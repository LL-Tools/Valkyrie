

module b17_C_gen_AntiSAT_k_256_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9805, n9807,
         n9808, n9809, n9810, n9811, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411;

  NOR2_X1 U11240 ( .A1(n15118), .A2(n15279), .ZN(n15072) );
  AND2_X1 U11241 ( .A1(n11063), .A2(n11051), .ZN(n13840) );
  NAND2_X1 U11242 ( .A1(n13170), .A2(n13169), .ZN(n13168) );
  NAND2_X1 U11243 ( .A1(n10921), .A2(n10920), .ZN(n13169) );
  CLKBUF_X1 U11244 ( .A(n10611), .Z(n11237) );
  NAND2_X2 U11245 ( .A1(n10896), .A2(n10895), .ZN(n11345) );
  BUF_X1 U11246 ( .A(n9811), .Z(n12683) );
  AND2_X1 U11247 ( .A1(n11709), .A2(n16412), .ZN(n12428) );
  AND2_X1 U11248 ( .A1(n12265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12113) );
  AND2_X1 U11249 ( .A1(n12300), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12414) );
  INV_X1 U11250 ( .A(n10197), .ZN(n12541) );
  AND2_X1 U11251 ( .A1(n11913), .A2(n11914), .ZN(n12809) );
  AND2_X1 U11252 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11915), .ZN(
        n12546) );
  CLKBUF_X1 U11253 ( .A(n10688), .Z(n11232) );
  INV_X1 U11254 ( .A(n12310), .ZN(n11783) );
  INV_X2 U11255 ( .A(n13852), .ZN(n17302) );
  CLKBUF_X1 U11256 ( .A(n10687), .Z(n10576) );
  CLKBUF_X2 U11257 ( .A(n10672), .Z(n13308) );
  CLKBUF_X2 U11258 ( .A(n10777), .Z(n12629) );
  INV_X2 U11259 ( .A(n17339), .ZN(n17223) );
  OR3_X1 U11260 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13851), .ZN(n13868) );
  NAND2_X2 U11261 ( .A1(n13848), .A2(n17041), .ZN(n17339) );
  NAND2_X2 U11262 ( .A1(n10301), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13901) );
  INV_X1 U11263 ( .A(n11861), .ZN(n11868) );
  NAND2_X1 U11264 ( .A1(n11696), .A2(n11695), .ZN(n11791) );
  CLKBUF_X2 U11265 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13837) );
  NAND3_X2 U11266 ( .A1(n10627), .A2(n10516), .A3(n10626), .ZN(n10694) );
  INV_X2 U11267 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10233) );
  AND2_X1 U11268 ( .A1(n10252), .A2(n13305), .ZN(n10672) );
  AND2_X1 U11269 ( .A1(n10527), .A2(n10529), .ZN(n10623) );
  AND2_X1 U11270 ( .A1(n10527), .A2(n13303), .ZN(n10733) );
  INV_X1 U11271 ( .A(n18867), .ZN(n9796) );
  INV_X1 U11272 ( .A(n9796), .ZN(n9797) );
  INV_X1 U11273 ( .A(n9796), .ZN(n9798) );
  BUF_X1 U11274 ( .A(n11198), .Z(n11625) );
  BUF_X1 U11275 ( .A(n11231), .Z(n11219) );
  NOR2_X1 U11276 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n15013), .ZN(n15083) );
  BUF_X1 U11277 ( .A(n11231), .Z(n9805) );
  AOI21_X1 U11278 ( .B1(n10256), .B2(n10258), .A(n9904), .ZN(n10253) );
  INV_X1 U11279 ( .A(n12403), .ZN(n13442) );
  INV_X2 U11280 ( .A(n17335), .ZN(n17349) );
  NOR2_X1 U11281 ( .A1(n12636), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12635) );
  INV_X2 U11283 ( .A(n12683), .ZN(n12404) );
  OR2_X1 U11284 ( .A1(n14773), .A2(n14767), .ZN(n14765) );
  INV_X1 U11286 ( .A(n13922), .ZN(n17329) );
  INV_X2 U11287 ( .A(n17275), .ZN(n9810) );
  NAND2_X1 U11288 ( .A1(n10203), .A2(n10202), .ZN(n10209) );
  INV_X2 U11289 ( .A(n13966), .ZN(n17176) );
  INV_X1 U11290 ( .A(n13146), .ZN(n21010) );
  INV_X2 U11291 ( .A(n11533), .ZN(n11531) );
  INV_X2 U11292 ( .A(n11531), .ZN(n14515) );
  INV_X1 U11293 ( .A(n15783), .ZN(n15789) );
  NAND2_X1 U11294 ( .A1(n12952), .A2(n11819), .ZN(n11817) );
  INV_X1 U11295 ( .A(n12581), .ZN(n12599) );
  AND2_X1 U11296 ( .A1(n14734), .A2(n14725), .ZN(n14727) );
  AND2_X1 U11297 ( .A1(n12790), .A2(n10350), .ZN(n14734) );
  XNOR2_X1 U11298 ( .A(n14692), .B(n14679), .ZN(n16120) );
  NOR2_X1 U11299 ( .A1(n15118), .A2(n15302), .ZN(n15102) );
  OAI21_X1 U11300 ( .B1(n19086), .B2(n15043), .A(n15211), .ZN(n15158) );
  NOR2_X1 U11301 ( .A1(n18226), .A2(n17932), .ZN(n17900) );
  NAND2_X1 U11302 ( .A1(n14143), .A2(n14126), .ZN(n14128) );
  OR2_X1 U11303 ( .A1(n14598), .A2(n11613), .ZN(n14578) );
  INV_X2 U11304 ( .A(n13868), .ZN(n17345) );
  INV_X1 U11305 ( .A(n18400), .ZN(n17445) );
  INV_X1 U11306 ( .A(n18028), .ZN(n17998) );
  INV_X1 U11307 ( .A(n17888), .ZN(n18226) );
  INV_X1 U11308 ( .A(n19268), .ZN(n19267) );
  INV_X1 U11309 ( .A(n20191), .ZN(n20184) );
  INV_X1 U11310 ( .A(n19250), .ZN(n13402) );
  INV_X1 U11311 ( .A(n17934), .ZN(n17893) );
  NAND2_X1 U11312 ( .A1(n17518), .A2(n18021), .ZN(n17938) );
  INV_X2 U11313 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18967) );
  OR2_X1 U11314 ( .A1(n9818), .A2(n15429), .ZN(n9799) );
  INV_X1 U11315 ( .A(n12604), .ZN(n11744) );
  NAND2_X2 U11316 ( .A1(n13446), .A2(n13447), .ZN(n13528) );
  AND2_X2 U11317 ( .A1(n13414), .A2(n13413), .ZN(n13447) );
  NAND2_X2 U11318 ( .A1(n11797), .A2(n12622), .ZN(n12813) );
  AND2_X1 U11319 ( .A1(n10529), .A2(n13305), .ZN(n9800) );
  AND2_X1 U11320 ( .A1(n10252), .A2(n13305), .ZN(n9801) );
  AND2_X1 U11321 ( .A1(n10252), .A2(n13305), .ZN(n9802) );
  AND2_X4 U11322 ( .A1(n13305), .A2(n10528), .ZN(n10723) );
  AND2_X4 U11323 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13305) );
  AND2_X2 U11324 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10528) );
  XNOR2_X2 U11325 ( .A(n12232), .B(n10512), .ZN(n14716) );
  NAND2_X2 U11326 ( .A1(n14723), .A2(n10514), .ZN(n12232) );
  INV_X2 U11327 ( .A(n13364), .ZN(n13401) );
  OR2_X2 U11328 ( .A1(n13364), .A2(n13367), .ZN(n13639) );
  OR3_X4 U11329 ( .A1(n18967), .A2(n18974), .A3(n13857), .ZN(n13933) );
  NAND2_X2 U11330 ( .A1(n11564), .A2(n12888), .ZN(n11657) );
  AND2_X2 U11331 ( .A1(n10365), .A2(n10364), .ZN(n11564) );
  NOR2_X2 U11333 ( .A1(n15140), .A2(n15331), .ZN(n15128) );
  AND2_X2 U11336 ( .A1(n10252), .A2(n14655), .ZN(n10842) );
  AND3_X2 U11337 ( .A1(n10287), .A2(n10289), .A3(n17990), .ZN(n17854) );
  BUF_X4 U11339 ( .A(n11231), .Z(n11627) );
  INV_X1 U11340 ( .A(n15618), .ZN(n13934) );
  XNOR2_X2 U11341 ( .A(n17550), .B(n15673), .ZN(n18019) );
  AND2_X1 U11342 ( .A1(n10527), .A2(n10529), .ZN(n9807) );
  AND2_X2 U11343 ( .A1(n11684), .A2(n13837), .ZN(n9808) );
  AND2_X1 U11344 ( .A1(n11684), .A2(n13837), .ZN(n12300) );
  NAND2_X4 U11345 ( .A1(n13849), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17293) );
  NOR2_X2 U11346 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17041) );
  NAND3_X2 U11347 ( .A1(n17042), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17144) );
  NAND2_X1 U11348 ( .A1(n10072), .A2(n9855), .ZN(n10326) );
  NAND2_X1 U11349 ( .A1(n9896), .A2(n10251), .ZN(n10250) );
  AOI211_X1 U11350 ( .C1(P2_EBX_REG_30__SCAN_IN), .C2(n19189), .A(n16122), .B(
        n16121), .ZN(n16123) );
  NAND2_X1 U11351 ( .A1(n15042), .A2(n14909), .ZN(n15044) );
  INV_X4 U11352 ( .A(n11531), .ZN(n15938) );
  AND2_X1 U11353 ( .A1(n10137), .A2(n13446), .ZN(n9823) );
  NAND2_X1 U11354 ( .A1(n10513), .A2(n11927), .ZN(n13104) );
  AND2_X1 U11355 ( .A1(n10312), .A2(n10311), .ZN(n17727) );
  AND2_X1 U11356 ( .A1(n10408), .A2(n10407), .ZN(n10513) );
  NOR2_X1 U11357 ( .A1(n15020), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15124) );
  OAI21_X1 U11358 ( .B1(n17738), .B2(n17722), .A(n15710), .ZN(n15711) );
  CLKBUF_X2 U11359 ( .A(n17822), .Z(n9847) );
  INV_X1 U11360 ( .A(n10209), .ZN(n15707) );
  AND2_X1 U11361 ( .A1(n10106), .A2(n13013), .ZN(n13006) );
  NAND2_X1 U11362 ( .A1(n13401), .A2(n9862), .ZN(n19478) );
  INV_X1 U11363 ( .A(n19576), .ZN(n9809) );
  CLKBUF_X1 U11364 ( .A(n13364), .Z(n13396) );
  XNOR2_X1 U11365 ( .A(n10134), .B(n11860), .ZN(n13363) );
  NAND2_X1 U11366 ( .A1(n20211), .A2(n10695), .ZN(n14318) );
  AOI21_X1 U11367 ( .B1(n19092), .B2(n19091), .A(n12675), .ZN(n19090) );
  OR2_X1 U11368 ( .A1(n14947), .A2(n14946), .ZN(n14964) );
  NOR2_X4 U11369 ( .A1(n18204), .A2(n18813), .ZN(n18261) );
  NAND2_X2 U11370 ( .A1(n13025), .A2(n13024), .ZN(n13023) );
  XNOR2_X1 U11371 ( .A(n12698), .B(n12696), .ZN(n12694) );
  AND2_X1 U11372 ( .A1(n11362), .A2(n11361), .ZN(n15783) );
  AND2_X1 U11373 ( .A1(n10275), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11888) );
  NOR2_X1 U11374 ( .A1(n16649), .A2(n19024), .ZN(n15572) );
  NAND2_X1 U11375 ( .A1(n16538), .A2(n15738), .ZN(n17811) );
  AND2_X1 U11376 ( .A1(n10218), .A2(n10217), .ZN(n18004) );
  AND2_X1 U11377 ( .A1(n10386), .A2(n11802), .ZN(n11820) );
  NOR2_X1 U11378 ( .A1(n17550), .A2(n17538), .ZN(n15746) );
  INV_X8 U11379 ( .A(n15043), .ZN(n15087) );
  NAND4_X2 U11380 ( .A1(n11799), .A2(n16440), .A3(n12956), .A4(n12622), .ZN(
        n16442) );
  BUF_X1 U11381 ( .A(n11817), .Z(n12936) );
  AOI211_X1 U11382 ( .C1(n15618), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n15608), .B(n15607), .ZN(n15736) );
  INV_X1 U11383 ( .A(n15684), .ZN(n17550) );
  AND3_X1 U11384 ( .A1(n11792), .A2(n19452), .A3(n11791), .ZN(n11799) );
  INV_X1 U11385 ( .A(n19452), .ZN(n10319) );
  INV_X2 U11386 ( .A(n13879), .ZN(n17324) );
  INV_X4 U11387 ( .A(n15538), .ZN(n15633) );
  CLKBUF_X3 U11388 ( .A(n11765), .Z(n9852) );
  INV_X2 U11389 ( .A(n12310), .ZN(n12299) );
  CLKBUF_X2 U11390 ( .A(n10646), .Z(n11632) );
  NOR2_X1 U11391 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18371), .ZN(n18715) );
  CLKBUF_X2 U11392 ( .A(n10734), .Z(n11229) );
  INV_X4 U11393 ( .A(n13901), .ZN(n17241) );
  CLKBUF_X2 U11394 ( .A(n10733), .Z(n11199) );
  INV_X1 U11395 ( .A(n13911), .ZN(n9813) );
  CLKBUF_X3 U11396 ( .A(n11198), .Z(n11144) );
  CLKBUF_X2 U11397 ( .A(n10800), .Z(n11230) );
  INV_X8 U11398 ( .A(n13933), .ZN(n17323) );
  INV_X4 U11399 ( .A(n11908), .ZN(n12265) );
  NOR2_X1 U11400 ( .A1(n12670), .A2(n19424), .ZN(n12667) );
  INV_X1 U11401 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18974) );
  INV_X1 U11402 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16415) );
  AOI21_X1 U11403 ( .B1(n14402), .B2(n15981), .A(n14401), .ZN(n14403) );
  XNOR2_X1 U11404 ( .A(n11654), .B(n11653), .ZN(n14106) );
  NAND2_X1 U11405 ( .A1(n14138), .A2(n10126), .ZN(n14408) );
  AND2_X1 U11406 ( .A1(n10368), .A2(n10366), .ZN(n14068) );
  AOI21_X1 U11407 ( .B1(n10125), .B2(n20298), .A(n14411), .ZN(n10124) );
  MUX2_X1 U11408 ( .A(n15420), .B(n9799), .S(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .Z(n15421) );
  AND2_X1 U11409 ( .A1(n11551), .A2(n10367), .ZN(n10366) );
  AOI21_X1 U11410 ( .B1(n15200), .B2(n15159), .A(n10239), .ZN(n15174) );
  NAND2_X1 U11411 ( .A1(n10326), .A2(n15008), .ZN(n15123) );
  AOI21_X1 U11412 ( .B1(n10283), .B2(n10282), .A(n10276), .ZN(n15213) );
  OR2_X1 U11413 ( .A1(n14392), .A2(n10377), .ZN(n14412) );
  NAND2_X1 U11414 ( .A1(n10241), .A2(n15158), .ZN(n15200) );
  OR2_X1 U11415 ( .A1(n15209), .A2(n15208), .ZN(n10241) );
  AND2_X1 U11416 ( .A1(n9824), .A2(n14404), .ZN(n14384) );
  NAND2_X1 U11417 ( .A1(n15196), .A2(n9892), .ZN(n15415) );
  NOR2_X1 U11418 ( .A1(n14716), .A2(n14715), .ZN(n14714) );
  NAND2_X1 U11419 ( .A1(n15480), .A2(n15435), .ZN(n15452) );
  AOI21_X1 U11420 ( .B1(n16530), .B2(n17934), .A(n16494), .ZN(n16495) );
  NAND2_X1 U11421 ( .A1(n13840), .A2(n13841), .ZN(n13844) );
  AOI21_X1 U11422 ( .B1(n16530), .B2(n18253), .A(n16529), .ZN(n16531) );
  AND2_X1 U11423 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15480) );
  OAI21_X1 U11424 ( .B1(n9896), .B2(n10244), .A(n10242), .ZN(n16224) );
  AND2_X1 U11425 ( .A1(n10271), .A2(n15495), .ZN(n9836) );
  INV_X1 U11426 ( .A(n13610), .ZN(n11012) );
  NAND2_X1 U11427 ( .A1(n10054), .A2(n10055), .ZN(n10141) );
  AND2_X1 U11428 ( .A1(n10056), .A2(n10057), .ZN(n10054) );
  OR2_X1 U11429 ( .A1(n16290), .A2(n16382), .ZN(n10075) );
  AOI21_X1 U11430 ( .B1(n10272), .B2(n16382), .A(n21411), .ZN(n10179) );
  INV_X1 U11431 ( .A(n10236), .ZN(n10142) );
  NAND2_X1 U11432 ( .A1(n10059), .A2(n10058), .ZN(n14873) );
  OR2_X1 U11433 ( .A1(n15939), .A2(n11535), .ZN(n14497) );
  INV_X1 U11434 ( .A(n16547), .ZN(n17676) );
  INV_X1 U11435 ( .A(n9826), .ZN(n10258) );
  AOI21_X1 U11436 ( .B1(n9826), .B2(n10257), .A(n9905), .ZN(n10256) );
  OR2_X1 U11437 ( .A1(n13674), .A2(n13673), .ZN(n10059) );
  AND2_X1 U11438 ( .A1(n11537), .A2(n9918), .ZN(n10148) );
  OR2_X1 U11439 ( .A1(n9833), .A2(n9834), .ZN(n16126) );
  AND2_X1 U11440 ( .A1(n9913), .A2(n11523), .ZN(n9826) );
  OR2_X1 U11441 ( .A1(n14515), .A2(n11536), .ZN(n14488) );
  OR2_X1 U11442 ( .A1(n15968), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11522) );
  OR2_X1 U11443 ( .A1(n9857), .A2(n15082), .ZN(n10070) );
  AND2_X1 U11444 ( .A1(n17707), .A2(n10506), .ZN(n15717) );
  AND2_X1 U11445 ( .A1(n13678), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15049) );
  NAND2_X1 U11446 ( .A1(n9856), .A2(n13451), .ZN(n13524) );
  AND2_X1 U11447 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  AND2_X1 U11448 ( .A1(n10324), .A2(n15008), .ZN(n9857) );
  NAND2_X1 U11449 ( .A1(n10081), .A2(n10086), .ZN(n10089) );
  XNOR2_X1 U11450 ( .A(n10434), .B(n12632), .ZN(n14527) );
  NAND3_X1 U11451 ( .A1(n17727), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17720), .ZN(n15716) );
  AND2_X1 U11452 ( .A1(n10325), .A2(n15113), .ZN(n10324) );
  AND2_X1 U11453 ( .A1(n12794), .A2(n12793), .ZN(n15354) );
  AND2_X1 U11454 ( .A1(n13528), .A2(n10085), .ZN(n10081) );
  NAND2_X1 U11455 ( .A1(n9823), .A2(n13667), .ZN(n14908) );
  INV_X1 U11456 ( .A(n12631), .ZN(n10434) );
  INV_X1 U11457 ( .A(n9823), .ZN(n10087) );
  AND2_X1 U11458 ( .A1(n10940), .A2(n10939), .ZN(n13345) );
  NAND2_X1 U11459 ( .A1(n13218), .A2(n10890), .ZN(n13170) );
  NOR2_X1 U11460 ( .A1(n17770), .A2(n15712), .ZN(n17721) );
  AND2_X1 U11461 ( .A1(n20161), .A2(n13495), .ZN(n20191) );
  NOR2_X1 U11462 ( .A1(n14841), .A2(n12769), .ZN(n12794) );
  OR2_X1 U11463 ( .A1(n10144), .A2(n10328), .ZN(n10066) );
  AND2_X1 U11464 ( .A1(n9985), .A2(n13666), .ZN(n13667) );
  INV_X1 U11465 ( .A(n15711), .ZN(n15712) );
  NAND2_X1 U11466 ( .A1(n10206), .A2(n10204), .ZN(n17770) );
  AND2_X1 U11467 ( .A1(n13184), .A2(n10347), .ZN(n13467) );
  OR2_X1 U11468 ( .A1(n9829), .A2(n9830), .ZN(n16189) );
  OR2_X1 U11469 ( .A1(n10207), .A2(n17933), .ZN(n10206) );
  AND2_X1 U11470 ( .A1(n16174), .A2(n15087), .ZN(n15020) );
  AND2_X1 U11471 ( .A1(n13087), .A2(n10474), .ZN(n10473) );
  AND2_X1 U11472 ( .A1(n10210), .A2(n18152), .ZN(n10207) );
  NAND2_X1 U11473 ( .A1(n10878), .A2(n10877), .ZN(n13087) );
  AOI22_X1 U11474 ( .A1(n17889), .A2(n18226), .B1(n18000), .B2(n18224), .ZN(
        n17920) );
  OR2_X1 U11475 ( .A1(n9885), .A2(n13109), .ZN(n13178) );
  AND3_X1 U11476 ( .A1(n13406), .A2(n13405), .A3(n9900), .ZN(n13407) );
  AND2_X1 U11477 ( .A1(n15706), .A2(n9945), .ZN(n10210) );
  NOR2_X1 U11478 ( .A1(n13395), .A2(n13394), .ZN(n13408) );
  OR2_X1 U11479 ( .A1(n13654), .A2(n13404), .ZN(n9900) );
  NOR2_X2 U11480 ( .A1(n15006), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15010) );
  OR2_X1 U11481 ( .A1(n15000), .A2(n14999), .ZN(n15006) );
  NAND2_X1 U11482 ( .A1(n13401), .A2(n13391), .ZN(n19624) );
  NAND2_X1 U11483 ( .A1(n13401), .A2(n13400), .ZN(n19576) );
  OR2_X1 U11484 ( .A1(n13403), .A2(n19250), .ZN(n19786) );
  AND2_X1 U11485 ( .A1(n13364), .A2(n13279), .ZN(n14880) );
  OR2_X1 U11486 ( .A1(n13078), .A2(n10887), .ZN(n13079) );
  OR2_X1 U11487 ( .A1(n11871), .A2(n11870), .ZN(n10396) );
  NAND2_X1 U11488 ( .A1(n10382), .A2(n11464), .ZN(n13094) );
  OAI21_X1 U11489 ( .B1(n13364), .B2(n10101), .A(n10103), .ZN(n13013) );
  NAND2_X1 U11490 ( .A1(n11605), .A2(n11604), .ZN(n20325) );
  OR2_X1 U11491 ( .A1(n13364), .A2(n13389), .ZN(n19542) );
  NAND2_X1 U11492 ( .A1(n12783), .A2(n12784), .ZN(n15000) );
  NOR2_X1 U11493 ( .A1(n13402), .A2(n13399), .ZN(n13391) );
  NOR2_X1 U11494 ( .A1(n13374), .A2(n13228), .ZN(n9862) );
  NAND2_X1 U11495 ( .A1(n12782), .A2(n15012), .ZN(n12783) );
  OR2_X1 U11496 ( .A1(n13374), .A2(n13373), .ZN(n13389) );
  AND2_X1 U11497 ( .A1(n14977), .A2(n14976), .ZN(n19096) );
  OR2_X1 U11498 ( .A1(n13339), .A2(n11488), .ZN(n10382) );
  AND2_X1 U11499 ( .A1(n14614), .A2(n14608), .ZN(n16055) );
  XNOR2_X1 U11500 ( .A(n13325), .B(n20477), .ZN(n20594) );
  XNOR2_X1 U11501 ( .A(n10859), .B(n10860), .ZN(n10873) );
  OR2_X1 U11502 ( .A1(n12691), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U11503 ( .A1(n11876), .A2(n11875), .ZN(n13792) );
  OAI21_X2 U11504 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19004), .A(n16650), 
        .ZN(n18028) );
  NOR2_X2 U11505 ( .A1(n19012), .A2(n16650), .ZN(n18021) );
  NOR2_X1 U11506 ( .A1(n19076), .A2(n19090), .ZN(n19075) );
  OR2_X1 U11507 ( .A1(n10859), .A2(n10860), .ZN(n10861) );
  BUF_X1 U11508 ( .A(n13363), .Z(n13374) );
  NAND2_X1 U11509 ( .A1(n11602), .A2(n15800), .ZN(n14614) );
  OR2_X1 U11510 ( .A1(n14975), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14976) );
  CLKBUF_X3 U11511 ( .A(n12675), .Z(n9835) );
  NAND2_X1 U11512 ( .A1(n10134), .A2(n11884), .ZN(n10346) );
  NOR2_X1 U11513 ( .A1(n20483), .A2(n20357), .ZN(n20864) );
  AND2_X1 U11514 ( .A1(n11571), .A2(n20107), .ZN(n11602) );
  NAND2_X1 U11515 ( .A1(n13200), .A2(n12839), .ZN(n11876) );
  NOR2_X1 U11516 ( .A1(n20483), .A2(n20266), .ZN(n20907) );
  NAND2_X1 U11517 ( .A1(n19005), .A2(n18805), .ZN(n16650) );
  NOR2_X1 U11518 ( .A1(n20483), .A2(n20376), .ZN(n20898) );
  NAND2_X1 U11519 ( .A1(n10261), .A2(n10833), .ZN(n10879) );
  NOR2_X1 U11520 ( .A1(n20483), .A2(n20367), .ZN(n20892) );
  NAND2_X1 U11521 ( .A1(n10073), .A2(n10176), .ZN(n10134) );
  CLKBUF_X2 U11522 ( .A(n12868), .Z(n19250) );
  INV_X1 U11523 ( .A(n10090), .ZN(n13200) );
  NOR2_X2 U11524 ( .A1(n19446), .A2(n19826), .ZN(n19447) );
  NOR2_X2 U11525 ( .A1(n19440), .A2(n19826), .ZN(n19441) );
  NOR2_X2 U11526 ( .A1(n19388), .A2(n19826), .ZN(n13231) );
  NOR2_X2 U11527 ( .A1(n19386), .A2(n19826), .ZN(n13210) );
  AND2_X1 U11528 ( .A1(n12704), .A2(n10355), .ZN(n10354) );
  NAND2_X1 U11529 ( .A1(n10163), .A2(n10162), .ZN(n20161) );
  OR2_X1 U11530 ( .A1(n13617), .A2(n13616), .ZN(n13735) );
  OAI22_X1 U11531 ( .A1(n19034), .A2(n15242), .B1(n15053), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U11532 ( .A1(n11873), .A2(n11872), .ZN(n10091) );
  OR2_X1 U11533 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  NAND3_X1 U11534 ( .A1(n11848), .A2(n11847), .A3(n11846), .ZN(n11872) );
  CLKBUF_X2 U11535 ( .A(n11891), .Z(n14685) );
  NOR2_X2 U11536 ( .A1(n15763), .A2(n15768), .ZN(n18353) );
  AOI21_X1 U11537 ( .B1(n11891), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11896), .ZN(n12696) );
  OR2_X1 U11538 ( .A1(n13360), .A2(n13359), .ZN(n16084) );
  NAND2_X2 U11539 ( .A1(n17589), .A2(n18848), .ZN(n17655) );
  OAI21_X1 U11540 ( .B1(n11839), .B2(n10502), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11847) );
  NOR2_X1 U11541 ( .A1(n15572), .A2(n15561), .ZN(n16665) );
  XNOR2_X1 U11542 ( .A(n15689), .B(n15688), .ZN(n17995) );
  NAND2_X1 U11543 ( .A1(n14915), .A2(n14913), .ZN(n14925) );
  BUF_X2 U11544 ( .A(n11892), .Z(n9986) );
  NAND2_X1 U11545 ( .A1(n10315), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10314) );
  NAND2_X1 U11546 ( .A1(n14915), .A2(n12404), .ZN(n15012) );
  AND3_X1 U11547 ( .A1(n10191), .A2(n10194), .A3(n13526), .ZN(n14917) );
  AND2_X1 U11548 ( .A1(n11796), .A2(n12962), .ZN(n11836) );
  NOR2_X1 U11549 ( .A1(n13448), .A2(n10195), .ZN(n10194) );
  AND2_X2 U11550 ( .A1(n12397), .A2(n11818), .ZN(n12965) );
  AND3_X1 U11551 ( .A1(n10780), .A2(n11596), .A3(n10779), .ZN(n10782) );
  INV_X1 U11552 ( .A(n9837), .ZN(n11807) );
  NOR2_X1 U11553 ( .A1(n15736), .A2(n15691), .ZN(n15694) );
  NAND2_X1 U11554 ( .A1(n12404), .A2(n10493), .ZN(n12577) );
  NOR2_X1 U11555 ( .A1(n17445), .A2(n18372), .ZN(n15564) );
  AND2_X1 U11556 ( .A1(n16442), .A2(n12931), .ZN(n9837) );
  NAND2_X1 U11557 ( .A1(n11745), .A2(n11744), .ZN(n12955) );
  NOR4_X2 U11558 ( .A1(n16997), .A2(n15765), .A3(n18393), .A4(n15552), .ZN(
        n17590) );
  INV_X1 U11559 ( .A(n12936), .ZN(n12364) );
  AND2_X2 U11560 ( .A1(n12553), .A2(n12552), .ZN(n15043) );
  NOR2_X1 U11561 ( .A1(n13138), .A2(n10757), .ZN(n10781) );
  INV_X1 U11562 ( .A(n11795), .ZN(n12444) );
  NAND2_X1 U11563 ( .A1(n10671), .A2(n10774), .ZN(n10754) );
  INV_X1 U11564 ( .A(n12354), .ZN(n14671) );
  OR2_X1 U11565 ( .A1(n12423), .A2(n12422), .ZN(n12684) );
  OR2_X1 U11566 ( .A1(n12505), .A2(n12506), .ZN(n13443) );
  OR2_X1 U11567 ( .A1(n12468), .A2(n12467), .ZN(n12847) );
  NAND2_X1 U11568 ( .A1(n11868), .A2(n11791), .ZN(n11795) );
  OR2_X1 U11569 ( .A1(n12485), .A2(n12484), .ZN(n12849) );
  NAND2_X1 U11570 ( .A1(n11453), .A2(n11584), .ZN(n11449) );
  AND2_X1 U11571 ( .A1(n10670), .A2(n10695), .ZN(n10774) );
  INV_X2 U11572 ( .A(n11791), .ZN(n9811) );
  NOR2_X1 U11573 ( .A1(n13496), .A2(n13599), .ZN(n12888) );
  INV_X1 U11574 ( .A(n13157), .ZN(n13579) );
  NOR2_X1 U11575 ( .A1(n10318), .A2(n10317), .ZN(n10316) );
  INV_X1 U11576 ( .A(n13599), .ZN(n10762) );
  OR2_X2 U11577 ( .A1(n16598), .A2(n16551), .ZN(n16601) );
  OR2_X1 U11578 ( .A1(n10821), .A2(n10820), .ZN(n11524) );
  OR2_X1 U11579 ( .A1(n10682), .A2(n10681), .ZN(n13589) );
  AND2_X1 U11580 ( .A1(n10515), .A2(n10517), .ZN(n13157) );
  NAND2_X1 U11581 ( .A1(n11788), .A2(n11787), .ZN(n19439) );
  NAND3_X1 U11582 ( .A1(n11736), .A2(n11735), .A3(n11734), .ZN(n11743) );
  AND4_X1 U11583 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10741) );
  AND4_X1 U11584 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(
        n10716) );
  AND4_X1 U11585 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10717) );
  AND4_X1 U11586 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10740) );
  NAND4_X1 U11587 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10668) );
  AND4_X1 U11588 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10518) );
  AND4_X1 U11589 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n10659) );
  AND4_X1 U11590 ( .A1(n10645), .A2(n10644), .A3(n10643), .A4(n10642), .ZN(
        n10658) );
  AND4_X1 U11591 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10657) );
  AND4_X1 U11592 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10715) );
  AND4_X1 U11593 ( .A1(n10702), .A2(n10701), .A3(n10700), .A4(n10699), .ZN(
        n10718) );
  AND4_X1 U11594 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10742) );
  AND3_X1 U11595 ( .A1(n11733), .A2(n16412), .A3(n11732), .ZN(n11736) );
  AND4_X1 U11596 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10616) );
  NAND2_X1 U11597 ( .A1(n12666), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12663) );
  AND2_X1 U11598 ( .A1(n11737), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11738) );
  AND2_X2 U11600 ( .A1(n12799), .A2(n19034), .ZN(n19412) );
  NAND2_X2 U11601 ( .A1(n20036), .A2(n19978), .ZN(n20042) );
  INV_X2 U11602 ( .A(n16634), .ZN(U215) );
  NAND2_X2 U11603 ( .A1(n18999), .A2(n18883), .ZN(n18935) );
  CLKBUF_X3 U11605 ( .A(n11721), .Z(n9848) );
  BUF_X2 U11606 ( .A(n10842), .Z(n11624) );
  BUF_X2 U11607 ( .A(n10623), .Z(n11626) );
  INV_X1 U11608 ( .A(n18956), .ZN(n18867) );
  CLKBUF_X1 U11609 ( .A(n10651), .Z(n11634) );
  BUF_X4 U11610 ( .A(n10723), .Z(n10698) );
  INV_X2 U11611 ( .A(n16637), .ZN(n16639) );
  AND2_X2 U11612 ( .A1(n13303), .A2(n10526), .ZN(n11198) );
  INV_X2 U11613 ( .A(n21023), .ZN(n20972) );
  NOR2_X1 U11614 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  AND2_X1 U11615 ( .A1(n10520), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U11616 ( .A1(n18974), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13855) );
  AND3_X4 U11617 ( .A1(n13801), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11709) );
  NAND2_X2 U11618 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13851) );
  NOR2_X2 U11619 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14655) );
  NAND2_X1 U11620 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18828) );
  INV_X1 U11621 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18988) );
  NOR2_X1 U11622 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11684) );
  NAND2_X2 U11623 ( .A1(n13176), .A2(n13175), .ZN(n13174) );
  AND2_X1 U11624 ( .A1(n9817), .A2(n13681), .ZN(n9814) );
  NAND4_X1 U11625 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n9815) );
  AND2_X1 U11626 ( .A1(n12403), .A2(n19439), .ZN(n9816) );
  AOI21_X1 U11627 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(n9817) );
  AND2_X1 U11628 ( .A1(n15430), .A2(n15419), .ZN(n9818) );
  AOI21_X1 U11629 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(n13680) );
  NAND2_X1 U11630 ( .A1(n10254), .A2(n10253), .ZN(n9819) );
  NAND2_X1 U11631 ( .A1(n11542), .A2(n15938), .ZN(n9820) );
  NAND2_X1 U11632 ( .A1(n10765), .A2(n10764), .ZN(n9821) );
  NAND2_X1 U11633 ( .A1(n10254), .A2(n10253), .ZN(n14518) );
  OAI21_X2 U11634 ( .B1(n10769), .B2(n10760), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10765) );
  NOR2_X2 U11635 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10529) );
  OR2_X1 U11636 ( .A1(n16290), .A2(n16382), .ZN(n9822) );
  XNOR2_X1 U11637 ( .A(n12635), .B(n11616), .ZN(n10369) );
  NOR2_X1 U11638 ( .A1(n14548), .A2(n14566), .ZN(n9824) );
  AOI21_X2 U11639 ( .B1(n15070), .B2(n10327), .A(n15034), .ZN(n15041) );
  AND2_X1 U11640 ( .A1(n10373), .A2(n10370), .ZN(n9825) );
  NOR3_X2 U11641 ( .A1(n10372), .A2(n10378), .A3(n10371), .ZN(n10370) );
  NAND2_X2 U11642 ( .A1(n12127), .A2(n12126), .ZN(n12162) );
  XNOR2_X2 U11643 ( .A(n12162), .B(n12186), .ZN(n14742) );
  NOR2_X1 U11644 ( .A1(n12162), .A2(n12163), .ZN(n12164) );
  INV_X1 U11645 ( .A(n14189), .ZN(n11264) );
  AOI211_X1 U11646 ( .C1(n10912), .C2(n21346), .A(n20716), .B(n20650), .ZN(
        n14653) );
  NAND2_X1 U11647 ( .A1(n9822), .A2(n10074), .ZN(n9827) );
  NAND2_X1 U11648 ( .A1(n10075), .A2(n10074), .ZN(n10271) );
  NOR2_X2 U11649 ( .A1(n9828), .A2(n15129), .ZN(n15103) );
  NAND2_X1 U11650 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U11651 ( .A1(n16112), .A2(n9835), .ZN(n9829) );
  AND2_X1 U11652 ( .A1(n9831), .A2(n16199), .ZN(n9830) );
  INV_X1 U11653 ( .A(n9835), .ZN(n9831) );
  NOR2_X1 U11655 ( .A1(n16152), .A2(n9835), .ZN(n9833) );
  AND2_X1 U11656 ( .A1(n9831), .A2(n16145), .ZN(n9834) );
  NAND2_X2 U11658 ( .A1(n14906), .A2(n14907), .ZN(n15042) );
  OR2_X1 U11659 ( .A1(n14392), .A2(n10377), .ZN(n9838) );
  AND2_X2 U11660 ( .A1(n10123), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13303) );
  NOR2_X1 U11661 ( .A1(n12636), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9840) );
  AND2_X4 U11662 ( .A1(n10529), .A2(n13305), .ZN(n10651) );
  NAND2_X1 U11663 ( .A1(n10473), .A2(n10472), .ZN(n13218) );
  XNOR2_X1 U11664 ( .A(n11527), .B(n10988), .ZN(n11515) );
  NAND2_X1 U11665 ( .A1(n10968), .A2(n10157), .ZN(n11527) );
  INV_X4 U11666 ( .A(n11908), .ZN(n11778) );
  OAI21_X2 U11667 ( .B1(n14716), .B2(n10097), .A(n10096), .ZN(n12258) );
  NAND4_X4 U11668 ( .A1(n10715), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n13599) );
  NAND2_X1 U11669 ( .A1(n15977), .A2(n9844), .ZN(n9841) );
  AND2_X2 U11670 ( .A1(n9841), .A2(n9842), .ZN(n15970) );
  OR2_X1 U11671 ( .A1(n9843), .A2(n13556), .ZN(n9842) );
  INV_X1 U11672 ( .A(n11514), .ZN(n9843) );
  AND2_X1 U11673 ( .A1(n11504), .A2(n11514), .ZN(n9844) );
  NOR2_X2 U11674 ( .A1(n9845), .A2(n10694), .ZN(n10669) );
  NOR2_X1 U11675 ( .A1(n15129), .A2(n15131), .ZN(n15115) );
  AND3_X1 U11676 ( .A1(n10619), .A2(n10618), .A3(n10617), .ZN(n10621) );
  INV_X4 U11678 ( .A(n9845), .ZN(n14043) );
  NAND2_X1 U11679 ( .A1(n9819), .A2(n11532), .ZN(n15960) );
  NAND2_X2 U11680 ( .A1(n13844), .A2(n11063), .ZN(n14246) );
  NAND2_X1 U11681 ( .A1(n20292), .A2(n11496), .ZN(n15979) );
  NAND2_X1 U11682 ( .A1(n20294), .A2(n20293), .ZN(n20292) );
  OAI21_X1 U11683 ( .B1(n11542), .B2(n10376), .A(n10149), .ZN(n14404) );
  OR2_X1 U11684 ( .A1(n10743), .A2(n10696), .ZN(n15797) );
  NAND2_X1 U11685 ( .A1(n12965), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9846) );
  NAND2_X2 U11686 ( .A1(n14154), .A2(n14153), .ZN(n14137) );
  AND2_X2 U11687 ( .A1(n11264), .A2(n10477), .ZN(n14154) );
  NAND2_X1 U11688 ( .A1(n13557), .A2(n13556), .ZN(n13555) );
  NOR2_X2 U11689 ( .A1(n12777), .A2(n15148), .ZN(n15138) );
  AND2_X1 U11690 ( .A1(n13303), .A2(n10526), .ZN(n9849) );
  XNOR2_X1 U11691 ( .A(n11484), .B(n20336), .ZN(n13248) );
  OAI21_X2 U11692 ( .B1(n10873), .B2(n11465), .A(n10861), .ZN(n10864) );
  NAND2_X1 U11693 ( .A1(n20346), .A2(n11475), .ZN(n11484) );
  XNOR2_X1 U11694 ( .A(n12695), .B(n12694), .ZN(n9850) );
  XNOR2_X1 U11695 ( .A(n12695), .B(n12694), .ZN(n9851) );
  NAND2_X1 U11696 ( .A1(n13132), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20346) );
  XNOR2_X1 U11697 ( .A(n13093), .B(n11473), .ZN(n13132) );
  AND2_X2 U11698 ( .A1(n10526), .A2(n10252), .ZN(n10646) );
  NOR2_X2 U11699 ( .A1(n12647), .A2(n15167), .ZN(n12648) );
  XNOR2_X2 U11700 ( .A(n11650), .B(n12626), .ZN(n14062) );
  NOR2_X4 U11701 ( .A1(n14137), .A2(n10486), .ZN(n11650) );
  NOR2_X2 U11703 ( .A1(n12665), .A2(n16299), .ZN(n12666) );
  NOR2_X2 U11704 ( .A1(n12663), .A2(n10338), .ZN(n12658) );
  NOR2_X2 U11705 ( .A1(n12655), .A2(n12672), .ZN(n12653) );
  NAND3_X1 U11706 ( .A1(n13594), .A2(n13599), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11349) );
  OR2_X1 U11707 ( .A1(n13594), .A2(n21012), .ZN(n10895) );
  NAND3_X1 U11708 ( .A1(n11868), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13442), 
        .ZN(n12227) );
  NAND2_X1 U11709 ( .A1(n10220), .A2(n10219), .ZN(n10218) );
  NAND2_X1 U11710 ( .A1(n17550), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10219) );
  NAND2_X1 U11711 ( .A1(n10769), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10784) );
  NOR2_X1 U11712 ( .A1(n12164), .A2(n12187), .ZN(n10400) );
  NAND2_X1 U11713 ( .A1(n10275), .A2(n9941), .ZN(n11806) );
  AND2_X1 U11714 ( .A1(n9815), .A2(n9946), .ZN(n10137) );
  NAND4_X1 U11715 ( .A1(n11802), .A2(n14671), .A3(n11819), .A4(n11801), .ZN(
        n12713) );
  NOR2_X1 U11716 ( .A1(n12956), .A2(n11817), .ZN(n11818) );
  NAND2_X1 U11717 ( .A1(n9811), .A2(n11868), .ZN(n11808) );
  INV_X1 U11718 ( .A(n14449), .ZN(n10372) );
  NAND2_X1 U11719 ( .A1(n14404), .A2(n11543), .ZN(n11544) );
  NAND2_X1 U11720 ( .A1(n10837), .A2(n10836), .ZN(n10859) );
  OAI21_X1 U11721 ( .B1(n10883), .B2(n10263), .A(n9901), .ZN(n10837) );
  INV_X1 U11722 ( .A(n10833), .ZN(n10263) );
  NAND2_X1 U11723 ( .A1(n10909), .A2(n14650), .ZN(n10943) );
  INV_X1 U11724 ( .A(n12227), .ZN(n12253) );
  NAND2_X1 U11725 ( .A1(n14742), .A2(n14743), .ZN(n10402) );
  NOR2_X1 U11726 ( .A1(n9935), .A2(n10109), .ZN(n10108) );
  INV_X1 U11727 ( .A(n13622), .ZN(n10109) );
  NOR2_X1 U11728 ( .A1(n9884), .A2(n10333), .ZN(n10332) );
  NAND2_X1 U11729 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10333) );
  INV_X1 U11730 ( .A(n13297), .ZN(n10349) );
  INV_X1 U11731 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U11732 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10341) );
  INV_X1 U11733 ( .A(n14741), .ZN(n10352) );
  NOR2_X1 U11734 ( .A1(n10067), .A2(n15363), .ZN(n10062) );
  NOR2_X1 U11735 ( .A1(n15175), .A2(n14995), .ZN(n10329) );
  INV_X1 U11736 ( .A(n13729), .ZN(n10356) );
  INV_X1 U11737 ( .A(n12713), .ZN(n14680) );
  NAND2_X1 U11738 ( .A1(n9915), .A2(n10273), .ZN(n10272) );
  INV_X1 U11739 ( .A(n15044), .ZN(n10273) );
  NOR2_X1 U11740 ( .A1(n15047), .A2(n9906), .ZN(n16290) );
  INV_X1 U11741 ( .A(n13459), .ZN(n10085) );
  AND2_X1 U11742 ( .A1(n12370), .A2(n12824), .ZN(n12371) );
  NOR2_X1 U11743 ( .A1(n19958), .A2(n14670), .ZN(n12978) );
  NAND2_X1 U11744 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18967), .ZN(
        n13856) );
  INV_X1 U11745 ( .A(n13965), .ZN(n15609) );
  AND2_X1 U11746 ( .A1(n10309), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10307) );
  INV_X1 U11747 ( .A(n17518), .ZN(n15738) );
  INV_X1 U11748 ( .A(n17964), .ZN(n10214) );
  AND2_X1 U11749 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15692), .ZN(
        n15693) );
  XNOR2_X1 U11750 ( .A(n15640), .B(n15684), .ZN(n15685) );
  NOR2_X1 U11751 ( .A1(n13488), .A2(n20317), .ZN(n10162) );
  NOR2_X1 U11752 ( .A1(n13507), .A2(n10762), .ZN(n13502) );
  NAND2_X1 U11753 ( .A1(n20161), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13507) );
  AND4_X1 U11754 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10739) );
  NOR2_X1 U11755 ( .A1(n11301), .A2(n10133), .ZN(n10132) );
  AOI21_X1 U11756 ( .B1(n10872), .B2(n11042), .A(n10476), .ZN(n10475) );
  INV_X1 U11757 ( .A(n10890), .ZN(n10476) );
  NAND2_X1 U11758 ( .A1(n11476), .A2(n10872), .ZN(n10472) );
  INV_X1 U11759 ( .A(n15829), .ZN(n20107) );
  AND3_X1 U11760 ( .A1(n11525), .A2(n10260), .A3(n11524), .ZN(n11526) );
  NAND2_X1 U11761 ( .A1(n10856), .A2(n21012), .ZN(n10858) );
  OAI21_X1 U11762 ( .B1(n10170), .B2(n11359), .A(n9910), .ZN(n11361) );
  AND2_X1 U11763 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  INV_X1 U11764 ( .A(n14812), .ZN(n10456) );
  AND2_X1 U11765 ( .A1(n13467), .A2(n13466), .ZN(n13478) );
  NOR2_X1 U11766 ( .A1(n11907), .A2(n10410), .ZN(n10409) );
  INV_X1 U11767 ( .A(n11904), .ZN(n10410) );
  INV_X1 U11768 ( .A(n16471), .ZN(n12992) );
  AND2_X1 U11769 ( .A1(n11903), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U11770 ( .A1(n11902), .A2(n10105), .ZN(n10104) );
  NAND2_X1 U11771 ( .A1(n15026), .A2(n10190), .ZN(n10143) );
  AND2_X1 U11772 ( .A1(n20065), .A2(n20072), .ZN(n20053) );
  INV_X1 U11773 ( .A(n15609), .ZN(n17326) );
  AOI21_X1 U11774 ( .B1(n16666), .B2(n15571), .A(n10122), .ZN(n15856) );
  NAND2_X1 U11775 ( .A1(n18799), .A2(n19013), .ZN(n10122) );
  XNOR2_X1 U11776 ( .A(n15685), .B(n18328), .ZN(n18005) );
  NAND2_X1 U11777 ( .A1(n15683), .A2(n18019), .ZN(n10220) );
  NAND2_X1 U11778 ( .A1(n15858), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18027) );
  INV_X1 U11779 ( .A(n20316), .ZN(n20344) );
  NAND2_X1 U11780 ( .A1(n12925), .A2(n12830), .ZN(n12835) );
  INV_X1 U11781 ( .A(n16294), .ZN(n19416) );
  AND4_X1 U11782 ( .A1(n14885), .A2(n14884), .A3(n14883), .A4(n14882), .ZN(
        n14902) );
  NAND2_X1 U11783 ( .A1(n11315), .A2(n11314), .ZN(n11322) );
  INV_X1 U11784 ( .A(n11820), .ZN(n11803) );
  NAND2_X1 U11785 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10120) );
  OR2_X1 U11786 ( .A1(n10978), .A2(n10977), .ZN(n11517) );
  NAND2_X1 U11787 ( .A1(n11449), .A2(n10416), .ZN(n10415) );
  NAND2_X1 U11788 ( .A1(n10153), .A2(n10753), .ZN(n10152) );
  NAND2_X1 U11789 ( .A1(n11798), .A2(n12939), .ZN(n11843) );
  NAND2_X1 U11790 ( .A1(n12955), .A2(n12957), .ZN(n11837) );
  INV_X1 U11791 ( .A(n15092), .ZN(n10322) );
  OAI21_X1 U11792 ( .B1(n9986), .B2(n13182), .A(n12726), .ZN(n10004) );
  NAND2_X1 U11793 ( .A1(n13664), .A2(n9898), .ZN(n9985) );
  AND4_X1 U11794 ( .A1(n13647), .A2(n13646), .A3(n13645), .A4(n13644), .ZN(
        n13664) );
  OAI21_X1 U11795 ( .B1(n11892), .B2(n11895), .A(n11893), .ZN(n9988) );
  AOI21_X1 U11796 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18369), .A(
        n13954), .ZN(n15567) );
  INV_X1 U11797 ( .A(n13703), .ZN(n11011) );
  NAND2_X1 U11798 ( .A1(n10489), .A2(n10487), .ZN(n10486) );
  NOR2_X1 U11799 ( .A1(n11310), .A2(n10490), .ZN(n10489) );
  INV_X1 U11800 ( .A(n14125), .ZN(n10490) );
  AND2_X1 U11801 ( .A1(n11275), .A2(n9956), .ZN(n10479) );
  NAND2_X1 U11802 ( .A1(n11248), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11261) );
  NAND2_X1 U11803 ( .A1(n9943), .A2(n10129), .ZN(n10128) );
  INV_X1 U11804 ( .A(n10130), .ZN(n10129) );
  NOR2_X1 U11805 ( .A1(n14271), .A2(n10482), .ZN(n10481) );
  INV_X1 U11806 ( .A(n9955), .ZN(n10482) );
  OR2_X1 U11807 ( .A1(n10131), .A2(n14289), .ZN(n10130) );
  INV_X1 U11808 ( .A(n14281), .ZN(n10131) );
  INV_X1 U11809 ( .A(n11646), .ZN(n11297) );
  NAND2_X1 U11810 ( .A1(n14656), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11646) );
  INV_X1 U11811 ( .A(n10375), .ZN(n10371) );
  NAND2_X1 U11812 ( .A1(n11531), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10375) );
  NAND2_X1 U11813 ( .A1(n14192), .A2(n14205), .ZN(n10423) );
  NAND2_X1 U11814 ( .A1(n14450), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10381) );
  NOR2_X1 U11815 ( .A1(n10421), .A2(n14294), .ZN(n10420) );
  INV_X1 U11816 ( .A(n14305), .ZN(n10421) );
  NAND2_X1 U11817 ( .A1(n15915), .A2(n13804), .ZN(n10427) );
  INV_X1 U11818 ( .A(n11449), .ZN(n11444) );
  INV_X1 U11819 ( .A(n11453), .ZN(n10777) );
  OR2_X1 U11820 ( .A1(n10831), .A2(n10830), .ZN(n11466) );
  NAND2_X1 U11821 ( .A1(n10854), .A2(n10853), .ZN(n20385) );
  NOR2_X1 U11822 ( .A1(n10806), .A2(n10805), .ZN(n11477) );
  AND2_X1 U11823 ( .A1(n10891), .A2(n20886), .ZN(n13573) );
  INV_X1 U11824 ( .A(n15797), .ZN(n14656) );
  AND2_X2 U11825 ( .A1(n10519), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10252) );
  CLKBUF_X1 U11826 ( .A(n11559), .Z(n13155) );
  INV_X1 U11827 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20723) );
  INV_X1 U11828 ( .A(n11476), .ZN(n14648) );
  NAND2_X1 U11829 ( .A1(n20594), .A2(n21012), .ZN(n10908) );
  INV_X1 U11830 ( .A(n13319), .ZN(n15808) );
  OR2_X1 U11831 ( .A1(n11353), .A2(n11318), .ZN(n11320) );
  NOR2_X1 U11832 ( .A1(n11349), .A2(n11488), .ZN(n11352) );
  INV_X1 U11833 ( .A(n11349), .ZN(n11357) );
  OR3_X1 U11834 ( .A1(n11353), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20353), .ZN(n11355) );
  OAI21_X1 U11835 ( .B1(n9986), .B2(n13058), .A(n12710), .ZN(n9994) );
  NOR2_X1 U11836 ( .A1(n9986), .A2(n14089), .ZN(n10052) );
  NOR2_X1 U11837 ( .A1(n9986), .A2(n12744), .ZN(n10034) );
  OAI21_X1 U11838 ( .B1(n9986), .B2(n12737), .A(n12735), .ZN(n10006) );
  NAND2_X1 U11839 ( .A1(n10102), .A2(n11902), .ZN(n11905) );
  NAND2_X1 U11840 ( .A1(n10454), .A2(n15507), .ZN(n10453) );
  INV_X1 U11841 ( .A(n16361), .ZN(n10454) );
  OAI21_X1 U11842 ( .B1(n9986), .B2(n15004), .A(n14082), .ZN(n10018) );
  OAI21_X1 U11843 ( .B1(n9986), .B2(n12733), .A(n12731), .ZN(n10000) );
  NOR2_X1 U11844 ( .A1(n9986), .A2(n13186), .ZN(n10031) );
  OAI21_X1 U11845 ( .B1(n9986), .B2(n15030), .A(n14100), .ZN(n10024) );
  INV_X1 U11846 ( .A(n14097), .ZN(n10047) );
  OAI21_X1 U11847 ( .B1(n9986), .B2(n15016), .A(n14094), .ZN(n10020) );
  INV_X1 U11848 ( .A(n14701), .ZN(n10362) );
  INV_X1 U11849 ( .A(n15124), .ZN(n10325) );
  OAI21_X1 U11850 ( .B1(n9986), .B2(n14092), .A(n14090), .ZN(n10022) );
  NOR2_X1 U11851 ( .A1(n9986), .A2(n14728), .ZN(n10049) );
  OR2_X1 U11852 ( .A1(n10507), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15008) );
  OR2_X1 U11853 ( .A1(n15021), .A2(n15331), .ZN(n15111) );
  NAND2_X1 U11854 ( .A1(n15003), .A2(n9929), .ZN(n15136) );
  OAI21_X1 U11855 ( .B1(n9986), .B2(n14998), .A(n14079), .ZN(n10014) );
  INV_X1 U11856 ( .A(n12787), .ZN(n10044) );
  OAI21_X1 U11857 ( .B1(n9986), .B2(n14760), .A(n12761), .ZN(n10016) );
  OAI21_X1 U11858 ( .B1(n9986), .B2(n14952), .A(n12758), .ZN(n10012) );
  OAI21_X1 U11859 ( .B1(n9986), .B2(n12755), .A(n12753), .ZN(n10010) );
  OAI21_X1 U11860 ( .B1(n9986), .B2(n14959), .A(n12748), .ZN(n10008) );
  NOR2_X1 U11861 ( .A1(n14866), .A2(n10463), .ZN(n10462) );
  INV_X1 U11862 ( .A(n13739), .ZN(n10463) );
  NAND2_X1 U11863 ( .A1(n9912), .A2(n12400), .ZN(n12582) );
  OAI21_X1 U11864 ( .B1(n9986), .B2(n14973), .A(n12745), .ZN(n10002) );
  INV_X1 U11865 ( .A(n13626), .ZN(n10357) );
  AND2_X1 U11866 ( .A1(n10248), .A2(n16244), .ZN(n10247) );
  INV_X1 U11867 ( .A(n14950), .ZN(n10246) );
  NAND2_X1 U11868 ( .A1(n10247), .A2(n16260), .ZN(n10243) );
  NOR2_X1 U11869 ( .A1(n10447), .A2(n16332), .ZN(n10446) );
  INV_X1 U11870 ( .A(n10449), .ZN(n10447) );
  OAI21_X1 U11871 ( .B1(n9986), .B2(n12724), .A(n12722), .ZN(n9998) );
  OAI21_X1 U11872 ( .B1(n9986), .B2(n12719), .A(n12717), .ZN(n9996) );
  NOR2_X1 U11873 ( .A1(n9986), .A2(n12716), .ZN(n10028) );
  INV_X1 U11874 ( .A(n13053), .ZN(n10353) );
  INV_X1 U11875 ( .A(n9992), .ZN(n9991) );
  AND2_X1 U11876 ( .A1(n10088), .A2(n10087), .ZN(n13531) );
  NAND2_X1 U11877 ( .A1(n10082), .A2(n10083), .ZN(n10086) );
  INV_X1 U11878 ( .A(n13447), .ZN(n10083) );
  NOR2_X1 U11879 ( .A1(n12551), .A2(n12550), .ZN(n12552) );
  NOR2_X1 U11880 ( .A1(n12540), .A2(n12539), .ZN(n12553) );
  NAND2_X1 U11881 ( .A1(n10319), .A2(n12604), .ZN(n11826) );
  NOR2_X1 U11882 ( .A1(n19250), .A2(n13399), .ZN(n13400) );
  NAND2_X1 U11883 ( .A1(n11689), .A2(n16412), .ZN(n11696) );
  AOI21_X1 U11884 ( .B1(n12816), .B2(n12348), .A(n12335), .ZN(n12342) );
  AND2_X1 U11885 ( .A1(n13837), .A2(n20078), .ZN(n12335) );
  NAND2_X1 U11886 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18988), .ZN(
        n13858) );
  NOR2_X1 U11887 ( .A1(n13858), .A2(n13855), .ZN(n13911) );
  AND2_X1 U11888 ( .A1(n10302), .A2(n18967), .ZN(n10301) );
  AND2_X1 U11889 ( .A1(n13852), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n15622) );
  AOI22_X1 U11890 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15613) );
  INV_X1 U11891 ( .A(n15620), .ZN(n10318) );
  NOR2_X1 U11892 ( .A1(n13868), .A2(n17210), .ZN(n10317) );
  NOR2_X1 U11893 ( .A1(n17144), .A2(n17361), .ZN(n10224) );
  NOR2_X1 U11894 ( .A1(n10296), .A2(n10300), .ZN(n10295) );
  INV_X1 U11895 ( .A(n10297), .ZN(n10296) );
  INV_X1 U11896 ( .A(n10295), .ZN(n10292) );
  INV_X1 U11897 ( .A(n18385), .ZN(n15559) );
  NAND2_X1 U11898 ( .A1(n18400), .A2(n18385), .ZN(n15765) );
  XNOR2_X1 U11899 ( .A(n15698), .B(n17955), .ZN(n15699) );
  NOR3_X1 U11900 ( .A1(n15557), .A2(n15556), .A3(n15555), .ZN(n15577) );
  NOR2_X1 U11901 ( .A1(n13877), .A2(n10115), .ZN(n10114) );
  NOR3_X1 U11902 ( .A1(n15765), .A2(n15551), .A3(n18809), .ZN(n15764) );
  NAND2_X1 U11903 ( .A1(n15572), .A2(n15729), .ZN(n17551) );
  NOR2_X1 U11904 ( .A1(n15785), .A2(n15786), .ZN(n12909) );
  NAND2_X1 U11905 ( .A1(n14310), .A2(n9940), .ZN(n14285) );
  NAND2_X1 U11906 ( .A1(n10694), .A2(n10695), .ZN(n11678) );
  AND2_X1 U11907 ( .A1(n20625), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11651) );
  NOR2_X1 U11908 ( .A1(n10491), .A2(n10486), .ZN(n10485) );
  INV_X1 U11909 ( .A(n12626), .ZN(n10491) );
  NAND2_X1 U11910 ( .A1(n11302), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U11911 ( .A1(n14123), .A2(n14125), .ZN(n14124) );
  AND2_X1 U11912 ( .A1(n11541), .A2(n10147), .ZN(n10145) );
  CLKBUF_X1 U11913 ( .A(n13610), .Z(n13611) );
  NAND2_X1 U11914 ( .A1(n10979), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10989) );
  AND2_X1 U11915 ( .A1(n13086), .A2(n10475), .ZN(n10474) );
  NAND2_X1 U11916 ( .A1(n13087), .A2(n13086), .ZN(n13220) );
  NOR2_X1 U11917 ( .A1(n14383), .A2(n11546), .ZN(n11547) );
  NAND2_X1 U11918 ( .A1(n11531), .A2(n11615), .ZN(n11546) );
  INV_X1 U11919 ( .A(n11522), .ZN(n10257) );
  OR2_X1 U11920 ( .A1(n20995), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U11921 ( .A1(n10855), .A2(n20385), .ZN(n13506) );
  INV_X1 U11922 ( .A(n20532), .ZN(n20560) );
  NOR2_X1 U11923 ( .A1(n20656), .A2(n20483), .ZN(n20810) );
  OR2_X1 U11924 ( .A1(n13332), .A2(n13339), .ZN(n20772) );
  NOR2_X2 U11925 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20848) );
  NAND2_X1 U11926 ( .A1(n14648), .A2(n14650), .ZN(n20857) );
  AOI21_X1 U11927 ( .B1(n20766), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20483), 
        .ZN(n20858) );
  NAND2_X1 U11928 ( .A1(n11752), .A2(n16412), .ZN(n11759) );
  NOR2_X1 U11929 ( .A1(n14822), .A2(n10458), .ZN(n10457) );
  INV_X1 U11930 ( .A(n15353), .ZN(n10458) );
  INV_X1 U11931 ( .A(n13448), .ZN(n10193) );
  NOR2_X1 U11932 ( .A1(n19248), .A2(n20079), .ZN(n19217) );
  NOR2_X1 U11933 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  INV_X1 U11934 ( .A(n12751), .ZN(n10038) );
  NAND2_X1 U11935 ( .A1(n12740), .A2(n10039), .ZN(n13466) );
  NOR2_X1 U11936 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  INV_X1 U11937 ( .A(n12739), .ZN(n10041) );
  NAND2_X1 U11938 ( .A1(n11987), .A2(n9939), .ZN(n10406) );
  AND2_X1 U11939 ( .A1(n9894), .A2(n10348), .ZN(n10347) );
  INV_X1 U11940 ( .A(n13347), .ZN(n10348) );
  NAND2_X1 U11941 ( .A1(n12258), .A2(n10390), .ZN(n10392) );
  NOR2_X1 U11942 ( .A1(n10391), .A2(n14699), .ZN(n10390) );
  NAND2_X1 U11943 ( .A1(n9866), .A2(n10094), .ZN(n10093) );
  INV_X1 U11944 ( .A(n14714), .ZN(n10094) );
  NAND2_X1 U11945 ( .A1(n10402), .A2(n10401), .ZN(n10397) );
  AND2_X1 U11946 ( .A1(n14742), .A2(n14743), .ZN(n14744) );
  INV_X1 U11947 ( .A(n10413), .ZN(n10411) );
  INV_X1 U11948 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12652) );
  INV_X1 U11949 ( .A(n15413), .ZN(n10268) );
  CLKBUF_X1 U11950 ( .A(n12659), .Z(n12660) );
  NAND2_X1 U11951 ( .A1(n10339), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10338) );
  NOR2_X1 U11952 ( .A1(n15482), .A2(n10140), .ZN(n10139) );
  INV_X1 U11953 ( .A(n15466), .ZN(n10140) );
  XNOR2_X1 U11954 ( .A(n11886), .B(n11859), .ZN(n11860) );
  INV_X1 U11955 ( .A(n10026), .ZN(n10025) );
  OAI21_X1 U11956 ( .B1(n9986), .B2(n14683), .A(n14681), .ZN(n10026) );
  INV_X1 U11957 ( .A(n14718), .ZN(n10358) );
  NOR2_X1 U11958 ( .A1(n14709), .A2(n14679), .ZN(n10359) );
  NAND2_X1 U11959 ( .A1(n10440), .A2(n15235), .ZN(n10435) );
  OR2_X1 U11960 ( .A1(n14804), .A2(n10438), .ZN(n10437) );
  AND2_X1 U11961 ( .A1(n9934), .A2(n10351), .ZN(n10350) );
  INV_X1 U11962 ( .A(n14735), .ZN(n10351) );
  AND2_X1 U11963 ( .A1(n10068), .A2(n10248), .ZN(n10067) );
  AND2_X1 U11964 ( .A1(n14943), .A2(n10249), .ZN(n10248) );
  INV_X1 U11965 ( .A(n15454), .ZN(n10249) );
  INV_X1 U11966 ( .A(n15452), .ZN(n16263) );
  NAND2_X1 U11967 ( .A1(n16290), .A2(n10272), .ZN(n10181) );
  AND2_X1 U11968 ( .A1(n10272), .A2(n21411), .ZN(n10074) );
  AND2_X1 U11969 ( .A1(n9959), .A2(n13023), .ZN(n13260) );
  NAND2_X1 U11970 ( .A1(n10086), .A2(n13528), .ZN(n13460) );
  NOR2_X1 U11971 ( .A1(n13794), .A2(n12939), .ZN(n16434) );
  AND2_X1 U11972 ( .A1(n12930), .A2(n12992), .ZN(n12967) );
  INV_X1 U11973 ( .A(n13792), .ZN(n13003) );
  NAND2_X1 U11974 ( .A1(n12918), .A2(n12375), .ZN(n16438) );
  NAND2_X1 U11975 ( .A1(n10102), .A2(n10100), .ZN(n10106) );
  NOR2_X1 U11976 ( .A1(n11903), .A2(n10101), .ZN(n10100) );
  AND2_X1 U11977 ( .A1(n15526), .A2(n20081), .ZN(n19623) );
  NOR2_X1 U11978 ( .A1(n15526), .A2(n20081), .ZN(n19820) );
  NAND2_X1 U11979 ( .A1(n20059), .A2(n20081), .ZN(n19790) );
  INV_X1 U11980 ( .A(n19659), .ZN(n19655) );
  NOR2_X1 U11981 ( .A1(n13858), .A2(n13856), .ZN(n13852) );
  NAND2_X1 U11982 ( .A1(n10308), .A2(n10303), .ZN(n16490) );
  AOI21_X1 U11983 ( .B1(n16547), .B2(n17811), .A(n10304), .ZN(n10303) );
  NOR2_X1 U11984 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10310) );
  AND2_X1 U11985 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10309) );
  NOR2_X1 U11986 ( .A1(n18080), .A2(n17795), .ZN(n10311) );
  NAND2_X1 U11987 ( .A1(n15559), .A2(n15727), .ZN(n18808) );
  NAND2_X1 U11988 ( .A1(n10214), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10213) );
  NAND2_X1 U11989 ( .A1(n15697), .A2(n10214), .ZN(n10212) );
  OR2_X1 U11990 ( .A1(n17974), .A2(n17973), .ZN(n10216) );
  OAI21_X1 U11991 ( .B1(n15722), .B2(n13958), .A(n15721), .ZN(n18803) );
  INV_X1 U11992 ( .A(n18005), .ZN(n10217) );
  INV_X1 U11993 ( .A(n13851), .ZN(n17042) );
  NAND2_X1 U11994 ( .A1(n15566), .A2(n15763), .ZN(n16666) );
  INV_X1 U11995 ( .A(n16997), .ZN(n18372) );
  NAND2_X1 U11996 ( .A1(n11580), .A2(n20107), .ZN(n10166) );
  AND2_X1 U11997 ( .A1(n14065), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13495) );
  AND2_X1 U11998 ( .A1(n13502), .A2(n13497), .ZN(n20186) );
  AND2_X1 U11999 ( .A1(n13502), .A2(n13500), .ZN(n20179) );
  NAND2_X1 U12000 ( .A1(n11368), .A2(n11367), .ZN(n14316) );
  AND2_X1 U12001 ( .A1(n11584), .A2(n20107), .ZN(n11367) );
  NAND2_X1 U12002 ( .A1(n11366), .A2(n11661), .ZN(n11368) );
  INV_X2 U12003 ( .A(n14316), .ZN(n20211) );
  NAND2_X2 U12004 ( .A1(n20211), .A2(n11664), .ZN(n14312) );
  INV_X1 U12005 ( .A(n14379), .ZN(n14375) );
  AND2_X1 U12006 ( .A1(n11663), .A2(n20107), .ZN(n14380) );
  OR2_X1 U12007 ( .A1(n13162), .A2(n11662), .ZN(n11663) );
  INV_X1 U12008 ( .A(n14062), .ZN(n10265) );
  NAND2_X1 U12009 ( .A1(n14137), .A2(n11301), .ZN(n10126) );
  NOR2_X1 U12010 ( .A1(n9840), .A2(n10266), .ZN(n14536) );
  AND2_X1 U12011 ( .A1(n12636), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10266) );
  OR2_X1 U12012 ( .A1(n16010), .A2(n11600), .ZN(n14592) );
  AND2_X1 U12013 ( .A1(n11602), .A2(n11576), .ZN(n20332) );
  NAND2_X1 U12014 ( .A1(n11655), .A2(n11657), .ZN(n11575) );
  OR2_X1 U12015 ( .A1(n12637), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20342) );
  AND2_X1 U12016 ( .A1(n11602), .A2(n11583), .ZN(n20316) );
  INV_X1 U12017 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20766) );
  CLKBUF_X1 U12018 ( .A(n13506), .Z(n20595) );
  NAND2_X1 U12019 ( .A1(n10383), .A2(n19249), .ZN(n13634) );
  NAND2_X1 U12020 ( .A1(n15212), .A2(n19420), .ZN(n10281) );
  NOR2_X1 U12021 ( .A1(n10280), .A2(n10278), .ZN(n10277) );
  INV_X1 U12022 ( .A(n10279), .ZN(n10278) );
  NOR2_X1 U12023 ( .A1(n16277), .A2(n19091), .ZN(n10280) );
  AOI21_X1 U12024 ( .B1(n16270), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15423), .ZN(n10279) );
  INV_X1 U12025 ( .A(n15210), .ZN(n10283) );
  OR2_X1 U12026 ( .A1(n12835), .A2(n12403), .ZN(n19415) );
  AND2_X1 U12027 ( .A1(n19423), .A2(n20071), .ZN(n19420) );
  NAND2_X1 U12028 ( .A1(n12835), .A2(n12831), .ZN(n19423) );
  AND2_X1 U12029 ( .A1(n19423), .A2(n12862), .ZN(n19411) );
  AND2_X1 U12030 ( .A1(n12832), .A2(n12403), .ZN(n16294) );
  XNOR2_X1 U12031 ( .A(n15070), .B(n15071), .ZN(n15290) );
  INV_X1 U12032 ( .A(n10241), .ZN(n15207) );
  AND2_X1 U12033 ( .A1(n12967), .A2(n20093), .ZN(n16393) );
  INV_X1 U12034 ( .A(n10383), .ZN(n13040) );
  INV_X1 U12035 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20086) );
  INV_X1 U12036 ( .A(n15526), .ZN(n20059) );
  NAND2_X1 U12037 ( .A1(n10396), .A2(n11883), .ZN(n12988) );
  AND2_X1 U12038 ( .A1(n19654), .A2(n20053), .ZN(n19599) );
  NAND2_X1 U12039 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17055), .ZN(n17019) );
  INV_X1 U12040 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17367) );
  NOR2_X1 U12041 ( .A1(n17613), .A2(n17425), .ZN(n17419) );
  NAND2_X1 U12042 ( .A1(n17514), .A2(n9965), .ZN(n17487) );
  NOR2_X1 U12043 ( .A1(n9897), .A2(n10222), .ZN(n10221) );
  INV_X1 U12044 ( .A(n15681), .ZN(n10225) );
  NAND2_X1 U12045 ( .A1(n10232), .A2(n16545), .ZN(n10231) );
  NAND2_X1 U12046 ( .A1(n16539), .A2(n17669), .ZN(n10232) );
  NAND2_X1 U12047 ( .A1(n10228), .A2(n17664), .ZN(n10227) );
  OR2_X1 U12048 ( .A1(n18043), .A2(n17674), .ZN(n10228) );
  INV_X1 U12049 ( .A(n18343), .ZN(n18361) );
  OR2_X1 U12050 ( .A1(n13648), .A2(n12052), .ZN(n13383) );
  OAI22_X1 U12051 ( .A1(n13388), .A2(n13387), .B1(n19478), .B2(n13386), .ZN(
        n13395) );
  NAND2_X1 U12052 ( .A1(n9809), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13405) );
  AND2_X1 U12053 ( .A1(n20766), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11331) );
  AND2_X1 U12054 ( .A1(n10168), .A2(n10167), .ZN(n11335) );
  AOI21_X1 U12055 ( .B1(n11357), .B2(n11553), .A(n11332), .ZN(n10167) );
  NAND2_X1 U12056 ( .A1(n11345), .A2(n13496), .ZN(n10168) );
  INV_X1 U12057 ( .A(n11345), .ZN(n11341) );
  AND2_X1 U12058 ( .A1(n14905), .A2(n14904), .ZN(n14907) );
  AOI22_X1 U12059 ( .A1(n14880), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10136), .B2(n10135), .ZN(n13425) );
  AND2_X1 U12060 ( .A1(n13364), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10135) );
  OAI21_X1 U12061 ( .B1(n13402), .B2(n10184), .A(n10183), .ZN(n10182) );
  INV_X1 U12062 ( .A(n13389), .ZN(n10136) );
  AOI21_X1 U12063 ( .B1(n12342), .B2(n12344), .A(n12343), .ZN(n12338) );
  NAND2_X1 U12064 ( .A1(n10833), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12065 ( .A1(n10747), .A2(n10746), .ZN(n10748) );
  NAND2_X1 U12066 ( .A1(n10768), .A2(n10767), .ZN(n10770) );
  OR2_X1 U12067 ( .A1(n10906), .A2(n10905), .ZN(n11490) );
  NAND2_X2 U12068 ( .A1(n11913), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12310) );
  NAND2_X1 U12069 ( .A1(n12721), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U12070 ( .A1(n11838), .A2(n12364), .ZN(n10274) );
  AND2_X1 U12071 ( .A1(n14671), .A2(n11801), .ZN(n10386) );
  NAND2_X1 U12072 ( .A1(n11795), .A2(n10319), .ZN(n10185) );
  AOI21_X1 U12073 ( .B1(n12570), .B2(n13443), .A(n9958), .ZN(n10189) );
  INV_X1 U12074 ( .A(n11774), .ZN(n11776) );
  INV_X1 U12075 ( .A(n13390), .ZN(n13399) );
  NAND2_X1 U12076 ( .A1(n10136), .A2(n9851), .ZN(n13424) );
  AND2_X1 U12077 ( .A1(n13363), .A2(n10090), .ZN(n13390) );
  NOR2_X1 U12078 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12079 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18822), .ZN(
        n15569) );
  NOR2_X1 U12080 ( .A1(n10119), .A2(n10118), .ZN(n10117) );
  NOR2_X1 U12081 ( .A1(n17349), .A2(n13874), .ZN(n10118) );
  NAND2_X1 U12082 ( .A1(n10120), .A2(n9899), .ZN(n10119) );
  NAND2_X1 U12083 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10116) );
  NOR2_X1 U12084 ( .A1(n13579), .A2(n13589), .ZN(n11365) );
  NOR2_X1 U12085 ( .A1(n11261), .A2(n14191), .ZN(n11271) );
  NAND2_X1 U12086 ( .A1(n11161), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U12087 ( .A1(n9868), .A2(n11539), .ZN(n10147) );
  NOR2_X1 U12088 ( .A1(n14237), .A2(n10484), .ZN(n10483) );
  INV_X1 U12089 ( .A(n14247), .ZN(n10484) );
  INV_X1 U12090 ( .A(n13790), .ZN(n10480) );
  AND2_X1 U12091 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10934), .ZN(
        n10956) );
  INV_X1 U12092 ( .A(n10694), .ZN(n10881) );
  INV_X1 U12093 ( .A(n14547), .ZN(n10379) );
  NAND2_X1 U12094 ( .A1(n10376), .A2(n15986), .ZN(n10374) );
  NOR2_X1 U12095 ( .A1(n14422), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10380) );
  NOR2_X1 U12096 ( .A1(n10986), .A2(n10158), .ZN(n10157) );
  INV_X1 U12097 ( .A(n10967), .ZN(n10158) );
  NOR2_X1 U12098 ( .A1(n14291), .A2(n10419), .ZN(n10418) );
  INV_X1 U12099 ( .A(n10420), .ZN(n10419) );
  INV_X1 U12100 ( .A(n11437), .ZN(n11441) );
  NAND2_X1 U12101 ( .A1(n10417), .A2(n10415), .ZN(n11371) );
  NAND2_X1 U12102 ( .A1(n11374), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n10417) );
  NAND2_X1 U12103 ( .A1(n9821), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10794) );
  INV_X1 U12104 ( .A(n11589), .ZN(n10751) );
  INV_X1 U12105 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12106 ( .A1(n10751), .A2(n10750), .ZN(n13139) );
  NOR2_X1 U12107 ( .A1(n13496), .A2(n14043), .ZN(n10750) );
  AOI22_X1 U12108 ( .A1(n10697), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10617) );
  CLKBUF_X1 U12109 ( .A(n13568), .Z(n14649) );
  OAI21_X1 U12110 ( .B1(n21018), .B2(n13329), .A(n20987), .ZN(n13578) );
  INV_X1 U12111 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20653) );
  OR3_X1 U12112 ( .A1(n13162), .A2(n13161), .A3(n13160), .ZN(n15795) );
  AOI22_X1 U12113 ( .A1(n11351), .A2(n11350), .B1(n11552), .B2(n11352), .ZN(
        n10170) );
  NAND2_X1 U12114 ( .A1(n21012), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10169) );
  OAI21_X1 U12115 ( .B1(n13443), .B2(n12936), .A(n10188), .ZN(n12820) );
  NAND2_X1 U12116 ( .A1(n12936), .A2(n12681), .ZN(n10188) );
  INV_X1 U12117 ( .A(n14966), .ZN(n10198) );
  AND2_X1 U12118 ( .A1(n10462), .A2(n14858), .ZN(n10461) );
  NOR2_X1 U12119 ( .A1(n12404), .A2(n12741), .ZN(n14962) );
  INV_X1 U12120 ( .A(n13449), .ZN(n10191) );
  NOR2_X1 U12121 ( .A1(n9986), .A2(n14955), .ZN(n10037) );
  NOR2_X1 U12122 ( .A1(n9986), .A2(n12741), .ZN(n10040) );
  CLKBUF_X1 U12123 ( .A(n11709), .Z(n12314) );
  NOR2_X1 U12124 ( .A1(n14699), .A2(n10395), .ZN(n10394) );
  INV_X1 U12125 ( .A(n14707), .ZN(n10395) );
  INV_X1 U12126 ( .A(n12233), .ZN(n10095) );
  NAND2_X1 U12127 ( .A1(n10399), .A2(n10398), .ZN(n12212) );
  NAND2_X1 U12128 ( .A1(n10404), .A2(n14730), .ZN(n10398) );
  NAND2_X1 U12129 ( .A1(n10400), .A2(n10402), .ZN(n10399) );
  NAND2_X1 U12130 ( .A1(n10414), .A2(n10505), .ZN(n10413) );
  INV_X1 U12131 ( .A(n13757), .ZN(n10414) );
  NOR2_X1 U12132 ( .A1(n16343), .A2(n10450), .ZN(n10449) );
  INV_X1 U12133 ( .A(n15458), .ZN(n10450) );
  INV_X1 U12134 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U12135 ( .A1(n11858), .A2(n11857), .ZN(n11885) );
  OR2_X1 U12136 ( .A1(n12443), .A2(n12442), .ZN(n12843) );
  NOR2_X1 U12137 ( .A1(n9855), .A2(n15302), .ZN(n10323) );
  NAND2_X1 U12138 ( .A1(n10326), .A2(n9857), .ZN(n15081) );
  INV_X1 U12139 ( .A(n15350), .ZN(n10187) );
  NAND2_X1 U12140 ( .A1(n12727), .A2(n10003), .ZN(n12728) );
  INV_X1 U12141 ( .A(n10004), .ZN(n10003) );
  NAND2_X1 U12142 ( .A1(n14875), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10057) );
  NAND2_X1 U12143 ( .A1(n14912), .A2(n9928), .ZN(n10238) );
  INV_X1 U12144 ( .A(n13667), .ZN(n9984) );
  INV_X1 U12145 ( .A(n13253), .ZN(n10443) );
  NAND2_X1 U12146 ( .A1(n11894), .A2(n9987), .ZN(n11896) );
  INV_X1 U12147 ( .A(n9988), .ZN(n9987) );
  NAND2_X1 U12148 ( .A1(n11808), .A2(n11774), .ZN(n12377) );
  NAND2_X1 U12149 ( .A1(n9851), .A2(n12839), .ZN(n10102) );
  NAND2_X1 U12150 ( .A1(n13401), .A2(n13369), .ZN(n13387) );
  INV_X1 U12151 ( .A(n13424), .ZN(n19757) );
  AOI22_X1 U12152 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11781) );
  NAND3_X1 U12153 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20057), .A3(n19863), 
        .ZN(n13213) );
  NAND2_X1 U12154 ( .A1(n12369), .A2(n12368), .ZN(n12824) );
  OR2_X1 U12155 ( .A1(n12367), .A2(n12366), .ZN(n12369) );
  AOI211_X1 U12156 ( .C1(n17242), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15602), .B(n15601), .ZN(n15603) );
  NOR2_X1 U12157 ( .A1(n18024), .A2(n10298), .ZN(n10297) );
  NOR2_X1 U12158 ( .A1(n10306), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10305) );
  INV_X1 U12159 ( .A(n10310), .ZN(n10306) );
  NOR2_X1 U12160 ( .A1(n17955), .A2(n15698), .ZN(n16538) );
  NOR2_X1 U12161 ( .A1(n18207), .A2(n18213), .ZN(n18183) );
  NOR2_X1 U12162 ( .A1(n15640), .A2(n15748), .ZN(n15745) );
  AOI21_X1 U12163 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(n15721) );
  AOI211_X1 U12164 ( .C1(n18389), .C2(n18817), .A(n15765), .B(n15575), .ZN(
        n15720) );
  OAI21_X1 U12165 ( .B1(n15559), .B2(n15558), .A(n15577), .ZN(n15766) );
  AOI221_X1 U12166 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18970), .C1(n18856), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18982), .ZN(n18371) );
  NAND2_X1 U12167 ( .A1(n10762), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U12168 ( .A1(n10175), .A2(n14052), .ZN(n10174) );
  INV_X1 U12169 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14191) );
  NOR2_X1 U12170 ( .A1(n9974), .A2(n21128), .ZN(n10175) );
  NOR2_X1 U12171 ( .A1(n14226), .A2(n21128), .ZN(n15861) );
  NAND2_X1 U12172 ( .A1(n11093), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11108) );
  AND2_X1 U12173 ( .A1(n13808), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n10172) );
  OR2_X1 U12174 ( .A1(n20179), .A2(n13810), .ZN(n20123) );
  INV_X1 U12175 ( .A(n10771), .ZN(n10772) );
  AND2_X1 U12176 ( .A1(n11434), .A2(n11433), .ZN(n14192) );
  NOR3_X1 U12177 ( .A1(n14276), .A2(n14218), .A3(n10424), .ZN(n14203) );
  AND2_X1 U12178 ( .A1(n11417), .A2(n11416), .ZN(n14294) );
  NAND2_X1 U12179 ( .A1(n14310), .A2(n14305), .ZN(n14304) );
  AND2_X1 U12180 ( .A1(n11411), .A2(n11410), .ZN(n14308) );
  INV_X1 U12181 ( .A(n11213), .ZN(n14271) );
  AND3_X1 U12182 ( .A1(n11010), .A2(n11009), .A3(n11008), .ZN(n13703) );
  NAND2_X1 U12183 ( .A1(n10912), .A2(n11117), .ZN(n10921) );
  AND2_X1 U12184 ( .A1(n13049), .A2(n15849), .ZN(n20212) );
  AND2_X1 U12185 ( .A1(n10666), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U12186 ( .A1(n11271), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11282) );
  AND2_X1 U12187 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  INV_X1 U12188 ( .A(n14165), .ZN(n10478) );
  AND2_X1 U12189 ( .A1(n11253), .A2(n11252), .ZN(n14199) );
  AND2_X1 U12190 ( .A1(n11160), .A2(n11159), .ZN(n14289) );
  NOR2_X1 U12191 ( .A1(n11108), .A2(n15900), .ZN(n11139) );
  CLKBUF_X1 U12192 ( .A(n14297), .Z(n14298) );
  INV_X1 U12193 ( .A(n14508), .ZN(n10160) );
  INV_X1 U12194 ( .A(n14505), .ZN(n10159) );
  NOR2_X1 U12195 ( .A1(n11074), .A2(n14250), .ZN(n11078) );
  AND2_X1 U12196 ( .A1(n11039), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U12197 ( .A1(n11044), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11074) );
  AND2_X1 U12198 ( .A1(n11117), .A2(n11062), .ZN(n13841) );
  NOR2_X1 U12199 ( .A1(n11013), .A2(n10664), .ZN(n11039) );
  INV_X1 U12200 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20142) );
  NOR2_X1 U12201 ( .A1(n10989), .A2(n20142), .ZN(n11007) );
  AOI21_X1 U12202 ( .B1(n11505), .B2(n11117), .A(n10982), .ZN(n13481) );
  AND2_X1 U12203 ( .A1(n10956), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10979) );
  OAI21_X1 U12204 ( .B1(n11295), .B2(n10962), .A(n10961), .ZN(n10963) );
  NAND2_X1 U12205 ( .A1(n14648), .A2(n10260), .ZN(n11483) );
  NAND2_X1 U12206 ( .A1(n14406), .A2(n11619), .ZN(n10367) );
  NAND2_X1 U12207 ( .A1(n10373), .A2(n10370), .ZN(n14383) );
  NAND2_X1 U12208 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  AND2_X1 U12209 ( .A1(n10375), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U12210 ( .A1(n11531), .A2(n10151), .ZN(n10150) );
  INV_X1 U12211 ( .A(n10376), .ZN(n10151) );
  INV_X1 U12212 ( .A(n10380), .ZN(n10377) );
  OR2_X1 U12213 ( .A1(n10423), .A2(n14178), .ZN(n10422) );
  NAND2_X1 U12214 ( .A1(n10381), .A2(n15938), .ZN(n14423) );
  NAND2_X1 U12215 ( .A1(n11542), .A2(n15938), .ZN(n14450) );
  NOR2_X1 U12216 ( .A1(n14276), .A2(n14218), .ZN(n14217) );
  NAND2_X1 U12217 ( .A1(n14481), .A2(n14480), .ZN(n14603) );
  OR3_X1 U12218 ( .A1(n14470), .A2(n15938), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U12219 ( .A1(n14310), .A2(n10420), .ZN(n14296) );
  NAND2_X1 U12220 ( .A1(n11538), .A2(n11537), .ZN(n14487) );
  OR3_X1 U12221 ( .A1(n16067), .A2(n10427), .A3(n11407), .ZN(n10426) );
  NAND2_X1 U12222 ( .A1(n14515), .A2(n16033), .ZN(n15951) );
  NOR3_X1 U12223 ( .A1(n16066), .A2(n16067), .A3(n10429), .ZN(n15916) );
  NOR2_X1 U12224 ( .A1(n16066), .A2(n16067), .ZN(n16065) );
  NAND2_X1 U12225 ( .A1(n13269), .A2(n11487), .ZN(n20294) );
  NAND2_X1 U12226 ( .A1(n11580), .A2(n13496), .ZN(n11655) );
  AND2_X1 U12227 ( .A1(n16055), .A2(n20323), .ZN(n14630) );
  INV_X1 U12228 ( .A(n20323), .ZN(n13561) );
  NAND2_X1 U12229 ( .A1(n10154), .A2(n10867), .ZN(n11582) );
  INV_X1 U12230 ( .A(n13139), .ZN(n10154) );
  NAND2_X1 U12231 ( .A1(n10863), .A2(n10862), .ZN(n10910) );
  NAND2_X1 U12232 ( .A1(n9821), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10894) );
  AND2_X1 U12233 ( .A1(n11564), .A2(n15776), .ZN(n15800) );
  INV_X1 U12234 ( .A(n15795), .ZN(n13327) );
  OR2_X1 U12235 ( .A1(n13332), .A2(n13570), .ZN(n20476) );
  NAND2_X1 U12236 ( .A1(n14649), .A2(n11476), .ZN(n20455) );
  NAND2_X1 U12237 ( .A1(n14648), .A2(n13569), .ZN(n20532) );
  OR2_X1 U12238 ( .A1(n14649), .A2(n14648), .ZN(n20695) );
  AND2_X1 U12239 ( .A1(n13332), .A2(n13570), .ZN(n20559) );
  AND2_X1 U12240 ( .A1(n13332), .A2(n13339), .ZN(n20799) );
  INV_X1 U12241 ( .A(n20857), .ZN(n20800) );
  NAND2_X1 U12242 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n16097) );
  AND4_X1 U12243 ( .A1(n19452), .A2(n19439), .A3(n11791), .A4(n12949), .ZN(
        n11797) );
  AND2_X1 U12244 ( .A1(n12594), .A2(n12593), .ZN(n14803) );
  AND3_X1 U12245 ( .A1(n10201), .A2(n10200), .A3(n15012), .ZN(n16174) );
  AND2_X1 U12246 ( .A1(n12590), .A2(n12589), .ZN(n14822) );
  AND2_X1 U12247 ( .A1(n16313), .A2(n10459), .ZN(n14842) );
  AND2_X1 U12248 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  INV_X1 U12249 ( .A(n14850), .ZN(n10460) );
  NAND2_X1 U12250 ( .A1(n14967), .A2(n9861), .ZN(n14969) );
  NAND2_X1 U12251 ( .A1(n16313), .A2(n10461), .ZN(n14857) );
  CLKBUF_X1 U12252 ( .A(n12655), .Z(n12656) );
  NOR2_X1 U12253 ( .A1(n19148), .A2(n19146), .ZN(n19133) );
  AND2_X1 U12254 ( .A1(n14929), .A2(n13182), .ZN(n14933) );
  NOR2_X1 U12255 ( .A1(n19168), .A2(n19166), .ZN(n19156) );
  NOR2_X2 U12256 ( .A1(n14925), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14929) );
  NOR2_X1 U12257 ( .A1(n19192), .A2(n19190), .ZN(n19176) );
  NOR2_X1 U12258 ( .A1(n19212), .A2(n19210), .ZN(n19200) );
  NAND2_X1 U12259 ( .A1(n12711), .A2(n9993), .ZN(n12712) );
  INV_X1 U12260 ( .A(n9994), .ZN(n9993) );
  NOR2_X1 U12261 ( .A1(n19410), .A2(n19237), .ZN(n19221) );
  NOR2_X1 U12262 ( .A1(n13630), .A2(n13761), .ZN(n13689) );
  NAND2_X1 U12263 ( .A1(n14088), .A2(n10051), .ZN(n14719) );
  NOR2_X1 U12264 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  INV_X1 U12265 ( .A(n14087), .ZN(n10053) );
  NAND2_X1 U12266 ( .A1(n12743), .A2(n10033), .ZN(n13477) );
  NOR2_X1 U12267 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U12268 ( .A(n12742), .ZN(n10035) );
  NAND2_X1 U12269 ( .A1(n12736), .A2(n10005), .ZN(n12738) );
  INV_X1 U12270 ( .A(n10006), .ZN(n10005) );
  NOR2_X1 U12271 ( .A1(n10391), .A2(n10389), .ZN(n10388) );
  INV_X1 U12272 ( .A(n10394), .ZN(n10389) );
  NAND2_X1 U12273 ( .A1(n10099), .A2(n10098), .ZN(n10097) );
  INV_X1 U12274 ( .A(n14715), .ZN(n10098) );
  NAND2_X1 U12275 ( .A1(n15354), .A2(n15353), .ZN(n15356) );
  NAND2_X1 U12276 ( .A1(n10412), .A2(n10505), .ZN(n13756) );
  INV_X1 U12277 ( .A(n13476), .ZN(n10405) );
  AND3_X1 U12278 ( .A1(n12573), .A2(n12572), .A3(n12571), .ZN(n16332) );
  NAND2_X1 U12279 ( .A1(n10448), .A2(n10449), .ZN(n16331) );
  AND3_X1 U12280 ( .A1(n12560), .A2(n12559), .A3(n12558), .ZN(n15489) );
  NOR2_X1 U12281 ( .A1(n16362), .A2(n10452), .ZN(n15488) );
  OR2_X1 U12282 ( .A1(n10453), .A2(n15489), .ZN(n10452) );
  OR2_X1 U12283 ( .A1(n16362), .A2(n10453), .ZN(n15508) );
  AND2_X1 U12284 ( .A1(n12409), .A2(n12408), .ZN(n16361) );
  NOR2_X1 U12285 ( .A1(n16362), .A2(n16361), .ZN(n16360) );
  AND2_X1 U12286 ( .A1(n12893), .A2(n19967), .ZN(n19334) );
  INV_X1 U12287 ( .A(n12615), .ZN(n19268) );
  OAI21_X1 U12288 ( .B1(n12614), .B2(n12613), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12615) );
  INV_X1 U12289 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15131) );
  CLKBUF_X1 U12290 ( .A(n15129), .Z(n15130) );
  NAND2_X1 U12291 ( .A1(n14083), .A2(n10017), .ZN(n14084) );
  INV_X1 U12292 ( .A(n10018), .ZN(n10017) );
  CLKBUF_X1 U12293 ( .A(n12777), .Z(n12778) );
  NAND2_X1 U12294 ( .A1(n12732), .A2(n9999), .ZN(n12734) );
  INV_X1 U12295 ( .A(n10000), .ZN(n9999) );
  NAND2_X1 U12296 ( .A1(n13184), .A2(n9894), .ZN(n13348) );
  NAND2_X1 U12297 ( .A1(n12730), .A2(n10030), .ZN(n13183) );
  NOR2_X1 U12298 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  INV_X1 U12299 ( .A(n12729), .ZN(n10032) );
  NAND2_X1 U12300 ( .A1(n13184), .A2(n13183), .ZN(n13298) );
  INV_X1 U12301 ( .A(n12663), .ZN(n10337) );
  AND2_X1 U12302 ( .A1(n15060), .A2(n15027), .ZN(n10327) );
  NAND2_X1 U12303 ( .A1(n14101), .A2(n10023), .ZN(n14102) );
  INV_X1 U12304 ( .A(n10024), .ZN(n10023) );
  NAND2_X1 U12305 ( .A1(n14098), .A2(n10045), .ZN(n14690) );
  NOR2_X1 U12306 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  NOR2_X1 U12307 ( .A1(n9986), .A2(n14099), .ZN(n10046) );
  AND3_X1 U12308 ( .A1(n16128), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15087), .ZN(n15068) );
  OR2_X1 U12309 ( .A1(n14789), .A2(n14788), .ZN(n15294) );
  NAND2_X1 U12310 ( .A1(n14095), .A2(n10019), .ZN(n14096) );
  INV_X1 U12311 ( .A(n10020), .ZN(n10019) );
  AND2_X1 U12312 ( .A1(n10363), .A2(n10362), .ZN(n14702) );
  NAND2_X1 U12313 ( .A1(n10071), .A2(n10070), .ZN(n15090) );
  NAND2_X1 U12314 ( .A1(n10072), .A2(n9903), .ZN(n10071) );
  NAND2_X1 U12315 ( .A1(n14091), .A2(n10021), .ZN(n14093) );
  INV_X1 U12316 ( .A(n10022), .ZN(n10021) );
  INV_X1 U12317 ( .A(n10363), .ZN(n14711) );
  NAND2_X1 U12318 ( .A1(n14086), .A2(n10048), .ZN(n14725) );
  NOR2_X1 U12319 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  INV_X1 U12320 ( .A(n14085), .ZN(n10050) );
  INV_X1 U12321 ( .A(n15111), .ZN(n15126) );
  NAND2_X1 U12322 ( .A1(n15195), .A2(n10186), .ZN(n15140) );
  AND2_X1 U12323 ( .A1(n9966), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10186) );
  AND2_X1 U12324 ( .A1(n15195), .A2(n9966), .ZN(n15146) );
  NAND2_X1 U12325 ( .A1(n14080), .A2(n10013), .ZN(n14081) );
  INV_X1 U12326 ( .A(n10014), .ZN(n10013) );
  NAND2_X1 U12327 ( .A1(n12790), .A2(n9934), .ZN(n14738) );
  AOI21_X1 U12328 ( .B1(n10066), .B2(n10062), .A(n10061), .ZN(n10060) );
  NAND2_X1 U12329 ( .A1(n10066), .A2(n10064), .ZN(n10063) );
  INV_X1 U12330 ( .A(n15364), .ZN(n10061) );
  NAND2_X1 U12331 ( .A1(n12788), .A2(n10042), .ZN(n12789) );
  NOR2_X1 U12332 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  NOR2_X1 U12333 ( .A1(n9986), .A2(n14754), .ZN(n10043) );
  NAND2_X1 U12334 ( .A1(n12790), .A2(n12789), .ZN(n14740) );
  NAND2_X1 U12335 ( .A1(n12762), .A2(n10015), .ZN(n12763) );
  INV_X1 U12336 ( .A(n10016), .ZN(n10015) );
  NAND2_X1 U12337 ( .A1(n15185), .A2(n10240), .ZN(n10239) );
  NAND2_X1 U12338 ( .A1(n12759), .A2(n10011), .ZN(n12760) );
  INV_X1 U12339 ( .A(n10012), .ZN(n10011) );
  NAND2_X1 U12340 ( .A1(n13478), .A2(n9865), .ZN(n14774) );
  NAND2_X1 U12341 ( .A1(n12754), .A2(n10009), .ZN(n12756) );
  INV_X1 U12342 ( .A(n10010), .ZN(n10009) );
  NAND2_X1 U12343 ( .A1(n12749), .A2(n10007), .ZN(n12750) );
  INV_X1 U12344 ( .A(n10008), .ZN(n10007) );
  AND2_X1 U12345 ( .A1(n12579), .A2(n12578), .ZN(n14866) );
  AND2_X1 U12346 ( .A1(n16313), .A2(n10462), .ZN(n14864) );
  NAND2_X1 U12347 ( .A1(n16313), .A2(n13739), .ZN(n14865) );
  NAND2_X1 U12348 ( .A1(n12746), .A2(n10001), .ZN(n12747) );
  INV_X1 U12349 ( .A(n10002), .ZN(n10001) );
  NAND2_X1 U12350 ( .A1(n13478), .A2(n9888), .ZN(n13730) );
  NAND2_X1 U12351 ( .A1(n13478), .A2(n13477), .ZN(n13625) );
  NOR2_X1 U12352 ( .A1(n16315), .A2(n16314), .ZN(n16313) );
  INV_X1 U12353 ( .A(n10247), .ZN(n10244) );
  AND2_X1 U12354 ( .A1(n10243), .A2(n10245), .ZN(n10242) );
  NAND2_X1 U12355 ( .A1(n10246), .A2(n16244), .ZN(n10245) );
  NAND2_X1 U12356 ( .A1(n10448), .A2(n10444), .ZN(n16314) );
  NOR2_X1 U12357 ( .A1(n10445), .A2(n10451), .ZN(n10444) );
  INV_X1 U12358 ( .A(n15437), .ZN(n10451) );
  INV_X1 U12359 ( .A(n10446), .ZN(n10445) );
  NOR2_X1 U12360 ( .A1(n16342), .A2(n16343), .ZN(n16341) );
  INV_X1 U12361 ( .A(n15482), .ZN(n10138) );
  NAND2_X1 U12362 ( .A1(n12723), .A2(n9997), .ZN(n12725) );
  INV_X1 U12363 ( .A(n9998), .ZN(n9997) );
  NAND2_X1 U12364 ( .A1(n12718), .A2(n9995), .ZN(n12720) );
  INV_X1 U12365 ( .A(n9996), .ZN(n9995) );
  NAND2_X1 U12366 ( .A1(n12715), .A2(n10027), .ZN(n13045) );
  NOR2_X1 U12367 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  INV_X1 U12368 ( .A(n12714), .ZN(n10029) );
  NAND2_X1 U12369 ( .A1(n13721), .A2(n12527), .ZN(n16375) );
  NAND2_X1 U12370 ( .A1(n12707), .A2(n9991), .ZN(n12709) );
  NAND2_X1 U12371 ( .A1(n12705), .A2(n10354), .ZN(n13054) );
  XNOR2_X1 U12372 ( .A(n14875), .B(n13672), .ZN(n14874) );
  OR2_X1 U12373 ( .A1(n19234), .A2(n13677), .ZN(n10058) );
  NAND2_X1 U12374 ( .A1(n10089), .A2(n10084), .ZN(n10080) );
  INV_X1 U12375 ( .A(n13532), .ZN(n10084) );
  NAND2_X1 U12376 ( .A1(n13023), .A2(n10441), .ZN(n13719) );
  AND2_X1 U12377 ( .A1(n12493), .A2(n10442), .ZN(n10441) );
  AND2_X1 U12378 ( .A1(n10443), .A2(n13261), .ZN(n10442) );
  NAND2_X1 U12379 ( .A1(n12702), .A2(n9989), .ZN(n12703) );
  INV_X1 U12380 ( .A(n9990), .ZN(n9989) );
  NAND2_X1 U12381 ( .A1(n10234), .A2(n10235), .ZN(n13523) );
  NAND2_X1 U12382 ( .A1(n13460), .A2(n13692), .ZN(n10234) );
  NOR3_X1 U12383 ( .A1(n11812), .A2(n11826), .A3(n12956), .ZN(n11813) );
  OR2_X1 U12384 ( .A1(n12943), .A2(n12942), .ZN(n12945) );
  NAND2_X1 U12385 ( .A1(n13023), .A2(n12493), .ZN(n13252) );
  NAND2_X1 U12386 ( .A1(n11862), .A2(n20079), .ZN(n11901) );
  XNOR2_X1 U12387 ( .A(n13792), .B(n11880), .ZN(n12997) );
  AND2_X1 U12388 ( .A1(n12981), .A2(n12980), .ZN(n16430) );
  INV_X1 U12389 ( .A(n13387), .ZN(n14881) );
  NAND2_X1 U12390 ( .A1(n9862), .A2(n13364), .ZN(n13434) );
  INV_X1 U12391 ( .A(n19477), .ZN(n19483) );
  OR3_X1 U12392 ( .A1(n19757), .A2(n19779), .A3(n19822), .ZN(n19761) );
  OR2_X1 U12393 ( .A1(n20065), .A2(n20072), .ZN(n19789) );
  NOR2_X1 U12394 ( .A1(n19268), .A2(n13213), .ZN(n19464) );
  NOR2_X1 U12395 ( .A1(n19267), .A2(n13213), .ZN(n19465) );
  INV_X1 U12396 ( .A(n19464), .ZN(n19466) );
  INV_X1 U12397 ( .A(n19465), .ZN(n19468) );
  OR2_X1 U12398 ( .A1(n20065), .A2(n13276), .ZN(n19659) );
  OR2_X1 U12399 ( .A1(n14880), .A2(n13280), .ZN(n13283) );
  NAND2_X1 U12400 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19863), .ZN(n19470) );
  XNOR2_X1 U12401 ( .A(n12347), .B(n12346), .ZN(n12804) );
  INV_X1 U12402 ( .A(n12387), .ZN(n16462) );
  NOR2_X1 U12403 ( .A1(n15727), .A2(n15560), .ZN(n15576) );
  AND2_X1 U12404 ( .A1(n16666), .A2(n16665), .ZN(n18800) );
  NOR2_X1 U12405 ( .A1(n17977), .A2(n10290), .ZN(n10289) );
  INV_X1 U12406 ( .A(n13855), .ZN(n10111) );
  INV_X1 U12407 ( .A(n15625), .ZN(n17275) );
  OAI211_X1 U12408 ( .C1(n13868), .C2(n17148), .A(n15661), .B(n15660), .ZN(
        n15740) );
  NOR2_X1 U12409 ( .A1(n15623), .A2(n15622), .ZN(n15624) );
  AOI21_X1 U12410 ( .B1(n17176), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n10224), .ZN(n10223) );
  NOR2_X1 U12411 ( .A1(n17588), .A2(n17551), .ZN(n17569) );
  AND3_X1 U12412 ( .A1(n10294), .A2(n10293), .A3(n10291), .ZN(n16977) );
  NAND2_X1 U12413 ( .A1(n10292), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10291) );
  OR2_X1 U12414 ( .A1(n16512), .A2(n10299), .ZN(n10294) );
  NAND2_X1 U12415 ( .A1(n16512), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16477) );
  NOR2_X1 U12416 ( .A1(n17662), .A2(n17663), .ZN(n16512) );
  AND2_X1 U12417 ( .A1(n17764), .A2(n9947), .ZN(n17688) );
  INV_X1 U12418 ( .A(n17703), .ZN(n10284) );
  NOR2_X1 U12419 ( .A1(n17703), .A2(n16679), .ZN(n17657) );
  NAND2_X1 U12420 ( .A1(n17764), .A2(n9873), .ZN(n17702) );
  NOR2_X1 U12421 ( .A1(n16680), .A2(n16681), .ZN(n17700) );
  NOR2_X1 U12422 ( .A1(n17746), .A2(n10286), .ZN(n10285) );
  NAND2_X1 U12423 ( .A1(n17764), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17745) );
  NOR2_X1 U12424 ( .A1(n17776), .A2(n17778), .ZN(n17764) );
  NOR2_X1 U12425 ( .A1(n17815), .A2(n17817), .ZN(n17803) );
  NOR2_X1 U12426 ( .A1(n10288), .A2(n16867), .ZN(n10287) );
  NAND2_X1 U12427 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10288) );
  NOR2_X1 U12428 ( .A1(n18008), .A2(n17018), .ZN(n17990) );
  NOR2_X1 U12429 ( .A1(n16524), .A2(n17659), .ZN(n16508) );
  NAND2_X1 U12430 ( .A1(n17706), .A2(n15762), .ZN(n18041) );
  NOR2_X1 U12431 ( .A1(n18076), .A2(n17725), .ZN(n17706) );
  NOR2_X1 U12432 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17758), .ZN(
        n17740) );
  NAND2_X1 U12433 ( .A1(n10209), .A2(n10205), .ZN(n10204) );
  NOR2_X1 U12434 ( .A1(n17933), .A2(n18164), .ZN(n10205) );
  NOR2_X1 U12435 ( .A1(n17887), .A2(n16534), .ZN(n18169) );
  NOR2_X1 U12436 ( .A1(n18174), .A2(n18173), .ZN(n18172) );
  NAND2_X1 U12437 ( .A1(n18226), .A2(n18183), .ZN(n18200) );
  INV_X1 U12438 ( .A(n17887), .ZN(n18224) );
  INV_X1 U12439 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17945) );
  INV_X1 U12440 ( .A(n17954), .ZN(n17955) );
  INV_X1 U12441 ( .A(n17988), .ZN(n10315) );
  NOR2_X1 U12442 ( .A1(n17995), .A2(n18317), .ZN(n17994) );
  INV_X1 U12443 ( .A(n18833), .ZN(n18804) );
  INV_X1 U12444 ( .A(n18389), .ZN(n15725) );
  NAND2_X1 U12445 ( .A1(n15733), .A2(n15720), .ZN(n18797) );
  NAND2_X1 U12446 ( .A1(n16665), .A2(n15565), .ZN(n15768) );
  NOR2_X1 U12447 ( .A1(n15766), .A2(n15560), .ZN(n15763) );
  NAND2_X1 U12448 ( .A1(n15764), .A2(n19024), .ZN(n18833) );
  INV_X1 U12449 ( .A(n13875), .ZN(n10121) );
  OAI211_X1 U12450 ( .C1(n9813), .C2(n15653), .A(n13921), .B(n13920), .ZN(
        n18393) );
  INV_X1 U12451 ( .A(n18685), .ZN(n18745) );
  OAI22_X1 U12452 ( .A1(n16474), .A2(n18797), .B1(n18803), .B2(n18332), .ZN(
        n18805) );
  AOI211_X1 U12453 ( .C1(n15764), .C2(n15582), .A(n15856), .B(n15581), .ZN(
        n18835) );
  INV_X1 U12454 ( .A(n12915), .ZN(n10164) );
  OAI21_X1 U12455 ( .B1(n14122), .B2(n21249), .A(n21178), .ZN(n10161) );
  AND2_X1 U12456 ( .A1(n20177), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n10433) );
  NOR3_X1 U12457 ( .A1(n14226), .A2(n10174), .A3(n14057), .ZN(n14151) );
  NOR2_X1 U12458 ( .A1(n14226), .A2(n10173), .ZN(n14222) );
  INV_X1 U12459 ( .A(n10175), .ZN(n10173) );
  NOR2_X1 U12460 ( .A1(n15905), .A2(n15886), .ZN(n15882) );
  INV_X1 U12461 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15900) );
  NOR2_X1 U12462 ( .A1(n21376), .A2(n14252), .ZN(n15906) );
  AND2_X1 U12463 ( .A1(n20179), .A2(n9971), .ZN(n15921) );
  INV_X1 U12464 ( .A(n14050), .ZN(n10171) );
  NAND2_X1 U12465 ( .A1(n20179), .A2(n9881), .ZN(n20129) );
  INV_X1 U12466 ( .A(n20170), .ZN(n20153) );
  AND2_X1 U12467 ( .A1(n20161), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20190) );
  INV_X1 U12468 ( .A(n20190), .ZN(n20172) );
  AND2_X1 U12469 ( .A1(n13502), .A2(n13501), .ZN(n20177) );
  INV_X1 U12470 ( .A(n20177), .ZN(n20201) );
  INV_X1 U12471 ( .A(n14312), .ZN(n20206) );
  OR3_X1 U12472 ( .A1(n14374), .A2(n11678), .A3(n14369), .ZN(n11676) );
  AND2_X1 U12473 ( .A1(n14380), .A2(n14044), .ZN(n14364) );
  INV_X1 U12474 ( .A(n14042), .ZN(n14361) );
  INV_X1 U12475 ( .A(n14380), .ZN(n14374) );
  NAND2_X1 U12476 ( .A1(n14380), .A2(n13083), .ZN(n14379) );
  BUF_X1 U12477 ( .A(n13128), .Z(n20241) );
  INV_X1 U12478 ( .A(n20245), .ZN(n20287) );
  XNOR2_X1 U12479 ( .A(n13491), .B(n13490), .ZN(n14065) );
  INV_X1 U12480 ( .A(n11652), .ZN(n11653) );
  NAND2_X1 U12481 ( .A1(n10488), .A2(n10485), .ZN(n11654) );
  NAND2_X1 U12482 ( .A1(n10472), .A2(n10475), .ZN(n13221) );
  NAND2_X1 U12483 ( .A1(n11602), .A2(n15788), .ZN(n20323) );
  NAND2_X1 U12484 ( .A1(n10255), .A2(n10256), .ZN(n13820) );
  OR2_X1 U12485 ( .A1(n15970), .A2(n10258), .ZN(n10255) );
  NAND2_X1 U12486 ( .A1(n10259), .A2(n11523), .ZN(n13748) );
  NAND2_X1 U12487 ( .A1(n15970), .A2(n11522), .ZN(n10259) );
  INV_X1 U12489 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20353) );
  INV_X1 U12490 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U12491 ( .A1(n16101), .A2(n20985), .ZN(n20995) );
  INV_X1 U12492 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16096) );
  INV_X1 U12493 ( .A(n20454), .ZN(n20472) );
  OAI21_X1 U12494 ( .B1(n20500), .B2(n20484), .A(n20810), .ZN(n20502) );
  OAI21_X1 U12495 ( .B1(n20680), .B2(n20985), .A(n20662), .ZN(n20683) );
  INV_X1 U12496 ( .A(n20715), .ZN(n20682) );
  AOI22_X1 U12497 ( .A1(n20728), .A2(n20725), .B1(n20722), .B2(n20721), .ZN(
        n20765) );
  NOR2_X1 U12498 ( .A1(n20483), .A2(n20255), .ZN(n20805) );
  INV_X1 U12499 ( .A(n20853), .ZN(n20806) );
  NOR2_X1 U12500 ( .A1(n20483), .A2(n20258), .ZN(n20816) );
  INV_X1 U12501 ( .A(n20871), .ZN(n20817) );
  INV_X1 U12502 ( .A(n20878), .ZN(n20823) );
  NOR2_X1 U12503 ( .A1(n20483), .A2(n20262), .ZN(n20828) );
  INV_X1 U12504 ( .A(n20887), .ZN(n20829) );
  OAI211_X1 U12505 ( .C1(n20840), .C2(n20811), .A(n20810), .B(n20809), .ZN(
        n20843) );
  NOR2_X2 U12506 ( .A1(n20857), .A2(n20772), .ZN(n20842) );
  INV_X1 U12507 ( .A(n20822), .ZN(n20877) );
  INV_X1 U12508 ( .A(n20752), .ZN(n20899) );
  NAND2_X1 U12509 ( .A1(n20800), .A2(n20799), .ZN(n20915) );
  INV_X1 U12510 ( .A(n20904), .ZN(n20911) );
  INV_X1 U12511 ( .A(n20758), .ZN(n20909) );
  NOR2_X1 U12512 ( .A1(n15783), .A2(n20985), .ZN(n15825) );
  INV_X1 U12513 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16101) );
  NAND2_X1 U12514 ( .A1(n16101), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20917) );
  INV_X1 U12515 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20985) );
  INV_X1 U12516 ( .A(n16132), .ZN(n16135) );
  NAND2_X1 U12517 ( .A1(n15354), .A2(n10457), .ZN(n14813) );
  INV_X1 U12518 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15167) );
  INV_X1 U12519 ( .A(n19189), .ZN(n19110) );
  INV_X1 U12520 ( .A(n10342), .ZN(n19054) );
  NOR2_X1 U12521 ( .A1(n19066), .A2(n19055), .ZN(n10343) );
  NOR2_X1 U12522 ( .A1(n19075), .A2(n9835), .ZN(n19065) );
  NOR2_X1 U12523 ( .A1(n19065), .A2(n19066), .ZN(n19064) );
  NOR2_X1 U12524 ( .A1(n19126), .A2(n19131), .ZN(n19117) );
  OR2_X1 U12525 ( .A1(n19032), .A2(n12679), .ZN(n19183) );
  AND2_X1 U12526 ( .A1(n19032), .A2(n16461), .ZN(n19251) );
  INV_X1 U12527 ( .A(n19110), .ZN(n19244) );
  INV_X1 U12528 ( .A(n19183), .ZN(n19248) );
  AND2_X1 U12529 ( .A1(n12768), .A2(n12767), .ZN(n19249) );
  NAND2_X1 U12530 ( .A1(n14694), .A2(n14693), .ZN(n14695) );
  OR2_X1 U12531 ( .A1(n11951), .A2(n11950), .ZN(n13175) );
  NOR2_X1 U12532 ( .A1(n11939), .A2(n11938), .ZN(n13108) );
  AND2_X1 U12533 ( .A1(n9874), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10407) );
  INV_X1 U12534 ( .A(n14779), .ZN(n14746) );
  INV_X1 U12535 ( .A(n20072), .ZN(n13276) );
  AND2_X1 U12536 ( .A1(n14782), .A2(n15234), .ZN(n16133) );
  NAND2_X1 U12537 ( .A1(n14708), .A2(n14707), .ZN(n14706) );
  NOR2_X1 U12538 ( .A1(n14744), .A2(n12164), .ZN(n14731) );
  NAND2_X1 U12539 ( .A1(n19282), .A2(n12605), .ZN(n14868) );
  AND2_X1 U12540 ( .A1(n12398), .A2(n12992), .ZN(n19282) );
  NAND2_X1 U12541 ( .A1(n12444), .A2(n19282), .ZN(n19269) );
  NAND2_X1 U12542 ( .A1(n13005), .A2(n11904), .ZN(n13016) );
  INV_X1 U12543 ( .A(n19282), .ZN(n19317) );
  INV_X1 U12544 ( .A(n19269), .ZN(n19319) );
  NOR2_X1 U12545 ( .A1(n13203), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19335) );
  NOR2_X1 U12546 ( .A1(n19383), .A2(n19405), .ZN(n12911) );
  CLKBUF_X2 U12547 ( .A(n12911), .Z(n19406) );
  INV_X1 U12548 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16252) );
  OAI21_X1 U12549 ( .B1(n16277), .B2(n16256), .A(n16255), .ZN(n10079) );
  INV_X1 U12550 ( .A(n19411), .ZN(n16277) );
  INV_X1 U12551 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19424) );
  INV_X1 U12552 ( .A(n19415), .ZN(n16293) );
  XNOR2_X1 U12553 ( .A(n14687), .B(n14686), .ZN(n16115) );
  NAND2_X1 U12554 ( .A1(n10358), .A2(n9930), .ZN(n14687) );
  NAND2_X1 U12555 ( .A1(n14682), .A2(n10025), .ZN(n14684) );
  NAND2_X1 U12556 ( .A1(n10065), .A2(n10066), .ZN(n15366) );
  NAND2_X1 U12557 ( .A1(n10250), .A2(n10067), .ZN(n10065) );
  NAND2_X1 U12558 ( .A1(n10250), .A2(n10248), .ZN(n16243) );
  NAND2_X1 U12559 ( .A1(n10250), .A2(n14943), .ZN(n15456) );
  NAND2_X1 U12560 ( .A1(n16241), .A2(n9907), .ZN(n16254) );
  INV_X1 U12561 ( .A(n15480), .ZN(n10270) );
  AND2_X1 U12562 ( .A1(n15251), .A2(n15250), .ZN(n15486) );
  NAND2_X1 U12563 ( .A1(n10141), .A2(n10142), .ZN(n15484) );
  NAND2_X1 U12564 ( .A1(n15224), .A2(n9827), .ZN(n15226) );
  INV_X1 U12565 ( .A(n16365), .ZN(n16407) );
  AND2_X1 U12566 ( .A1(n12967), .A2(n12941), .ZN(n16399) );
  NAND2_X1 U12567 ( .A1(n13003), .A2(n13002), .ZN(n20081) );
  INV_X1 U12568 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20069) );
  INV_X1 U12569 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16427) );
  NAND2_X1 U12570 ( .A1(n12995), .A2(n12998), .ZN(n20072) );
  OR2_X1 U12571 ( .A1(n12997), .A2(n12996), .ZN(n12998) );
  AND2_X1 U12572 ( .A1(n16438), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16465) );
  AOI21_X1 U12573 ( .B1(n10383), .B2(n15524), .A(n13779), .ZN(n16414) );
  NAND2_X1 U12574 ( .A1(n13005), .A2(n13008), .ZN(n15526) );
  OR2_X1 U12575 ( .A1(n19516), .A2(n19826), .ZN(n19533) );
  INV_X1 U12576 ( .A(n19582), .ZN(n19600) );
  OR3_X1 U12577 ( .A1(n19631), .A2(n19826), .A3(n19630), .ZN(n19650) );
  NOR2_X2 U12578 ( .A1(n13287), .A2(n19483), .ZN(n19751) );
  NOR2_X2 U12579 ( .A1(n19790), .A2(n19537), .ZN(n19781) );
  NAND2_X1 U12580 ( .A1(n19820), .A2(n20053), .ZN(n19819) );
  OAI22_X1 U12581 ( .A1(n19451), .A2(n19468), .B1(n19450), .B2(n19466), .ZN(
        n19879) );
  INV_X1 U12582 ( .A(n19886), .ZN(n19892) );
  OAI21_X1 U12583 ( .B1(n19868), .B2(n19867), .A(n19866), .ZN(n19894) );
  INV_X1 U12584 ( .A(n19942), .ZN(n19926) );
  NOR2_X1 U12585 ( .A1(n19790), .A2(n19659), .ZN(n19931) );
  OR2_X1 U12586 ( .A1(n19956), .A2(n19822), .ZN(n16471) );
  NOR2_X1 U12587 ( .A1(n17590), .A2(n15576), .ZN(n16649) );
  NAND2_X1 U12588 ( .A1(n19005), .A2(n18799), .ZN(n17588) );
  NOR2_X1 U12589 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16789), .ZN(n16775) );
  NOR2_X1 U12590 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16814), .ZN(n16796) );
  NAND2_X1 U12591 ( .A1(n18849), .A2(n16668), .ZN(n17045) );
  NOR2_X1 U12592 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16858), .ZN(n16844) );
  NOR2_X1 U12593 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16981), .ZN(n16965) );
  INV_X1 U12594 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17018) );
  NOR2_X1 U12595 ( .A1(n18970), .A2(n18865), .ZN(n17014) );
  OAI211_X1 U12596 ( .C1(n18857), .C2(n18858), .A(n16667), .B(n19023), .ZN(
        n17055) );
  NOR2_X1 U12597 ( .A1(n17061), .A2(n17120), .ZN(n17125) );
  OAI211_X1 U12598 ( .C1(n17339), .C2(n17367), .A(n13867), .B(n13866), .ZN(
        n18400) );
  AOI211_X1 U12599 ( .C1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(n17176), .A(
        n13865), .B(n13864), .ZN(n13866) );
  NOR2_X1 U12600 ( .A1(n16940), .A2(n17321), .ZN(n17343) );
  NOR2_X1 U12601 ( .A1(n16960), .A2(n17368), .ZN(n17344) );
  NOR3_X1 U12602 ( .A1(n16989), .A2(n17384), .A3(n17371), .ZN(n17375) );
  INV_X1 U12603 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17383) );
  INV_X1 U12604 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17389) );
  INV_X1 U12605 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17391) );
  NAND2_X1 U12606 ( .A1(n17438), .A2(n9879), .ZN(n17425) );
  NAND2_X1 U12607 ( .A1(n17438), .A2(n17445), .ZN(n17433) );
  NAND2_X1 U12608 ( .A1(n17438), .A2(n9877), .ZN(n17434) );
  NOR2_X1 U12609 ( .A1(n17606), .A2(n17439), .ZN(n17438) );
  INV_X1 U12610 ( .A(n17455), .ZN(n17473) );
  NOR2_X1 U12611 ( .A1(n17487), .A2(n17656), .ZN(n17480) );
  AND2_X1 U12612 ( .A1(n17401), .A2(n10112), .ZN(n17514) );
  AND2_X1 U12613 ( .A1(n17400), .A2(n9972), .ZN(n10112) );
  INV_X1 U12614 ( .A(n17514), .ZN(n17513) );
  AOI211_X2 U12615 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n15672), .B(n15671), .ZN(n17518) );
  NOR2_X1 U12616 ( .A1(n17445), .A2(n17542), .ZN(n17530) );
  INV_X1 U12617 ( .A(n17528), .ZN(n17549) );
  OAI21_X1 U12618 ( .B1(n15856), .B2(n15855), .A(n19005), .ZN(n17542) );
  NOR3_X1 U12619 ( .A1(n15854), .A2(n18372), .A3(n10113), .ZN(n15855) );
  INV_X1 U12620 ( .A(n17542), .ZN(n17401) );
  NOR2_X2 U12621 ( .A1(n18817), .A2(n17542), .ZN(n17528) );
  INV_X1 U12622 ( .A(n17541), .ZN(n17543) );
  NOR2_X1 U12623 ( .A1(n19012), .A2(n17652), .ZN(n17644) );
  OAI211_X1 U12624 ( .C1(n19012), .C2(n19013), .A(n17590), .B(n17589), .ZN(
        n17647) );
  BUF_X1 U12625 ( .A(n17647), .Z(n17652) );
  INV_X1 U12627 ( .A(n16977), .ZN(n17006) );
  AND2_X1 U12628 ( .A1(n16528), .A2(n18000), .ZN(n16494) );
  NOR2_X1 U12629 ( .A1(n18041), .A2(n16524), .ZN(n16506) );
  OAI21_X1 U12630 ( .B1(n17675), .B2(n17811), .A(n16547), .ZN(n17670) );
  NAND2_X1 U12631 ( .A1(n17845), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18174) );
  INV_X1 U12632 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17858) );
  INV_X1 U12633 ( .A(n17872), .ZN(n17857) );
  INV_X1 U12634 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17868) );
  NOR2_X2 U12635 ( .A1(n18970), .A2(n17953), .ZN(n17872) );
  NOR2_X2 U12636 ( .A1(n17518), .A2(n18032), .ZN(n17934) );
  INV_X1 U12637 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17977) );
  NAND2_X1 U12638 ( .A1(n17990), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17976) );
  NAND2_X1 U12639 ( .A1(n17802), .A2(n17857), .ZN(n17996) );
  INV_X1 U12640 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18008) );
  NAND2_X1 U12641 ( .A1(n18715), .A2(n16476), .ZN(n18685) );
  INV_X1 U12642 ( .A(n17996), .ZN(n18025) );
  INV_X1 U12643 ( .A(n18021), .ZN(n18032) );
  INV_X1 U12644 ( .A(n18000), .ZN(n18033) );
  INV_X1 U12645 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18970) );
  NAND2_X1 U12646 ( .A1(n16490), .A2(n16489), .ZN(n16491) );
  AND2_X1 U12647 ( .A1(n16528), .A2(n18356), .ZN(n16529) );
  NAND2_X1 U12648 ( .A1(n17675), .A2(n10309), .ZN(n15840) );
  NAND2_X1 U12649 ( .A1(n17676), .A2(n10310), .ZN(n15841) );
  NOR2_X1 U12650 ( .A1(n18357), .A2(n17661), .ZN(n10230) );
  INV_X1 U12651 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18856) );
  NAND2_X1 U12652 ( .A1(n10208), .A2(n10210), .ZN(n17801) );
  NAND2_X1 U12653 ( .A1(n10209), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10208) );
  INV_X1 U12654 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18173) );
  INV_X1 U12655 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18285) );
  NAND2_X1 U12656 ( .A1(n10212), .A2(n10211), .ZN(n17963) );
  NAND2_X2 U12657 ( .A1(n19012), .A2(n18261), .ZN(n18332) );
  INV_X1 U12658 ( .A(n10218), .ZN(n18006) );
  NOR2_X1 U12659 ( .A1(n18797), .A2(n18351), .ZN(n18343) );
  INV_X1 U12660 ( .A(n10220), .ZN(n18016) );
  NOR2_X1 U12661 ( .A1(n18332), .A2(n18351), .ZN(n18356) );
  INV_X1 U12662 ( .A(n18334), .ZN(n18351) );
  INV_X1 U12663 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18822) );
  AND2_X1 U12664 ( .A1(n19022), .A2(n16644), .ZN(n19004) );
  INV_X1 U12665 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18823) );
  INV_X1 U12666 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18369) );
  OAI211_X1 U12667 ( .C1(n18847), .C2(n18835), .A(n18370), .B(n15583), .ZN(
        n18986) );
  INV_X1 U12668 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18415) );
  NOR2_X1 U12669 ( .A1(n18857), .A2(n18856), .ZN(n19005) );
  INV_X1 U12670 ( .A(n17014), .ZN(n18863) );
  NAND2_X1 U12671 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18970), .ZN(n18857) );
  INV_X1 U12672 ( .A(n14369), .ZN(n13577) );
  OAI21_X1 U12674 ( .B1(n14527), .B2(n20174), .A(n10430), .ZN(P1_U2810) );
  INV_X1 U12675 ( .A(n10431), .ZN(n10430) );
  OAI21_X1 U12676 ( .B1(n14062), .B2(n20133), .A(n10432), .ZN(n10431) );
  AOI211_X1 U12677 ( .C1(n10161), .C2(n14061), .A(n10433), .B(n14049), .ZN(
        n10432) );
  NAND2_X1 U12678 ( .A1(n20179), .A2(n13808), .ZN(n20146) );
  AND2_X1 U12679 ( .A1(n11457), .A2(n10495), .ZN(n11458) );
  OR2_X1 U12680 ( .A1(n14114), .A2(n14312), .ZN(n11457) );
  OAI211_X1 U12681 ( .C1(n14536), .C2(n20108), .A(n12641), .B(n10264), .ZN(
        P1_U2969) );
  NAND2_X1 U12682 ( .A1(n10265), .A2(n20296), .ZN(n10264) );
  INV_X1 U12683 ( .A(n14560), .ZN(n10125) );
  OAI21_X1 U12684 ( .B1(n14068), .B2(n20340), .A(n11622), .ZN(P1_U3000) );
  OAI21_X1 U12685 ( .B1(n14560), .B2(n20340), .A(n10155), .ZN(P1_U3004) );
  NOR2_X1 U12686 ( .A1(n14561), .A2(n10156), .ZN(n10155) );
  NOR2_X1 U12687 ( .A1(n14545), .A2(n14556), .ZN(n10156) );
  NOR2_X1 U12688 ( .A1(n13040), .A2(n14776), .ZN(n10385) );
  NAND2_X1 U12689 ( .A1(n10281), .A2(n10277), .ZN(n10276) );
  AOI21_X1 U12690 ( .B1(n15415), .B2(n15211), .A(n19416), .ZN(n10282) );
  OAI21_X1 U12691 ( .B1(n16254), .B2(n19416), .A(n10076), .ZN(P2_U3002) );
  INV_X1 U12692 ( .A(n10077), .ZN(n10076) );
  OAI21_X1 U12693 ( .B1(n16253), .B2(n19415), .A(n10078), .ZN(n10077) );
  AOI21_X1 U12694 ( .B1(n19150), .B2(n19420), .A(n10079), .ZN(n10078) );
  AND2_X1 U12695 ( .A1(n19420), .A2(n10383), .ZN(n10384) );
  AOI21_X1 U12696 ( .B1(n15273), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15272), .ZN(n15274) );
  AOI21_X1 U12697 ( .B1(n15308), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15285), .ZN(n15286) );
  AOI21_X1 U12698 ( .B1(n16548), .B2(n17661), .A(n10227), .ZN(n10226) );
  NAND2_X1 U12699 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  AND2_X1 U12700 ( .A1(n11709), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U12701 ( .A1(n17041), .A2(n10111), .ZN(n15538) );
  NOR2_X1 U12702 ( .A1(n13363), .A2(n13200), .ZN(n9854) );
  NAND3_X2 U12703 ( .A1(n13801), .A2(n10233), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U12704 ( .A1(n10507), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9855) );
  NAND2_X1 U12705 ( .A1(n14246), .A2(n14247), .ZN(n14236) );
  NAND2_X1 U12706 ( .A1(n11194), .A2(n9955), .ZN(n14224) );
  AND2_X1 U12707 ( .A1(n10069), .A2(n13692), .ZN(n9856) );
  NOR2_X4 U12708 ( .A1(n13851), .A2(n13855), .ZN(n15618) );
  INV_X1 U12709 ( .A(n12429), .ZN(n11964) );
  AND2_X1 U12710 ( .A1(n12313), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11954) );
  AND2_X1 U12711 ( .A1(n11012), .A2(n9936), .ZN(n13789) );
  INV_X1 U12712 ( .A(n12258), .ZN(n10092) );
  NAND2_X1 U12713 ( .A1(n14200), .A2(n10479), .ZN(n14164) );
  NAND2_X1 U12714 ( .A1(n10337), .A2(n10339), .ZN(n12662) );
  NAND2_X1 U12715 ( .A1(n14200), .A2(n9956), .ZN(n14175) );
  OR2_X1 U12716 ( .A1(n12659), .A2(n9884), .ZN(n9858) );
  AND2_X1 U12717 ( .A1(n14246), .A2(n10483), .ZN(n9859) );
  NAND2_X1 U12718 ( .A1(n11194), .A2(n9925), .ZN(n9860) );
  NOR2_X1 U12720 ( .A1(n12688), .A2(n10198), .ZN(n9861) );
  NAND2_X1 U12721 ( .A1(n10055), .A2(n10057), .ZN(n16291) );
  AND2_X1 U12722 ( .A1(n9861), .A2(n9942), .ZN(n9863) );
  INV_X1 U12723 ( .A(n15136), .ZN(n10072) );
  AND2_X1 U12724 ( .A1(n9888), .A2(n10356), .ZN(n9864) );
  AND2_X1 U12725 ( .A1(n9864), .A2(n13759), .ZN(n9865) );
  NAND2_X2 U12726 ( .A1(n15494), .A2(n15051), .ZN(n15195) );
  AND2_X1 U12727 ( .A1(n10095), .A2(n12256), .ZN(n9866) );
  AND2_X1 U12728 ( .A1(n14480), .A2(n9975), .ZN(n9867) );
  AND2_X1 U12729 ( .A1(n11531), .A2(n9976), .ZN(n9868) );
  AND2_X1 U12730 ( .A1(n9863), .A2(n14952), .ZN(n9869) );
  AND2_X1 U12731 ( .A1(n9857), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U12732 ( .A1(n10108), .A2(n9961), .ZN(n9871) );
  INV_X2 U12733 ( .A(n12580), .ZN(n12510) );
  NAND2_X1 U12734 ( .A1(n10408), .A2(n13011), .ZN(n13014) );
  INV_X1 U12735 ( .A(n16648), .ZN(n18799) );
  INV_X1 U12736 ( .A(n15198), .ZN(n10240) );
  AND2_X1 U12737 ( .A1(n15103), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15095) );
  AND2_X1 U12738 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9872) );
  AND2_X1 U12739 ( .A1(n10285), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9873) );
  NAND2_X1 U12740 ( .A1(n10107), .A2(n10108), .ZN(n13621) );
  AND2_X1 U12741 ( .A1(n13011), .A2(n9969), .ZN(n9874) );
  AND2_X1 U12742 ( .A1(n14307), .A2(n10483), .ZN(n9875) );
  AND2_X1 U12743 ( .A1(n9872), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9876) );
  AND2_X1 U12744 ( .A1(n17445), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n9877) );
  AND2_X1 U12745 ( .A1(n9877), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n9878) );
  INV_X1 U12746 ( .A(n11301), .ZN(n10487) );
  AND2_X1 U12747 ( .A1(n9878), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n9879) );
  AND2_X1 U12748 ( .A1(n10439), .A2(n10438), .ZN(n9880) );
  AND2_X1 U12749 ( .A1(n10172), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n9881) );
  NAND2_X2 U12750 ( .A1(n10758), .A2(n13599), .ZN(n11374) );
  INV_X1 U12751 ( .A(n12434), .ZN(n12009) );
  INV_X1 U12752 ( .A(n15611), .ZN(n13879) );
  INV_X1 U12753 ( .A(n12428), .ZN(n11963) );
  OR3_X1 U12754 ( .A1(n14276), .A2(n14218), .A3(n10422), .ZN(n9882) );
  NOR3_X1 U12755 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13858), .ZN(n13870) );
  INV_X1 U12756 ( .A(n10113), .ZN(n19012) );
  AND2_X1 U12757 ( .A1(n15195), .A2(n15252), .ZN(n9883) );
  AND2_X1 U12758 ( .A1(n14154), .A2(n10132), .ZN(n14123) );
  OR2_X1 U12759 ( .A1(n16252), .A2(n10335), .ZN(n9884) );
  OR2_X1 U12760 ( .A1(n13101), .A2(n13100), .ZN(n9885) );
  AND2_X1 U12761 ( .A1(n14908), .A2(n9983), .ZN(n13678) );
  NAND2_X1 U12762 ( .A1(n14246), .A2(n9875), .ZN(n14301) );
  NOR2_X1 U12763 ( .A1(n12663), .A2(n10341), .ZN(n12661) );
  INV_X1 U12764 ( .A(n10312), .ZN(n17796) );
  NOR2_X1 U12765 ( .A1(n12663), .A2(n19186), .ZN(n12664) );
  AND2_X1 U12766 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12669) );
  OR2_X1 U12767 ( .A1(n10748), .A2(n10749), .ZN(n9886) );
  OR3_X1 U12768 ( .A1(n16118), .A2(n15043), .A3(n15269), .ZN(n9887) );
  AND2_X1 U12769 ( .A1(n13477), .A2(n10357), .ZN(n9888) );
  AND2_X1 U12770 ( .A1(n10354), .A2(n10353), .ZN(n9889) );
  NOR2_X1 U12771 ( .A1(n14288), .A2(n14289), .ZN(n9890) );
  INV_X1 U12772 ( .A(n10127), .ZN(n11194) );
  OR2_X1 U12773 ( .A1(n14288), .A2(n10130), .ZN(n10127) );
  AND2_X1 U12774 ( .A1(n11194), .A2(n10481), .ZN(n9891) );
  AND2_X1 U12775 ( .A1(n15195), .A2(n10268), .ZN(n9892) );
  OR3_X1 U12776 ( .A1(n14276), .A2(n14218), .A3(n10423), .ZN(n9893) );
  AND2_X1 U12777 ( .A1(n13183), .A2(n10349), .ZN(n9894) );
  OR3_X1 U12778 ( .A1(n17671), .A2(n18270), .A3(n16547), .ZN(n9895) );
  AND3_X1 U12779 ( .A1(n10141), .A2(n10142), .A3(n10139), .ZN(n9896) );
  INV_X1 U12780 ( .A(n13496), .ZN(n20355) );
  AND2_X2 U12781 ( .A1(n10233), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11913) );
  AND2_X1 U12782 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n9897) );
  AND3_X1 U12783 ( .A1(n13662), .A2(n13663), .A3(n13661), .ZN(n9898) );
  NAND2_X1 U12784 ( .A1(n13202), .A2(n13363), .ZN(n13368) );
  OR2_X1 U12785 ( .A1(n17339), .A2(n17391), .ZN(n9899) );
  AND2_X1 U12786 ( .A1(n10262), .A2(n10880), .ZN(n9901) );
  INV_X1 U12787 ( .A(n10269), .ZN(n16281) );
  OAI21_X1 U12788 ( .B1(n15195), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10270), .ZN(n10269) );
  INV_X2 U12789 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16412) );
  AND2_X1 U12790 ( .A1(n11360), .A2(n10169), .ZN(n9902) );
  AND2_X1 U12791 ( .A1(n10190), .A2(n9855), .ZN(n9903) );
  NOR2_X1 U12792 ( .A1(n14515), .A2(n16075), .ZN(n9904) );
  NOR2_X1 U12793 ( .A1(n13746), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9905) );
  AND2_X1 U12794 ( .A1(n15049), .A2(n15048), .ZN(n9906) );
  OR2_X1 U12795 ( .A1(n16263), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9907) );
  NAND2_X1 U12796 ( .A1(n10182), .A2(n13396), .ZN(n9908) );
  AND2_X1 U12797 ( .A1(n11782), .A2(n16412), .ZN(n9909) );
  AND2_X1 U12798 ( .A1(n11358), .A2(n9902), .ZN(n9910) );
  NAND2_X1 U12799 ( .A1(n14967), .A2(n9863), .ZN(n10199) );
  AND2_X1 U12800 ( .A1(n15162), .A2(n15159), .ZN(n9911) );
  AND2_X1 U12801 ( .A1(n9811), .A2(n12403), .ZN(n9912) );
  INV_X1 U12802 ( .A(n17041), .ZN(n13857) );
  NAND2_X1 U12803 ( .A1(n13746), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9913) );
  AND2_X1 U12804 ( .A1(n17676), .A2(n10305), .ZN(n9914) );
  OR2_X1 U12805 ( .A1(n9814), .A2(n15049), .ZN(n9915) );
  INV_X1 U12806 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17883) );
  INV_X1 U12807 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19186) );
  AND2_X1 U12808 ( .A1(n15682), .A2(n15679), .ZN(n9916) );
  AND2_X1 U12809 ( .A1(n12507), .A2(n10189), .ZN(n9917) );
  AND2_X1 U12810 ( .A1(n11532), .A2(n11539), .ZN(n9918) );
  INV_X1 U12811 ( .A(n15082), .ZN(n10190) );
  AND3_X1 U12812 ( .A1(n10141), .A2(n10142), .A3(n10138), .ZN(n9919) );
  AND2_X1 U12813 ( .A1(n10756), .A2(n14043), .ZN(n11572) );
  OR2_X1 U12814 ( .A1(n13368), .A2(n13433), .ZN(n9920) );
  AND2_X1 U12815 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9921) );
  AND2_X1 U12816 ( .A1(n9889), .A2(n13045), .ZN(n9922) );
  INV_X1 U12817 ( .A(n10328), .ZN(n10068) );
  NAND2_X1 U12818 ( .A1(n9911), .A2(n10329), .ZN(n10328) );
  OR2_X1 U12819 ( .A1(n15699), .A2(n18285), .ZN(n9923) );
  INV_X1 U12820 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19034) );
  INV_X1 U12821 ( .A(n12453), .ZN(n12581) );
  AND2_X1 U12822 ( .A1(n13442), .A2(n20079), .ZN(n12453) );
  NAND2_X1 U12823 ( .A1(n10107), .A2(n11987), .ZN(n13295) );
  INV_X1 U12824 ( .A(n16342), .ZN(n10448) );
  INV_X1 U12825 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20079) );
  INV_X1 U12826 ( .A(n11902), .ZN(n10101) );
  AND2_X1 U12827 ( .A1(n16373), .A2(n12554), .ZN(n16362) );
  INV_X1 U12828 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20078) );
  NOR2_X1 U12829 ( .A1(n13174), .A2(n9871), .ZN(n14762) );
  NOR2_X1 U12830 ( .A1(n13621), .A2(n10413), .ZN(n13755) );
  NAND2_X1 U12831 ( .A1(n11012), .A2(n11011), .ZN(n13702) );
  INV_X1 U12832 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13850) );
  NOR3_X1 U12833 ( .A1(n12659), .A2(n9884), .A3(n19109), .ZN(n12654) );
  NOR2_X1 U12834 ( .A1(n12651), .A2(n12652), .ZN(n12650) );
  NOR2_X1 U12835 ( .A1(n12659), .A2(n16252), .ZN(n12657) );
  AND2_X1 U12836 ( .A1(n17438), .A2(n9878), .ZN(n9924) );
  AND2_X1 U12837 ( .A1(n10481), .A2(n14214), .ZN(n9925) );
  OR2_X1 U12838 ( .A1(n13448), .A2(n13449), .ZN(n9926) );
  OR2_X1 U12839 ( .A1(n13449), .A2(n10192), .ZN(n9927) );
  AND2_X1 U12840 ( .A1(n15501), .A2(n15498), .ZN(n9928) );
  OR3_X1 U12841 ( .A1(n16201), .A2(n15043), .A3(n15352), .ZN(n9929) );
  AND2_X1 U12842 ( .A1(n10360), .A2(n10359), .ZN(n9930) );
  AND2_X1 U12843 ( .A1(n14310), .A2(n10418), .ZN(n9931) );
  AND2_X1 U12844 ( .A1(n13478), .A2(n9864), .ZN(n9932) );
  AND2_X1 U12845 ( .A1(n10448), .A2(n10446), .ZN(n9933) );
  INV_X1 U12846 ( .A(n15363), .ZN(n10064) );
  AND2_X1 U12847 ( .A1(n12789), .A2(n10352), .ZN(n9934) );
  OR2_X1 U12848 ( .A1(n10406), .A2(n10405), .ZN(n9935) );
  AND2_X1 U12849 ( .A1(n10480), .A2(n11011), .ZN(n9936) );
  INV_X1 U12850 ( .A(n19066), .ZN(n10345) );
  NAND2_X1 U12851 ( .A1(n12997), .A2(n12996), .ZN(n12995) );
  OR2_X1 U12852 ( .A1(n14226), .A2(n10174), .ZN(n9937) );
  AND2_X1 U12853 ( .A1(n10397), .A2(n10403), .ZN(n9938) );
  INV_X1 U12854 ( .A(n13621), .ZN(n10412) );
  AND2_X1 U12855 ( .A1(n13346), .A2(n12574), .ZN(n9939) );
  INV_X1 U12856 ( .A(n10425), .ZN(n15918) );
  NOR3_X1 U12857 ( .A1(n16066), .A2(n16067), .A3(n10427), .ZN(n10425) );
  AND2_X1 U12858 ( .A1(n10418), .A2(n14283), .ZN(n9940) );
  AND2_X1 U12859 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13837), .ZN(n9941) );
  OR2_X1 U12860 ( .A1(n12404), .A2(n12689), .ZN(n9942) );
  NAND2_X1 U12861 ( .A1(n10908), .A2(n10907), .ZN(n14650) );
  NOR2_X1 U12862 ( .A1(n16066), .A2(n10426), .ZN(n10428) );
  NOR2_X1 U12863 ( .A1(n14774), .A2(n14775), .ZN(n12757) );
  INV_X1 U12864 ( .A(n16260), .ZN(n10251) );
  AND2_X1 U12865 ( .A1(n14937), .A2(n16265), .ZN(n16260) );
  NAND2_X1 U12866 ( .A1(n12752), .A2(n10036), .ZN(n13759) );
  AND2_X1 U12867 ( .A1(n14199), .A2(n9925), .ZN(n9943) );
  INV_X1 U12868 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10520) );
  AND2_X1 U12869 ( .A1(n9936), .A2(n13803), .ZN(n9944) );
  OR2_X1 U12870 ( .A1(n17811), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9945) );
  AND2_X1 U12871 ( .A1(n13413), .A2(n13529), .ZN(n9946) );
  AND2_X1 U12872 ( .A1(n9873), .A2(n10284), .ZN(n9947) );
  AND2_X1 U12873 ( .A1(n10208), .A2(n10207), .ZN(n9948) );
  AND2_X1 U12874 ( .A1(n9875), .A2(n11124), .ZN(n9949) );
  AND2_X1 U12875 ( .A1(n9876), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U12876 ( .A(n11916), .ZN(n13773) );
  INV_X2 U12877 ( .A(n13773), .ZN(n11917) );
  INV_X1 U12878 ( .A(n10165), .ZN(n13060) );
  NOR2_X1 U12879 ( .A1(n15783), .A2(n10166), .ZN(n10165) );
  INV_X1 U12880 ( .A(n13174), .ZN(n10107) );
  NOR2_X1 U12881 ( .A1(n16086), .A2(n16085), .ZN(n9951) );
  INV_X1 U12882 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10286) );
  INV_X1 U12883 ( .A(n20108), .ZN(n20298) );
  INV_X1 U12884 ( .A(n14693), .ZN(n10391) );
  INV_X1 U12885 ( .A(n14749), .ZN(n14769) );
  INV_X1 U12886 ( .A(n14769), .ZN(n14776) );
  NOR2_X1 U12887 ( .A1(n13174), .A2(n10406), .ZN(n13469) );
  AND2_X1 U12888 ( .A1(n10408), .A2(n9874), .ZN(n13044) );
  NAND2_X1 U12889 ( .A1(n13397), .A2(n9854), .ZN(n19507) );
  AND2_X1 U12890 ( .A1(n12705), .A2(n12704), .ZN(n9952) );
  INV_X1 U12891 ( .A(n10163), .ZN(n21006) );
  NOR2_X1 U12892 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  INV_X1 U12893 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21012) );
  NAND2_X1 U12894 ( .A1(n15103), .A2(n9872), .ZN(n15074) );
  INV_X1 U12895 ( .A(n13041), .ZN(n10355) );
  INV_X1 U12896 ( .A(n11488), .ZN(n10260) );
  AND2_X1 U12897 ( .A1(n14795), .A2(n14787), .ZN(n9953) );
  INV_X1 U12898 ( .A(n14153), .ZN(n10133) );
  INV_X1 U12899 ( .A(n13668), .ZN(n10195) );
  INV_X1 U12900 ( .A(n17811), .ZN(n17933) );
  INV_X1 U12901 ( .A(n14730), .ZN(n10403) );
  INV_X1 U12902 ( .A(n12256), .ZN(n10099) );
  AND2_X1 U12903 ( .A1(n20179), .A2(n10172), .ZN(n9954) );
  INV_X1 U12904 ( .A(n14205), .ZN(n10424) );
  AND2_X1 U12905 ( .A1(n11193), .A2(n11192), .ZN(n9955) );
  AND2_X1 U12906 ( .A1(n11263), .A2(n11262), .ZN(n9956) );
  AND2_X1 U12907 ( .A1(n12705), .A2(n9889), .ZN(n9957) );
  AND2_X1 U12908 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n9958) );
  OAI21_X1 U12909 ( .B1(n10305), .B2(n17933), .A(n16523), .ZN(n10304) );
  AND2_X1 U12910 ( .A1(n12493), .A2(n10443), .ZN(n9959) );
  NOR2_X1 U12911 ( .A1(n12994), .A2(n10385), .ZN(n9960) );
  AND2_X1 U12912 ( .A1(n10411), .A2(n14772), .ZN(n9961) );
  AND2_X1 U12913 ( .A1(n10216), .A2(n10215), .ZN(n9962) );
  INV_X1 U12914 ( .A(n10185), .ZN(n12376) );
  INV_X1 U12915 ( .A(n10361), .ZN(n10360) );
  NAND2_X1 U12916 ( .A1(n10362), .A2(n14690), .ZN(n10361) );
  OR2_X1 U12917 ( .A1(n12867), .A2(n10384), .ZN(P2_U3012) );
  INV_X1 U12918 ( .A(n10888), .ZN(n11045) );
  NOR2_X1 U12919 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10888) );
  AND2_X1 U12920 ( .A1(n16512), .A2(n10297), .ZN(n9964) );
  INV_X1 U12921 ( .A(n16534), .ZN(n10202) );
  AND2_X1 U12922 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13768) );
  AND3_X1 U12923 ( .A1(n17484), .A2(n17485), .A3(P3_EAX_REG_14__SCAN_IN), .ZN(
        n9965) );
  AND2_X1 U12924 ( .A1(n15252), .A2(n10187), .ZN(n9966) );
  AND2_X1 U12925 ( .A1(n17990), .A2(n10289), .ZN(n9967) );
  NOR2_X1 U12926 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13827) );
  INV_X1 U12927 ( .A(n15235), .ZN(n10438) );
  NOR2_X1 U12928 ( .A1(n17994), .A2(n15690), .ZN(n9968) );
  AND2_X1 U12929 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9969) );
  INV_X1 U12930 ( .A(n10440), .ZN(n10439) );
  NAND2_X1 U12931 ( .A1(n9953), .A2(n14781), .ZN(n10440) );
  AND2_X1 U12932 ( .A1(n15103), .A2(n9876), .ZN(n9970) );
  AND2_X1 U12933 ( .A1(n9881), .A2(n10171), .ZN(n9971) );
  AND2_X1 U12934 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .ZN(n9972) );
  INV_X1 U12935 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n10416) );
  INV_X1 U12936 ( .A(n13826), .ZN(n20296) );
  AND2_X1 U12937 ( .A1(n17764), .A2(n10285), .ZN(n9973) );
  AND2_X1 U12938 ( .A1(n13334), .A2(n21008), .ZN(n15981) );
  AND2_X1 U12939 ( .A1(n19034), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12839) );
  INV_X1 U12940 ( .A(n12839), .ZN(n10105) );
  NAND2_X1 U12941 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n9974) );
  AND3_X1 U12942 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9975) );
  OR2_X1 U12943 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12944 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10376) );
  INV_X1 U12945 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10299) );
  INV_X1 U12946 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10290) );
  INV_X1 U12947 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10298) );
  INV_X1 U12948 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10110) );
  INV_X1 U12949 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10300) );
  INV_X1 U12950 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10336) );
  INV_X1 U12951 ( .A(n9977), .ZN(n20889) );
  NOR2_X1 U12952 ( .A1(n21101), .A2(n20379), .ZN(n9978) );
  NOR2_X1 U12953 ( .A1(n16565), .A2(n20377), .ZN(n9979) );
  NOR2_X1 U12954 ( .A1(n9978), .A2(n9979), .ZN(n9977) );
  NAND2_X1 U12955 ( .A1(n20296), .A2(n14369), .ZN(n20379) );
  OAI22_X2 U12956 ( .A1(n20372), .A2(n20377), .B1(n21054), .B2(n20379), .ZN(
        n20900) );
  NOR4_X2 U12957 ( .A1(n17812), .A2(n17930), .A3(n17811), .A4(n17945), .ZN(
        n17909) );
  AND3_X1 U12958 ( .A1(n10211), .A2(n10212), .A3(n9923), .ZN(n17812) );
  INV_X1 U12959 ( .A(n9980), .ZN(n20830) );
  NOR2_X1 U12960 ( .A1(n21369), .A2(n20379), .ZN(n9981) );
  NOR2_X1 U12961 ( .A1(n19451), .A2(n20377), .ZN(n9982) );
  NOR2_X1 U12962 ( .A1(n9981), .A2(n9982), .ZN(n9980) );
  NAND2_X1 U12963 ( .A1(n13270), .A2(n13271), .ZN(n13269) );
  NAND2_X1 U12964 ( .A1(n13248), .A2(n13247), .ZN(n13246) );
  OAI21_X1 U12965 ( .B1(n14408), .B2(n13826), .A(n10124), .ZN(P1_U2972) );
  XNOR2_X1 U12966 ( .A(n14407), .B(n14556), .ZN(n14560) );
  NAND2_X1 U12967 ( .A1(n10334), .A2(n10332), .ZN(n12655) );
  NOR2_X1 U12968 ( .A1(n16126), .A2(n16125), .ZN(n16127) );
  NOR2_X1 U12969 ( .A1(n16199), .A2(n16198), .ZN(n16197) );
  NOR2_X1 U12970 ( .A1(n15169), .A2(n12676), .ZN(n12779) );
  NOR2_X1 U12971 ( .A1(n16154), .A2(n16153), .ZN(n16152) );
  NOR2_X1 U12972 ( .A1(n16165), .A2(n16164), .ZN(n16163) );
  NOR2_X1 U12973 ( .A1(n16190), .A2(n16189), .ZN(n16188) );
  XNOR2_X1 U12974 ( .A(n10331), .B(n15064), .ZN(n16124) );
  NOR2_X1 U12975 ( .A1(n16127), .A2(n9835), .ZN(n10331) );
  NOR2_X4 U12976 ( .A1(n14964), .A2(n14962), .ZN(n14967) );
  AND2_X1 U12977 ( .A1(n10330), .A2(n14950), .ZN(n10144) );
  OR2_X2 U12978 ( .A1(n15314), .A2(n16402), .ZN(n15324) );
  OR3_X1 U12979 ( .A1(n14979), .A2(n15198), .A3(n15214), .ZN(n14980) );
  INV_X1 U12980 ( .A(n13526), .ZN(n10196) );
  NAND2_X1 U12981 ( .A1(n15145), .A2(n15144), .ZN(n15003) );
  NAND2_X1 U12982 ( .A1(n14932), .A2(n12686), .ZN(n14947) );
  NAND2_X1 U12983 ( .A1(n11806), .A2(n11805), .ZN(n11850) );
  NAND2_X2 U12984 ( .A1(n17695), .A2(n18048), .ZN(n17694) );
  NOR2_X4 U12985 ( .A1(n15708), .A2(n15707), .ZN(n17738) );
  INV_X1 U12986 ( .A(n17900), .ZN(n10203) );
  NAND2_X2 U12987 ( .A1(n17686), .A2(n16546), .ZN(n16547) );
  NOR2_X1 U12988 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13859), .ZN(
        n13965) );
  OAI22_X1 U12989 ( .A1(n13434), .A2(n13435), .B1(n9851), .B2(n9920), .ZN(
        n13436) );
  NAND2_X1 U12990 ( .A1(n9984), .A2(n10087), .ZN(n9983) );
  OAI21_X1 U12991 ( .B1(n9986), .B2(n13019), .A(n12701), .ZN(n9990) );
  OAI21_X1 U12992 ( .B1(n9986), .B2(n12708), .A(n12706), .ZN(n9992) );
  INV_X1 U12993 ( .A(n10238), .ZN(n10056) );
  NAND2_X1 U12994 ( .A1(n14873), .A2(n14874), .ZN(n10055) );
  OAI21_X2 U12995 ( .B1(n10063), .B2(n10250), .A(n10060), .ZN(n15145) );
  NAND3_X1 U12996 ( .A1(n10086), .A2(n13528), .A3(n15043), .ZN(n10069) );
  NAND2_X1 U12997 ( .A1(n10091), .A2(n11877), .ZN(n10073) );
  XNOR2_X1 U12998 ( .A(n11849), .B(n11850), .ZN(n11877) );
  INV_X1 U12999 ( .A(n13446), .ZN(n10082) );
  NOR2_X1 U13000 ( .A1(n13531), .A2(n10080), .ZN(n13675) );
  INV_X1 U13001 ( .A(n10089), .ZN(n13533) );
  NAND2_X1 U13002 ( .A1(n13528), .A2(n12509), .ZN(n10088) );
  NAND2_X1 U13003 ( .A1(n11874), .A2(n10091), .ZN(n10090) );
  XNOR2_X1 U13004 ( .A(n13277), .B(n10091), .ZN(n12868) );
  NAND2_X1 U13005 ( .A1(n12233), .A2(n10099), .ZN(n10096) );
  AND2_X2 U13006 ( .A1(n10093), .A2(n10092), .ZN(n14708) );
  NOR2_X1 U13007 ( .A1(n13174), .A2(n9935), .ZN(n13623) );
  NAND2_X1 U13008 ( .A1(n14762), .A2(n14764), .ZN(n14750) );
  NAND4_X1 U13009 ( .A1(n10121), .A2(n10114), .A3(n13876), .A4(n13873), .ZN(
        n10113) );
  NAND3_X1 U13010 ( .A1(n13872), .A2(n10117), .A3(n10116), .ZN(n10115) );
  AND2_X4 U13011 ( .A1(n13303), .A2(n13305), .ZN(n11633) );
  NAND2_X1 U13012 ( .A1(n14246), .A2(n9949), .ZN(n14297) );
  INV_X1 U13013 ( .A(n14297), .ZN(n11143) );
  OR2_X2 U13014 ( .A1(n14288), .A2(n10128), .ZN(n14189) );
  NAND2_X1 U13015 ( .A1(n13445), .A2(n13444), .ZN(n13446) );
  OR2_X2 U13016 ( .A1(n15024), .A2(n10143), .ZN(n15070) );
  NAND2_X2 U13017 ( .A1(n10146), .A2(n10145), .ZN(n14481) );
  NAND3_X1 U13018 ( .A1(n11538), .A2(n10148), .A3(n14518), .ZN(n10146) );
  NAND4_X1 U13019 ( .A1(n11655), .A2(n10152), .A3(n11582), .A4(n11657), .ZN(
        n10769) );
  INV_X1 U13020 ( .A(n10752), .ZN(n10153) );
  NAND2_X1 U13021 ( .A1(n10968), .A2(n10967), .ZN(n10985) );
  NAND3_X1 U13022 ( .A1(n10160), .A2(n10159), .A3(n15951), .ZN(n15939) );
  NAND2_X1 U13023 ( .A1(n11849), .A2(n10177), .ZN(n10176) );
  INV_X1 U13024 ( .A(n11850), .ZN(n10177) );
  AND2_X1 U13025 ( .A1(n9827), .A2(n10178), .ZN(n15496) );
  NAND2_X1 U13026 ( .A1(n15224), .A2(n16358), .ZN(n10178) );
  NAND2_X1 U13027 ( .A1(n10181), .A2(n10179), .ZN(n15224) );
  NAND3_X1 U13028 ( .A1(n9851), .A2(n9854), .A3(n13402), .ZN(n19691) );
  NAND2_X1 U13029 ( .A1(n9854), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10184) );
  NAND3_X1 U13030 ( .A1(n19250), .A2(n9854), .A3(n9851), .ZN(n14893) );
  NAND3_X1 U13031 ( .A1(n13402), .A2(n9854), .A3(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10183) );
  NAND3_X1 U13032 ( .A1(n11808), .A2(n11774), .A3(n19452), .ZN(n12382) );
  NAND3_X1 U13033 ( .A1(n10185), .A2(n12382), .A3(n12604), .ZN(n12947) );
  AND4_X2 U13034 ( .A1(n10191), .A2(n10194), .A3(n12685), .A4(n13526), .ZN(
        n14915) );
  NAND2_X1 U13035 ( .A1(n13526), .A2(n10193), .ZN(n10192) );
  NAND2_X1 U13036 ( .A1(n16412), .A2(n11778), .ZN(n10197) );
  NAND2_X1 U13037 ( .A1(n14967), .A2(n9869), .ZN(n12691) );
  NAND2_X1 U13038 ( .A1(n14967), .A2(n14966), .ZN(n14975) );
  INV_X1 U13039 ( .A(n10199), .ZN(n14954) );
  NAND2_X1 U13040 ( .A1(n15010), .A2(n14728), .ZN(n10200) );
  OR2_X1 U13041 ( .A1(n15010), .A2(n15009), .ZN(n10201) );
  OR2_X2 U13042 ( .A1(n17974), .A2(n10213), .ZN(n10211) );
  INV_X1 U13043 ( .A(n10216), .ZN(n17972) );
  INV_X1 U13044 ( .A(n15697), .ZN(n10215) );
  NOR2_X2 U13045 ( .A1(n18004), .A2(n15686), .ZN(n15689) );
  NAND3_X1 U13046 ( .A1(n10225), .A2(n9916), .A3(n10221), .ZN(n15858) );
  NAND3_X1 U13047 ( .A1(n15678), .A2(n15680), .A3(n10223), .ZN(n10222) );
  NAND3_X1 U13048 ( .A1(n10229), .A2(n10226), .A3(n9895), .ZN(P3_U2834) );
  AOI21_X1 U13049 ( .B1(n13692), .B2(n15087), .A(n13451), .ZN(n10235) );
  OAI21_X1 U13050 ( .B1(n16292), .B2(n10238), .A(n14924), .ZN(n10236) );
  NAND2_X1 U13051 ( .A1(n10237), .A2(n14912), .ZN(n15227) );
  NAND2_X1 U13052 ( .A1(n16291), .A2(n16292), .ZN(n10237) );
  NAND2_X1 U13053 ( .A1(n11888), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11852) );
  NAND3_X1 U13054 ( .A1(n10274), .A2(n11843), .A3(n11836), .ZN(n10275) );
  NAND2_X1 U13055 ( .A1(n10252), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13302) );
  AND2_X2 U13056 ( .A1(n10527), .A2(n10252), .ZN(n10697) );
  NOR2_X1 U13057 ( .A1(n13304), .A2(n10252), .ZN(n13311) );
  NAND2_X1 U13058 ( .A1(n15970), .A2(n10256), .ZN(n10254) );
  INV_X1 U13059 ( .A(n10864), .ZN(n10862) );
  MUX2_X1 U13060 ( .A(n20443), .B(n20856), .S(n11476), .Z(n13335) );
  NAND2_X1 U13061 ( .A1(n10883), .A2(n21012), .ZN(n10261) );
  XNOR2_X2 U13062 ( .A(n10811), .B(n10810), .ZN(n10883) );
  OAI21_X2 U13063 ( .B1(n14481), .B2(n10267), .A(n11531), .ZN(n14449) );
  NAND3_X1 U13064 ( .A1(n10494), .A2(n11545), .A3(n14461), .ZN(n10267) );
  NAND3_X1 U13065 ( .A1(n17990), .A2(n10289), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17922) );
  NAND3_X1 U13066 ( .A1(n16512), .A2(n10299), .A3(n10295), .ZN(n10293) );
  AND2_X2 U13067 ( .A1(n10302), .A2(n9921), .ZN(n17335) );
  NAND2_X1 U13068 ( .A1(n17675), .A2(n10307), .ZN(n10308) );
  INV_X1 U13069 ( .A(n10308), .ZN(n16486) );
  NAND2_X1 U13070 ( .A1(n17888), .A2(n17826), .ZN(n17937) );
  AND3_X2 U13071 ( .A1(n17826), .A2(n17888), .A3(n17811), .ZN(n17932) );
  OR2_X2 U13072 ( .A1(n15702), .A2(n17930), .ZN(n17888) );
  OR2_X2 U13073 ( .A1(n17770), .A2(n17757), .ZN(n10312) );
  NAND2_X1 U13074 ( .A1(n15690), .A2(n10315), .ZN(n10313) );
  OAI21_X2 U13075 ( .B1(n17995), .B2(n10314), .A(n10313), .ZN(n17987) );
  NAND3_X1 U13076 ( .A1(n15619), .A2(n15624), .A3(n10316), .ZN(n15684) );
  NAND2_X1 U13077 ( .A1(n12403), .A2(n10319), .ZN(n12385) );
  NAND2_X1 U13078 ( .A1(n10320), .A2(n10321), .ZN(n15025) );
  NAND2_X1 U13079 ( .A1(n15136), .A2(n9870), .ZN(n10320) );
  AOI21_X1 U13080 ( .B1(n9857), .B2(n10323), .A(n10322), .ZN(n10321) );
  NOR2_X2 U13081 ( .A1(n15123), .A2(n15124), .ZN(n15122) );
  AOI21_X2 U13082 ( .B1(n15070), .B2(n15027), .A(n15068), .ZN(n15062) );
  OAI21_X2 U13083 ( .B1(n15044), .B2(n15087), .A(n19208), .ZN(n14911) );
  NOR3_X1 U13084 ( .A1(n15161), .A2(n14980), .A3(n15177), .ZN(n10330) );
  INV_X1 U13085 ( .A(n12659), .ZN(n10334) );
  NAND2_X1 U13086 ( .A1(n15103), .A2(n9950), .ZN(n12649) );
  NAND3_X1 U13087 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12670) );
  AOI21_X1 U13088 ( .B1(n19075), .B2(n10345), .A(n9835), .ZN(n10344) );
  AOI22_X1 U13089 ( .A1(n19075), .A2(n10343), .B1(n9835), .B2(n15180), .ZN(
        n10342) );
  NAND2_X2 U13090 ( .A1(n10346), .A2(n11887), .ZN(n12695) );
  NAND2_X1 U13091 ( .A1(n9922), .A2(n12705), .ZN(n13101) );
  NOR2_X1 U13092 ( .A1(n14718), .A2(n14709), .ZN(n10363) );
  OR3_X1 U13093 ( .A1(n14718), .A2(n10361), .A3(n14709), .ZN(n14692) );
  NOR2_X1 U13094 ( .A1(n10748), .A2(n11586), .ZN(n10365) );
  INV_X1 U13095 ( .A(n10749), .ZN(n10364) );
  NAND2_X1 U13096 ( .A1(n10369), .A2(n11531), .ZN(n10368) );
  NAND2_X1 U13097 ( .A1(n9820), .A2(n10374), .ZN(n10373) );
  NAND2_X2 U13098 ( .A1(n10381), .A2(n14449), .ZN(n14392) );
  NAND2_X1 U13099 ( .A1(n14481), .A2(n9867), .ZN(n11542) );
  XNOR2_X2 U13100 ( .A(n10879), .B(n10880), .ZN(n13339) );
  NAND2_X1 U13101 ( .A1(n13363), .A2(n12839), .ZN(n11867) );
  CLKBUF_X1 U13102 ( .A(n13363), .Z(n10383) );
  NAND2_X1 U13103 ( .A1(n14708), .A2(n10394), .ZN(n10393) );
  NAND2_X1 U13104 ( .A1(n10392), .A2(n10387), .ZN(n12323) );
  AOI21_X1 U13105 ( .B1(n14708), .B2(n10388), .A(n12296), .ZN(n10387) );
  OAI21_X1 U13106 ( .B1(n10092), .B2(n14699), .A(n10393), .ZN(n14694) );
  NAND3_X1 U13107 ( .A1(n10396), .A2(n11882), .A3(n11883), .ZN(n12990) );
  NAND2_X1 U13108 ( .A1(n11871), .A2(n11870), .ZN(n11883) );
  INV_X1 U13109 ( .A(n12164), .ZN(n10401) );
  INV_X1 U13110 ( .A(n12187), .ZN(n10404) );
  NAND2_X1 U13111 ( .A1(n13005), .A2(n10409), .ZN(n10408) );
  NAND4_X4 U13112 ( .A1(n10741), .A2(n10739), .A3(n10742), .A4(n10740), .ZN(
        n13496) );
  AND2_X2 U13113 ( .A1(n13496), .A2(n13599), .ZN(n11584) );
  INV_X1 U13114 ( .A(n10428), .ZN(n14309) );
  INV_X1 U13115 ( .A(n13804), .ZN(n10429) );
  INV_X2 U13116 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13801) );
  INV_X2 U13117 ( .A(n12582), .ZN(n12567) );
  NAND2_X1 U13118 ( .A1(n14804), .A2(n10439), .ZN(n15234) );
  NAND2_X1 U13119 ( .A1(n14804), .A2(n9880), .ZN(n10436) );
  AND2_X1 U13120 ( .A1(n14804), .A2(n9953), .ZN(n14789) );
  AND2_X1 U13121 ( .A1(n14804), .A2(n14795), .ZN(n14797) );
  NAND3_X1 U13122 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(n16119) );
  NAND2_X1 U13123 ( .A1(n15354), .A2(n10455), .ZN(n14815) );
  NOR2_X1 U13124 ( .A1(n10464), .A2(n10744), .ZN(n11559) );
  NOR2_X1 U13125 ( .A1(n11565), .A2(n10464), .ZN(n11573) );
  NAND2_X1 U13126 ( .A1(n10693), .A2(n11468), .ZN(n10464) );
  INV_X1 U13127 ( .A(n10795), .ZN(n10471) );
  NAND2_X1 U13128 ( .A1(n10465), .A2(n10795), .ZN(n13325) );
  NAND2_X1 U13129 ( .A1(n10855), .A2(n10788), .ZN(n10465) );
  NAND3_X1 U13130 ( .A1(n10470), .A2(n10468), .A3(n10466), .ZN(n13137) );
  NAND2_X1 U13131 ( .A1(n10795), .A2(n10467), .ZN(n10466) );
  INV_X1 U13132 ( .A(n10788), .ZN(n10467) );
  NAND2_X1 U13133 ( .A1(n10469), .A2(n10795), .ZN(n10468) );
  INV_X1 U13134 ( .A(n10855), .ZN(n10469) );
  NAND3_X1 U13135 ( .A1(n10471), .A2(n10855), .A3(n10788), .ZN(n10470) );
  OAI22_X2 U13136 ( .A1(n13137), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11477), 
        .B2(n10895), .ZN(n10808) );
  NAND2_X1 U13137 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U13138 ( .A1(n11012), .A2(n9944), .ZN(n11050) );
  INV_X1 U13139 ( .A(n14137), .ZN(n10488) );
  INV_X1 U13140 ( .A(n13017), .ZN(n12705) );
  NAND2_X1 U13141 ( .A1(n12700), .A2(n12699), .ZN(n13017) );
  NAND2_X1 U13142 ( .A1(n15236), .A2(n10438), .ZN(n15240) );
  NAND2_X1 U13143 ( .A1(n14727), .A2(n14719), .ZN(n14718) );
  NAND2_X1 U13144 ( .A1(n13007), .A2(n13006), .ZN(n13005) );
  AND2_X1 U13145 ( .A1(n9885), .A2(n13102), .ZN(n19193) );
  NAND2_X1 U13146 ( .A1(n16133), .A2(n19251), .ZN(n16134) );
  NAND2_X1 U13147 ( .A1(n12990), .A2(n11883), .ZN(n13007) );
  AND2_X1 U13148 ( .A1(n13348), .A2(n13299), .ZN(n19150) );
  CLKBUF_X1 U13149 ( .A(n14750), .Z(n14763) );
  AND2_X2 U13150 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13828) );
  NAND2_X1 U13151 ( .A1(n11771), .A2(n16412), .ZN(n11772) );
  NAND2_X1 U13152 ( .A1(n11764), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11773) );
  AOI22_X1 U13153 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U13154 ( .A1(n12990), .A2(n12989), .ZN(n20065) );
  OR2_X1 U13155 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  OAI21_X1 U13156 ( .B1(n14321), .B2(n14318), .A(n11458), .ZN(P1_U2843) );
  NOR2_X1 U13157 ( .A1(n11453), .A2(n13089), .ZN(n11437) );
  AOI21_X2 U13158 ( .B1(n11310), .B2(n14124), .A(n11650), .ZN(n14390) );
  INV_X1 U13159 ( .A(n10668), .ZN(n10756) );
  NAND2_X1 U13160 ( .A1(n11791), .A2(n11861), .ZN(n11774) );
  XNOR2_X1 U13161 ( .A(n10966), .B(n10967), .ZN(n11497) );
  XNOR2_X1 U13162 ( .A(n12323), .B(n12322), .ZN(n14105) );
  NAND2_X1 U13163 ( .A1(n15488), .A2(n15472), .ZN(n16342) );
  NAND2_X1 U13164 ( .A1(n9846), .A2(n13801), .ZN(n11833) );
  INV_X1 U13165 ( .A(n13612), .ZN(n13613) );
  NAND2_X1 U13166 ( .A1(n10943), .A2(n10911), .ZN(n13568) );
  XNOR2_X1 U13167 ( .A(n10943), .B(n10941), .ZN(n11489) );
  NAND2_X1 U13168 ( .A1(n11586), .A2(n13579), .ZN(n10747) );
  AOI21_X1 U13169 ( .B1(n14106), .B2(n15981), .A(n14066), .ZN(n14067) );
  NAND2_X1 U13170 ( .A1(n14106), .A2(n11665), .ZN(n11683) );
  NAND2_X2 U13171 ( .A1(n14380), .A2(n13082), .ZN(n14382) );
  NOR2_X1 U13172 ( .A1(n20654), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10492) );
  INV_X1 U13173 ( .A(n12399), .ZN(n12580) );
  INV_X1 U13174 ( .A(n12494), .ZN(n12131) );
  AND2_X1 U13175 ( .A1(n17399), .A2(n18400), .ZN(n17396) );
  AND2_X1 U13176 ( .A1(n12403), .A2(n20079), .ZN(n10493) );
  AND2_X1 U13177 ( .A1(n16001), .A2(n14613), .ZN(n10494) );
  OR2_X1 U13178 ( .A1(n21191), .A2(n20211), .ZN(n10495) );
  OR2_X1 U13179 ( .A1(n20211), .A2(n21195), .ZN(n10496) );
  OR2_X1 U13180 ( .A1(n13868), .A2(n15630), .ZN(n10497) );
  NOR2_X1 U13181 ( .A1(n20140), .A2(n20160), .ZN(n10498) );
  AND3_X1 U13182 ( .A1(n11920), .A2(n11919), .A3(n11918), .ZN(n10499) );
  NOR2_X1 U13183 ( .A1(n13857), .A2(n13856), .ZN(n15611) );
  INV_X1 U13184 ( .A(n10868), .ZN(n11295) );
  INV_X2 U13185 ( .A(n19020), .ZN(n18999) );
  INV_X2 U13186 ( .A(n13821), .ZN(n20291) );
  INV_X1 U13187 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13451) );
  AND3_X1 U13188 ( .A1(n15632), .A2(n10497), .A3(n15631), .ZN(n10500) );
  INV_X2 U13189 ( .A(n20100), .ZN(n20036) );
  NAND2_X1 U13190 ( .A1(n11917), .A2(n16412), .ZN(n10501) );
  AND2_X1 U13191 ( .A1(n11838), .A2(n11837), .ZN(n10502) );
  OR2_X1 U13192 ( .A1(n15848), .A2(n16507), .ZN(n10503) );
  INV_X1 U13193 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15673) );
  INV_X1 U13194 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12668) );
  OR2_X1 U13195 ( .A1(n19334), .A2(n19366), .ZN(n19333) );
  AND2_X1 U13196 ( .A1(n16484), .A2(n16487), .ZN(n10504) );
  OR2_X1 U13197 ( .A1(n12060), .A2(n12059), .ZN(n10505) );
  INV_X1 U13198 ( .A(n15640), .ZN(n17538) );
  INV_X1 U13199 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13200 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17480), .ZN(n17475) );
  INV_X1 U13201 ( .A(n17475), .ZN(n17444) );
  OR2_X1 U13202 ( .A1(n17811), .A2(n15762), .ZN(n10506) );
  AND2_X1 U13203 ( .A1(n16185), .A2(n15087), .ZN(n10507) );
  NAND2_X1 U13204 ( .A1(n10881), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11042) );
  AND3_X1 U13205 ( .A1(n12330), .A2(n12329), .A3(n12328), .ZN(n10508) );
  INV_X1 U13206 ( .A(n13558), .ZN(n20322) );
  INV_X4 U13207 ( .A(n17302), .ZN(n17351) );
  INV_X1 U13208 ( .A(n12435), .ZN(n12415) );
  INV_X1 U13209 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19257) );
  OR2_X1 U13210 ( .A1(n18970), .A2(n18029), .ZN(n19006) );
  OR2_X1 U13211 ( .A1(n18029), .A2(n17998), .ZN(n17802) );
  AND2_X1 U13212 ( .A1(n11715), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10509) );
  AND2_X1 U13213 ( .A1(n11777), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10510) );
  AND2_X1 U13214 ( .A1(n13426), .A2(n13425), .ZN(n10511) );
  AND2_X1 U13215 ( .A1(n12229), .A2(n12252), .ZN(n10512) );
  OR2_X1 U13216 ( .A1(n12212), .A2(n12211), .ZN(n10514) );
  AND4_X1 U13217 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10515) );
  AND2_X1 U13218 ( .A1(n10625), .A2(n10624), .ZN(n10516) );
  AND4_X1 U13219 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10517) );
  INV_X1 U13220 ( .A(n11558), .ZN(n10753) );
  NOR3_X1 U13221 ( .A1(n13438), .A2(n13437), .A3(n13436), .ZN(n13439) );
  OR2_X1 U13222 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11313), .ZN(
        n11312) );
  OR2_X1 U13223 ( .A1(n10931), .A2(n10930), .ZN(n11507) );
  AOI22_X1 U13224 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U13225 ( .A1(n13443), .A2(n12403), .ZN(n13444) );
  AND2_X1 U13226 ( .A1(n16415), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12343) );
  XNOR2_X1 U13227 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11321) );
  BUF_X1 U13228 ( .A(n10697), .Z(n11623) );
  OR2_X1 U13229 ( .A1(n10586), .A2(n10585), .ZN(n11287) );
  INV_X1 U13230 ( .A(n14300), .ZN(n11142) );
  OR2_X1 U13231 ( .A1(n10953), .A2(n10952), .ZN(n11506) );
  NAND2_X1 U13232 ( .A1(n11365), .A2(n10762), .ZN(n11589) );
  NAND2_X1 U13233 ( .A1(n10745), .A2(n13157), .ZN(n10746) );
  NAND2_X1 U13234 ( .A1(n11678), .A2(n10696), .ZN(n10744) );
  NOR2_X1 U13235 ( .A1(n16482), .A2(n15837), .ZN(n16483) );
  OR2_X1 U13236 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20353), .ZN(
        n11319) );
  INV_X1 U13237 ( .A(n14177), .ZN(n11275) );
  AND2_X1 U13238 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11214), .ZN(
        n11248) );
  INV_X1 U13239 ( .A(n14302), .ZN(n11124) );
  INV_X1 U13240 ( .A(n10993), .ZN(n10994) );
  OR2_X1 U13241 ( .A1(n10848), .A2(n10847), .ZN(n11467) );
  INV_X1 U13242 ( .A(n10895), .ZN(n11525) );
  AND4_X1 U13243 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  AND2_X1 U13244 ( .A1(n16427), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U13245 ( .A1(n13589), .A2(n13157), .ZN(n11363) );
  AND2_X1 U13246 ( .A1(n11320), .A2(n11319), .ZN(n11557) );
  INV_X1 U13247 ( .A(n11295), .ZN(n11258) );
  AND2_X1 U13248 ( .A1(n10665), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11284) );
  NOR2_X1 U13249 ( .A1(n11155), .A2(n11156), .ZN(n11161) );
  INV_X1 U13250 ( .A(n10963), .ZN(n10964) );
  AND2_X1 U13251 ( .A1(n10811), .A2(n10809), .ZN(n10852) );
  AND2_X1 U13252 ( .A1(n12232), .A2(n10512), .ZN(n12233) );
  AND2_X1 U13253 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  INV_X1 U13254 ( .A(n12577), .ZN(n12570) );
  NAND2_X1 U13255 ( .A1(n12253), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11880) );
  INV_X1 U13256 ( .A(n17144), .ZN(n15612) );
  NAND2_X1 U13257 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n15631) );
  INV_X1 U13258 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14023) );
  INV_X1 U13259 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17128) );
  NOR2_X1 U13260 ( .A1(n15797), .A2(n11363), .ZN(n13148) );
  OAI211_X1 U13261 ( .C1(n13581), .C2(n12637), .A(n10794), .B(n10793), .ZN(
        n10795) );
  NOR2_X1 U13262 ( .A1(n10695), .A2(n20625), .ZN(n10868) );
  OR2_X1 U13263 ( .A1(n13489), .A2(n14048), .ZN(n13491) );
  OR2_X1 U13264 ( .A1(n11648), .A2(n14116), .ZN(n13489) );
  NAND2_X1 U13265 ( .A1(n11284), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11299) );
  INV_X1 U13266 ( .A(n11196), .ZN(n11214) );
  INV_X1 U13267 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U13268 ( .A1(n10965), .A2(n10964), .ZN(n13353) );
  INV_X1 U13269 ( .A(n11042), .ZN(n11117) );
  NAND2_X1 U13270 ( .A1(n10894), .A2(n10893), .ZN(n20477) );
  INV_X1 U13271 ( .A(n20365), .ZN(n20373) );
  INV_X1 U13272 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15148) );
  INV_X1 U13273 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12672) );
  INV_X1 U13274 ( .A(n13018), .ZN(n12704) );
  OR2_X1 U13275 ( .A1(n12020), .A2(n12019), .ZN(n12574) );
  NOR2_X1 U13276 ( .A1(n13294), .A2(n13293), .ZN(n11987) );
  INV_X1 U13277 ( .A(n13103), .ZN(n11927) );
  OR2_X1 U13278 ( .A1(n12252), .A2(n12257), .ZN(n12291) );
  AND2_X1 U13279 ( .A1(n12206), .A2(n12205), .ZN(n12209) );
  AND2_X1 U13280 ( .A1(n12584), .A2(n12583), .ZN(n12769) );
  AND3_X1 U13281 ( .A1(n16433), .A2(n12920), .A3(n12802), .ZN(n12393) );
  INV_X1 U13282 ( .A(n15103), .ZN(n15116) );
  INV_X1 U13283 ( .A(n15089), .ZN(n15088) );
  NOR2_X1 U13284 ( .A1(n16390), .A2(n15246), .ZN(n15439) );
  AND2_X1 U13285 ( .A1(n12923), .A2(n12386), .ZN(n16431) );
  AOI21_X1 U13286 ( .B1(n12868), .B2(n12839), .A(n11879), .ZN(n12996) );
  INV_X1 U13287 ( .A(n19542), .ZN(n19546) );
  AOI22_X1 U13288 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18823), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n13850), .ZN(n15570) );
  AOI21_X1 U13289 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15723) );
  OR2_X1 U13290 ( .A1(n18808), .A2(n15573), .ZN(n15562) );
  NOR2_X1 U13291 ( .A1(n13851), .A2(n13856), .ZN(n15625) );
  OR2_X1 U13292 ( .A1(n9914), .A2(n16482), .ZN(n16485) );
  NAND2_X1 U13293 ( .A1(n17933), .A2(n18058), .ZN(n15713) );
  NOR2_X1 U13294 ( .A1(n17738), .A2(n18140), .ZN(n17757) );
  NOR2_X1 U13295 ( .A1(n18200), .A2(n17866), .ZN(n17845) );
  NAND2_X1 U13296 ( .A1(n18353), .A2(n18833), .ZN(n18204) );
  OR2_X1 U13297 ( .A1(n17533), .A2(n15745), .ZN(n15742) );
  INV_X1 U13298 ( .A(n15768), .ZN(n15566) );
  INV_X2 U13299 ( .A(n15609), .ZN(n17352) );
  NOR2_X1 U13300 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13848) );
  INV_X1 U13301 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14232) );
  INV_X1 U13302 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14250) );
  INV_X1 U13303 ( .A(n20123), .ZN(n20160) );
  AND2_X1 U13304 ( .A1(n13494), .A2(n21346), .ZN(n13500) );
  AND2_X2 U13305 ( .A1(n13589), .A2(n13496), .ZN(n11453) );
  NOR2_X1 U13306 ( .A1(n11191), .A2(n14232), .ZN(n11195) );
  AND2_X1 U13307 ( .A1(n11078), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U13308 ( .A1(n11007), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U13309 ( .A1(n20108), .A2(n12638), .ZN(n13821) );
  AOI21_X1 U13310 ( .B1(n20303), .B2(n20322), .A(n13561), .ZN(n16081) );
  AND2_X1 U13311 ( .A1(n20448), .A2(n20447), .ZN(n20452) );
  INV_X1 U13312 ( .A(n20799), .ZN(n20531) );
  INV_X1 U13313 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20625) );
  INV_X1 U13314 ( .A(n20559), .ZN(n20694) );
  INV_X1 U13315 ( .A(n13339), .ZN(n13570) );
  NAND2_X1 U13316 ( .A1(n20296), .A2(n13577), .ZN(n20377) );
  OR2_X1 U13317 ( .A1(n11558), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21011) );
  AND2_X1 U13318 ( .A1(n12392), .A2(n12824), .ZN(n12920) );
  AND2_X1 U13319 ( .A1(n12592), .A2(n12591), .ZN(n14812) );
  INV_X1 U13320 ( .A(n13762), .ZN(n12675) );
  XNOR2_X1 U13321 ( .A(n12649), .B(n15054), .ZN(n15053) );
  INV_X1 U13322 ( .A(n12987), .ZN(n11882) );
  NAND2_X1 U13323 ( .A1(n19282), .A2(n12622), .ZN(n13264) );
  NAND2_X1 U13324 ( .A1(n15033), .A2(n9887), .ZN(n15034) );
  AND2_X1 U13325 ( .A1(n19056), .A2(n14982), .ZN(n15175) );
  AND3_X1 U13326 ( .A1(n12407), .A2(n12406), .A3(n12405), .ZN(n16315) );
  NOR2_X1 U13327 ( .A1(n15042), .A2(n15043), .ZN(n15050) );
  INV_X1 U13328 ( .A(n16399), .ZN(n16364) );
  AND2_X1 U13329 ( .A1(n13542), .A2(n13541), .ZN(n16390) );
  NAND2_X1 U13330 ( .A1(n16465), .A2(n19034), .ZN(n13205) );
  INV_X1 U13331 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13767) );
  INV_X1 U13332 ( .A(n20057), .ZN(n19861) );
  INV_X1 U13333 ( .A(n20053), .ZN(n19537) );
  INV_X1 U13334 ( .A(n19820), .ZN(n13287) );
  NOR2_X1 U13335 ( .A1(n15721), .A2(n15723), .ZN(n16648) );
  NOR2_X1 U13336 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16881), .ZN(n16868) );
  NOR2_X1 U13337 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16909), .ZN(n16890) );
  INV_X1 U13338 ( .A(n17051), .ZN(n17044) );
  INV_X1 U13339 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17221) );
  INV_X1 U13340 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17148) );
  NAND2_X1 U13341 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17688), .ZN(
        n17662) );
  NOR2_X1 U13342 ( .A1(n10286), .A2(n16807), .ZN(n16682) );
  NOR2_X1 U13343 ( .A1(n16830), .A2(n16843), .ZN(n17775) );
  NAND2_X1 U13344 ( .A1(n16485), .A2(n10504), .ZN(n16492) );
  AOI21_X1 U13345 ( .B1(n10202), .B2(n16536), .A(n16535), .ZN(n18097) );
  AOI21_X1 U13346 ( .B1(n15767), .B2(n10113), .A(n15766), .ZN(n18807) );
  INV_X1 U13347 ( .A(n18813), .ZN(n18818) );
  INV_X1 U13348 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17930) );
  NOR2_X1 U13349 ( .A1(n15579), .A2(n15578), .ZN(n15735) );
  INV_X1 U13350 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U13351 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17241), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13867) );
  NOR2_X1 U13352 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21018) );
  NOR2_X1 U13353 ( .A1(n14065), .A2(n16101), .ZN(n13492) );
  INV_X1 U13354 ( .A(n20133), .ZN(n20155) );
  INV_X1 U13355 ( .A(n13145), .ZN(n15776) );
  OAI21_X1 U13356 ( .B1(n14527), .B2(n14312), .A(n10496), .ZN(n12633) );
  INV_X1 U13357 ( .A(n11676), .ZN(n14362) );
  INV_X1 U13358 ( .A(n20289), .ZN(n20283) );
  NAND2_X1 U13359 ( .A1(n11195), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11196) );
  NAND2_X1 U13360 ( .A1(n11139), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11155) );
  AND2_X1 U13361 ( .A1(n13845), .A2(n13844), .ZN(n15964) );
  NOR2_X1 U13362 ( .A1(n10913), .A2(n10663), .ZN(n10934) );
  NOR2_X1 U13363 ( .A1(n16081), .A2(n13560), .ZN(n16044) );
  INV_X2 U13364 ( .A(n20342), .ZN(n20317) );
  INV_X1 U13365 ( .A(n16055), .ZN(n20327) );
  NAND2_X1 U13366 ( .A1(n21012), .A2(n13578), .ZN(n20483) );
  INV_X1 U13367 ( .A(n15825), .ZN(n20987) );
  OAI22_X1 U13368 ( .A1(n13584), .A2(n13583), .B1(n20479), .B2(n20598), .ZN(
        n20380) );
  NOR2_X2 U13369 ( .A1(n20455), .A2(n20476), .ZN(n20407) );
  OAI21_X1 U13370 ( .B1(n20426), .B2(n20985), .A(n20415), .ZN(n20439) );
  NOR2_X2 U13371 ( .A1(n20455), .A2(n20531), .ZN(n20471) );
  NOR2_X2 U13372 ( .A1(n20455), .A2(n20694), .ZN(n20501) );
  NOR2_X2 U13373 ( .A1(n20532), .A2(n20772), .ZN(n20554) );
  NOR2_X2 U13374 ( .A1(n20532), .A2(n20531), .ZN(n20589) );
  INV_X1 U13375 ( .A(n20599), .ZN(n20621) );
  INV_X1 U13376 ( .A(n20476), .ZN(n20593) );
  NOR2_X2 U13377 ( .A1(n20695), .A2(n20772), .ZN(n20681) );
  INV_X1 U13378 ( .A(n20695), .ZN(n20650) );
  NOR2_X2 U13379 ( .A1(n20695), .A2(n20694), .ZN(n20760) );
  NOR2_X1 U13380 ( .A1(n20483), .A2(n20260), .ZN(n20822) );
  AND2_X1 U13381 ( .A1(n15782), .A2(n15789), .ZN(n15817) );
  INV_X1 U13382 ( .A(n21011), .ZN(n15849) );
  AND2_X1 U13383 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20972), .ZN(n20951) );
  OAI21_X1 U13384 ( .B1(n20092), .B2(n12829), .A(n12828), .ZN(n12925) );
  NAND2_X1 U13385 ( .A1(n16135), .A2(n16134), .ZN(n16136) );
  INV_X1 U13386 ( .A(n19247), .ZN(n19233) );
  INV_X1 U13387 ( .A(n19217), .ZN(n19185) );
  AND2_X1 U13388 ( .A1(n12768), .A2(n12693), .ZN(n19247) );
  OAI21_X1 U13389 ( .B1(n12878), .B2(n12677), .A(n16104), .ZN(n19189) );
  INV_X1 U13390 ( .A(n19953), .ZN(n19226) );
  INV_X1 U13391 ( .A(n19185), .ZN(n19245) );
  OR2_X1 U13392 ( .A1(n12034), .A2(n12033), .ZN(n13476) );
  AND3_X1 U13393 ( .A1(n11974), .A2(n11973), .A3(n11972), .ZN(n13294) );
  OR2_X1 U13394 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  OR2_X1 U13395 ( .A1(n12084), .A2(n12083), .ZN(n14772) );
  OR2_X1 U13396 ( .A1(n12046), .A2(n12045), .ZN(n13622) );
  INV_X1 U13397 ( .A(n19289), .ZN(n19294) );
  AND2_X1 U13398 ( .A1(n19282), .A2(n11744), .ZN(n19318) );
  INV_X1 U13399 ( .A(n12403), .ZN(n13000) );
  INV_X1 U13400 ( .A(n19408), .ZN(n19383) );
  INV_X1 U13401 ( .A(n15474), .ZN(n19170) );
  INV_X1 U13402 ( .A(n19423), .ZN(n16270) );
  INV_X1 U13403 ( .A(n15436), .ZN(n19128) );
  NOR2_X2 U13404 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U13405 ( .A1(n13205), .A2(n13204), .ZN(n19863) );
  NOR2_X1 U13406 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13836) );
  INV_X1 U13407 ( .A(n19486), .ZN(n19503) );
  AND2_X1 U13408 ( .A1(n20065), .A2(n13276), .ZN(n19477) );
  AND2_X1 U13409 ( .A1(n19623), .A2(n20053), .ZN(n19562) );
  AND2_X1 U13410 ( .A1(n19623), .A2(n19830), .ZN(n19618) );
  AND2_X1 U13411 ( .A1(n19654), .A2(n19830), .ZN(n19649) );
  INV_X1 U13412 ( .A(n19653), .ZN(n19680) );
  AND2_X1 U13413 ( .A1(n15526), .A2(n19322), .ZN(n19654) );
  INV_X1 U13414 ( .A(n19724), .ZN(n19728) );
  INV_X1 U13415 ( .A(n19863), .ZN(n19826) );
  OAI21_X1 U13416 ( .B1(n19814), .B2(n20079), .A(n19795), .ZN(n19816) );
  INV_X1 U13417 ( .A(n19789), .ZN(n19830) );
  NOR2_X2 U13418 ( .A1(n13287), .A2(n19659), .ZN(n19942) );
  XOR2_X1 U13419 ( .A(n10113), .B(n16997), .Z(n19024) );
  NOR2_X1 U13420 ( .A1(n18800), .A2(n17588), .ZN(n19009) );
  NOR2_X1 U13421 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16771), .ZN(n16755) );
  NOR2_X1 U13422 ( .A1(n18921), .A2(n16799), .ZN(n16800) );
  NOR2_X1 U13423 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16838), .ZN(n16818) );
  NOR2_X1 U13424 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16915), .ZN(n16914) );
  NOR2_X1 U13425 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16959), .ZN(n16927) );
  INV_X1 U13426 ( .A(n17045), .ZN(n17023) );
  INV_X1 U13427 ( .A(n17019), .ZN(n17037) );
  NOR2_X1 U13428 ( .A1(n16790), .A2(n17158), .ZN(n17126) );
  INV_X1 U13429 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16910) );
  AOI21_X1 U13430 ( .B1(n15764), .B2(n15582), .A(n13959), .ZN(n15854) );
  NOR2_X1 U13431 ( .A1(n17596), .A2(n17469), .ZN(n17464) );
  INV_X1 U13432 ( .A(n17530), .ZN(n17537) );
  INV_X1 U13433 ( .A(n17588), .ZN(n17589) );
  INV_X1 U13434 ( .A(n18095), .ZN(n18100) );
  NOR2_X1 U13435 ( .A1(n17920), .A2(n16534), .ZN(n17822) );
  NOR2_X1 U13436 ( .A1(n17868), .A2(n17858), .ZN(n17852) );
  NOR2_X1 U13437 ( .A1(n15761), .A2(n17929), .ZN(n17887) );
  NAND2_X1 U13438 ( .A1(n18028), .A2(n17989), .ZN(n17953) );
  NOR2_X1 U13439 ( .A1(n18097), .A2(n18351), .ZN(n18110) );
  INV_X1 U13440 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18164) );
  OAI21_X2 U13441 ( .B1(n18808), .B2(n15768), .A(n18807), .ZN(n18813) );
  INV_X1 U13442 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18237) );
  NOR2_X2 U13443 ( .A1(n17518), .A2(n18361), .ZN(n18253) );
  INV_X1 U13444 ( .A(n18339), .ZN(n18297) );
  AOI21_X2 U13445 ( .B1(n15735), .B2(n15734), .A(n18847), .ZN(n18334) );
  INV_X1 U13446 ( .A(n18715), .ZN(n18455) );
  NOR2_X1 U13447 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18960), .ZN(
        n18982) );
  INV_X1 U13448 ( .A(n19005), .ZN(n18847) );
  INV_X1 U13449 ( .A(n18743), .ZN(n18738) );
  INV_X1 U13450 ( .A(n18407), .ZN(n18473) );
  INV_X1 U13451 ( .A(n18477), .ZN(n18541) );
  INV_X1 U13452 ( .A(n18523), .ZN(n18585) );
  INV_X1 U13453 ( .A(n18545), .ZN(n18609) );
  INV_X1 U13454 ( .A(n18567), .ZN(n18633) );
  INV_X1 U13455 ( .A(n18589), .ZN(n18655) );
  INV_X1 U13456 ( .A(n18614), .ZN(n18677) );
  INV_X1 U13457 ( .A(n18637), .ZN(n18706) );
  AND2_X1 U13458 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18745), .ZN(n18774) );
  AND2_X1 U13459 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18745), .ZN(n18789) );
  INV_X1 U13460 ( .A(n19013), .ZN(n19007) );
  INV_X1 U13461 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18883) );
  NAND2_X2 U13462 ( .A1(n11675), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14369)
         );
  INV_X1 U13463 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21346) );
  INV_X1 U13464 ( .A(n20186), .ZN(n20174) );
  NAND2_X1 U13465 ( .A1(n20161), .A2(n13492), .ZN(n20133) );
  INV_X1 U13466 ( .A(n12633), .ZN(n12634) );
  INV_X1 U13467 ( .A(n20212), .ZN(n20243) );
  AND2_X1 U13468 ( .A1(n13115), .A2(n13114), .ZN(n20357) );
  OR2_X1 U13469 ( .A1(n20286), .A2(n13496), .ZN(n20245) );
  OR2_X1 U13470 ( .A1(n13060), .A2(n13059), .ZN(n20289) );
  OR2_X2 U13471 ( .A1(n20291), .A2(n13096), .ZN(n20302) );
  NAND2_X2 U13472 ( .A1(n15817), .A2(n20107), .ZN(n20108) );
  INV_X1 U13473 ( .A(n20332), .ZN(n20340) );
  OAI21_X1 U13474 ( .B1(n13331), .B2(n13330), .A(n20483), .ZN(n20352) );
  AOI21_X1 U13475 ( .B1(n13576), .B2(n13583), .A(n13575), .ZN(n20384) );
  OR2_X1 U13476 ( .A1(n20455), .A2(n20772), .ZN(n20437) );
  AOI22_X1 U13477 ( .A1(n20414), .A2(n20412), .B1(n20656), .B2(n10492), .ZN(
        n20442) );
  AOI22_X1 U13478 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20450), .B1(n20453), 
        .B2(n20449), .ZN(n20475) );
  NAND2_X1 U13479 ( .A1(n20560), .A2(n20593), .ZN(n20529) );
  AOI22_X1 U13480 ( .A1(n20537), .A2(n20534), .B1(n10492), .B2(n20722), .ZN(
        n20558) );
  NAND2_X1 U13481 ( .A1(n20560), .A2(n20559), .ZN(n20599) );
  NAND2_X1 U13482 ( .A1(n20650), .A2(n20593), .ZN(n20649) );
  AOI22_X1 U13483 ( .A1(n20661), .A2(n20657), .B1(n20656), .B2(n20655), .ZN(
        n20686) );
  NAND2_X1 U13484 ( .A1(n20650), .A2(n20799), .ZN(n20715) );
  INV_X1 U13485 ( .A(n20805), .ZN(n20852) );
  INV_X1 U13486 ( .A(n20892), .ZN(n20751) );
  NAND2_X1 U13487 ( .A1(n20716), .A2(n13339), .ZN(n20798) );
  INV_X1 U13488 ( .A(n20880), .ZN(n20827) );
  INV_X1 U13489 ( .A(n20910), .ZN(n20846) );
  NAND2_X1 U13490 ( .A1(n20800), .A2(n20559), .ZN(n20904) );
  OR2_X1 U13491 ( .A1(n20917), .A2(n21012), .ZN(n15829) );
  INV_X1 U13492 ( .A(n20984), .ZN(n20980) );
  INV_X1 U13493 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20936) );
  NAND2_X1 U13494 ( .A1(n12921), .A2(n12830), .ZN(n12878) );
  INV_X1 U13495 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19627) );
  INV_X1 U13496 ( .A(n19251), .ZN(n19232) );
  INV_X1 U13497 ( .A(n19249), .ZN(n19230) );
  NAND2_X1 U13498 ( .A1(n12993), .A2(n12992), .ZN(n14749) );
  AND2_X1 U13499 ( .A1(n19270), .A2(n19269), .ZN(n19289) );
  INV_X1 U13500 ( .A(n19285), .ZN(n19325) );
  NAND2_X1 U13501 ( .A1(n19334), .A2(n14671), .ZN(n19327) );
  INV_X1 U13502 ( .A(n19334), .ZN(n19368) );
  OR2_X1 U13503 ( .A1(n12878), .A2(n13000), .ZN(n12914) );
  OR2_X1 U13504 ( .A1(n12878), .A2(n12877), .ZN(n19408) );
  INV_X1 U13505 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19109) );
  INV_X1 U13506 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16269) );
  INV_X1 U13507 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16299) );
  INV_X1 U13508 ( .A(n19420), .ZN(n16284) );
  INV_X1 U13509 ( .A(n16393), .ZN(n16404) );
  NAND2_X1 U13510 ( .A1(n12967), .A2(n12935), .ZN(n16365) );
  INV_X1 U13511 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20062) );
  AOI21_X1 U13512 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19034), .A(n12983), 
        .ZN(n15527) );
  NAND2_X1 U13513 ( .A1(n19477), .A2(n19623), .ZN(n19486) );
  NAND2_X1 U13514 ( .A1(n19477), .A2(n19654), .ZN(n19536) );
  INV_X1 U13515 ( .A(n19562), .ZN(n19573) );
  INV_X1 U13516 ( .A(n19618), .ZN(n19611) );
  INV_X1 U13517 ( .A(n19649), .ZN(n19646) );
  NAND2_X1 U13518 ( .A1(n19655), .A2(n19654), .ZN(n19715) );
  OR2_X1 U13519 ( .A1(n19790), .A2(n19483), .ZN(n19724) );
  NOR2_X1 U13520 ( .A1(n13516), .A2(n19826), .ZN(n19755) );
  INV_X1 U13521 ( .A(n19900), .ZN(n19801) );
  INV_X1 U13522 ( .A(n19910), .ZN(n19806) );
  INV_X1 U13523 ( .A(n19832), .ZN(n19871) );
  NAND2_X1 U13524 ( .A1(n19820), .A2(n19830), .ZN(n19886) );
  INV_X1 U13525 ( .A(n19838), .ZN(n19908) );
  INV_X1 U13526 ( .A(n19931), .ZN(n19946) );
  INV_X1 U13527 ( .A(n16468), .ZN(n19949) );
  INV_X1 U13528 ( .A(n20052), .ZN(n19957) );
  NAND2_X1 U13529 ( .A1(n19959), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20100) );
  INV_X1 U13530 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19011) );
  INV_X1 U13531 ( .A(n17052), .ZN(n17026) );
  NOR2_X1 U13532 ( .A1(n16750), .A2(n17110), .ZN(n17114) );
  NOR2_X1 U13533 ( .A1(n16910), .A2(n17318), .ZN(n17306) );
  INV_X1 U13534 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17381) );
  NOR4_X2 U13535 ( .A1(n19012), .A2(n16997), .A3(n15854), .A4(n18847), .ZN(
        n17399) );
  NAND2_X1 U13536 ( .A1(n17530), .A2(n18397), .ZN(n17455) );
  NOR3_X1 U13537 ( .A1(n17625), .A2(n17545), .A3(n17544), .ZN(n17540) );
  NAND2_X1 U13538 ( .A1(n17569), .A2(n18372), .ZN(n17568) );
  INV_X1 U13539 ( .A(n17569), .ZN(n17587) );
  INV_X1 U13540 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18213) );
  INV_X1 U13541 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18248) );
  INV_X1 U13542 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18024) );
  INV_X1 U13543 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18198) );
  INV_X1 U13544 ( .A(n18253), .ZN(n18270) );
  INV_X1 U13545 ( .A(n18356), .ZN(n18349) );
  INV_X1 U13546 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18839) );
  INV_X1 U13547 ( .A(n18986), .ZN(n18989) );
  INV_X1 U13548 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18412) );
  INV_X1 U13549 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18689) );
  NAND2_X1 U13550 ( .A1(n18401), .A2(n18372), .ZN(n18749) );
  NAND2_X1 U13551 ( .A1(n18401), .A2(n18381), .ZN(n18761) );
  NAND2_X1 U13552 ( .A1(n18401), .A2(n18397), .ZN(n18785) );
  INV_X1 U13553 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18960) );
  INV_X1 U13554 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18880) );
  NAND2_X1 U13555 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18880), .ZN(n19020) );
  NOR2_X1 U13556 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12646), .ZN(n16631)
         );
  INV_X1 U13557 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19326) );
  INV_X1 U13558 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19983) );
  OAI21_X1 U13559 ( .B1(n14062), .B2(n14318), .A(n12634), .ZN(P1_U2842) );
  NAND2_X1 U13560 ( .A1(n11683), .A2(n11682), .ZN(P1_U2873) );
  OR4_X1 U13561 ( .A1(n12798), .A2(n12797), .A3(n12796), .A4(n12795), .ZN(
        P2_U2833) );
  AND2_X2 U13562 ( .A1(n13303), .A2(n14655), .ZN(n10734) );
  INV_X1 U13563 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13564 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10525) );
  INV_X1 U13565 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10521) );
  AND2_X2 U13566 ( .A1(n10521), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10526) );
  AND2_X4 U13567 ( .A1(n10526), .A2(n10528), .ZN(n11231) );
  AOI22_X1 U13568 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11199), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13569 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11626), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10523) );
  BUF_X4 U13570 ( .A(n11633), .Z(n10728) );
  AND2_X2 U13571 ( .A1(n14655), .A2(n10528), .ZN(n10688) );
  AOI22_X1 U13572 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10522) );
  NAND4_X1 U13573 ( .A1(n10525), .A2(n10524), .A3(n10523), .A4(n10522), .ZN(
        n10535) );
  AOI22_X1 U13574 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10533) );
  AND2_X2 U13575 ( .A1(n10526), .A2(n10529), .ZN(n10687) );
  AOI22_X1 U13576 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11632), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10532) );
  AND2_X2 U13577 ( .A1(n10527), .A2(n10528), .ZN(n10800) );
  AOI22_X1 U13578 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10531) );
  AND2_X2 U13579 ( .A1(n14655), .A2(n10529), .ZN(n10611) );
  AOI22_X1 U13580 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13581 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  NOR2_X1 U13582 ( .A1(n10535), .A2(n10534), .ZN(n11292) );
  AOI22_X1 U13583 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13584 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13585 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13586 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10536) );
  NAND4_X1 U13587 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10545) );
  AOI22_X1 U13588 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13589 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13590 ( .A1(n9805), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13591 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13592 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  NOR2_X1 U13593 ( .A1(n10545), .A2(n10544), .ZN(n11276) );
  AOI22_X1 U13594 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13595 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13596 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13597 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13598 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10555) );
  AOI22_X1 U13599 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13600 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13601 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13602 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10550) );
  NAND4_X1 U13603 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10554) );
  NOR2_X1 U13604 ( .A1(n10555), .A2(n10554), .ZN(n11255) );
  AOI22_X1 U13605 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11626), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13606 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13607 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13608 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10556) );
  NAND4_X1 U13609 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10565) );
  AOI22_X1 U13610 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13611 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13612 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13613 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10560) );
  NAND4_X1 U13614 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10564) );
  NOR2_X1 U13615 ( .A1(n10565), .A2(n10564), .ZN(n11254) );
  NOR2_X1 U13616 ( .A1(n11255), .A2(n11254), .ZN(n11267) );
  AOI22_X1 U13617 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13618 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13619 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10567) );
  INV_X1 U13620 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20362) );
  AOI22_X1 U13621 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13622 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10575) );
  AOI22_X1 U13623 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13624 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13625 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13626 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10570) );
  NAND4_X1 U13627 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10574) );
  OR2_X1 U13628 ( .A1(n10575), .A2(n10574), .ZN(n11265) );
  NAND2_X1 U13629 ( .A1(n11267), .A2(n11265), .ZN(n11277) );
  NOR2_X1 U13630 ( .A1(n11276), .A2(n11277), .ZN(n11288) );
  AOI22_X1 U13631 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13632 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13633 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13634 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10577) );
  NAND4_X1 U13635 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10586) );
  AOI22_X1 U13636 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13637 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13638 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13639 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10581) );
  NAND4_X1 U13640 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n10585) );
  NAND2_X1 U13641 ( .A1(n11288), .A2(n11287), .ZN(n11293) );
  NOR2_X1 U13642 ( .A1(n11292), .A2(n11293), .ZN(n11306) );
  AOI22_X1 U13643 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13644 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13645 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10588) );
  INV_X1 U13646 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20371) );
  AOI22_X1 U13647 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10587) );
  NAND4_X1 U13648 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10596) );
  AOI22_X1 U13649 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13650 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13651 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13652 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10591) );
  NAND4_X1 U13653 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10595) );
  OR2_X1 U13654 ( .A1(n10596), .A2(n10595), .ZN(n11305) );
  NAND2_X1 U13655 ( .A1(n11306), .A2(n11305), .ZN(n11641) );
  AOI22_X1 U13656 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13657 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11626), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13658 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13659 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10597) );
  NAND4_X1 U13660 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .ZN(
        n10606) );
  AOI22_X1 U13661 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13662 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13663 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13664 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10601) );
  NAND4_X1 U13665 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .ZN(
        n10605) );
  NOR2_X1 U13666 ( .A1(n10606), .A2(n10605), .ZN(n11642) );
  XOR2_X1 U13667 ( .A(n11641), .B(n11642), .Z(n10662) );
  AOI22_X1 U13668 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10697), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13669 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9807), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13670 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13671 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13672 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13673 ( .A1(n10687), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9802), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13674 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13675 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13676 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13677 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9800), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13678 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9801), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13679 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13681 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10623), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13682 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13683 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10626) );
  INV_X1 U13684 ( .A(n10669), .ZN(n10743) );
  AOI22_X1 U13685 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13686 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13687 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10672), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13688 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10628) );
  NAND4_X1 U13689 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10637) );
  AOI22_X1 U13690 ( .A1(n11198), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10697), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13691 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13692 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13693 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10632) );
  NAND4_X1 U13694 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n10636) );
  OR2_X2 U13695 ( .A1(n10637), .A2(n10636), .ZN(n10695) );
  NAND2_X1 U13696 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13697 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10640) );
  NAND2_X1 U13698 ( .A1(n10697), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10639) );
  NAND2_X1 U13699 ( .A1(n10723), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U13700 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10645) );
  NAND2_X1 U13701 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10644) );
  NAND2_X1 U13702 ( .A1(n10687), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10643) );
  NAND2_X1 U13703 ( .A1(n10672), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10642) );
  NAND2_X1 U13704 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10650) );
  NAND2_X1 U13705 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13706 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10648) );
  NAND2_X1 U13707 ( .A1(n10688), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10647) );
  NAND2_X1 U13708 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10655) );
  NAND2_X1 U13709 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13710 ( .A1(n10611), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10653) );
  NAND2_X1 U13711 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10652) );
  NAND2_X1 U13712 ( .A1(n10695), .A2(n13594), .ZN(n10696) );
  INV_X1 U13713 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n10660) );
  INV_X1 U13714 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14116) );
  OAI22_X1 U13715 ( .A1(n11295), .A2(n10660), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14116), .ZN(n10661) );
  AOI21_X1 U13716 ( .B1(n10662), .B2(n11297), .A(n10661), .ZN(n10667) );
  NAND2_X1 U13717 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10913) );
  INV_X1 U13718 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10663) );
  INV_X1 U13719 ( .A(n11282), .ZN(n10665) );
  INV_X1 U13720 ( .A(n11299), .ZN(n10666) );
  XNOR2_X1 U13721 ( .A(n11648), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14386) );
  INV_X1 U13722 ( .A(n11045), .ZN(n10916) );
  MUX2_X1 U13723 ( .A(n10667), .B(n14386), .S(n10916), .Z(n11310) );
  NAND2_X1 U13724 ( .A1(n10669), .A2(n10756), .ZN(n10671) );
  NAND2_X1 U13725 ( .A1(n9845), .A2(n10694), .ZN(n10670) );
  INV_X1 U13726 ( .A(n10754), .ZN(n10693) );
  AOI22_X1 U13727 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13728 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13729 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10672), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13730 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10673) );
  NAND4_X1 U13731 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n10682) );
  AOI22_X1 U13732 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10697), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13733 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13734 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13735 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10677) );
  NAND4_X1 U13736 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  AOI22_X1 U13737 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13738 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13739 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10697), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13740 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13741 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13742 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13743 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10672), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13744 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10689) );
  INV_X1 U13745 ( .A(n11363), .ZN(n11468) );
  NAND2_X1 U13746 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10702) );
  NAND2_X1 U13747 ( .A1(n11198), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10701) );
  NAND2_X1 U13748 ( .A1(n10697), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10700) );
  NAND2_X1 U13749 ( .A1(n10698), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10699) );
  NAND2_X1 U13750 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10706) );
  NAND2_X1 U13751 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10705) );
  NAND2_X1 U13752 ( .A1(n10687), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U13753 ( .A1(n10672), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10703) );
  NAND2_X1 U13754 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13755 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10709) );
  NAND2_X1 U13756 ( .A1(n9805), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10708) );
  NAND2_X1 U13757 ( .A1(n10688), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13758 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10714) );
  NAND2_X1 U13759 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10713) );
  NAND2_X1 U13760 ( .A1(n10611), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U13761 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13762 ( .A1(n11559), .A2(n13599), .ZN(n10752) );
  INV_X1 U13763 ( .A(n10752), .ZN(n11580) );
  NAND2_X1 U13764 ( .A1(n10687), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13765 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13766 ( .A1(n10672), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U13767 ( .A1(n10688), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U13768 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10727) );
  NAND2_X1 U13769 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10726) );
  NAND2_X1 U13770 ( .A1(n10697), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10725) );
  NAND2_X1 U13771 ( .A1(n10723), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U13772 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13773 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13774 ( .A1(n10646), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13775 ( .A1(n10842), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10729) );
  NAND2_X1 U13776 ( .A1(n10733), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10738) );
  NAND2_X1 U13777 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13778 ( .A1(n10611), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10736) );
  NAND2_X1 U13779 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13780 ( .A1(n10743), .A2(n13589), .ZN(n10778) );
  NAND2_X1 U13781 ( .A1(n10778), .A2(n10744), .ZN(n10749) );
  INV_X1 U13782 ( .A(n11572), .ZN(n11586) );
  AND2_X1 U13783 ( .A1(n14043), .A2(n10694), .ZN(n10745) );
  INV_X1 U13784 ( .A(n11678), .ZN(n10867) );
  NAND2_X1 U13785 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20925) );
  OAI21_X1 U13786 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20925), .ZN(n11558) );
  OR2_X1 U13787 ( .A1(n10754), .A2(n13594), .ZN(n11567) );
  NAND2_X1 U13788 ( .A1(n11567), .A2(n15797), .ZN(n10759) );
  NAND2_X1 U13789 ( .A1(n11572), .A2(n11453), .ZN(n11594) );
  NAND2_X1 U13790 ( .A1(n13579), .A2(n13599), .ZN(n10755) );
  NAND2_X1 U13791 ( .A1(n11594), .A2(n10755), .ZN(n13138) );
  NAND2_X1 U13792 ( .A1(n20355), .A2(n13599), .ZN(n13146) );
  NOR2_X1 U13793 ( .A1(n13146), .A2(n10756), .ZN(n10757) );
  INV_X1 U13794 ( .A(n13589), .ZN(n10758) );
  NAND2_X2 U13795 ( .A1(n11374), .A2(n10777), .ZN(n13165) );
  NAND2_X1 U13796 ( .A1(n13165), .A2(n11363), .ZN(n11588) );
  NAND3_X1 U13797 ( .A1(n10759), .A2(n10781), .A3(n11588), .ZN(n10760) );
  INV_X1 U13798 ( .A(n11365), .ZN(n10761) );
  NAND2_X1 U13799 ( .A1(n10761), .A2(n20355), .ZN(n10763) );
  INV_X1 U13800 ( .A(n10896), .ZN(n21016) );
  OAI21_X1 U13801 ( .B1(n9886), .B2(n10763), .A(n21016), .ZN(n10764) );
  NAND2_X1 U13802 ( .A1(n10765), .A2(n10764), .ZN(n10792) );
  NAND2_X1 U13803 ( .A1(n10792), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10768) );
  NAND2_X1 U13804 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10790) );
  OAI21_X1 U13805 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10790), .ZN(n20654) );
  NAND2_X1 U13806 ( .A1(n20917), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10785) );
  OAI21_X1 U13807 ( .B1(n12637), .B2(n20654), .A(n10785), .ZN(n10766) );
  INV_X1 U13808 ( .A(n10766), .ZN(n10767) );
  XNOR2_X2 U13809 ( .A(n10770), .B(n10784), .ZN(n20445) );
  NAND2_X1 U13810 ( .A1(n10792), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10773) );
  INV_X1 U13811 ( .A(n12637), .ZN(n10892) );
  MUX2_X1 U13812 ( .A(n20917), .B(n10892), .S(n20766), .Z(n10771) );
  NAND2_X1 U13813 ( .A1(n10773), .A2(n10772), .ZN(n10811) );
  NAND2_X1 U13814 ( .A1(n9886), .A2(n12888), .ZN(n11592) );
  NAND3_X1 U13815 ( .A1(n11567), .A2(n13496), .A3(n15797), .ZN(n10783) );
  INV_X1 U13816 ( .A(n10774), .ZN(n10776) );
  NAND2_X1 U13817 ( .A1(n10762), .A2(n13496), .ZN(n13145) );
  INV_X1 U13818 ( .A(n20995), .ZN(n16093) );
  NAND3_X1 U13819 ( .A1(n13145), .A2(n16093), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10775) );
  AOI21_X1 U13820 ( .B1(n21010), .B2(n10776), .A(n10775), .ZN(n10780) );
  OR2_X1 U13821 ( .A1(n11589), .A2(n10694), .ZN(n11596) );
  INV_X1 U13822 ( .A(n12888), .ZN(n13493) );
  AND2_X1 U13823 ( .A1(n13493), .A2(n12629), .ZN(n12917) );
  NAND2_X1 U13824 ( .A1(n12917), .A2(n10778), .ZN(n10779) );
  NAND4_X1 U13825 ( .A1(n11592), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10809) );
  NAND2_X2 U13826 ( .A1(n20445), .A2(n10852), .ZN(n10855) );
  INV_X1 U13827 ( .A(n10784), .ZN(n10787) );
  NAND2_X1 U13828 ( .A1(n10785), .A2(n10521), .ZN(n10786) );
  NAND2_X1 U13829 ( .A1(n10787), .A2(n10786), .ZN(n10788) );
  INV_X1 U13830 ( .A(n10790), .ZN(n10789) );
  NAND2_X1 U13831 ( .A1(n10789), .A2(n11313), .ZN(n20687) );
  NAND2_X1 U13832 ( .A1(n10790), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10791) );
  AND2_X1 U13833 ( .A1(n20687), .A2(n10791), .ZN(n13581) );
  NAND2_X1 U13834 ( .A1(n20917), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10793) );
  AOI22_X1 U13835 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13836 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U13837 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13838 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10796) );
  NAND4_X1 U13839 ( .A1(n10799), .A2(n10798), .A3(n10797), .A4(n10796), .ZN(
        n10806) );
  AOI22_X1 U13840 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13841 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13842 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13843 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10801) );
  NAND4_X1 U13844 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10805) );
  INV_X1 U13845 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13587) );
  OAI22_X1 U13846 ( .A1(n10896), .A2(n11477), .B1(n11349), .B2(n13587), .ZN(
        n10807) );
  XNOR2_X1 U13847 ( .A(n10808), .B(n10807), .ZN(n10865) );
  INV_X1 U13848 ( .A(n10865), .ZN(n10863) );
  INV_X1 U13849 ( .A(n10809), .ZN(n10810) );
  AOI22_X1 U13850 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13851 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10623), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13852 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13853 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13854 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10821) );
  AOI22_X1 U13855 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10842), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13856 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13857 ( .A1(n13308), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13858 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10816) );
  NAND4_X1 U13859 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10820) );
  INV_X1 U13860 ( .A(n11524), .ZN(n11528) );
  AOI22_X1 U13861 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13862 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13863 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13864 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13865 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10831) );
  AOI22_X1 U13866 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13867 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13868 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13869 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13870 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  XNOR2_X1 U13871 ( .A(n11528), .B(n11466), .ZN(n10832) );
  NAND2_X1 U13872 ( .A1(n10832), .A2(n11525), .ZN(n10833) );
  INV_X1 U13873 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13603) );
  AOI21_X1 U13874 ( .B1(n10756), .B2(n11524), .A(n21012), .ZN(n10835) );
  NAND2_X1 U13875 ( .A1(n10762), .A2(n11466), .ZN(n10834) );
  OAI211_X1 U13876 ( .C1(n11349), .C2(n13603), .A(n10835), .B(n10834), .ZN(
        n10880) );
  NAND2_X1 U13877 ( .A1(n11525), .A2(n11524), .ZN(n10836) );
  AOI22_X1 U13878 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10697), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13879 ( .A1(n9805), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13880 ( .A1(n10623), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13881 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10838) );
  NAND4_X1 U13882 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10848) );
  AOI22_X1 U13883 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13884 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13885 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13886 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U13887 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10847) );
  INV_X1 U13888 ( .A(n11467), .ZN(n10849) );
  OR2_X1 U13889 ( .A1(n10896), .A2(n10849), .ZN(n10851) );
  NAND2_X1 U13890 ( .A1(n11357), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10850) );
  OAI211_X1 U13891 ( .C1(n11524), .C2(n10895), .A(n10851), .B(n10850), .ZN(
        n10860) );
  INV_X1 U13892 ( .A(n20445), .ZN(n10854) );
  INV_X1 U13893 ( .A(n10852), .ZN(n10853) );
  INV_X1 U13894 ( .A(n13506), .ZN(n10856) );
  NAND2_X1 U13895 ( .A1(n11525), .A2(n11467), .ZN(n10857) );
  NAND2_X2 U13896 ( .A1(n10858), .A2(n10857), .ZN(n11465) );
  NAND2_X1 U13897 ( .A1(n10865), .A2(n10864), .ZN(n10866) );
  NAND2_X1 U13898 ( .A1(n10910), .A2(n10866), .ZN(n11476) );
  NAND2_X1 U13899 ( .A1(n10867), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10937) );
  XNOR2_X1 U13900 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14071) );
  AOI21_X1 U13901 ( .B1(n10916), .B2(n14071), .A(n11651), .ZN(n10870) );
  NAND2_X1 U13902 ( .A1(n10868), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10869) );
  OAI211_X1 U13903 ( .C1(n10937), .C2(n13320), .A(n10870), .B(n10869), .ZN(
        n10871) );
  INV_X1 U13904 ( .A(n10871), .ZN(n10872) );
  NAND2_X1 U13905 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10890) );
  XNOR2_X2 U13906 ( .A(n11465), .B(n10873), .ZN(n13332) );
  NAND2_X1 U13907 ( .A1(n13332), .A2(n11117), .ZN(n10878) );
  AOI22_X1 U13908 ( .A1(n10868), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20625), .ZN(n10876) );
  INV_X1 U13909 ( .A(n10937), .ZN(n10874) );
  NAND2_X1 U13910 ( .A1(n10874), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10875) );
  AND2_X1 U13911 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  NAND2_X1 U13912 ( .A1(n13339), .A2(n10881), .ZN(n10882) );
  NAND2_X1 U13913 ( .A1(n10882), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13078) );
  NAND2_X1 U13914 ( .A1(n20625), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U13915 ( .A1(n10868), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10884) );
  OAI211_X1 U13916 ( .C1(n10937), .C2(n10520), .A(n10885), .B(n10884), .ZN(
        n10886) );
  AOI21_X1 U13917 ( .B1(n10883), .B2(n11117), .A(n10886), .ZN(n10887) );
  INV_X1 U13918 ( .A(n10887), .ZN(n13080) );
  OR2_X1 U13919 ( .A1(n13080), .A2(n11045), .ZN(n10889) );
  NAND2_X1 U13920 ( .A1(n13079), .A2(n10889), .ZN(n13086) );
  INV_X1 U13921 ( .A(n10910), .ZN(n10909) );
  NOR3_X1 U13922 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11313), .A3(
        n20723), .ZN(n20567) );
  NAND2_X1 U13923 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20567), .ZN(
        n20579) );
  NAND2_X1 U13924 ( .A1(n20653), .A2(n20579), .ZN(n10891) );
  NAND3_X1 U13925 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20855) );
  INV_X1 U13926 ( .A(n20855), .ZN(n20847) );
  NAND2_X1 U13927 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20847), .ZN(
        n20886) );
  AOI22_X1 U13928 ( .A1(n10892), .A2(n13573), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20917), .ZN(n10893) );
  AOI22_X1 U13929 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13930 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13931 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13932 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U13933 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10906) );
  AOI22_X1 U13934 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13935 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10611), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13936 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13937 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10901) );
  NAND4_X1 U13938 ( .A1(n10904), .A2(n10903), .A3(n10902), .A4(n10901), .ZN(
        n10905) );
  AOI22_X1 U13939 ( .A1(n11345), .A2(n11490), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11357), .ZN(n10907) );
  INV_X1 U13940 ( .A(n14650), .ZN(n13569) );
  NAND2_X1 U13941 ( .A1(n10910), .A2(n13569), .ZN(n10911) );
  INV_X1 U13942 ( .A(n13568), .ZN(n10912) );
  INV_X1 U13943 ( .A(n10913), .ZN(n10915) );
  INV_X1 U13944 ( .A(n10934), .ZN(n10914) );
  OAI21_X1 U13945 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10915), .A(
        n10914), .ZN(n20189) );
  AOI22_X1 U13946 ( .A1(n10916), .A2(n20189), .B1(n11651), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U13947 ( .A1(n11258), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10917) );
  OAI211_X1 U13948 ( .C1(n10937), .C2(n10519), .A(n10918), .B(n10917), .ZN(
        n10919) );
  INV_X1 U13949 ( .A(n10919), .ZN(n10920) );
  AOI22_X1 U13950 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9805), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13951 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10728), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13952 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11626), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13953 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11632), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U13954 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10931) );
  AOI22_X1 U13955 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13956 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11229), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13957 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13958 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13959 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  NAND2_X1 U13960 ( .A1(n11345), .A2(n11507), .ZN(n10933) );
  NAND2_X1 U13961 ( .A1(n11357), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10932) );
  NAND2_X1 U13962 ( .A1(n10933), .A2(n10932), .ZN(n10941) );
  NAND2_X1 U13963 ( .A1(n11489), .A2(n11117), .ZN(n10940) );
  XNOR2_X1 U13964 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n10934), .ZN(
        n20301) );
  OAI21_X1 U13965 ( .B1(n21346), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20625), .ZN(n10936) );
  NAND2_X1 U13966 ( .A1(n11258), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10935) );
  OAI211_X1 U13967 ( .C1(n10937), .C2(n16096), .A(n10936), .B(n10935), .ZN(
        n10938) );
  OAI21_X1 U13968 ( .B1(n11045), .B2(n20301), .A(n10938), .ZN(n10939) );
  NOR2_X2 U13969 ( .A1(n13168), .A2(n13345), .ZN(n13354) );
  INV_X1 U13970 ( .A(n10941), .ZN(n10942) );
  OR2_X2 U13971 ( .A1(n10943), .A2(n10942), .ZN(n10966) );
  AOI22_X1 U13972 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13973 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13974 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13975 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10944) );
  NAND4_X1 U13976 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(
        n10953) );
  AOI22_X1 U13977 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13978 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13979 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13980 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10948) );
  NAND4_X1 U13981 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n10952) );
  NAND2_X1 U13982 ( .A1(n11345), .A2(n11506), .ZN(n10955) );
  NAND2_X1 U13983 ( .A1(n11357), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10954) );
  NAND2_X1 U13984 ( .A1(n10955), .A2(n10954), .ZN(n10967) );
  NAND2_X1 U13985 ( .A1(n11497), .A2(n11117), .ZN(n10965) );
  INV_X1 U13986 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10962) );
  INV_X1 U13987 ( .A(n10979), .ZN(n10960) );
  INV_X1 U13988 ( .A(n10956), .ZN(n10958) );
  INV_X1 U13989 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U13990 ( .A1(n10958), .A2(n10957), .ZN(n10959) );
  NAND2_X1 U13991 ( .A1(n10960), .A2(n10959), .ZN(n20169) );
  AOI22_X1 U13992 ( .A1(n20169), .A2(n10916), .B1(n11651), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13993 ( .A1(n13354), .A2(n13353), .ZN(n13352) );
  INV_X1 U13994 ( .A(n13352), .ZN(n10984) );
  INV_X1 U13995 ( .A(n10966), .ZN(n10968) );
  AOI22_X1 U13996 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13997 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13998 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13999 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U14000 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10978) );
  AOI22_X1 U14001 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U14002 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14003 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14004 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10973) );
  NAND4_X1 U14005 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10977) );
  AOI22_X1 U14006 ( .A1(n11345), .A2(n11517), .B1(n11357), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U14007 ( .A1(n10985), .A2(n10986), .ZN(n11505) );
  INV_X1 U14008 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10981) );
  OAI21_X1 U14009 ( .B1(n10979), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10989), .ZN(n20159) );
  AOI22_X1 U14010 ( .A1(n20159), .A2(n10916), .B1(n11651), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10980) );
  OAI21_X1 U14011 ( .B1(n11295), .B2(n10981), .A(n10980), .ZN(n10982) );
  INV_X1 U14012 ( .A(n13481), .ZN(n10983) );
  NAND2_X1 U14013 ( .A1(n10984), .A2(n10983), .ZN(n13614) );
  INV_X1 U14014 ( .A(n13614), .ZN(n10996) );
  INV_X1 U14015 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U14016 ( .A1(n11345), .A2(n11524), .ZN(n10987) );
  OAI21_X1 U14017 ( .B1(n13609), .B2(n11349), .A(n10987), .ZN(n10988) );
  NAND2_X1 U14018 ( .A1(n11515), .A2(n11117), .ZN(n10995) );
  NAND2_X1 U14019 ( .A1(n10989), .A2(n20142), .ZN(n10991) );
  INV_X1 U14020 ( .A(n11007), .ZN(n10990) );
  NAND2_X1 U14021 ( .A1(n10991), .A2(n10990), .ZN(n20150) );
  AOI22_X1 U14022 ( .A1(n20150), .A2(n10916), .B1(n11651), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10992) );
  OAI21_X1 U14023 ( .B1(n11295), .B2(n20230), .A(n10992), .ZN(n10993) );
  NAND2_X1 U14024 ( .A1(n10995), .A2(n10994), .ZN(n13612) );
  NAND2_X1 U14025 ( .A1(n10996), .A2(n13612), .ZN(n13610) );
  AOI22_X1 U14026 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14027 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14028 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14029 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U14030 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11006) );
  AOI22_X1 U14031 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14032 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14033 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14034 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11001) );
  NAND4_X1 U14035 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11005) );
  OAI21_X1 U14036 ( .B1(n11006), .B2(n11005), .A(n11117), .ZN(n11010) );
  NAND2_X1 U14037 ( .A1(n11258), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11009) );
  XNOR2_X1 U14038 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11007), .ZN(
        n20132) );
  AOI22_X1 U14039 ( .A1(n10916), .A2(n20132), .B1(n11651), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11008) );
  XNOR2_X1 U14040 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11013), .ZN(
        n20126) );
  INV_X1 U14041 ( .A(n20126), .ZN(n11028) );
  AOI22_X1 U14042 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14043 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14044 ( .A1(n11627), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14045 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11014) );
  NAND4_X1 U14046 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11023) );
  AOI22_X1 U14047 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14048 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14049 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14050 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11018) );
  NAND4_X1 U14051 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11022) );
  OAI21_X1 U14052 ( .B1(n11023), .B2(n11022), .A(n11117), .ZN(n11026) );
  NAND2_X1 U14053 ( .A1(n11258), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U14054 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11024) );
  NAND3_X1 U14055 ( .A1(n11026), .A2(n11025), .A3(n11024), .ZN(n11027) );
  AOI21_X1 U14056 ( .B1(n11028), .B2(n10916), .A(n11027), .ZN(n13790) );
  AOI22_X1 U14057 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14058 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9805), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U14059 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14060 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11029) );
  NAND4_X1 U14061 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11038) );
  AOI22_X1 U14062 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14063 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14064 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14065 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11033) );
  NAND4_X1 U14066 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n11037) );
  NOR2_X1 U14067 ( .A1(n11038), .A2(n11037), .ZN(n11043) );
  XNOR2_X1 U14068 ( .A(n11039), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14522) );
  NAND2_X1 U14069 ( .A1(n14522), .A2(n10916), .ZN(n11041) );
  AOI22_X1 U14070 ( .A1(n11258), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11651), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11040) );
  OAI211_X1 U14071 ( .C1(n11043), .C2(n11042), .A(n11041), .B(n11040), .ZN(
        n13803) );
  INV_X1 U14072 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11047) );
  INV_X1 U14073 ( .A(n11651), .ZN(n11157) );
  OAI21_X1 U14074 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11044), .A(
        n11074), .ZN(n15967) );
  NAND2_X1 U14075 ( .A1(n15967), .A2(n10888), .ZN(n11046) );
  OAI21_X1 U14076 ( .B1(n11047), .B2(n11157), .A(n11046), .ZN(n11048) );
  AOI21_X1 U14077 ( .B1(n11258), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11048), .ZN(
        n11049) );
  OR2_X2 U14078 ( .A1(n11050), .A2(n11049), .ZN(n11063) );
  AOI22_X1 U14079 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14080 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14081 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14082 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U14083 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11061) );
  AOI22_X1 U14084 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14085 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14086 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14087 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14088 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11060) );
  OR2_X1 U14089 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  INV_X1 U14090 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14381) );
  AOI22_X1 U14091 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14092 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10728), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14093 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14094 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11624), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11064) );
  NAND4_X1 U14095 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11073) );
  AOI22_X1 U14096 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14097 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11626), .B1(
        n9805), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14098 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14099 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11068) );
  NAND4_X1 U14100 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11072) );
  OAI21_X1 U14101 ( .B1(n11073), .B2(n11072), .A(n11117), .ZN(n11077) );
  XNOR2_X1 U14102 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11074), .ZN(
        n15955) );
  INV_X1 U14103 ( .A(n15955), .ZN(n11075) );
  AOI22_X1 U14104 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n10916), .B2(n11075), .ZN(n11076) );
  OAI211_X1 U14105 ( .C1(n11295), .C2(n14381), .A(n11077), .B(n11076), .ZN(
        n14247) );
  XNOR2_X1 U14106 ( .A(n11078), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14510) );
  AOI22_X1 U14107 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14108 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9805), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14109 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14110 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11079) );
  NAND4_X1 U14111 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11088) );
  AOI22_X1 U14112 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14113 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14114 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14115 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U14116 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11087) );
  OAI21_X1 U14117 ( .B1(n11088), .B2(n11087), .A(n11117), .ZN(n11091) );
  NAND2_X1 U14118 ( .A1(n11258), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11090) );
  NAND2_X1 U14119 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11089) );
  NAND3_X1 U14120 ( .A1(n11091), .A2(n11090), .A3(n11089), .ZN(n11092) );
  AOI21_X1 U14121 ( .B1(n14510), .B2(n10916), .A(n11092), .ZN(n14237) );
  XOR2_X1 U14122 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11093), .Z(
        n15943) );
  AOI22_X1 U14123 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14124 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14125 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14126 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11094) );
  NAND4_X1 U14127 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n11103) );
  AOI22_X1 U14128 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9805), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14129 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14130 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14131 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11098) );
  NAND4_X1 U14132 ( .A1(n11101), .A2(n11100), .A3(n11099), .A4(n11098), .ZN(
        n11102) );
  OAI21_X1 U14133 ( .B1(n11103), .B2(n11102), .A(n11117), .ZN(n11106) );
  NAND2_X1 U14134 ( .A1(n11258), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14135 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11104) );
  AND3_X1 U14136 ( .A1(n11106), .A2(n11105), .A3(n11104), .ZN(n11107) );
  OAI21_X1 U14137 ( .B1(n15943), .B2(n11045), .A(n11107), .ZN(n14307) );
  XNOR2_X1 U14138 ( .A(n11108), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15897) );
  INV_X1 U14139 ( .A(n15897), .ZN(n14502) );
  AOI22_X1 U14140 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14141 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14142 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14143 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11109) );
  NAND4_X1 U14144 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        n11119) );
  AOI22_X1 U14145 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14146 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14147 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14148 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11113) );
  NAND4_X1 U14149 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n11118) );
  OAI21_X1 U14150 ( .B1(n11119), .B2(n11118), .A(n11117), .ZN(n11122) );
  NAND2_X1 U14151 ( .A1(n11258), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14152 ( .A1(n11651), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11120) );
  NAND3_X1 U14153 ( .A1(n11122), .A2(n11121), .A3(n11120), .ZN(n11123) );
  AOI21_X1 U14154 ( .B1(n14502), .B2(n10888), .A(n11123), .ZN(n14302) );
  AOI22_X1 U14155 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14156 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11626), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14157 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14158 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11125) );
  NAND4_X1 U14159 ( .A1(n11128), .A2(n11127), .A3(n11126), .A4(n11125), .ZN(
        n11134) );
  AOI22_X1 U14160 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14161 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14162 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14163 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11129) );
  NAND4_X1 U14164 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n11133) );
  NOR2_X1 U14165 ( .A1(n11134), .A2(n11133), .ZN(n11138) );
  OAI21_X1 U14166 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21346), .A(
        n20625), .ZN(n11135) );
  INV_X1 U14167 ( .A(n11135), .ZN(n11136) );
  AOI21_X1 U14168 ( .B1(n11258), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11136), .ZN(
        n11137) );
  OAI21_X1 U14169 ( .B1(n11646), .B2(n11138), .A(n11137), .ZN(n11141) );
  OAI21_X1 U14170 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11139), .A(
        n11155), .ZN(n15937) );
  OR2_X1 U14171 ( .A1(n11045), .A2(n15937), .ZN(n11140) );
  NAND2_X1 U14172 ( .A1(n11141), .A2(n11140), .ZN(n14300) );
  NAND2_X1 U14173 ( .A1(n11143), .A2(n11142), .ZN(n14288) );
  AOI22_X1 U14174 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14175 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14176 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14177 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11145) );
  NAND4_X1 U14178 ( .A1(n11148), .A2(n11147), .A3(n11146), .A4(n11145), .ZN(
        n11154) );
  AOI22_X1 U14179 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14180 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U14181 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11150) );
  AOI22_X1 U14182 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11149) );
  NAND4_X1 U14183 ( .A1(n11152), .A2(n11151), .A3(n11150), .A4(n11149), .ZN(
        n11153) );
  OAI21_X1 U14184 ( .B1(n11154), .B2(n11153), .A(n11297), .ZN(n11160) );
  XNOR2_X1 U14185 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11155), .ZN(
        n15877) );
  INV_X1 U14186 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11156) );
  OAI22_X1 U14187 ( .A1(n15877), .A2(n11045), .B1(n11157), .B2(n11156), .ZN(
        n11158) );
  AOI21_X1 U14188 ( .B1(n11258), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11158), .ZN(
        n11159) );
  INV_X1 U14189 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11163) );
  INV_X1 U14190 ( .A(n11161), .ZN(n11162) );
  NAND2_X1 U14191 ( .A1(n11163), .A2(n11162), .ZN(n11164) );
  AND2_X1 U14192 ( .A1(n11164), .A2(n11191), .ZN(n15868) );
  INV_X1 U14193 ( .A(n15868), .ZN(n14483) );
  AOI22_X1 U14194 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14195 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14196 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14197 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11165) );
  NAND4_X1 U14198 ( .A1(n11168), .A2(n11167), .A3(n11166), .A4(n11165), .ZN(
        n11174) );
  AOI22_X1 U14199 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14200 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14201 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14202 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11169) );
  NAND4_X1 U14203 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11173) );
  NOR2_X1 U14204 ( .A1(n11174), .A2(n11173), .ZN(n11176) );
  AOI22_X1 U14205 ( .A1(n11258), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20625), .ZN(n11175) );
  OAI21_X1 U14206 ( .B1(n11646), .B2(n11176), .A(n11175), .ZN(n11177) );
  MUX2_X1 U14207 ( .A(n14483), .B(n11177), .S(n11045), .Z(n14281) );
  AOI22_X1 U14208 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14209 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11626), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14210 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14211 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11178) );
  NAND4_X1 U14212 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11187) );
  AOI22_X1 U14213 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11627), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14214 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14215 ( .A1(n13308), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14216 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11182) );
  NAND4_X1 U14217 ( .A1(n11185), .A2(n11184), .A3(n11183), .A4(n11182), .ZN(
        n11186) );
  NOR2_X1 U14218 ( .A1(n11187), .A2(n11186), .ZN(n11190) );
  AOI21_X1 U14219 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14232), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11188) );
  AOI21_X1 U14220 ( .B1(n11258), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11188), .ZN(
        n11189) );
  OAI21_X1 U14221 ( .B1(n11646), .B2(n11190), .A(n11189), .ZN(n11193) );
  XNOR2_X1 U14222 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11191), .ZN(
        n14474) );
  NAND2_X1 U14223 ( .A1(n14474), .A2(n10888), .ZN(n11192) );
  OR2_X1 U14224 ( .A1(n11195), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11197) );
  NAND2_X1 U14225 ( .A1(n11197), .A2(n11196), .ZN(n15932) );
  AOI22_X1 U14226 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14227 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11199), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14228 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10728), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14229 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11200) );
  NAND4_X1 U14230 ( .A1(n11203), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n11209) );
  AOI22_X1 U14231 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11626), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14232 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11231), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14233 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11632), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14234 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U14235 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11208) );
  NOR2_X1 U14236 ( .A1(n11209), .A2(n11208), .ZN(n11211) );
  AOI22_X1 U14237 ( .A1(n11258), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20625), .ZN(n11210) );
  OAI21_X1 U14238 ( .B1(n11646), .B2(n11211), .A(n11210), .ZN(n11212) );
  MUX2_X1 U14239 ( .A(n15932), .B(n11212), .S(n11045), .Z(n11213) );
  XNOR2_X1 U14240 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11214), .ZN(
        n14466) );
  AOI22_X1 U14241 ( .A1(n11229), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14242 ( .A1(n10728), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14243 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14244 ( .A1(n11632), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11215) );
  NAND4_X1 U14245 ( .A1(n11218), .A2(n11217), .A3(n11216), .A4(n11215), .ZN(
        n11225) );
  AOI22_X1 U14246 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14247 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14248 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10698), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14249 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11220) );
  NAND4_X1 U14250 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11224) );
  NOR2_X1 U14251 ( .A1(n11225), .A2(n11224), .ZN(n11227) );
  AOI22_X1 U14252 ( .A1(n11258), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20625), .ZN(n11226) );
  OAI21_X1 U14253 ( .B1(n11646), .B2(n11227), .A(n11226), .ZN(n11228) );
  MUX2_X1 U14254 ( .A(n14466), .B(n11228), .S(n11045), .Z(n14214) );
  AOI22_X1 U14255 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11229), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14256 ( .A1(n11624), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11231), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14257 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14258 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11232), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14259 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11243) );
  AOI22_X1 U14260 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14261 ( .A1(n9849), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11237), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14262 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14263 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11238) );
  NAND4_X1 U14264 ( .A1(n11241), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11242) );
  NOR2_X1 U14265 ( .A1(n11243), .A2(n11242), .ZN(n11247) );
  OAI21_X1 U14266 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21346), .A(
        n20625), .ZN(n11244) );
  INV_X1 U14267 ( .A(n11244), .ZN(n11245) );
  AOI21_X1 U14268 ( .B1(n11258), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11245), .ZN(
        n11246) );
  OAI21_X1 U14269 ( .B1(n11646), .B2(n11247), .A(n11246), .ZN(n11253) );
  INV_X1 U14270 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11250) );
  INV_X1 U14271 ( .A(n11248), .ZN(n11249) );
  NAND2_X1 U14272 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  AND2_X1 U14273 ( .A1(n11261), .A2(n11251), .ZN(n14452) );
  NAND2_X1 U14274 ( .A1(n14452), .A2(n10888), .ZN(n11252) );
  XOR2_X1 U14275 ( .A(n11255), .B(n11254), .Z(n11256) );
  NAND2_X1 U14276 ( .A1(n11256), .A2(n11297), .ZN(n11260) );
  AOI21_X1 U14277 ( .B1(n14191), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11257) );
  AOI21_X1 U14278 ( .B1(n11258), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11257), .ZN(
        n11259) );
  NAND2_X1 U14279 ( .A1(n11260), .A2(n11259), .ZN(n11263) );
  XNOR2_X1 U14280 ( .A(n11261), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14190) );
  NAND2_X1 U14281 ( .A1(n14190), .A2(n10888), .ZN(n11262) );
  INV_X1 U14282 ( .A(n11265), .ZN(n11266) );
  XNOR2_X1 U14283 ( .A(n11267), .B(n11266), .ZN(n11270) );
  INV_X1 U14284 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11268) );
  INV_X1 U14285 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14181) );
  OAI22_X1 U14286 ( .A1(n11295), .A2(n11268), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14181), .ZN(n11269) );
  AOI21_X1 U14287 ( .B1(n11270), .B2(n11297), .A(n11269), .ZN(n11274) );
  INV_X1 U14288 ( .A(n11271), .ZN(n11272) );
  NAND2_X1 U14289 ( .A1(n11272), .A2(n14181), .ZN(n11273) );
  AND2_X1 U14290 ( .A1(n11282), .A2(n11273), .ZN(n14180) );
  MUX2_X1 U14291 ( .A(n11274), .B(n14180), .S(n10916), .Z(n14177) );
  XOR2_X1 U14292 ( .A(n11277), .B(n11276), .Z(n11281) );
  INV_X1 U14293 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n11279) );
  INV_X1 U14294 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11278) );
  OAI22_X1 U14295 ( .A1(n11295), .A2(n11279), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11278), .ZN(n11280) );
  AOI21_X1 U14296 ( .B1(n11281), .B2(n11297), .A(n11280), .ZN(n11283) );
  XNOR2_X1 U14297 ( .A(n11282), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14427) );
  MUX2_X1 U14298 ( .A(n11283), .B(n14427), .S(n10888), .Z(n14165) );
  INV_X1 U14299 ( .A(n11284), .ZN(n11285) );
  INV_X1 U14300 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14157) );
  NAND2_X1 U14301 ( .A1(n11285), .A2(n14157), .ZN(n11286) );
  NAND2_X1 U14302 ( .A1(n11299), .A2(n11286), .ZN(n14418) );
  XNOR2_X1 U14303 ( .A(n11288), .B(n11287), .ZN(n11290) );
  AOI22_X1 U14304 ( .A1(n11258), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20625), .ZN(n11289) );
  OAI21_X1 U14305 ( .B1(n11290), .B2(n11646), .A(n11289), .ZN(n11291) );
  MUX2_X1 U14306 ( .A(n14418), .B(n11291), .S(n11045), .Z(n14153) );
  XOR2_X1 U14307 ( .A(n11293), .B(n11292), .Z(n11298) );
  INV_X1 U14308 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n11294) );
  INV_X1 U14309 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14146) );
  OAI22_X1 U14310 ( .A1(n11295), .A2(n11294), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14146), .ZN(n11296) );
  AOI21_X1 U14311 ( .B1(n11298), .B2(n11297), .A(n11296), .ZN(n11300) );
  XNOR2_X1 U14312 ( .A(n11299), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14145) );
  MUX2_X1 U14313 ( .A(n11300), .B(n14145), .S(n10888), .Z(n11301) );
  INV_X1 U14314 ( .A(n11302), .ZN(n11303) );
  INV_X1 U14315 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14129) );
  NAND2_X1 U14316 ( .A1(n11303), .A2(n14129), .ZN(n11304) );
  NAND2_X1 U14317 ( .A1(n11648), .A2(n11304), .ZN(n14400) );
  XNOR2_X1 U14318 ( .A(n11306), .B(n11305), .ZN(n11308) );
  AOI22_X1 U14319 ( .A1(n11258), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20625), .ZN(n11307) );
  OAI21_X1 U14320 ( .B1(n11308), .B2(n11646), .A(n11307), .ZN(n11309) );
  MUX2_X1 U14321 ( .A(n14400), .B(n11309), .S(n11045), .Z(n14125) );
  INV_X1 U14322 ( .A(n14390), .ZN(n14321) );
  NAND2_X1 U14323 ( .A1(n14043), .A2(n13496), .ZN(n11488) );
  XNOR2_X1 U14324 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14325 ( .A1(n11331), .A2(n11330), .ZN(n11329) );
  NAND2_X1 U14326 ( .A1(n20723), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14327 ( .A1(n11329), .A2(n11311), .ZN(n11340) );
  NAND2_X1 U14328 ( .A1(n11340), .A2(n11312), .ZN(n11315) );
  NAND2_X1 U14329 ( .A1(n11313), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U14330 ( .A1(n11322), .A2(n11321), .ZN(n11317) );
  NAND2_X1 U14331 ( .A1(n20653), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14332 ( .A1(n11317), .A2(n11316), .ZN(n11353) );
  NOR2_X1 U14333 ( .A1(n16096), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U14334 ( .A1(n11352), .A2(n11557), .ZN(n11362) );
  NAND2_X1 U14335 ( .A1(n11557), .A2(n11345), .ZN(n11360) );
  XNOR2_X1 U14336 ( .A(n11322), .B(n11321), .ZN(n11552) );
  AND2_X1 U14337 ( .A1(n10520), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11323) );
  NOR2_X1 U14338 ( .A1(n11331), .A2(n11323), .ZN(n11326) );
  INV_X1 U14339 ( .A(n11326), .ZN(n11324) );
  NOR2_X1 U14340 ( .A1(n11341), .A2(n11324), .ZN(n11328) );
  AND2_X1 U14341 ( .A1(n14043), .A2(n20355), .ZN(n11325) );
  NOR2_X1 U14342 ( .A1(n12888), .A2(n11325), .ZN(n11343) );
  OAI211_X1 U14343 ( .C1(n10762), .C2(n11586), .A(n11343), .B(n11326), .ZN(
        n11327) );
  OAI21_X1 U14344 ( .B1(n11352), .B2(n11328), .A(n11327), .ZN(n11334) );
  INV_X1 U14345 ( .A(n11334), .ZN(n11338) );
  OAI21_X1 U14346 ( .B1(n11331), .B2(n11330), .A(n11329), .ZN(n11553) );
  NOR2_X1 U14347 ( .A1(n21012), .A2(n14043), .ZN(n11332) );
  INV_X1 U14348 ( .A(n11335), .ZN(n11337) );
  INV_X1 U14349 ( .A(n11332), .ZN(n11333) );
  NAND3_X1 U14350 ( .A1(n11341), .A2(n13496), .A3(n11333), .ZN(n11354) );
  AOI22_X1 U14351 ( .A1(n11335), .A2(n11334), .B1(n11553), .B2(n11354), .ZN(
        n11336) );
  AOI21_X1 U14352 ( .B1(n11338), .B2(n11337), .A(n11336), .ZN(n11348) );
  MUX2_X1 U14353 ( .A(n11313), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11339) );
  XNOR2_X1 U14354 ( .A(n11340), .B(n11339), .ZN(n11554) );
  OAI21_X1 U14355 ( .B1(n11341), .B2(n11554), .A(n11343), .ZN(n11342) );
  AOI21_X1 U14356 ( .B1(n11357), .B2(n11554), .A(n11342), .ZN(n11347) );
  INV_X1 U14357 ( .A(n11343), .ZN(n11344) );
  NAND2_X1 U14358 ( .A1(n11345), .A2(n11344), .ZN(n11346) );
  OAI22_X1 U14359 ( .A1(n11348), .A2(n11347), .B1(n11554), .B2(n11346), .ZN(
        n11351) );
  NAND2_X1 U14360 ( .A1(n11349), .A2(n11552), .ZN(n11350) );
  NOR2_X1 U14361 ( .A1(n11357), .A2(n11355), .ZN(n11359) );
  INV_X1 U14362 ( .A(n11354), .ZN(n11356) );
  INV_X1 U14363 ( .A(n11355), .ZN(n11555) );
  NAND3_X1 U14364 ( .A1(n11357), .A2(n11356), .A3(n11555), .ZN(n11358) );
  NAND2_X1 U14365 ( .A1(n15783), .A2(n13148), .ZN(n11366) );
  INV_X1 U14366 ( .A(n10695), .ZN(n11664) );
  NOR2_X1 U14367 ( .A1(n14043), .A2(n13594), .ZN(n11364) );
  NAND4_X1 U14368 ( .A1(n11365), .A2(n11664), .A3(n11364), .A4(n10694), .ZN(
        n11661) );
  INV_X2 U14369 ( .A(n11584), .ZN(n13089) );
  NAND2_X1 U14370 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11369) );
  OR2_X1 U14371 ( .A1(n11584), .A2(n11374), .ZN(n11414) );
  AND2_X1 U14372 ( .A1(n11369), .A2(n11414), .ZN(n11370) );
  NAND2_X1 U14373 ( .A1(n11371), .A2(n11370), .ZN(n11373) );
  NAND2_X1 U14374 ( .A1(n11374), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11372) );
  OAI21_X1 U14375 ( .B1(n11453), .B2(P1_EBX_REG_0__SCAN_IN), .A(n11372), .ZN(
        n13167) );
  XNOR2_X1 U14376 ( .A(n11373), .B(n13167), .ZN(n13088) );
  NAND2_X1 U14377 ( .A1(n13088), .A2(n11584), .ZN(n13091) );
  NAND2_X1 U14378 ( .A1(n13091), .A2(n11373), .ZN(n13223) );
  INV_X1 U14379 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21243) );
  NAND2_X1 U14380 ( .A1(n11444), .A2(n21243), .ZN(n11378) );
  INV_X1 U14381 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20336) );
  NAND2_X1 U14382 ( .A1(n11374), .A2(n20336), .ZN(n11376) );
  NAND2_X1 U14383 ( .A1(n11584), .A2(n21243), .ZN(n11375) );
  NAND3_X1 U14384 ( .A1(n11376), .A2(n12629), .A3(n11375), .ZN(n11377) );
  AND2_X1 U14385 ( .A1(n11378), .A2(n11377), .ZN(n13222) );
  NOR2_X1 U14386 ( .A1(n13223), .A2(n13222), .ZN(n13224) );
  INV_X1 U14387 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20202) );
  NAND2_X1 U14388 ( .A1(n11437), .A2(n20202), .ZN(n11381) );
  INV_X1 U14389 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20320) );
  NAND2_X1 U14390 ( .A1(n11584), .A2(n20202), .ZN(n11379) );
  OAI211_X1 U14391 ( .C1(n11453), .C2(n20320), .A(n11379), .B(n11374), .ZN(
        n11380) );
  AND2_X1 U14392 ( .A1(n11381), .A2(n11380), .ZN(n13171) );
  NAND2_X1 U14393 ( .A1(n13224), .A2(n13171), .ZN(n13360) );
  MUX2_X1 U14394 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11384) );
  NAND2_X1 U14395 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11382) );
  AND2_X1 U14396 ( .A1(n11382), .A2(n11414), .ZN(n11383) );
  AND2_X1 U14397 ( .A1(n11384), .A2(n11383), .ZN(n13359) );
  INV_X1 U14398 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13559) );
  INV_X1 U14399 ( .A(n13165), .ZN(n11418) );
  NAND2_X1 U14400 ( .A1(n13559), .A2(n11418), .ZN(n11386) );
  MUX2_X1 U14401 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11385) );
  NAND2_X1 U14402 ( .A1(n11386), .A2(n11385), .ZN(n16083) );
  NOR2_X1 U14403 ( .A1(n16084), .A2(n16083), .ZN(n16086) );
  INV_X1 U14404 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14405 ( .A1(n11374), .A2(n11585), .ZN(n11388) );
  INV_X1 U14406 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21334) );
  NAND2_X1 U14407 ( .A1(n11584), .A2(n21334), .ZN(n11387) );
  NAND3_X1 U14408 ( .A1(n11388), .A2(n12629), .A3(n11387), .ZN(n11389) );
  OAI21_X1 U14409 ( .B1(n11449), .B2(P1_EBX_REG_6__SCAN_IN), .A(n11389), .ZN(
        n13482) );
  NAND2_X1 U14410 ( .A1(n16086), .A2(n13482), .ZN(n13617) );
  MUX2_X1 U14411 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n11390) );
  OAI21_X1 U14412 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13165), .A(
        n11390), .ZN(n13616) );
  INV_X1 U14413 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21250) );
  NAND2_X1 U14414 ( .A1(n11444), .A2(n21250), .ZN(n11394) );
  INV_X1 U14415 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13751) );
  NAND2_X1 U14416 ( .A1(n11374), .A2(n13751), .ZN(n11392) );
  NAND2_X1 U14417 ( .A1(n11584), .A2(n21250), .ZN(n11391) );
  NAND3_X1 U14418 ( .A1(n11392), .A2(n12629), .A3(n11391), .ZN(n11393) );
  AND2_X1 U14419 ( .A1(n11394), .A2(n11393), .ZN(n13734) );
  OR2_X2 U14420 ( .A1(n13735), .A2(n13734), .ZN(n16066) );
  INV_X1 U14421 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16075) );
  NAND2_X1 U14422 ( .A1(n16075), .A2(n11418), .ZN(n11396) );
  MUX2_X1 U14423 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11395) );
  NAND2_X1 U14424 ( .A1(n11396), .A2(n11395), .ZN(n16067) );
  INV_X1 U14425 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16064) );
  NAND2_X1 U14426 ( .A1(n11374), .A2(n16064), .ZN(n11398) );
  INV_X1 U14427 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21347) );
  NAND2_X1 U14428 ( .A1(n11584), .A2(n21347), .ZN(n11397) );
  NAND3_X1 U14429 ( .A1(n11398), .A2(n12629), .A3(n11397), .ZN(n11399) );
  OAI21_X1 U14430 ( .B1(n11449), .B2(P1_EBX_REG_10__SCAN_IN), .A(n11399), .ZN(
        n13804) );
  MUX2_X1 U14431 ( .A(n11437), .B(n11453), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11401) );
  NOR2_X1 U14432 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11400) );
  NOR2_X1 U14433 ( .A1(n11401), .A2(n11400), .ZN(n15915) );
  MUX2_X1 U14434 ( .A(n11437), .B(n11453), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11403) );
  NOR2_X1 U14435 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11402) );
  NOR2_X1 U14436 ( .A1(n11403), .A2(n11402), .ZN(n14239) );
  MUX2_X1 U14437 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11406) );
  NAND2_X1 U14438 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11404) );
  AND2_X1 U14439 ( .A1(n11404), .A2(n11414), .ZN(n11405) );
  NAND2_X1 U14440 ( .A1(n11406), .A2(n11405), .ZN(n14248) );
  NAND2_X1 U14441 ( .A1(n14239), .A2(n14248), .ZN(n11407) );
  INV_X1 U14442 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15908) );
  NAND2_X1 U14443 ( .A1(n11444), .A2(n15908), .ZN(n11411) );
  INV_X1 U14444 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16025) );
  NAND2_X1 U14445 ( .A1(n11374), .A2(n16025), .ZN(n11409) );
  NAND2_X1 U14446 ( .A1(n11584), .A2(n15908), .ZN(n11408) );
  NAND3_X1 U14447 ( .A1(n11409), .A2(n12629), .A3(n11408), .ZN(n11410) );
  NOR2_X2 U14448 ( .A1(n14309), .A2(n14308), .ZN(n14310) );
  MUX2_X1 U14449 ( .A(n11437), .B(n11453), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11413) );
  NOR2_X1 U14450 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11412) );
  NOR2_X1 U14451 ( .A1(n11413), .A2(n11412), .ZN(n14305) );
  MUX2_X1 U14452 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11417) );
  INV_X1 U14453 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14643) );
  OAI21_X1 U14454 ( .B1(n11584), .B2(n14643), .A(n11414), .ZN(n11415) );
  INV_X1 U14455 ( .A(n11415), .ZN(n11416) );
  INV_X1 U14456 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14622) );
  NAND2_X1 U14457 ( .A1(n14622), .A2(n11418), .ZN(n11420) );
  MUX2_X1 U14458 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11419) );
  NAND2_X1 U14459 ( .A1(n11420), .A2(n11419), .ZN(n14291) );
  INV_X1 U14460 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16001) );
  NAND2_X1 U14461 ( .A1(n11374), .A2(n16001), .ZN(n11422) );
  INV_X1 U14462 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21379) );
  NAND2_X1 U14463 ( .A1(n11584), .A2(n21379), .ZN(n11421) );
  NAND3_X1 U14464 ( .A1(n11422), .A2(n12629), .A3(n11421), .ZN(n11423) );
  OAI21_X1 U14465 ( .B1(n11449), .B2(P1_EBX_REG_18__SCAN_IN), .A(n11423), .ZN(
        n14283) );
  MUX2_X1 U14466 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11424) );
  OAI21_X1 U14467 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13165), .A(
        n11424), .ZN(n14229) );
  OR2_X2 U14468 ( .A1(n14285), .A2(n14229), .ZN(n14274) );
  INV_X1 U14469 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21353) );
  NAND2_X1 U14470 ( .A1(n11444), .A2(n21353), .ZN(n11428) );
  INV_X1 U14471 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U14472 ( .A1(n11374), .A2(n14461), .ZN(n11426) );
  NAND2_X1 U14473 ( .A1(n11584), .A2(n21353), .ZN(n11425) );
  NAND3_X1 U14474 ( .A1(n11426), .A2(n12629), .A3(n11425), .ZN(n11427) );
  AND2_X1 U14475 ( .A1(n11428), .A2(n11427), .ZN(n14273) );
  OR2_X2 U14476 ( .A1(n14274), .A2(n14273), .ZN(n14276) );
  MUX2_X1 U14477 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11429) );
  OAI21_X1 U14478 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13165), .A(
        n11429), .ZN(n14218) );
  MUX2_X1 U14479 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11431) );
  NAND2_X1 U14480 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11430) );
  NAND2_X1 U14481 ( .A1(n11431), .A2(n11430), .ZN(n14205) );
  INV_X1 U14482 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21229) );
  NAND2_X1 U14483 ( .A1(n11437), .A2(n21229), .ZN(n11434) );
  INV_X1 U14484 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U14485 ( .A1(n11584), .A2(n21229), .ZN(n11432) );
  OAI211_X1 U14486 ( .C1(n11453), .C2(n14596), .A(n11432), .B(n11374), .ZN(
        n11433) );
  MUX2_X1 U14487 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11436) );
  NAND2_X1 U14488 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11435) );
  AND2_X1 U14489 ( .A1(n11436), .A2(n11435), .ZN(n14178) );
  INV_X1 U14490 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21159) );
  NAND2_X1 U14491 ( .A1(n11437), .A2(n21159), .ZN(n11440) );
  INV_X1 U14492 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U14493 ( .A1(n11584), .A2(n21159), .ZN(n11438) );
  OAI211_X1 U14494 ( .C1(n11453), .C2(n14563), .A(n11438), .B(n11374), .ZN(
        n11439) );
  NAND2_X1 U14495 ( .A1(n11440), .A2(n11439), .ZN(n14167) );
  NOR2_X2 U14496 ( .A1(n9882), .A2(n14167), .ZN(n14166) );
  MUX2_X1 U14497 ( .A(n11441), .B(n12629), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11443) );
  OR2_X1 U14498 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U14499 ( .A1(n11443), .A2(n11442), .ZN(n14140) );
  INV_X1 U14500 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U14501 ( .A1(n11444), .A2(n21132), .ZN(n11447) );
  INV_X1 U14502 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14415) );
  NAND2_X1 U14503 ( .A1(n11374), .A2(n14415), .ZN(n11445) );
  OAI211_X1 U14504 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n13089), .A(n11445), .B(
        n12629), .ZN(n11446) );
  AND2_X1 U14505 ( .A1(n11447), .A2(n11446), .ZN(n14139) );
  NOR2_X1 U14506 ( .A1(n14140), .A2(n14139), .ZN(n11448) );
  AND2_X2 U14507 ( .A1(n14166), .A2(n11448), .ZN(n14143) );
  MUX2_X1 U14508 ( .A(n11449), .B(n11374), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11451) );
  NAND2_X1 U14509 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11450) );
  NAND2_X1 U14510 ( .A1(n11451), .A2(n11450), .ZN(n14126) );
  OR2_X1 U14511 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11452) );
  INV_X1 U14512 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n21191) );
  NAND2_X1 U14513 ( .A1(n11584), .A2(n21191), .ZN(n11454) );
  NAND2_X1 U14514 ( .A1(n11452), .A2(n11454), .ZN(n12628) );
  MUX2_X1 U14515 ( .A(n12628), .B(n11454), .S(n11453), .Z(n11455) );
  OR2_X2 U14516 ( .A1(n14128), .A2(n11455), .ZN(n12627) );
  NAND2_X1 U14517 ( .A1(n14128), .A2(n11455), .ZN(n11456) );
  NAND2_X1 U14518 ( .A1(n12627), .A2(n11456), .ZN(n14114) );
  OR2_X1 U14519 ( .A1(n13568), .A2(n11488), .ZN(n11462) );
  NAND2_X1 U14520 ( .A1(n11466), .A2(n11467), .ZN(n11478) );
  NAND2_X1 U14521 ( .A1(n11478), .A2(n11477), .ZN(n11491) );
  INV_X1 U14522 ( .A(n11490), .ZN(n11459) );
  XNOR2_X1 U14523 ( .A(n11491), .B(n11459), .ZN(n11460) );
  NAND2_X1 U14524 ( .A1(n11460), .A2(n21010), .ZN(n11461) );
  NAND2_X1 U14525 ( .A1(n11462), .A2(n11461), .ZN(n11486) );
  XNOR2_X1 U14526 ( .A(n11486), .B(n20320), .ZN(n13271) );
  NAND2_X1 U14527 ( .A1(n10762), .A2(n13589), .ZN(n11479) );
  OAI21_X1 U14528 ( .B1(n13146), .B2(n11466), .A(n11479), .ZN(n11463) );
  INV_X1 U14529 ( .A(n11463), .ZN(n11464) );
  NAND2_X1 U14530 ( .A1(n13094), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13093) );
  OR2_X1 U14531 ( .A1(n11465), .A2(n20355), .ZN(n11472) );
  OAI21_X1 U14532 ( .B1(n11467), .B2(n11466), .A(n11478), .ZN(n11469) );
  OAI211_X1 U14533 ( .C1(n11469), .C2(n13146), .A(n11468), .B(n14043), .ZN(
        n11470) );
  INV_X1 U14534 ( .A(n11470), .ZN(n11471) );
  NAND2_X1 U14535 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  INV_X1 U14536 ( .A(n11473), .ZN(n11474) );
  OR2_X1 U14537 ( .A1(n13093), .A2(n11474), .ZN(n11475) );
  XNOR2_X1 U14538 ( .A(n11478), .B(n11477), .ZN(n11481) );
  INV_X1 U14539 ( .A(n11479), .ZN(n11480) );
  AOI21_X1 U14540 ( .B1(n11481), .B2(n21010), .A(n11480), .ZN(n11482) );
  NAND2_X1 U14541 ( .A1(n11483), .A2(n11482), .ZN(n13247) );
  NAND2_X1 U14542 ( .A1(n11484), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11485) );
  NAND2_X1 U14543 ( .A1(n13246), .A2(n11485), .ZN(n13270) );
  NAND2_X1 U14544 ( .A1(n11486), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11487) );
  NAND2_X1 U14545 ( .A1(n11489), .A2(n10260), .ZN(n11494) );
  NAND2_X1 U14546 ( .A1(n11491), .A2(n11490), .ZN(n11509) );
  XNOR2_X1 U14547 ( .A(n11509), .B(n11507), .ZN(n11492) );
  NAND2_X1 U14548 ( .A1(n11492), .A2(n21010), .ZN(n11493) );
  NAND2_X1 U14549 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  INV_X1 U14550 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20312) );
  XNOR2_X1 U14551 ( .A(n11495), .B(n20312), .ZN(n20293) );
  NAND2_X1 U14552 ( .A1(n11495), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14553 ( .A1(n11497), .A2(n10260), .ZN(n11502) );
  INV_X1 U14554 ( .A(n11507), .ZN(n11498) );
  OR2_X1 U14555 ( .A1(n11509), .A2(n11498), .ZN(n11499) );
  XNOR2_X1 U14556 ( .A(n11499), .B(n11506), .ZN(n11500) );
  NAND2_X1 U14557 ( .A1(n11500), .A2(n21010), .ZN(n11501) );
  NAND2_X1 U14558 ( .A1(n11502), .A2(n11501), .ZN(n11503) );
  XNOR2_X1 U14559 ( .A(n11503), .B(n13559), .ZN(n15978) );
  NAND2_X1 U14560 ( .A1(n15979), .A2(n15978), .ZN(n15977) );
  NAND2_X1 U14561 ( .A1(n11503), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11504) );
  NAND2_X1 U14562 ( .A1(n15977), .A2(n11504), .ZN(n13557) );
  NAND3_X1 U14563 ( .A1(n11527), .A2(n10260), .A3(n11505), .ZN(n11512) );
  NAND2_X1 U14564 ( .A1(n11507), .A2(n11506), .ZN(n11508) );
  OR2_X1 U14565 ( .A1(n11509), .A2(n11508), .ZN(n11516) );
  XNOR2_X1 U14566 ( .A(n11516), .B(n11517), .ZN(n11510) );
  NAND2_X1 U14567 ( .A1(n11510), .A2(n21010), .ZN(n11511) );
  NAND2_X1 U14568 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  XNOR2_X1 U14569 ( .A(n11513), .B(n11585), .ZN(n13556) );
  NAND2_X1 U14570 ( .A1(n11513), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U14571 ( .A1(n11515), .A2(n10260), .ZN(n11521) );
  INV_X1 U14572 ( .A(n11516), .ZN(n11518) );
  NAND2_X1 U14573 ( .A1(n11518), .A2(n11517), .ZN(n11529) );
  XNOR2_X1 U14574 ( .A(n11529), .B(n11524), .ZN(n11519) );
  NAND2_X1 U14575 ( .A1(n11519), .A2(n21010), .ZN(n11520) );
  NAND2_X1 U14576 ( .A1(n11521), .A2(n11520), .ZN(n15968) );
  NAND2_X1 U14577 ( .A1(n15968), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11523) );
  NAND2_X2 U14578 ( .A1(n11527), .A2(n11526), .ZN(n11533) );
  OR3_X1 U14579 ( .A1(n11529), .A2(n11528), .A3(n13146), .ZN(n11530) );
  NAND2_X1 U14580 ( .A1(n11533), .A2(n11530), .ZN(n13746) );
  NAND2_X1 U14581 ( .A1(n15938), .A2(n16075), .ZN(n11532) );
  XNOR2_X1 U14582 ( .A(n11533), .B(n16031), .ZN(n14508) );
  NAND2_X1 U14583 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11534) );
  AND2_X1 U14584 ( .A1(n14515), .A2(n11534), .ZN(n14505) );
  INV_X1 U14585 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16033) );
  AND2_X1 U14586 ( .A1(n14515), .A2(n16025), .ZN(n11535) );
  NOR2_X1 U14587 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14496) );
  INV_X1 U14588 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14636) );
  AND2_X1 U14589 ( .A1(n14496), .A2(n14636), .ZN(n11536) );
  NAND2_X1 U14590 ( .A1(n14497), .A2(n14488), .ZN(n11538) );
  XNOR2_X1 U14591 ( .A(n15938), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14634) );
  NAND2_X1 U14592 ( .A1(n15938), .A2(n14636), .ZN(n14631) );
  AND2_X1 U14593 ( .A1(n14634), .A2(n14631), .ZN(n11537) );
  NAND2_X1 U14594 ( .A1(n15938), .A2(n14622), .ZN(n11539) );
  NOR2_X1 U14595 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11540) );
  OR2_X1 U14596 ( .A1(n14515), .A2(n11540), .ZN(n15947) );
  OR2_X1 U14597 ( .A1(n14515), .A2(n16033), .ZN(n15950) );
  NAND2_X1 U14598 ( .A1(n15947), .A2(n15950), .ZN(n14506) );
  INV_X1 U14599 ( .A(n14488), .ZN(n14632) );
  NOR2_X1 U14600 ( .A1(n14506), .A2(n14632), .ZN(n11541) );
  XNOR2_X1 U14601 ( .A(n15938), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14480) );
  AND2_X1 U14602 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U14603 ( .A1(n14564), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14566) );
  INV_X1 U14604 ( .A(n14566), .ZN(n11543) );
  NOR2_X1 U14605 ( .A1(n11544), .A2(n11531), .ZN(n14406) );
  NAND2_X1 U14606 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14548) );
  INV_X1 U14607 ( .A(n14548), .ZN(n14528) );
  AND2_X1 U14608 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11549) );
  INV_X1 U14609 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11616) );
  AND3_X1 U14610 ( .A1(n14528), .A2(n11549), .A3(n11616), .ZN(n11619) );
  INV_X1 U14611 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11615) );
  NOR2_X1 U14612 ( .A1(n11531), .A2(n11615), .ZN(n11548) );
  INV_X1 U14613 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11545) );
  INV_X1 U14614 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U14615 ( .A1(n14596), .A2(n14436), .ZN(n14422) );
  INV_X1 U14616 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14556) );
  INV_X1 U14617 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U14618 ( .A1(n14556), .A2(n14396), .ZN(n14547) );
  AOI21_X1 U14619 ( .B1(n14384), .B2(n11548), .A(n11547), .ZN(n12636) );
  AOI21_X1 U14620 ( .B1(n14384), .B2(n11549), .A(n11616), .ZN(n11550) );
  NAND2_X1 U14621 ( .A1(n11550), .A2(n14515), .ZN(n11551) );
  NOR4_X1 U14622 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11556) );
  NOR2_X1 U14623 ( .A1(n11557), .A2(n11556), .ZN(n12887) );
  NAND2_X1 U14624 ( .A1(n13496), .A2(n21011), .ZN(n21009) );
  NAND3_X1 U14625 ( .A1(n12887), .A2(n16097), .A3(n21009), .ZN(n11563) );
  NAND2_X1 U14626 ( .A1(n13496), .A2(n16097), .ZN(n13059) );
  NAND2_X1 U14627 ( .A1(n15849), .A2(n16097), .ZN(n13154) );
  NAND2_X1 U14628 ( .A1(n13059), .A2(n13154), .ZN(n13494) );
  NAND2_X1 U14629 ( .A1(n13155), .A2(n13494), .ZN(n11560) );
  NAND3_X1 U14630 ( .A1(n11560), .A2(n13599), .A3(n11678), .ZN(n11561) );
  NAND2_X1 U14631 ( .A1(n11561), .A2(n15789), .ZN(n11562) );
  MUX2_X1 U14632 ( .A(n11563), .B(n11562), .S(n13157), .Z(n11570) );
  NAND2_X1 U14633 ( .A1(n11564), .A2(n10762), .ZN(n15785) );
  AND2_X1 U14634 ( .A1(n10743), .A2(n10762), .ZN(n11565) );
  OAI21_X1 U14635 ( .B1(n10669), .B2(n10762), .A(n13146), .ZN(n11566) );
  NAND2_X1 U14636 ( .A1(n11567), .A2(n11566), .ZN(n11593) );
  NAND2_X1 U14637 ( .A1(n11573), .A2(n11593), .ZN(n11568) );
  NAND2_X1 U14638 ( .A1(n15785), .A2(n11568), .ZN(n13159) );
  NAND3_X1 U14639 ( .A1(n15783), .A2(n10669), .A3(n13496), .ZN(n11569) );
  NAND3_X1 U14640 ( .A1(n11570), .A2(n13159), .A3(n11569), .ZN(n11571) );
  AND2_X1 U14641 ( .A1(n11573), .A2(n11572), .ZN(n15782) );
  NAND2_X1 U14642 ( .A1(n13148), .A2(n12888), .ZN(n15780) );
  OAI21_X1 U14643 ( .B1(n10756), .B2(n11582), .A(n15780), .ZN(n11574) );
  OR3_X1 U14644 ( .A1(n11575), .A2(n15782), .A3(n11574), .ZN(n11576) );
  AOI22_X1 U14645 ( .A1(n13165), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13089), .ZN(n11579) );
  AND2_X1 U14646 ( .A1(n13089), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11577) );
  AOI21_X1 U14647 ( .B1(n13165), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11577), .ZN(
        n12632) );
  MUX2_X1 U14648 ( .A(n12632), .B(n12629), .S(n12627), .Z(n11578) );
  XOR2_X1 U14649 ( .A(n11579), .B(n11578), .Z(n14265) );
  NAND2_X1 U14650 ( .A1(n10153), .A2(n20355), .ZN(n11581) );
  OAI21_X1 U14651 ( .B1(n11582), .B2(n13594), .A(n11581), .ZN(n11583) );
  NAND2_X1 U14652 ( .A1(n14265), .A2(n20316), .ZN(n11621) );
  AND2_X1 U14653 ( .A1(n13148), .A2(n11584), .ZN(n15788) );
  INV_X1 U14654 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16043) );
  NAND2_X1 U14655 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16061) );
  NOR2_X1 U14656 ( .A1(n11585), .A2(n16061), .ZN(n16053) );
  NAND3_X1 U14657 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16053), .ZN(n16051) );
  NOR2_X1 U14658 ( .A1(n16043), .A2(n16051), .ZN(n16039) );
  NAND2_X1 U14659 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16039), .ZN(
        n11598) );
  NOR2_X1 U14660 ( .A1(n20312), .A2(n20320), .ZN(n20307) );
  INV_X1 U14661 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20324) );
  INV_X1 U14662 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20350) );
  OAI21_X1 U14663 ( .B1(n20324), .B2(n20350), .A(n20336), .ZN(n20304) );
  NAND3_X1 U14664 ( .A1(n20307), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n20304), .ZN(n13560) );
  NOR3_X1 U14665 ( .A1(n20323), .A2(n11598), .A3(n13560), .ZN(n14609) );
  NAND2_X1 U14666 ( .A1(n11586), .A2(n15776), .ZN(n11587) );
  AND2_X1 U14667 ( .A1(n11588), .A2(n11587), .ZN(n11591) );
  OAI21_X1 U14668 ( .B1(n10751), .B2(n10754), .A(n13496), .ZN(n11590) );
  AND4_X1 U14669 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n13142) );
  MUX2_X1 U14670 ( .A(n11594), .B(n13157), .S(n13599), .Z(n11595) );
  NAND3_X1 U14671 ( .A1(n13142), .A2(n11596), .A3(n11595), .ZN(n11597) );
  NAND2_X1 U14672 ( .A1(n11602), .A2(n11597), .ZN(n14608) );
  NAND2_X1 U14673 ( .A1(n20324), .A2(n14614), .ZN(n20338) );
  NAND2_X1 U14674 ( .A1(n20327), .A2(n20338), .ZN(n13558) );
  NOR2_X1 U14675 ( .A1(n20336), .A2(n20350), .ZN(n20303) );
  AND2_X1 U14676 ( .A1(n20303), .A2(n20307), .ZN(n13562) );
  NAND2_X1 U14677 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13562), .ZN(
        n16037) );
  INV_X1 U14678 ( .A(n11598), .ZN(n11609) );
  NAND2_X1 U14679 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11609), .ZN(
        n11608) );
  OR2_X1 U14680 ( .A1(n16037), .A2(n11608), .ZN(n14624) );
  NOR2_X1 U14681 ( .A1(n13558), .A2(n14624), .ZN(n14586) );
  AOI21_X1 U14682 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14609), .A(
        n14586), .ZN(n16010) );
  NAND2_X1 U14683 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14639) );
  NOR3_X1 U14684 ( .A1(n16025), .A2(n14622), .A3(n14639), .ZN(n16002) );
  NAND2_X1 U14685 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16002), .ZN(
        n11607) );
  NAND4_X1 U14686 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11599) );
  OR2_X1 U14687 ( .A1(n11607), .A2(n11599), .ZN(n11600) );
  NAND2_X1 U14688 ( .A1(n11543), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11601) );
  NOR2_X1 U14689 ( .A1(n14592), .A2(n11601), .ZN(n14557) );
  AND2_X1 U14690 ( .A1(n20317), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14063) );
  INV_X1 U14691 ( .A(n14630), .ZN(n20339) );
  INV_X1 U14692 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14531) );
  OR2_X1 U14693 ( .A1(n14608), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11605) );
  INV_X1 U14694 ( .A(n11602), .ZN(n11603) );
  NAND2_X1 U14695 ( .A1(n11603), .A2(n20342), .ZN(n11604) );
  INV_X1 U14696 ( .A(n20325), .ZN(n11606) );
  NAND2_X1 U14697 ( .A1(n14630), .A2(n11606), .ZN(n16057) );
  INV_X1 U14698 ( .A(n16057), .ZN(n11617) );
  INV_X1 U14699 ( .A(n11607), .ZN(n11611) );
  NOR2_X1 U14700 ( .A1(n13560), .A2(n11608), .ZN(n16021) );
  INV_X1 U14701 ( .A(n16037), .ZN(n16054) );
  NAND2_X1 U14702 ( .A1(n16054), .A2(n11609), .ZN(n14611) );
  NAND2_X1 U14703 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11611), .ZN(
        n14607) );
  AOI221_X1 U14704 ( .B1(n14611), .B2(n20327), .C1(n14607), .C2(n20327), .A(
        n20325), .ZN(n11610) );
  OAI221_X1 U14705 ( .B1(n20323), .B2(n11611), .C1(n20323), .C2(n16021), .A(
        n11610), .ZN(n15994) );
  NAND2_X1 U14706 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15831) );
  OAI21_X1 U14707 ( .B1(n15994), .B2(n15831), .A(n16057), .ZN(n15985) );
  INV_X1 U14708 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15986) );
  NOR2_X1 U14709 ( .A1(n11545), .A2(n15986), .ZN(n15993) );
  OR2_X1 U14710 ( .A1(n14630), .A2(n15993), .ZN(n11612) );
  NAND2_X1 U14711 ( .A1(n15985), .A2(n11612), .ZN(n14598) );
  NOR2_X1 U14712 ( .A1(n14630), .A2(n14564), .ZN(n11613) );
  NAND2_X1 U14713 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11614) );
  OAI21_X1 U14714 ( .B1(n14578), .B2(n11614), .A(n16057), .ZN(n14545) );
  OAI21_X1 U14715 ( .B1(n14528), .B2(n11617), .A(n14545), .ZN(n14541) );
  AOI211_X1 U14716 ( .C1(n11615), .C2(n20339), .A(n14531), .B(n14541), .ZN(
        n14529) );
  NOR3_X1 U14717 ( .A1(n14529), .A2(n11617), .A3(n11616), .ZN(n11618) );
  AOI211_X1 U14718 ( .C1(n11619), .C2(n14557), .A(n14063), .B(n11618), .ZN(
        n11620) );
  AOI22_X1 U14719 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14720 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11624), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14721 ( .A1(n11626), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10687), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14722 ( .A1(n11231), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10688), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11628) );
  NAND4_X1 U14723 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11640) );
  AOI22_X1 U14724 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11632), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14725 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13308), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14726 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10723), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14727 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14728 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  NOR2_X1 U14729 ( .A1(n11640), .A2(n11639), .ZN(n11644) );
  NOR2_X1 U14730 ( .A1(n11642), .A2(n11641), .ZN(n11643) );
  XOR2_X1 U14731 ( .A(n11644), .B(n11643), .Z(n11647) );
  AOI22_X1 U14732 ( .A1(n11258), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20625), .ZN(n11645) );
  OAI21_X1 U14733 ( .B1(n11647), .B2(n11646), .A(n11645), .ZN(n11649) );
  INV_X1 U14734 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14048) );
  XNOR2_X1 U14735 ( .A(n13489), .B(n14048), .ZN(n14047) );
  MUX2_X1 U14736 ( .A(n11649), .B(n14047), .S(n10888), .Z(n12626) );
  AOI22_X1 U14737 ( .A1(n11258), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11651), .ZN(n11652) );
  INV_X1 U14738 ( .A(n16097), .ZN(n21005) );
  OAI21_X1 U14739 ( .B1(n11655), .B2(n21005), .A(n15780), .ZN(n11656) );
  NAND2_X1 U14740 ( .A1(n11656), .A2(n15789), .ZN(n11660) );
  INV_X1 U14741 ( .A(n11657), .ZN(n11658) );
  NAND3_X1 U14742 ( .A1(n11658), .A2(n12887), .A3(n16097), .ZN(n11659) );
  NAND2_X1 U14743 ( .A1(n11660), .A2(n11659), .ZN(n13162) );
  NOR2_X1 U14744 ( .A1(n11661), .A2(n13493), .ZN(n11662) );
  AND2_X1 U14745 ( .A1(n14380), .A2(n11664), .ZN(n11665) );
  NOR4_X1 U14746 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11669) );
  NOR4_X1 U14747 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11668) );
  NOR4_X1 U14748 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11667) );
  NOR4_X1 U14749 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11666) );
  AND4_X1 U14750 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11674) );
  NOR4_X1 U14751 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11672) );
  NOR4_X1 U14752 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11671) );
  NOR4_X1 U14753 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11670) );
  AND4_X1 U14754 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n20936), .ZN(
        n11673) );
  NAND2_X1 U14755 ( .A1(n11674), .A2(n11673), .ZN(n11675) );
  AOI22_X1 U14756 ( .A1(n14362), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n14374), .ZN(n11677) );
  INV_X1 U14757 ( .A(n11677), .ZN(n11681) );
  OR3_X1 U14758 ( .A1(n14374), .A2(n13577), .A3(n11678), .ZN(n14042) );
  INV_X1 U14759 ( .A(DATAI_31_), .ZN(n11679) );
  NOR2_X1 U14760 ( .A1(n14042), .A2(n11679), .ZN(n11680) );
  NOR2_X1 U14761 ( .A1(n11681), .A2(n11680), .ZN(n11682) );
  AND2_X4 U14762 ( .A1(n11913), .A2(n16415), .ZN(n11765) );
  AOI22_X1 U14763 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11687) );
  AND2_X4 U14764 ( .A1(n13827), .A2(n16415), .ZN(n11721) );
  AOI22_X1 U14765 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11686) );
  AND2_X4 U14766 ( .A1(n13828), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11916) );
  AND2_X4 U14767 ( .A1(n13828), .A2(n16415), .ZN(n12313) );
  AOI22_X1 U14768 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11685) );
  NAND4_X1 U14769 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11689) );
  AOI22_X1 U14770 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14771 ( .A1(n12300), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11765), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14772 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14773 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11690) );
  NAND4_X1 U14774 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11694) );
  NAND2_X1 U14775 ( .A1(n11694), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11695) );
  AOI22_X1 U14776 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14777 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14778 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14779 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14780 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  NAND2_X1 U14781 ( .A1(n11701), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11708) );
  AOI22_X1 U14782 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14783 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14784 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14785 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14786 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NAND2_X1 U14787 ( .A1(n11706), .A2(n16412), .ZN(n11707) );
  NAND2_X2 U14788 ( .A1(n11708), .A2(n11707), .ZN(n11861) );
  AOI22_X1 U14789 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14790 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14791 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14792 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11710) );
  AND4_X1 U14793 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11714) );
  NAND2_X1 U14794 ( .A1(n11714), .A2(n16412), .ZN(n11720) );
  AOI22_X1 U14795 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14796 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14797 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14798 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U14799 ( .A1(n10509), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11719) );
  NAND2_X2 U14800 ( .A1(n11720), .A2(n11719), .ZN(n19452) );
  AOI22_X1 U14801 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14802 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14803 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14804 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14805 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11731) );
  AOI22_X1 U14806 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14807 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14808 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9808), .ZN(n11726) );
  NAND4_X1 U14809 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11730) );
  MUX2_X2 U14810 ( .A(n11731), .B(n11730), .S(n16412), .Z(n12604) );
  AOI22_X1 U14811 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14812 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14813 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14814 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14815 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14816 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14817 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14818 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U14819 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11742) );
  NAND2_X2 U14820 ( .A1(n11743), .A2(n11742), .ZN(n11792) );
  INV_X2 U14821 ( .A(n11792), .ZN(n12949) );
  NAND2_X1 U14822 ( .A1(n12947), .A2(n12949), .ZN(n11747) );
  NAND3_X1 U14823 ( .A1(n19452), .A2(n9811), .A3(n11861), .ZN(n11775) );
  INV_X1 U14824 ( .A(n11775), .ZN(n11745) );
  NAND2_X1 U14825 ( .A1(n12955), .A2(n11792), .ZN(n11746) );
  NAND2_X1 U14826 ( .A1(n11747), .A2(n11746), .ZN(n11838) );
  AOI22_X1 U14827 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14828 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14829 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14830 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U14831 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  AOI22_X1 U14832 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14833 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14834 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14835 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U14836 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11757) );
  NAND2_X1 U14837 ( .A1(n11757), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11758) );
  NAND2_X2 U14838 ( .A1(n11759), .A2(n11758), .ZN(n12952) );
  AOI22_X1 U14839 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14840 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14841 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14842 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11760) );
  NAND4_X1 U14843 ( .A1(n11762), .A2(n11763), .A3(n11761), .A4(n11760), .ZN(
        n11764) );
  AOI22_X1 U14844 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14845 ( .A1(n9803), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14846 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14847 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11767) );
  NAND4_X1 U14848 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11771) );
  NAND2_X2 U14849 ( .A1(n11773), .A2(n11772), .ZN(n11819) );
  OAI21_X1 U14850 ( .B1(n11826), .B2(n11776), .A(n11775), .ZN(n11790) );
  AOI22_X1 U14851 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14852 ( .A1(n11778), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14853 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14854 ( .A1(n11781), .A2(n10510), .A3(n11780), .A4(n11779), .ZN(
        n11788) );
  AOI22_X1 U14855 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12313), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14856 ( .A1(n11765), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14857 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11709), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14858 ( .A1(n12299), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11721), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14859 ( .A1(n9909), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11787) );
  NAND2_X1 U14860 ( .A1(n11795), .A2(n12949), .ZN(n11789) );
  NAND3_X1 U14861 ( .A1(n11790), .A2(n19439), .A3(n11789), .ZN(n11794) );
  INV_X2 U14862 ( .A(n12952), .ZN(n16440) );
  AND2_X2 U14863 ( .A1(n12604), .A2(n11861), .ZN(n12622) );
  NAND2_X2 U14864 ( .A1(n19439), .A2(n11792), .ZN(n12956) );
  NAND3_X1 U14865 ( .A1(n11799), .A2(n12622), .A3(n12956), .ZN(n11793) );
  NAND3_X1 U14866 ( .A1(n11794), .A2(n16440), .A3(n11793), .ZN(n12962) );
  INV_X4 U14867 ( .A(n11819), .ZN(n12403) );
  AND2_X1 U14868 ( .A1(n11795), .A2(n12403), .ZN(n12957) );
  NAND2_X1 U14869 ( .A1(n11837), .A2(n16440), .ZN(n11796) );
  NAND3_X1 U14870 ( .A1(n12813), .A2(n19439), .A3(n13442), .ZN(n12939) );
  AND4_X2 U14871 ( .A1(n19452), .A2(n19439), .A3(n12604), .A4(n12949), .ZN(
        n11802) );
  INV_X1 U14872 ( .A(n11808), .ZN(n11801) );
  NAND2_X1 U14873 ( .A1(n11802), .A2(n11801), .ZN(n12387) );
  NAND2_X1 U14874 ( .A1(n12952), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12354) );
  AND2_X1 U14875 ( .A1(n12387), .A2(n14671), .ZN(n11798) );
  NAND2_X1 U14876 ( .A1(n12403), .A2(n19439), .ZN(n12394) );
  NOR2_X1 U14877 ( .A1(n11791), .A2(n12949), .ZN(n11800) );
  NAND4_X1 U14878 ( .A1(n9816), .A2(n16440), .A3(n12622), .A4(n11800), .ZN(
        n12931) );
  NAND2_X1 U14879 ( .A1(n19034), .A2(n13767), .ZN(n16459) );
  OAI21_X1 U14880 ( .B1(n16459), .B2(n20078), .A(n11803), .ZN(n11804) );
  AOI21_X1 U14881 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n11807), .A(n11804), 
        .ZN(n11805) );
  NOR2_X1 U14882 ( .A1(n11808), .A2(n11819), .ZN(n11809) );
  NAND2_X1 U14883 ( .A1(n11809), .A2(n11792), .ZN(n11811) );
  NAND2_X1 U14884 ( .A1(n12444), .A2(n12949), .ZN(n11810) );
  NAND2_X1 U14885 ( .A1(n11811), .A2(n11810), .ZN(n11825) );
  OAI21_X2 U14886 ( .B1(n11819), .B2(n12952), .A(n11817), .ZN(n14674) );
  INV_X1 U14887 ( .A(n14674), .ZN(n11812) );
  NAND2_X1 U14888 ( .A1(n11825), .A2(n11813), .ZN(n12933) );
  NAND2_X1 U14889 ( .A1(n9837), .A2(n12933), .ZN(n11814) );
  NAND2_X1 U14890 ( .A1(n11814), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U14891 ( .A1(n11820), .A2(n12403), .ZN(n11815) );
  NAND2_X2 U14892 ( .A1(n11816), .A2(n11815), .ZN(n11891) );
  INV_X1 U14893 ( .A(n12955), .ZN(n12397) );
  NAND2_X2 U14894 ( .A1(n12965), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11892) );
  INV_X1 U14895 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U14896 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11821) );
  OAI211_X1 U14897 ( .C1(n11892), .C2(n11823), .A(n11822), .B(n11821), .ZN(
        n11824) );
  AOI21_X2 U14898 ( .B1(n11891), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11824), .ZN(n11849) );
  NAND2_X1 U14899 ( .A1(n11833), .A2(n12364), .ZN(n11829) );
  INV_X1 U14900 ( .A(n11826), .ZN(n11827) );
  AND2_X1 U14901 ( .A1(n14674), .A2(n11827), .ZN(n11828) );
  NAND2_X1 U14902 ( .A1(n11825), .A2(n11828), .ZN(n13794) );
  NAND2_X1 U14903 ( .A1(n11829), .A2(n13794), .ZN(n11832) );
  NOR2_X1 U14904 ( .A1(n12956), .A2(n19034), .ZN(n11831) );
  NOR2_X1 U14905 ( .A1(n16459), .A2(n20086), .ZN(n11830) );
  AOI21_X1 U14906 ( .B1(n11832), .B2(n11831), .A(n11830), .ZN(n11835) );
  NAND2_X1 U14907 ( .A1(n11888), .A2(n11833), .ZN(n11834) );
  NAND2_X1 U14908 ( .A1(n11835), .A2(n11834), .ZN(n11873) );
  NAND2_X1 U14909 ( .A1(n11891), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11848) );
  INV_X1 U14910 ( .A(n11836), .ZN(n11839) );
  INV_X1 U14911 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11841) );
  INV_X1 U14912 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11840) );
  OAI22_X1 U14913 ( .A1(n11892), .A2(n11841), .B1(n12713), .B2(n11840), .ZN(
        n11845) );
  NAND2_X1 U14914 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11842) );
  NAND3_X1 U14915 ( .A1(n11843), .A2(n16459), .A3(n11842), .ZN(n11844) );
  NOR2_X1 U14916 ( .A1(n11845), .A2(n11844), .ZN(n11846) );
  AOI21_X1 U14917 ( .B1(n19034), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U14918 ( .A1(n11852), .A2(n11851), .ZN(n11886) );
  INV_X1 U14919 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11855) );
  INV_X2 U14920 ( .A(n12713), .ZN(n12721) );
  NAND2_X1 U14921 ( .A1(n12721), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11854) );
  NAND2_X1 U14922 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11853) );
  OAI211_X1 U14923 ( .C1(n11892), .C2(n11855), .A(n11854), .B(n11853), .ZN(
        n11856) );
  INV_X1 U14924 ( .A(n11856), .ZN(n11858) );
  NAND2_X1 U14925 ( .A1(n11891), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11857) );
  INV_X1 U14926 ( .A(n11885), .ZN(n11859) );
  NAND2_X1 U14927 ( .A1(n11861), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U14928 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19756) );
  NAND2_X1 U14929 ( .A1(n19756), .A2(n20069), .ZN(n11864) );
  NAND2_X1 U14930 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19855) );
  INV_X1 U14931 ( .A(n19855), .ZN(n11863) );
  NAND2_X1 U14932 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11863), .ZN(
        n11897) );
  NAND2_X1 U14933 ( .A1(n11864), .A2(n11897), .ZN(n19575) );
  NOR2_X1 U14934 ( .A1(n19861), .A2(n19575), .ZN(n11865) );
  AOI21_X1 U14935 ( .B1(n11901), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11865), .ZN(n11866) );
  NAND2_X1 U14936 ( .A1(n11867), .A2(n11866), .ZN(n11871) );
  INV_X1 U14937 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11869) );
  NOR2_X1 U14938 ( .A1(n12227), .A2(n11869), .ZN(n11870) );
  AOI22_X1 U14939 ( .A1(n11901), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20057), .B2(n20086), .ZN(n11875) );
  NAND2_X1 U14940 ( .A1(n11901), .A2(n13837), .ZN(n11878) );
  NAND2_X1 U14941 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20078), .ZN(
        n19479) );
  NAND2_X1 U14942 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20086), .ZN(
        n19508) );
  NAND2_X1 U14943 ( .A1(n19479), .A2(n19508), .ZN(n19574) );
  NAND2_X1 U14944 ( .A1(n20057), .A2(n19574), .ZN(n19509) );
  NAND2_X1 U14945 ( .A1(n11878), .A2(n19509), .ZN(n11879) );
  NAND2_X1 U14946 ( .A1(n13003), .A2(n11880), .ZN(n11881) );
  NAND2_X1 U14947 ( .A1(n12995), .A2(n11881), .ZN(n12987) );
  NAND2_X1 U14948 ( .A1(n11886), .A2(n11885), .ZN(n11884) );
  NAND2_X1 U14949 ( .A1(n11888), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11890) );
  OR2_X1 U14950 ( .A1(n16459), .A2(n20062), .ZN(n11889) );
  NAND2_X1 U14951 ( .A1(n11890), .A2(n11889), .ZN(n12698) );
  INV_X1 U14952 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U14953 ( .A1(n12721), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11894) );
  NAND2_X1 U14954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11893) );
  XNOR2_X2 U14955 ( .A(n12695), .B(n12694), .ZN(n13364) );
  INV_X1 U14956 ( .A(n11897), .ZN(n11898) );
  NAND2_X1 U14957 ( .A1(n11898), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19427) );
  OAI211_X1 U14958 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n11898), .A(
        n19427), .B(n20057), .ZN(n11899) );
  INV_X1 U14959 ( .A(n11899), .ZN(n11900) );
  AOI21_X1 U14960 ( .B1(n11901), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11900), .ZN(n11902) );
  INV_X1 U14961 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13418) );
  NOR2_X1 U14962 ( .A1(n12227), .A2(n13418), .ZN(n11903) );
  NAND2_X1 U14963 ( .A1(n11861), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11904) );
  AND2_X1 U14964 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11907) );
  INV_X1 U14965 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11906) );
  NOR2_X1 U14966 ( .A1(n12227), .A2(n11906), .ZN(n13011) );
  AND2_X2 U14967 ( .A1(n9848), .A2(n16412), .ZN(n12429) );
  AOI22_X1 U14968 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11912) );
  AND2_X2 U14969 ( .A1(n9852), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12427) );
  AOI22_X1 U14970 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11911) );
  AND2_X2 U14971 ( .A1(n9848), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12135) );
  AOI22_X1 U14972 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11910) );
  AND2_X2 U14973 ( .A1(n12313), .A2(n16412), .ZN(n12014) );
  AOI22_X1 U14974 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12014), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11909) );
  NAND4_X1 U14975 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11926) );
  NAND2_X1 U14976 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12145) );
  INV_X1 U14977 ( .A(n12145), .ZN(n11914) );
  NAND3_X1 U14978 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13837), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12807) );
  INV_X1 U14979 ( .A(n12807), .ZN(n11915) );
  AOI22_X1 U14980 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11920) );
  INV_X2 U14981 ( .A(n10501), .ZN(n12534) );
  NAND2_X1 U14982 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11919) );
  AND2_X1 U14983 ( .A1(n9808), .A2(n16412), .ZN(n12435) );
  NAND2_X1 U14984 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11918) );
  AOI22_X1 U14985 ( .A1(n12494), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11924) );
  AND2_X2 U14986 ( .A1(n11783), .A2(n16412), .ZN(n12434) );
  NAND2_X1 U14987 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11923) );
  AND2_X2 U14988 ( .A1(n9852), .A2(n16412), .ZN(n12426) );
  NAND2_X1 U14989 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U14990 ( .A1(n10499), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11925) );
  NOR2_X1 U14991 ( .A1(n11926), .A2(n11925), .ZN(n13103) );
  AOI22_X1 U14992 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14993 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14994 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U14995 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U14996 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11939) );
  AOI22_X1 U14997 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12414), .ZN(n11937) );
  AOI22_X1 U14998 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12546), .ZN(n11934) );
  NAND2_X1 U14999 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U15000 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11932) );
  AND3_X1 U15001 ( .A1(n11934), .A2(n11933), .A3(n11932), .ZN(n11936) );
  INV_X1 U15002 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15003 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11935) );
  NAND3_X1 U15004 ( .A1(n11937), .A2(n11936), .A3(n11935), .ZN(n11938) );
  NOR2_X2 U15005 ( .A1(n13104), .A2(n13108), .ZN(n13176) );
  AOI22_X1 U15006 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15007 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12546), .ZN(n11942) );
  NAND2_X1 U15008 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U15009 ( .A1(n12414), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11940) );
  AND3_X1 U15010 ( .A1(n11942), .A2(n11941), .A3(n11940), .ZN(n11944) );
  AOI22_X1 U15011 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n12435), .ZN(n11943) );
  NAND3_X1 U15012 ( .A1(n11945), .A2(n11944), .A3(n11943), .ZN(n11951) );
  AOI22_X1 U15013 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15014 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15015 ( .A1(n12113), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15016 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U15017 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11950) );
  INV_X1 U15018 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13429) );
  INV_X1 U15019 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13432) );
  INV_X1 U15020 ( .A(n12414), .ZN(n11992) );
  OAI22_X1 U15021 ( .A1(n12009), .A2(n13429), .B1(n13432), .B2(n11992), .ZN(
        n11953) );
  INV_X1 U15022 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13415) );
  OAI22_X1 U15023 ( .A1(n13415), .A2(n10197), .B1(n12131), .B2(n13418), .ZN(
        n11952) );
  OR2_X1 U15024 ( .A1(n11953), .A2(n11952), .ZN(n11959) );
  AOI22_X1 U15025 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12546), .ZN(n11957) );
  NAND2_X1 U15026 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11956) );
  NAND2_X1 U15027 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11955) );
  NAND3_X1 U15028 ( .A1(n11957), .A2(n11956), .A3(n11955), .ZN(n11958) );
  NOR2_X1 U15029 ( .A1(n11959), .A2(n11958), .ZN(n11974) );
  INV_X1 U15030 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13430) );
  INV_X1 U15031 ( .A(n12426), .ZN(n11962) );
  INV_X1 U15032 ( .A(n12427), .ZN(n11961) );
  INV_X1 U15033 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11960) );
  OAI22_X1 U15034 ( .A1(n13430), .A2(n11962), .B1(n11961), .B2(n11960), .ZN(
        n11966) );
  INV_X1 U15035 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13417) );
  INV_X1 U15036 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13428) );
  OAI22_X1 U15037 ( .A1(n13417), .A2(n11964), .B1(n11963), .B2(n13428), .ZN(
        n11965) );
  NOR2_X1 U15038 ( .A1(n11966), .A2(n11965), .ZN(n11973) );
  INV_X1 U15039 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13427) );
  INV_X1 U15040 ( .A(n12135), .ZN(n11968) );
  INV_X1 U15041 ( .A(n12113), .ZN(n11967) );
  INV_X1 U15042 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13431) );
  OAI22_X1 U15043 ( .A1(n13427), .A2(n11968), .B1(n11967), .B2(n13431), .ZN(
        n11971) );
  INV_X1 U15044 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13433) );
  INV_X1 U15045 ( .A(n12014), .ZN(n11969) );
  INV_X1 U15046 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13435) );
  OAI22_X1 U15047 ( .A1(n13433), .A2(n11969), .B1(n10501), .B2(n13435), .ZN(
        n11970) );
  NOR2_X1 U15048 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  AOI22_X1 U15049 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12541), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15050 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15051 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15052 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15053 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11986) );
  AOI22_X1 U15054 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n12435), .ZN(n11984) );
  AOI22_X1 U15055 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15056 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12546), .ZN(n11981) );
  NAND2_X1 U15057 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11980) );
  NAND2_X1 U15058 ( .A1(n12414), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11979) );
  AND3_X1 U15059 ( .A1(n11981), .A2(n11980), .A3(n11979), .ZN(n11982) );
  NAND3_X1 U15060 ( .A1(n11984), .A2(n11983), .A3(n11982), .ZN(n11985) );
  NOR2_X1 U15061 ( .A1(n11986), .A2(n11985), .ZN(n13293) );
  NAND2_X1 U15062 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U15063 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U15064 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U15065 ( .A1(n12428), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11988) );
  AND4_X1 U15066 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n12005) );
  INV_X1 U15067 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13640) );
  INV_X1 U15068 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13658) );
  OAI22_X1 U15069 ( .A1(n12009), .A2(n13640), .B1(n11992), .B2(n13658), .ZN(
        n11994) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13650) );
  INV_X1 U15071 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12103) );
  OAI22_X1 U15072 ( .A1(n10197), .A2(n13650), .B1(n12131), .B2(n12103), .ZN(
        n11993) );
  NOR2_X1 U15073 ( .A1(n11994), .A2(n11993), .ZN(n12004) );
  AOI22_X1 U15074 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U15075 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U15076 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11995) );
  AND3_X1 U15077 ( .A1(n11997), .A2(n11996), .A3(n11995), .ZN(n12003) );
  NAND2_X1 U15078 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U15079 ( .A1(n12113), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12000) );
  NAND2_X1 U15080 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U15081 ( .A1(n12014), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11998) );
  AND4_X1 U15082 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12002) );
  NAND4_X1 U15083 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n13346) );
  AOI22_X1 U15084 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12546), .ZN(n12008) );
  NAND2_X1 U15085 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12007) );
  NAND2_X1 U15086 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12006) );
  AND3_X1 U15087 ( .A1(n12008), .A2(n12007), .A3(n12006), .ZN(n12013) );
  AOI22_X1 U15088 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12494), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15089 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U15090 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12010) );
  NAND4_X1 U15091 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12020) );
  AOI22_X1 U15092 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12541), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15093 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15094 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15095 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U15096 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12019) );
  AOI22_X1 U15097 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n12414), .ZN(n12028) );
  AOI22_X1 U15098 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12546), .ZN(n12023) );
  NAND2_X1 U15099 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12022) );
  NAND2_X1 U15100 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12021) );
  AND3_X1 U15101 ( .A1(n12023), .A2(n12022), .A3(n12021), .ZN(n12027) );
  INV_X1 U15102 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12306) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12024) );
  OAI22_X1 U15104 ( .A1(n12306), .A2(n10197), .B1(n12131), .B2(n12024), .ZN(
        n12025) );
  INV_X1 U15105 ( .A(n12025), .ZN(n12026) );
  NAND3_X1 U15106 ( .A1(n12028), .A2(n12027), .A3(n12026), .ZN(n12034) );
  AOI22_X1 U15107 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15108 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15109 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15110 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15111 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12033) );
  AOI22_X1 U15112 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15113 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U15114 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12036) );
  NAND2_X1 U15115 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12035) );
  AND3_X1 U15116 ( .A1(n12037), .A2(n12036), .A3(n12035), .ZN(n12039) );
  AOI22_X1 U15117 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12038) );
  NAND3_X1 U15118 ( .A1(n12040), .A2(n12039), .A3(n12038), .ZN(n12046) );
  AOI22_X1 U15119 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12426), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15120 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15121 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15122 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12014), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12041) );
  NAND4_X1 U15123 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12045) );
  AOI22_X1 U15124 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15125 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15126 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15127 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15128 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12060) );
  AOI22_X1 U15129 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n12414), .ZN(n12058) );
  INV_X1 U15130 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13388) );
  NOR2_X1 U15131 ( .A1(n12415), .A2(n13388), .ZN(n12054) );
  INV_X1 U15132 ( .A(n12809), .ZN(n12104) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12051) );
  INV_X1 U15134 ( .A(n12546), .ZN(n12102) );
  OAI22_X1 U15135 ( .A1(n12104), .A2(n12052), .B1(n12051), .B2(n12102), .ZN(
        n12053) );
  NOR2_X1 U15136 ( .A1(n12054), .A2(n12053), .ZN(n12057) );
  AOI22_X1 U15137 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15138 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12055) );
  NAND4_X1 U15139 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12059) );
  AOI22_X1 U15140 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15141 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15142 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15143 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12061) );
  NAND4_X1 U15144 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12072) );
  AOI22_X1 U15145 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n12414), .ZN(n12070) );
  AOI22_X1 U15146 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12546), .ZN(n12067) );
  NAND2_X1 U15147 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12066) );
  NAND2_X1 U15148 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12065) );
  AND3_X1 U15149 ( .A1(n12067), .A2(n12066), .A3(n12065), .ZN(n12069) );
  AOI22_X1 U15150 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12068) );
  NAND3_X1 U15151 ( .A1(n12070), .A2(n12069), .A3(n12068), .ZN(n12071) );
  NOR2_X1 U15152 ( .A1(n12072), .A2(n12071), .ZN(n13757) );
  AOI22_X1 U15153 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15154 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15155 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15156 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U15157 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12084) );
  AOI22_X1 U15158 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n12414), .ZN(n12082) );
  NOR2_X1 U15159 ( .A1(n12415), .A2(n13433), .ZN(n12078) );
  OAI22_X1 U15160 ( .A1(n12104), .A2(n13418), .B1(n13417), .B2(n12102), .ZN(
        n12077) );
  NOR2_X1 U15161 ( .A1(n12078), .A2(n12077), .ZN(n12081) );
  AOI22_X1 U15162 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U15163 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12079) );
  NAND4_X1 U15164 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12083) );
  AOI22_X1 U15165 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n12414), .ZN(n12090) );
  AOI22_X1 U15166 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12546), .ZN(n12087) );
  NAND2_X1 U15167 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12086) );
  NAND2_X1 U15168 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12085) );
  AND3_X1 U15169 ( .A1(n12087), .A2(n12086), .A3(n12085), .ZN(n12089) );
  AOI22_X1 U15170 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12088) );
  NAND3_X1 U15171 ( .A1(n12090), .A2(n12089), .A3(n12088), .ZN(n12096) );
  AOI22_X1 U15172 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15173 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15174 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15175 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15176 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12095) );
  OR2_X1 U15177 ( .A1(n12096), .A2(n12095), .ZN(n14764) );
  INV_X1 U15178 ( .A(n14750), .ZN(n12127) );
  AOI22_X1 U15179 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12426), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15180 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15181 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15182 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12014), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12097) );
  NAND4_X1 U15183 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12112) );
  AOI22_X1 U15184 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12110) );
  INV_X1 U15185 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12101) );
  NOR2_X1 U15186 ( .A1(n12415), .A2(n12101), .ZN(n12106) );
  INV_X1 U15187 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13649) );
  OAI22_X1 U15188 ( .A1(n12104), .A2(n12103), .B1(n12102), .B2(n13649), .ZN(
        n12105) );
  NOR2_X1 U15189 ( .A1(n12106), .A2(n12105), .ZN(n12109) );
  AOI22_X1 U15190 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U15191 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12107) );
  NAND4_X1 U15192 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12111) );
  NOR2_X1 U15193 ( .A1(n12112), .A2(n12111), .ZN(n14757) );
  AOI22_X1 U15194 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15195 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15196 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15197 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U15198 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12125) );
  AOI22_X1 U15199 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n12414), .ZN(n12123) );
  AOI22_X1 U15200 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12546), .ZN(n12120) );
  NAND2_X1 U15201 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12119) );
  NAND2_X1 U15202 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12118) );
  AND3_X1 U15203 ( .A1(n12120), .A2(n12119), .A3(n12118), .ZN(n12122) );
  AOI22_X1 U15204 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12121) );
  NAND3_X1 U15205 ( .A1(n12123), .A2(n12122), .A3(n12121), .ZN(n12124) );
  NOR2_X1 U15206 ( .A1(n12125), .A2(n12124), .ZN(n14751) );
  NOR2_X1 U15207 ( .A1(n14757), .A2(n14751), .ZN(n12126) );
  AOI22_X1 U15208 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n12414), .ZN(n12134) );
  AOI22_X1 U15209 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12546), .ZN(n12130) );
  NAND2_X1 U15210 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U15211 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12128) );
  AND3_X1 U15212 ( .A1(n12130), .A2(n12129), .A3(n12128), .ZN(n12133) );
  AOI22_X1 U15213 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12132) );
  NAND3_X1 U15214 ( .A1(n12134), .A2(n12133), .A3(n12132), .ZN(n12141) );
  AOI22_X1 U15215 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15216 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15217 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15218 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15219 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  OR2_X1 U15220 ( .A1(n12141), .A2(n12140), .ZN(n12166) );
  AOI22_X1 U15221 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11783), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12151) );
  INV_X1 U15222 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12143) );
  INV_X1 U15223 ( .A(n12313), .ZN(n12304) );
  INV_X1 U15224 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12142) );
  OAI22_X1 U15225 ( .A1(n11908), .A2(n12143), .B1(n12304), .B2(n12142), .ZN(
        n12148) );
  INV_X1 U15226 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19552) );
  INV_X1 U15227 ( .A(n12300), .ZN(n12307) );
  INV_X1 U15228 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12144) );
  OR2_X1 U15229 ( .A1(n12307), .A2(n12144), .ZN(n12146) );
  OAI21_X1 U15230 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n12145), .ZN(n12305) );
  OAI211_X1 U15231 ( .C1(n13773), .C2(n19552), .A(n12146), .B(n12305), .ZN(
        n12147) );
  NOR2_X1 U15232 ( .A1(n12148), .A2(n12147), .ZN(n12150) );
  AOI22_X1 U15233 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12149) );
  NAND3_X1 U15234 ( .A1(n12151), .A2(n12150), .A3(n12149), .ZN(n12160) );
  AOI22_X1 U15235 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15236 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15237 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12156) );
  INV_X1 U15238 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13292) );
  INV_X1 U15239 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12152) );
  OR2_X1 U15240 ( .A1(n12307), .A2(n12152), .ZN(n12153) );
  INV_X1 U15241 ( .A(n12305), .ZN(n12275) );
  OAI211_X1 U15242 ( .C1(n12304), .C2(n13292), .A(n12153), .B(n12275), .ZN(
        n12154) );
  INV_X1 U15243 ( .A(n12154), .ZN(n12155) );
  NAND4_X1 U15244 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12159) );
  AND2_X1 U15245 ( .A1(n12160), .A2(n12159), .ZN(n12165) );
  NAND2_X1 U15246 ( .A1(n13000), .A2(n12165), .ZN(n12161) );
  XNOR2_X1 U15247 ( .A(n12166), .B(n12161), .ZN(n12186) );
  INV_X1 U15248 ( .A(n12165), .ZN(n12184) );
  NOR2_X1 U15249 ( .A1(n13000), .A2(n12184), .ZN(n14743) );
  INV_X1 U15250 ( .A(n12186), .ZN(n12163) );
  AND2_X1 U15251 ( .A1(n12166), .A2(n12165), .ZN(n12182) );
  AOI22_X1 U15252 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9848), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15253 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15254 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12170) );
  INV_X1 U15255 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13371) );
  INV_X1 U15256 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13392) );
  OR2_X1 U15257 ( .A1(n12307), .A2(n13392), .ZN(n12167) );
  OAI211_X1 U15258 ( .C1(n12304), .C2(n13371), .A(n12167), .B(n12305), .ZN(
        n12168) );
  INV_X1 U15259 ( .A(n12168), .ZN(n12169) );
  NAND4_X1 U15260 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12181) );
  AOI22_X1 U15261 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9848), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15262 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15263 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12177) );
  INV_X1 U15264 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12174) );
  INV_X1 U15265 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13404) );
  OR2_X1 U15266 ( .A1(n12307), .A2(n13404), .ZN(n12173) );
  OAI211_X1 U15267 ( .C1(n12304), .C2(n12174), .A(n12173), .B(n12275), .ZN(
        n12175) );
  INV_X1 U15268 ( .A(n12175), .ZN(n12176) );
  NAND4_X1 U15269 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12180) );
  AND2_X1 U15270 ( .A1(n12181), .A2(n12180), .ZN(n12183) );
  NAND2_X1 U15271 ( .A1(n12182), .A2(n12183), .ZN(n12188) );
  OAI211_X1 U15272 ( .C1(n12182), .C2(n12183), .A(n12253), .B(n12188), .ZN(
        n14730) );
  NAND2_X1 U15273 ( .A1(n12403), .A2(n12183), .ZN(n14733) );
  NOR2_X1 U15274 ( .A1(n14733), .A2(n12184), .ZN(n12185) );
  INV_X1 U15275 ( .A(n12188), .ZN(n12207) );
  AOI22_X1 U15276 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9848), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15277 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15278 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12194) );
  INV_X1 U15279 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12191) );
  INV_X1 U15280 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12189) );
  OR2_X1 U15281 ( .A1(n12307), .A2(n12189), .ZN(n12190) );
  OAI211_X1 U15282 ( .C1(n12304), .C2(n12191), .A(n12190), .B(n12305), .ZN(
        n12192) );
  INV_X1 U15283 ( .A(n12192), .ZN(n12193) );
  NAND4_X1 U15284 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12206) );
  AOI22_X1 U15285 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9848), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15286 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15287 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12202) );
  INV_X1 U15288 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12199) );
  INV_X1 U15289 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12197) );
  OR2_X1 U15290 ( .A1(n12307), .A2(n12197), .ZN(n12198) );
  OAI211_X1 U15291 ( .C1(n12304), .C2(n12199), .A(n12198), .B(n12275), .ZN(
        n12200) );
  INV_X1 U15292 ( .A(n12200), .ZN(n12201) );
  NAND4_X1 U15293 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12205) );
  NAND2_X1 U15294 ( .A1(n12207), .A2(n12209), .ZN(n12228) );
  OAI211_X1 U15295 ( .C1(n12207), .C2(n12209), .A(n12228), .B(n12253), .ZN(
        n12211) );
  INV_X1 U15296 ( .A(n12211), .ZN(n12208) );
  XNOR2_X1 U15297 ( .A(n12212), .B(n12208), .ZN(n14722) );
  INV_X1 U15298 ( .A(n12209), .ZN(n12210) );
  NOR2_X1 U15299 ( .A1(n13000), .A2(n12210), .ZN(n14724) );
  NAND2_X1 U15300 ( .A1(n14722), .A2(n14724), .ZN(n14723) );
  AOI22_X1 U15301 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9848), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15302 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15303 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12216) );
  OR2_X1 U15304 ( .A1(n12307), .A2(n13415), .ZN(n12213) );
  OAI211_X1 U15305 ( .C1(n12304), .C2(n13429), .A(n12213), .B(n12305), .ZN(
        n12214) );
  INV_X1 U15306 ( .A(n12214), .ZN(n12215) );
  NAND4_X1 U15307 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12226) );
  AOI22_X1 U15308 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9848), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15309 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15310 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12222) );
  INV_X1 U15311 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19914) );
  OR2_X1 U15312 ( .A1(n12307), .A2(n13431), .ZN(n12219) );
  OAI211_X1 U15313 ( .C1(n12304), .C2(n19914), .A(n12219), .B(n12275), .ZN(
        n12220) );
  INV_X1 U15314 ( .A(n12220), .ZN(n12221) );
  NAND4_X1 U15315 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12225) );
  NAND2_X1 U15316 ( .A1(n12226), .A2(n12225), .ZN(n12230) );
  AOI21_X1 U15317 ( .B1(n12228), .B2(n12230), .A(n12227), .ZN(n12229) );
  OR2_X1 U15318 ( .A1(n12228), .A2(n12230), .ZN(n12252) );
  INV_X1 U15319 ( .A(n12230), .ZN(n12231) );
  NAND2_X1 U15320 ( .A1(n12403), .A2(n12231), .ZN(n14715) );
  AOI22_X1 U15321 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9848), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15322 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15323 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12239) );
  INV_X1 U15324 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12236) );
  INV_X1 U15325 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12234) );
  OR2_X1 U15326 ( .A1(n12307), .A2(n12234), .ZN(n12235) );
  OAI211_X1 U15327 ( .C1(n12304), .C2(n12236), .A(n12235), .B(n12305), .ZN(
        n12237) );
  INV_X1 U15328 ( .A(n12237), .ZN(n12238) );
  NAND4_X1 U15329 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12251) );
  AOI22_X1 U15330 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9848), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15331 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15332 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12247) );
  INV_X1 U15333 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12244) );
  INV_X1 U15334 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12242) );
  OR2_X1 U15335 ( .A1(n12307), .A2(n12242), .ZN(n12243) );
  OAI211_X1 U15336 ( .C1(n12304), .C2(n12244), .A(n12243), .B(n12275), .ZN(
        n12245) );
  INV_X1 U15337 ( .A(n12245), .ZN(n12246) );
  NAND4_X1 U15338 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12250) );
  NAND2_X1 U15339 ( .A1(n12251), .A2(n12250), .ZN(n12257) );
  INV_X1 U15340 ( .A(n12257), .ZN(n12255) );
  INV_X1 U15341 ( .A(n12252), .ZN(n12254) );
  OAI211_X1 U15342 ( .C1(n12255), .C2(n12254), .A(n12291), .B(n12253), .ZN(
        n12256) );
  NOR2_X1 U15343 ( .A1(n13000), .A2(n12257), .ZN(n14707) );
  AOI22_X1 U15344 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9848), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15345 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15346 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12262) );
  OR2_X1 U15347 ( .A1(n12307), .A2(n13650), .ZN(n12259) );
  OAI211_X1 U15348 ( .C1(n12304), .C2(n13640), .A(n12259), .B(n12305), .ZN(
        n12260) );
  INV_X1 U15349 ( .A(n12260), .ZN(n12261) );
  NAND4_X1 U15350 ( .A1(n12264), .A2(n12263), .A3(n12262), .A4(n12261), .ZN(
        n12274) );
  AOI22_X1 U15351 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9848), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15352 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15353 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12270) );
  INV_X1 U15354 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12267) );
  INV_X1 U15355 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13655) );
  OR2_X1 U15356 ( .A1(n12307), .A2(n13655), .ZN(n12266) );
  OAI211_X1 U15357 ( .C1(n12304), .C2(n12267), .A(n12266), .B(n12275), .ZN(
        n12268) );
  INV_X1 U15358 ( .A(n12268), .ZN(n12269) );
  NAND4_X1 U15359 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(
        n12273) );
  NAND2_X1 U15360 ( .A1(n12274), .A2(n12273), .ZN(n14699) );
  AOI22_X1 U15361 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11783), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12282) );
  INV_X1 U15362 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14892) );
  INV_X1 U15363 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19935) );
  OAI22_X1 U15364 ( .A1(n11908), .A2(n14892), .B1(n12304), .B2(n19935), .ZN(
        n12279) );
  INV_X1 U15365 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12277) );
  INV_X1 U15366 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14896) );
  OR2_X1 U15367 ( .A1(n12307), .A2(n14896), .ZN(n12276) );
  OAI211_X1 U15368 ( .C1(n13773), .C2(n12277), .A(n12276), .B(n12275), .ZN(
        n12278) );
  NOR2_X1 U15369 ( .A1(n12279), .A2(n12278), .ZN(n12281) );
  AOI22_X1 U15370 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12280) );
  NAND3_X1 U15371 ( .A1(n12282), .A2(n12281), .A3(n12280), .ZN(n12290) );
  AOI22_X1 U15372 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11778), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15373 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15374 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12286) );
  INV_X1 U15375 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14877) );
  INV_X1 U15376 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14888) );
  OR2_X1 U15377 ( .A1(n12307), .A2(n14888), .ZN(n12283) );
  OAI211_X1 U15378 ( .C1(n12304), .C2(n14877), .A(n12283), .B(n12305), .ZN(
        n12284) );
  INV_X1 U15379 ( .A(n12284), .ZN(n12285) );
  NAND4_X1 U15380 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12289) );
  NAND2_X1 U15381 ( .A1(n12290), .A2(n12289), .ZN(n12295) );
  INV_X1 U15382 ( .A(n12291), .ZN(n14698) );
  INV_X1 U15383 ( .A(n14699), .ZN(n12292) );
  AND2_X1 U15384 ( .A1(n13000), .A2(n12292), .ZN(n12293) );
  NAND2_X1 U15385 ( .A1(n14698), .A2(n12293), .ZN(n12294) );
  NOR2_X1 U15386 ( .A1(n12294), .A2(n12295), .ZN(n12296) );
  AOI21_X1 U15387 ( .B1(n12295), .B2(n12294), .A(n12296), .ZN(n14693) );
  AOI22_X1 U15388 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15389 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U15390 ( .A1(n12298), .A2(n12297), .ZN(n12320) );
  INV_X1 U15391 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15392 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11916), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12302) );
  AOI21_X1 U15393 ( .B1(n9808), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12305), .ZN(n12301) );
  OAI211_X1 U15394 ( .C1(n12304), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12319) );
  OAI21_X1 U15395 ( .B1(n12307), .B2(n12306), .A(n12305), .ZN(n12312) );
  INV_X1 U15396 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12309) );
  INV_X1 U15397 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12308) );
  OAI22_X1 U15398 ( .A1(n12310), .A2(n12309), .B1(n13773), .B2(n12308), .ZN(
        n12311) );
  AOI211_X1 U15399 ( .C1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n12313), .A(
        n12312), .B(n12311), .ZN(n12317) );
  AOI22_X1 U15400 ( .A1(n9852), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12314), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15401 ( .A1(n9848), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12315) );
  NAND3_X1 U15402 ( .A1(n12317), .A2(n12316), .A3(n12315), .ZN(n12318) );
  OAI21_X1 U15403 ( .B1(n12320), .B2(n12319), .A(n12318), .ZN(n12321) );
  INV_X1 U15404 ( .A(n12321), .ZN(n12322) );
  AOI22_X1 U15405 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12113), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15406 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15407 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15408 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12014), .B1(
        n11954), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12324) );
  NAND4_X1 U15409 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12334) );
  AOI22_X1 U15410 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n12414), .ZN(n12332) );
  AOI22_X1 U15411 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12546), .ZN(n12330) );
  NAND2_X1 U15412 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12329) );
  NAND2_X1 U15413 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12328) );
  AOI22_X1 U15414 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12331) );
  NAND3_X1 U15415 ( .A1(n12332), .A2(n10508), .A3(n12331), .ZN(n12333) );
  NOR2_X1 U15416 ( .A1(n12334), .A2(n12333), .ZN(n12509) );
  MUX2_X1 U15417 ( .A(n20078), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n13837), .Z(n12816) );
  NAND2_X1 U15418 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20086), .ZN(
        n12349) );
  INV_X1 U15419 ( .A(n12349), .ZN(n12348) );
  NAND2_X1 U15420 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20069), .ZN(
        n12344) );
  XNOR2_X1 U15421 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12339) );
  NOR2_X1 U15422 ( .A1(n16412), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12336) );
  AOI21_X1 U15423 ( .B1(n12338), .B2(n12339), .A(n12336), .ZN(n12365) );
  NOR2_X1 U15424 ( .A1(n16427), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12337) );
  AND2_X1 U15425 ( .A1(n12365), .A2(n12337), .ZN(n12361) );
  MUX2_X1 U15426 ( .A(n12509), .B(n12361), .S(n12936), .Z(n12682) );
  INV_X1 U15427 ( .A(n12338), .ZN(n12341) );
  INV_X1 U15428 ( .A(n12339), .ZN(n12340) );
  XNOR2_X1 U15429 ( .A(n12341), .B(n12340), .ZN(n12681) );
  OAI21_X1 U15430 ( .B1(n12682), .B2(n12681), .A(n11817), .ZN(n12360) );
  INV_X1 U15431 ( .A(n12342), .ZN(n12347) );
  INV_X1 U15432 ( .A(n12343), .ZN(n12345) );
  NAND2_X1 U15433 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  INV_X1 U15434 ( .A(n12804), .ZN(n12351) );
  AOI21_X1 U15435 ( .B1(n13801), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12348), .ZN(n12815) );
  XNOR2_X1 U15436 ( .A(n12816), .B(n12349), .ZN(n12390) );
  OAI21_X1 U15437 ( .B1(n13000), .B2(n12815), .A(n12390), .ZN(n12350) );
  OAI21_X1 U15438 ( .B1(n12351), .B2(n13000), .A(n12350), .ZN(n12353) );
  NAND2_X1 U15439 ( .A1(n12816), .A2(n12815), .ZN(n12352) );
  AOI22_X1 U15440 ( .A1(n12353), .A2(n16440), .B1(n12364), .B2(n12352), .ZN(
        n12358) );
  NAND2_X1 U15441 ( .A1(n12354), .A2(n13000), .ZN(n12355) );
  MUX2_X1 U15442 ( .A(n12355), .B(n12936), .S(n12804), .Z(n12356) );
  INV_X1 U15443 ( .A(n12356), .ZN(n12357) );
  NOR2_X1 U15444 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  NAND2_X1 U15445 ( .A1(n12360), .A2(n12359), .ZN(n12372) );
  INV_X1 U15446 ( .A(n12361), .ZN(n12363) );
  INV_X1 U15447 ( .A(n12681), .ZN(n12362) );
  NAND2_X1 U15448 ( .A1(n12363), .A2(n12362), .ZN(n12389) );
  NAND2_X1 U15449 ( .A1(n12389), .A2(n12364), .ZN(n12370) );
  INV_X1 U15450 ( .A(n12365), .ZN(n12367) );
  INV_X1 U15451 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12808) );
  NAND2_X1 U15452 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12808), .ZN(
        n12368) );
  NAND2_X1 U15453 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  MUX2_X1 U15454 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12373), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12918) );
  INV_X1 U15455 ( .A(n12824), .ZN(n12374) );
  NAND2_X1 U15456 ( .A1(n12374), .A2(n14671), .ZN(n12375) );
  INV_X1 U15457 ( .A(n19439), .ZN(n12951) );
  OAI21_X1 U15458 ( .B1(n12376), .B2(n12951), .A(n16442), .ZN(n12384) );
  NAND2_X1 U15459 ( .A1(n12377), .A2(n12604), .ZN(n12378) );
  AND2_X1 U15460 ( .A1(n12403), .A2(n12952), .ZN(n12826) );
  NAND2_X1 U15461 ( .A1(n12378), .A2(n12826), .ZN(n12948) );
  NAND2_X1 U15462 ( .A1(n12385), .A2(n16440), .ZN(n12379) );
  NAND2_X1 U15463 ( .A1(n12379), .A2(n12604), .ZN(n12380) );
  NAND2_X1 U15464 ( .A1(n12380), .A2(n19439), .ZN(n12381) );
  AND4_X1 U15465 ( .A1(n12382), .A2(n12948), .A3(n12956), .A4(n12381), .ZN(
        n12383) );
  AND2_X1 U15466 ( .A1(n12384), .A2(n12383), .ZN(n12923) );
  INV_X1 U15467 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U15468 ( .A1(n16462), .A2(n12952), .ZN(n12388) );
  NAND2_X1 U15469 ( .A1(n16442), .A2(n12388), .ZN(n16433) );
  INV_X1 U15470 ( .A(n12389), .ZN(n12805) );
  AND2_X1 U15471 ( .A1(n12804), .A2(n12390), .ZN(n12391) );
  NAND2_X1 U15472 ( .A1(n12805), .A2(n12391), .ZN(n12392) );
  NAND2_X1 U15473 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19950) );
  AND2_X1 U15474 ( .A1(n14674), .A2(n19950), .ZN(n12802) );
  AOI21_X1 U15475 ( .B1(n16438), .B2(n16431), .A(n12393), .ZN(n12976) );
  NAND2_X1 U15476 ( .A1(n16440), .A2(n11792), .ZN(n12395) );
  NOR2_X1 U15477 ( .A1(n12394), .A2(n12395), .ZN(n12396) );
  NAND2_X1 U15478 ( .A1(n12397), .A2(n12396), .ZN(n12959) );
  NAND2_X1 U15479 ( .A1(n12976), .A2(n12959), .ZN(n12398) );
  NAND2_X1 U15480 ( .A1(n13767), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19956) );
  NOR2_X1 U15481 ( .A1(n12604), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15482 ( .A1(n12399), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12402) );
  AND2_X1 U15483 ( .A1(n12604), .A2(n20079), .ZN(n12400) );
  NAND2_X1 U15484 ( .A1(n12567), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U15485 ( .A1(n12402), .A2(n12401), .ZN(n14843) );
  AOI222_X1 U15486 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n12567), .B1(n12510), 
        .B2(P2_EAX_REG_19__SCAN_IN), .C1(n12599), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U15487 ( .A1(n12399), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15488 ( .A1(n12567), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15489 ( .A1(n12570), .A2(n13476), .ZN(n12405) );
  AOI22_X1 U15490 ( .A1(n12510), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12599), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U15491 ( .A1(n12567), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15492 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12426), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15493 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15494 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15495 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12014), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12410) );
  NAND4_X1 U15496 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n12410), .ZN(
        n12423) );
  AOI22_X1 U15497 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15498 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15499 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12416) );
  AND2_X1 U15500 ( .A1(n12417), .A2(n12416), .ZN(n12420) );
  AOI22_X1 U15501 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15502 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12418) );
  NAND4_X1 U15503 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12422) );
  INV_X1 U15504 ( .A(n12684), .ZN(n13665) );
  AOI22_X1 U15505 ( .A1(n12510), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12453), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12425) );
  NAND2_X1 U15506 ( .A1(n12567), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12424) );
  OAI211_X1 U15507 ( .C1(n13665), .C2(n12577), .A(n12425), .B(n12424), .ZN(
        n13718) );
  AOI22_X1 U15508 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12426), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15509 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15510 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15511 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12014), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U15512 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12443) );
  AOI22_X1 U15513 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15514 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12437) );
  NAND2_X1 U15515 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12436) );
  AND2_X1 U15516 ( .A1(n12437), .A2(n12436), .ZN(n12440) );
  AOI22_X1 U15517 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12439) );
  NAND2_X1 U15518 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12438) );
  NAND4_X1 U15519 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n12438), .ZN(
        n12442) );
  INV_X1 U15520 ( .A(n12843), .ZN(n12447) );
  NAND2_X1 U15521 ( .A1(n12444), .A2(n12453), .ZN(n12487) );
  AND2_X1 U15522 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12445) );
  NOR2_X1 U15523 ( .A1(n12399), .A2(n12445), .ZN(n12446) );
  OAI211_X1 U15524 ( .C1(n12447), .C2(n12577), .A(n12487), .B(n12446), .ZN(
        n13256) );
  NAND2_X1 U15525 ( .A1(n12567), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12452) );
  INV_X1 U15526 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12449) );
  NAND2_X1 U15527 ( .A1(n13442), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12448) );
  OAI211_X1 U15528 ( .C1(n12604), .C2(n12449), .A(n12448), .B(n20079), .ZN(
        n12450) );
  INV_X1 U15529 ( .A(n12450), .ZN(n12451) );
  NAND2_X1 U15530 ( .A1(n12452), .A2(n12451), .ZN(n13257) );
  NAND2_X1 U15531 ( .A1(n13256), .A2(n13257), .ZN(n12471) );
  AOI22_X1 U15532 ( .A1(n12399), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12453), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U15533 ( .A1(n12567), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12454) );
  AND2_X1 U15534 ( .A1(n12455), .A2(n12454), .ZN(n12472) );
  XNOR2_X1 U15535 ( .A(n12471), .B(n12472), .ZN(n12943) );
  NAND2_X1 U15536 ( .A1(n11795), .A2(n12604), .ZN(n12456) );
  MUX2_X1 U15537 ( .A(n12456), .B(n20078), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12470) );
  AOI22_X1 U15538 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15539 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15540 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12113), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15541 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15542 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12468) );
  AOI22_X1 U15543 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n12414), .ZN(n12466) );
  AOI22_X1 U15544 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12546), .ZN(n12462) );
  NAND2_X1 U15545 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12461) );
  AND2_X1 U15546 ( .A1(n12462), .A2(n12461), .ZN(n12465) );
  AOI22_X1 U15547 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U15548 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12463) );
  NAND4_X1 U15549 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12467) );
  NAND2_X1 U15550 ( .A1(n12570), .A2(n12847), .ZN(n12469) );
  NAND2_X1 U15551 ( .A1(n12470), .A2(n12469), .ZN(n12942) );
  NAND2_X1 U15552 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  NAND2_X1 U15553 ( .A1(n12945), .A2(n12473), .ZN(n12491) );
  AOI22_X1 U15554 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12429), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15555 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15556 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12428), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15557 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12014), .B1(
        n11954), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15558 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12485) );
  AOI22_X1 U15559 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15560 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n12414), .ZN(n12482) );
  AOI22_X1 U15561 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12546), .ZN(n12479) );
  NAND2_X1 U15562 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12478) );
  AND2_X1 U15563 ( .A1(n12479), .A2(n12478), .ZN(n12481) );
  NAND2_X1 U15564 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12480) );
  NAND4_X1 U15565 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12484) );
  INV_X1 U15566 ( .A(n12849), .ZN(n13411) );
  NAND2_X1 U15567 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12486) );
  OAI211_X1 U15568 ( .C1(n13411), .C2(n12577), .A(n12487), .B(n12486), .ZN(
        n12490) );
  XNOR2_X1 U15569 ( .A(n12491), .B(n12490), .ZN(n13025) );
  AOI22_X1 U15570 ( .A1(n12510), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12453), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U15571 ( .A1(n12567), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12488) );
  AND2_X1 U15572 ( .A1(n12489), .A2(n12488), .ZN(n13024) );
  INV_X1 U15573 ( .A(n12490), .ZN(n12492) );
  NAND2_X1 U15574 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  INV_X1 U15575 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U15576 ( .A1(n12567), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12599), .ZN(n12508) );
  AOI22_X1 U15577 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15578 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12135), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15579 ( .A1(n12113), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15580 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15581 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12506) );
  AOI22_X1 U15582 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15583 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12546), .ZN(n12500) );
  NAND2_X1 U15584 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12499) );
  AND2_X1 U15585 ( .A1(n12500), .A2(n12499), .ZN(n12503) );
  AOI22_X1 U15586 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15587 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12501) );
  NAND4_X1 U15588 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12505) );
  NAND2_X1 U15589 ( .A1(n12510), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12507) );
  AND2_X1 U15590 ( .A1(n12508), .A2(n9917), .ZN(n13253) );
  INV_X1 U15591 ( .A(n12509), .ZN(n13529) );
  AOI22_X1 U15592 ( .A1(n12567), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n12570), 
        .B2(n13529), .ZN(n12512) );
  AOI22_X1 U15593 ( .A1(n12510), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12599), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U15594 ( .A1(n12512), .A2(n12511), .ZN(n13261) );
  INV_X1 U15595 ( .A(n13719), .ZN(n12513) );
  NAND2_X1 U15596 ( .A1(n13718), .A2(n12513), .ZN(n13721) );
  AOI22_X1 U15597 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12426), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15598 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12428), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15599 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12135), .B1(
        n12113), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15600 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12014), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U15601 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n12525) );
  AOI22_X1 U15602 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15603 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12546), .ZN(n12519) );
  NAND2_X1 U15604 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12518) );
  AND2_X1 U15605 ( .A1(n12519), .A2(n12518), .ZN(n12522) );
  AOI22_X1 U15606 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12494), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15607 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12520) );
  NAND4_X1 U15608 ( .A1(n12523), .A2(n12522), .A3(n12521), .A4(n12520), .ZN(
        n12524) );
  NOR2_X1 U15609 ( .A1(n12525), .A2(n12524), .ZN(n14903) );
  INV_X1 U15610 ( .A(n14903), .ZN(n12526) );
  NAND2_X1 U15611 ( .A1(n12570), .A2(n12526), .ZN(n12527) );
  AOI22_X1 U15612 ( .A1(n12399), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12599), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U15613 ( .A1(n12567), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15614 ( .A1(n12529), .A2(n12528), .ZN(n16374) );
  NAND2_X1 U15615 ( .A1(n16375), .A2(n16374), .ZN(n16373) );
  NAND2_X1 U15616 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12533) );
  NAND2_X1 U15617 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15618 ( .A1(n12429), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15619 ( .A1(n12428), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12530) );
  NAND4_X1 U15620 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12540) );
  NAND2_X1 U15621 ( .A1(n12135), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U15622 ( .A1(n12113), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12537) );
  NAND2_X1 U15623 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U15624 ( .A1(n12014), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12535) );
  NAND4_X1 U15625 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12539) );
  NAND2_X1 U15626 ( .A1(n12434), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12545) );
  NAND2_X1 U15627 ( .A1(n12414), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12544) );
  NAND2_X1 U15628 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12543) );
  NAND2_X1 U15629 ( .A1(n12494), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12542) );
  NAND4_X1 U15630 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        n12551) );
  AOI22_X1 U15631 ( .A1(n12809), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12546), .ZN(n12549) );
  NAND2_X1 U15632 ( .A1(n11954), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U15633 ( .A1(n12435), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12547) );
  NAND3_X1 U15634 ( .A1(n12549), .A2(n12548), .A3(n12547), .ZN(n12550) );
  NAND2_X1 U15635 ( .A1(n12570), .A2(n15087), .ZN(n12554) );
  AOI22_X1 U15636 ( .A1(n12510), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12599), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15637 ( .A1(n12567), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12555) );
  OAI211_X1 U15638 ( .C1(n13103), .C2(n12577), .A(n12556), .B(n12555), .ZN(
        n15507) );
  AOI22_X1 U15639 ( .A1(n12399), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12453), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U15640 ( .A1(n12567), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12559) );
  INV_X1 U15641 ( .A(n13108), .ZN(n12557) );
  NAND2_X1 U15642 ( .A1(n12570), .A2(n12557), .ZN(n12558) );
  INV_X1 U15643 ( .A(n13175), .ZN(n12563) );
  AOI22_X1 U15644 ( .A1(n12399), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U15645 ( .A1(n12567), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12561) );
  OAI211_X1 U15646 ( .C1(n12563), .C2(n12577), .A(n12562), .B(n12561), .ZN(
        n15472) );
  NOR2_X1 U15647 ( .A1(n12577), .A2(n13294), .ZN(n12566) );
  INV_X1 U15648 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n12564) );
  INV_X1 U15649 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16265) );
  OAI22_X1 U15650 ( .A1(n12580), .A2(n12564), .B1(n12581), .B2(n16265), .ZN(
        n12565) );
  AOI211_X1 U15651 ( .C1(n12567), .C2(P2_REIP_REG_11__SCAN_IN), .A(n12566), 
        .B(n12565), .ZN(n16343) );
  AOI22_X1 U15652 ( .A1(n12510), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U15653 ( .A1(n12567), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12568) );
  OAI211_X1 U15654 ( .C1(n13293), .C2(n12577), .A(n12569), .B(n12568), .ZN(
        n15458) );
  AOI22_X1 U15655 ( .A1(n12399), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15656 ( .A1(n12567), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15657 ( .A1(n12570), .A2(n13346), .ZN(n12571) );
  INV_X1 U15658 ( .A(n12574), .ZN(n13470) );
  AOI22_X1 U15659 ( .A1(n12399), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U15660 ( .A1(n12567), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12575) );
  OAI211_X1 U15661 ( .C1(n13470), .C2(n12577), .A(n12576), .B(n12575), .ZN(
        n15437) );
  INV_X1 U15662 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15430) );
  INV_X1 U15663 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13740) );
  INV_X1 U15664 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20009) );
  OAI222_X1 U15665 ( .A1(n12581), .A2(n15430), .B1(n12580), .B2(n13740), .C1(
        n12582), .C2(n20009), .ZN(n13739) );
  AOI22_X1 U15666 ( .A1(n12399), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U15667 ( .A1(n12567), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12578) );
  INV_X1 U15668 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20013) );
  INV_X1 U15669 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16300) );
  INV_X1 U15670 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14859) );
  OAI222_X1 U15671 ( .A1(n12582), .A2(n20013), .B1(n12581), .B2(n16300), .C1(
        n12580), .C2(n14859), .ZN(n14858) );
  NAND2_X1 U15672 ( .A1(n14843), .A2(n14842), .ZN(n14841) );
  AOI22_X1 U15673 ( .A1(n12510), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12584) );
  NAND2_X1 U15674 ( .A1(n12567), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15675 ( .A1(n12510), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15676 ( .A1(n12567), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15677 ( .A1(n12586), .A2(n12585), .ZN(n12793) );
  AOI22_X1 U15678 ( .A1(n12510), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12588) );
  NAND2_X1 U15679 ( .A1(n12567), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U15680 ( .A1(n12588), .A2(n12587), .ZN(n15353) );
  AOI22_X1 U15681 ( .A1(n12510), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U15682 ( .A1(n12567), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15683 ( .A1(n12510), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U15684 ( .A1(n12567), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15685 ( .A1(n12510), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12594) );
  NAND2_X1 U15686 ( .A1(n12567), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12593) );
  NOR2_X2 U15687 ( .A1(n14815), .A2(n14803), .ZN(n14804) );
  AOI22_X1 U15688 ( .A1(n12510), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U15689 ( .A1(n12567), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12595) );
  NAND2_X1 U15690 ( .A1(n12596), .A2(n12595), .ZN(n14795) );
  AOI22_X1 U15691 ( .A1(n12510), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U15692 ( .A1(n12567), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U15693 ( .A1(n12598), .A2(n12597), .ZN(n14787) );
  AOI22_X1 U15694 ( .A1(n12510), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12599), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U15695 ( .A1(n12567), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U15696 ( .A1(n12601), .A2(n12600), .ZN(n14781) );
  AOI22_X1 U15697 ( .A1(n12510), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U15698 ( .A1(n12567), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12602) );
  AND2_X1 U15699 ( .A1(n12603), .A2(n12602), .ZN(n15235) );
  INV_X1 U15700 ( .A(n16119), .ZN(n12621) );
  AND2_X1 U15701 ( .A1(n9853), .A2(n12604), .ZN(n12605) );
  NOR4_X1 U15702 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12609) );
  NOR4_X1 U15703 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12608) );
  NOR4_X1 U15704 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12607) );
  NOR4_X1 U15705 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12606) );
  NAND4_X1 U15706 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12614) );
  NOR4_X1 U15707 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12612) );
  NOR4_X1 U15708 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12611) );
  NOR4_X1 U15709 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12610) );
  NAND4_X1 U15710 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n19983), .ZN(
        n12613) );
  NAND2_X1 U15711 ( .A1(n19267), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12617) );
  INV_X1 U15712 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16575) );
  OR2_X1 U15713 ( .A1(n19267), .A2(n16575), .ZN(n12616) );
  NAND2_X1 U15714 ( .A1(n12617), .A2(n12616), .ZN(n19382) );
  INV_X1 U15715 ( .A(n19382), .ZN(n12619) );
  INV_X1 U15716 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12618) );
  OAI22_X1 U15717 ( .A1(n14868), .A2(n12619), .B1(n19282), .B2(n12618), .ZN(
        n12620) );
  AOI21_X1 U15718 ( .B1(n12621), .B2(n19318), .A(n12620), .ZN(n12624) );
  NOR2_X2 U15719 ( .A1(n13264), .A2(n19267), .ZN(n19262) );
  NOR2_X2 U15720 ( .A1(n13264), .A2(n19268), .ZN(n19264) );
  AOI22_X1 U15721 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19262), .B1(n19264), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n12623) );
  AND2_X1 U15722 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  OAI21_X1 U15723 ( .B1(n14105), .B2(n19269), .A(n12625), .ZN(P2_U2889) );
  INV_X1 U15724 ( .A(n12627), .ZN(n12630) );
  OAI22_X1 U15725 ( .A1(n12630), .A2(n12629), .B1(n12628), .B2(n14128), .ZN(
        n12631) );
  INV_X1 U15726 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21195) );
  AND2_X1 U15727 ( .A1(n20848), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13334) );
  AND2_X1 U15728 ( .A1(n21012), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21008) );
  INV_X1 U15729 ( .A(n15981), .ZN(n13826) );
  INV_X1 U15730 ( .A(n20848), .ZN(n20804) );
  NAND2_X1 U15731 ( .A1(n20804), .A2(n12637), .ZN(n21007) );
  NAND2_X1 U15732 ( .A1(n21007), .A2(n21012), .ZN(n12638) );
  INV_X1 U15733 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21178) );
  NOR2_X1 U15734 ( .A1(n20342), .A2(n21178), .ZN(n14533) );
  NAND2_X1 U15735 ( .A1(n21012), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U15736 ( .A1(n21346), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12639) );
  AND2_X1 U15737 ( .A1(n15819), .A2(n12639), .ZN(n13096) );
  NOR2_X1 U15738 ( .A1(n20302), .A2(n14047), .ZN(n12640) );
  AOI211_X1 U15739 ( .C1(n20291), .C2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14533), .B(n12640), .ZN(n12641) );
  NOR2_X1 U15740 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12643) );
  NOR4_X1 U15741 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12642) );
  NAND4_X1 U15742 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12643), .A4(n12642), .ZN(n12646) );
  INV_X1 U15743 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21104) );
  INV_X1 U15744 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21140) );
  NOR4_X1 U15745 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21104), .A4(n21140), .ZN(n12645) );
  NOR4_X1 U15746 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12644)
         );
  NAND3_X1 U15747 ( .A1(n13577), .A2(n12645), .A3(n12644), .ZN(U214) );
  NOR2_X1 U15748 ( .A1(n19267), .A2(n12646), .ZN(n16551) );
  NAND2_X1 U15749 ( .A1(n16551), .A2(U214), .ZN(U212) );
  NAND2_X1 U15750 ( .A1(n12667), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12665) );
  NAND2_X1 U15751 ( .A1(n12658), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12659) );
  NAND2_X1 U15752 ( .A1(n12653), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12651) );
  NAND2_X1 U15753 ( .A1(n12650), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12647) );
  AOI21_X1 U15754 ( .B1(n15167), .B2(n12647), .A(n12648), .ZN(n15169) );
  INV_X1 U15755 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15242) );
  NAND2_X1 U15756 ( .A1(n12648), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12777) );
  NAND2_X1 U15757 ( .A1(n15138), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15129) );
  INV_X1 U15758 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15076) );
  INV_X1 U15759 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15054) );
  OAI21_X1 U15760 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12650), .A(
        n12647), .ZN(n15180) );
  INV_X1 U15761 ( .A(n15180), .ZN(n19055) );
  AOI21_X1 U15762 ( .B1(n12652), .B2(n12651), .A(n12650), .ZN(n19066) );
  OAI21_X1 U15763 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12653), .A(
        n12651), .ZN(n15202) );
  INV_X1 U15764 ( .A(n15202), .ZN(n19076) );
  OAI21_X1 U15765 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12654), .A(
        n12656), .ZN(n19104) );
  INV_X1 U15766 ( .A(n19104), .ZN(n19098) );
  OAI21_X1 U15767 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12657), .A(
        n9858), .ZN(n16238) );
  INV_X1 U15768 ( .A(n16238), .ZN(n19126) );
  OAI21_X1 U15769 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12658), .A(
        n12660), .ZN(n16256) );
  INV_X1 U15770 ( .A(n16256), .ZN(n19148) );
  OAI21_X1 U15771 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12661), .A(
        n12662), .ZN(n16276) );
  INV_X1 U15772 ( .A(n16276), .ZN(n19168) );
  AOI21_X1 U15773 ( .B1(n19186), .B2(n12663), .A(n12664), .ZN(n19192) );
  AOI21_X1 U15774 ( .B1(n16299), .B2(n12665), .A(n12666), .ZN(n19212) );
  AOI21_X1 U15775 ( .B1(n19424), .B2(n12670), .A(n12667), .ZN(n19410) );
  AOI21_X1 U15776 ( .B1(n19257), .B2(n12668), .A(n12669), .ZN(n13630) );
  AOI22_X1 U15777 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19034), .ZN(n13764) );
  AOI22_X1 U15778 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19257), .B2(n19034), .ZN(
        n13763) );
  NAND2_X1 U15779 ( .A1(n13764), .A2(n13763), .ZN(n13761) );
  OAI21_X1 U15780 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12669), .A(
        n12670), .ZN(n13690) );
  NAND2_X1 U15781 ( .A1(n13689), .A2(n13690), .ZN(n19237) );
  OAI21_X1 U15782 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12667), .A(
        n12665), .ZN(n19223) );
  NAND2_X1 U15783 ( .A1(n19221), .A2(n19223), .ZN(n19210) );
  OAI21_X1 U15784 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12666), .A(
        n12663), .ZN(n19201) );
  NAND2_X1 U15785 ( .A1(n19200), .A2(n19201), .ZN(n19190) );
  INV_X1 U15786 ( .A(n12661), .ZN(n12671) );
  OAI21_X1 U15787 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n12664), .A(
        n12671), .ZN(n19177) );
  NAND2_X1 U15788 ( .A1(n19176), .A2(n19177), .ZN(n19166) );
  AOI21_X1 U15789 ( .B1(n16269), .B2(n12662), .A(n12658), .ZN(n16257) );
  INV_X1 U15790 ( .A(n16257), .ZN(n19157) );
  NAND2_X1 U15791 ( .A1(n19156), .A2(n19157), .ZN(n19146) );
  AOI21_X1 U15792 ( .B1(n16252), .B2(n12660), .A(n12657), .ZN(n16239) );
  INV_X1 U15793 ( .A(n16239), .ZN(n19142) );
  NAND2_X1 U15794 ( .A1(n19133), .A2(n19142), .ZN(n19131) );
  AOI21_X1 U15795 ( .B1(n19109), .B2(n9858), .A(n12654), .ZN(n19112) );
  INV_X1 U15796 ( .A(n19112), .ZN(n19116) );
  NAND2_X1 U15797 ( .A1(n19117), .A2(n19116), .ZN(n19097) );
  NOR2_X1 U15798 ( .A1(n19098), .A2(n19097), .ZN(n19092) );
  NAND2_X1 U15799 ( .A1(n12656), .A2(n12672), .ZN(n12674) );
  INV_X1 U15800 ( .A(n12653), .ZN(n12673) );
  NAND2_X1 U15801 ( .A1(n12674), .A2(n12673), .ZN(n19091) );
  NOR2_X1 U15802 ( .A1(n9835), .A2(n19054), .ZN(n12676) );
  NOR3_X1 U15803 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15853) );
  NAND2_X1 U15804 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15853), .ZN(n19953) );
  AOI211_X1 U15805 ( .C1(n15169), .C2(n12676), .A(n12779), .B(n19953), .ZN(
        n12776) );
  AND2_X1 U15806 ( .A1(n12920), .A2(n16462), .ZN(n12921) );
  AND2_X1 U15807 ( .A1(n12952), .A2(n12992), .ZN(n12830) );
  INV_X1 U15808 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14683) );
  NAND2_X1 U15809 ( .A1(n19950), .A2(n19627), .ZN(n12766) );
  NAND2_X1 U15810 ( .A1(n14683), .A2(n12766), .ZN(n12677) );
  INV_X2 U15811 ( .A(n12914), .ZN(n19405) );
  INV_X1 U15812 ( .A(n19950), .ZN(n19958) );
  INV_X1 U15813 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19959) );
  NAND2_X2 U15814 ( .A1(n20036), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20038) );
  NOR2_X1 U15815 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19036) );
  INV_X1 U15816 ( .A(n19036), .ZN(n19971) );
  NAND3_X1 U15817 ( .A1(n19959), .A2(n20038), .A3(n19971), .ZN(n14670) );
  NAND2_X1 U15818 ( .A1(n19627), .A2(n12978), .ZN(n12771) );
  NAND2_X1 U15819 ( .A1(n19405), .A2(n12771), .ZN(n16104) );
  INV_X1 U15820 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14760) );
  INV_X1 U15821 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20019) );
  NOR2_X1 U15822 ( .A1(n16442), .A2(n16471), .ZN(n12891) );
  NAND2_X1 U15823 ( .A1(n12891), .A2(n12920), .ZN(n13710) );
  NAND2_X1 U15824 ( .A1(n13710), .A2(n12878), .ZN(n19032) );
  NAND2_X1 U15825 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19822), .ZN(n19948) );
  NOR2_X1 U15826 ( .A1(n19956), .A2(n19948), .ZN(n16455) );
  NAND2_X1 U15827 ( .A1(n13836), .A2(n19822), .ZN(n19033) );
  INV_X1 U15828 ( .A(n19033), .ZN(n12799) );
  NOR2_X1 U15829 ( .A1(n16455), .A2(n19412), .ZN(n12678) );
  NAND2_X1 U15830 ( .A1(n19953), .A2(n12678), .ZN(n12679) );
  OAI22_X1 U15831 ( .A1(n19110), .A2(n14760), .B1(n20019), .B2(n19183), .ZN(
        n12775) );
  MUX2_X1 U15832 ( .A(n12849), .B(n12804), .S(n12936), .Z(n12817) );
  MUX2_X1 U15833 ( .A(n12817), .B(n11855), .S(n12683), .Z(n12852) );
  NOR2_X1 U15834 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n12680) );
  MUX2_X1 U15835 ( .A(n12847), .B(n12680), .S(n12683), .Z(n12855) );
  NAND2_X1 U15836 ( .A1(n12852), .A2(n12855), .ZN(n13449) );
  MUX2_X1 U15837 ( .A(n12820), .B(P2_EBX_REG_3__SCAN_IN), .S(n9853), .Z(n13448) );
  INV_X1 U15838 ( .A(n12682), .ZN(n12822) );
  INV_X1 U15839 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13019) );
  MUX2_X1 U15840 ( .A(n12822), .B(n13019), .S(n9853), .Z(n13526) );
  INV_X1 U15841 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12708) );
  MUX2_X1 U15842 ( .A(n12684), .B(n12708), .S(n9853), .Z(n13668) );
  MUX2_X1 U15843 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n14903), .S(n12404), .Z(
        n14910) );
  MUX2_X1 U15844 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n15043), .S(n12404), .Z(
        n14918) );
  NOR2_X1 U15845 ( .A1(n14910), .A2(n14918), .ZN(n12685) );
  INV_X1 U15846 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U15847 ( .A1(n12683), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14913) );
  INV_X1 U15848 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U15849 ( .A1(n13186), .A2(n14933), .ZN(n14944) );
  NAND2_X1 U15850 ( .A1(n15012), .A2(n14944), .ZN(n14932) );
  NAND2_X1 U15851 ( .A1(n12683), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12686) );
  INV_X1 U15852 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12737) );
  NOR2_X1 U15853 ( .A1(n12404), .A2(n12737), .ZN(n14946) );
  INV_X1 U15854 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U15855 ( .A1(n9853), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14966) );
  NOR2_X1 U15856 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n12687) );
  NOR2_X1 U15857 ( .A1(n12404), .A2(n12687), .ZN(n12688) );
  NOR2_X1 U15858 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n12689) );
  INV_X1 U15859 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14952) );
  NOR2_X1 U15860 ( .A1(n12404), .A2(n14760), .ZN(n12690) );
  AND2_X1 U15861 ( .A1(n12691), .A2(n12690), .ZN(n12692) );
  OR2_X1 U15862 ( .A1(n12783), .A2(n12692), .ZN(n14951) );
  NOR2_X1 U15863 ( .A1(n12878), .A2(n12403), .ZN(n12768) );
  AND2_X1 U15864 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12766), .ZN(n12693) );
  OAI22_X1 U15865 ( .A1(n15167), .A2(n19185), .B1(n14951), .B2(n19233), .ZN(
        n12774) );
  NAND2_X1 U15866 ( .A1(n12695), .A2(n12694), .ZN(n12700) );
  INV_X1 U15867 ( .A(n12696), .ZN(n12697) );
  OR2_X1 U15868 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  NAND2_X1 U15869 ( .A1(n12721), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U15870 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12701) );
  AOI21_X1 U15871 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12703), .ZN(n13018) );
  NAND2_X1 U15872 ( .A1(n12721), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U15873 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12706) );
  AOI21_X1 U15874 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12709), .ZN(n13041) );
  INV_X1 U15875 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13058) );
  NAND2_X1 U15876 ( .A1(n12721), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U15877 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12710) );
  AOI21_X1 U15878 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12712), .ZN(n13053) );
  INV_X1 U15879 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U15880 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12715) );
  AOI22_X1 U15881 ( .A1(n14680), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12714) );
  INV_X1 U15882 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15883 ( .A1(n12721), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U15884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12717) );
  AOI21_X1 U15885 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12720), .ZN(n13100) );
  INV_X1 U15886 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U15887 ( .A1(n12721), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15888 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12722) );
  AOI21_X1 U15889 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12725), .ZN(n13109) );
  NAND2_X1 U15890 ( .A1(n14680), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15891 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12726) );
  AOI21_X1 U15892 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12728), .ZN(n13177) );
  NOR2_X2 U15893 ( .A1(n13178), .A2(n13177), .ZN(n13184) );
  NAND2_X1 U15894 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12730) );
  AOI22_X1 U15895 ( .A1(n14680), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12729) );
  INV_X1 U15896 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U15897 ( .A1(n14680), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U15898 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12731) );
  AOI21_X1 U15899 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12734), .ZN(n13297) );
  NAND2_X1 U15900 ( .A1(n14680), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U15901 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12735) );
  AOI21_X1 U15902 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12738), .ZN(n13347) );
  NAND2_X1 U15903 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12740) );
  AOI22_X1 U15904 ( .A1(n14680), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12739) );
  INV_X1 U15905 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U15906 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12743) );
  AOI22_X1 U15907 ( .A1(n14680), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12742) );
  INV_X1 U15908 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14973) );
  NAND2_X1 U15909 ( .A1(n14680), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15910 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12745) );
  AOI21_X1 U15911 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12747), .ZN(n13626) );
  INV_X1 U15912 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n14959) );
  NAND2_X1 U15913 ( .A1(n14680), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U15914 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12748) );
  AOI21_X1 U15915 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12750), .ZN(n13729) );
  INV_X1 U15916 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14955) );
  NAND2_X1 U15917 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12752) );
  AOI22_X1 U15918 ( .A1(n14680), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12751) );
  INV_X1 U15919 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15920 ( .A1(n14680), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U15921 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12753) );
  AOI21_X1 U15922 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12756), .ZN(n14775) );
  INV_X1 U15923 ( .A(n12757), .ZN(n14773) );
  NAND2_X1 U15924 ( .A1(n14680), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U15925 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12758) );
  AOI21_X1 U15926 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12760), .ZN(n14767) );
  NAND2_X1 U15927 ( .A1(n14680), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12762) );
  NAND2_X1 U15928 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12761) );
  AOI21_X1 U15929 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12763), .ZN(n12764) );
  AND2_X1 U15930 ( .A1(n14765), .A2(n12764), .ZN(n12765) );
  NOR2_X2 U15931 ( .A1(n14765), .A2(n12764), .ZN(n12790) );
  OR2_X1 U15932 ( .A1(n12765), .A2(n12790), .ZN(n15385) );
  INV_X1 U15933 ( .A(n12766), .ZN(n12767) );
  AND2_X1 U15934 ( .A1(n14841), .A2(n12769), .ZN(n12770) );
  NOR2_X1 U15935 ( .A1(n12794), .A2(n12770), .ZN(n14837) );
  INV_X1 U15936 ( .A(n14837), .ZN(n15381) );
  INV_X1 U15937 ( .A(n12771), .ZN(n12772) );
  AND2_X1 U15938 ( .A1(n12826), .A2(n12772), .ZN(n16461) );
  OAI22_X1 U15939 ( .A1(n15385), .A2(n19230), .B1(n15381), .B2(n19232), .ZN(
        n12773) );
  OR4_X1 U15940 ( .A1(n12776), .A2(n12775), .A3(n12774), .A4(n12773), .ZN(
        P2_U2834) );
  OAI21_X1 U15941 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12648), .A(
        n12778), .ZN(n16219) );
  INV_X1 U15942 ( .A(n16219), .ZN(n12781) );
  NOR2_X1 U15943 ( .A1(n9835), .A2(n12779), .ZN(n12780) );
  NOR2_X1 U15944 ( .A1(n12781), .A2(n12780), .ZN(n16112) );
  AOI211_X1 U15945 ( .C1(n12781), .C2(n12780), .A(n16112), .B(n19953), .ZN(
        n12798) );
  INV_X1 U15946 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14754) );
  INV_X1 U15947 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20021) );
  OAI22_X1 U15948 ( .A1(n19110), .A2(n14754), .B1(n20021), .B2(n19183), .ZN(
        n12797) );
  INV_X1 U15949 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12786) );
  INV_X1 U15950 ( .A(n12782), .ZN(n12785) );
  NAND2_X1 U15951 ( .A1(n12683), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12784) );
  OAI21_X1 U15952 ( .B1(n12785), .B2(n12784), .A(n15000), .ZN(n14996) );
  OAI22_X1 U15953 ( .A1(n12786), .A2(n19185), .B1(n14996), .B2(n19233), .ZN(
        n12796) );
  NAND2_X1 U15954 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12788) );
  AOI22_X1 U15955 ( .A1(n14680), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12787) );
  OR2_X1 U15956 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  AND2_X1 U15957 ( .A1(n12791), .A2(n14740), .ZN(n16216) );
  INV_X1 U15958 ( .A(n16216), .ZN(n14755) );
  INV_X1 U15959 ( .A(n15354), .ZN(n12792) );
  OAI21_X1 U15960 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(n15373) );
  OAI22_X1 U15961 ( .A1(n14755), .A2(n19230), .B1(n15373), .B2(n19232), .ZN(
        n12795) );
  INV_X1 U15962 ( .A(n13710), .ZN(n19258) );
  INV_X1 U15963 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20102) );
  OAI211_X1 U15964 ( .C1(n19258), .C2(n20102), .A(n19033), .B(n12878), .ZN(
        P2_U2814) );
  INV_X1 U15965 ( .A(n14674), .ZN(n12954) );
  INV_X1 U15966 ( .A(n19032), .ZN(n12801) );
  OAI21_X1 U15967 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n12799), .A(n12801), 
        .ZN(n12800) );
  OAI21_X1 U15968 ( .B1(n12954), .B2(n12801), .A(n12800), .ZN(P2_U3612) );
  INV_X1 U15969 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12982) );
  NOR2_X1 U15970 ( .A1(n12802), .A2(n12978), .ZN(n12803) );
  NAND3_X1 U15971 ( .A1(n16433), .A2(n12920), .A3(n12803), .ZN(n16446) );
  AND2_X1 U15972 ( .A1(n16446), .A2(n12992), .ZN(n20089) );
  NAND3_X1 U15973 ( .A1(n12805), .A2(n12815), .A3(n12804), .ZN(n12806) );
  NAND3_X1 U15974 ( .A1(n12920), .A2(n13767), .A3(n12806), .ZN(n12812) );
  NAND2_X1 U15975 ( .A1(n12808), .A2(n12807), .ZN(n16439) );
  OAI21_X1 U15976 ( .B1(n12809), .B2(n16439), .A(n12982), .ZN(n12810) );
  AND2_X1 U15977 ( .A1(n12810), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20083) );
  INV_X1 U15978 ( .A(n20083), .ZN(n12811) );
  AND2_X1 U15979 ( .A1(n12812), .A2(n12811), .ZN(n20092) );
  INV_X1 U15980 ( .A(n12813), .ZN(n12814) );
  NAND2_X1 U15981 ( .A1(n12814), .A2(n13000), .ZN(n12829) );
  MUX2_X1 U15982 ( .A(n12843), .B(n12815), .S(n12936), .Z(n12836) );
  NAND2_X1 U15983 ( .A1(n12836), .A2(n12816), .ZN(n12819) );
  INV_X1 U15984 ( .A(n12817), .ZN(n12818) );
  NAND2_X1 U15985 ( .A1(n12819), .A2(n12818), .ZN(n12823) );
  INV_X1 U15986 ( .A(n12820), .ZN(n12821) );
  NAND3_X1 U15987 ( .A1(n12823), .A2(n12822), .A3(n12821), .ZN(n12825) );
  AND2_X1 U15988 ( .A1(n12825), .A2(n12824), .ZN(n20090) );
  INV_X1 U15989 ( .A(n12826), .ZN(n12827) );
  NOR2_X1 U15990 ( .A1(n12813), .A2(n12827), .ZN(n20093) );
  NAND2_X1 U15991 ( .A1(n20090), .A2(n20093), .ZN(n12828) );
  OAI21_X1 U15992 ( .B1(n12982), .B2(n20089), .A(n12835), .ZN(P2_U2819) );
  OR2_X1 U15993 ( .A1(n20057), .A2(n13836), .ZN(n20070) );
  NAND2_X1 U15994 ( .A1(n20070), .A2(n19034), .ZN(n12831) );
  AND2_X1 U15995 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20071) );
  INV_X1 U15996 ( .A(n12835), .ZN(n12832) );
  AND2_X1 U15997 ( .A1(n12403), .A2(n12843), .ZN(n12848) );
  INV_X1 U15998 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12833) );
  AND2_X1 U15999 ( .A1(n12848), .A2(n12833), .ZN(n12834) );
  NOR2_X1 U16000 ( .A1(n12848), .A2(n12833), .ZN(n12845) );
  OR2_X1 U16001 ( .A1(n12834), .A2(n12845), .ZN(n16403) );
  INV_X1 U16002 ( .A(n16403), .ZN(n12838) );
  AND2_X1 U16003 ( .A1(n19412), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16406) );
  MUX2_X1 U16004 ( .A(n12836), .B(P2_EBX_REG_0__SCAN_IN), .S(n9853), .Z(n13706) );
  NAND2_X1 U16005 ( .A1(n13706), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12874) );
  OAI21_X1 U16006 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13706), .A(
        n12874), .ZN(n16401) );
  NOR2_X1 U16007 ( .A1(n19415), .A2(n16401), .ZN(n12837) );
  AOI211_X1 U16008 ( .C1(n16294), .C2(n12838), .A(n16406), .B(n12837), .ZN(
        n12842) );
  NAND2_X1 U16009 ( .A1(n19627), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U16010 ( .A1(n10105), .A2(n12840), .ZN(n12862) );
  OAI21_X1 U16011 ( .B1(n16270), .B2(n12862), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U16012 ( .C1(n16284), .C2(n10090), .A(n12842), .B(n12841), .ZN(
        P2_U3014) );
  INV_X1 U16013 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13537) );
  XOR2_X1 U16014 ( .A(n12843), .B(n12847), .Z(n12844) );
  AND2_X1 U16015 ( .A1(n12845), .A2(n12844), .ZN(n12846) );
  INV_X1 U16016 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13765) );
  XNOR2_X1 U16017 ( .A(n12845), .B(n12844), .ZN(n12870) );
  NOR2_X1 U16018 ( .A1(n13765), .A2(n12870), .ZN(n12869) );
  NOR2_X1 U16019 ( .A1(n12846), .A2(n12869), .ZN(n13456) );
  XNOR2_X1 U16020 ( .A(n13537), .B(n13456), .ZN(n12850) );
  NAND2_X1 U16021 ( .A1(n12848), .A2(n12847), .ZN(n13412) );
  XNOR2_X1 U16022 ( .A(n13412), .B(n12849), .ZN(n12851) );
  NAND2_X1 U16023 ( .A1(n12850), .A2(n12851), .ZN(n13030) );
  NOR2_X1 U16024 ( .A1(n12851), .A2(n12850), .ZN(n13457) );
  INV_X1 U16025 ( .A(n13457), .ZN(n13029) );
  NAND3_X1 U16026 ( .A1(n13030), .A2(n16294), .A3(n13029), .ZN(n12866) );
  INV_X1 U16027 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19982) );
  NOR2_X1 U16028 ( .A1(n19982), .A2(n16334), .ZN(n13027) );
  AOI21_X1 U16029 ( .B1(n16270), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13027), .ZN(n12865) );
  OAI21_X1 U16030 ( .B1(n12852), .B2(n12855), .A(n13449), .ZN(n13631) );
  XNOR2_X1 U16031 ( .A(n13631), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12861) );
  INV_X1 U16032 ( .A(n12861), .ZN(n12859) );
  NAND2_X1 U16033 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12853) );
  NOR2_X1 U16034 ( .A1(n12404), .A2(n12853), .ZN(n12854) );
  NOR2_X1 U16035 ( .A1(n12855), .A2(n12854), .ZN(n19246) );
  NAND2_X1 U16036 ( .A1(n19246), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12857) );
  INV_X1 U16037 ( .A(n19246), .ZN(n12856) );
  AOI22_X1 U16038 ( .A1(n12874), .A2(n12857), .B1(n13765), .B2(n12856), .ZN(
        n12860) );
  INV_X1 U16039 ( .A(n12860), .ZN(n12858) );
  NAND2_X1 U16040 ( .A1(n12859), .A2(n12858), .ZN(n13022) );
  NAND2_X1 U16041 ( .A1(n12861), .A2(n12860), .ZN(n13454) );
  NAND3_X1 U16042 ( .A1(n13022), .A2(n16293), .A3(n13454), .ZN(n12864) );
  NAND2_X1 U16043 ( .A1(n19411), .A2(n13630), .ZN(n12863) );
  NAND4_X1 U16044 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  AOI21_X1 U16045 ( .B1(n13765), .B2(n12870), .A(n12869), .ZN(n12946) );
  NAND2_X1 U16046 ( .A1(n16294), .A2(n12946), .ZN(n12871) );
  NAND2_X1 U16047 ( .A1(n19412), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12938) );
  OAI211_X1 U16048 ( .C1(n19423), .C2(n19257), .A(n12871), .B(n12938), .ZN(
        n12872) );
  INV_X1 U16049 ( .A(n12872), .ZN(n12876) );
  XNOR2_X1 U16050 ( .A(n19246), .B(n13765), .ZN(n12873) );
  XNOR2_X1 U16051 ( .A(n12874), .B(n12873), .ZN(n12972) );
  AOI22_X1 U16052 ( .A1(n19411), .A2(n19257), .B1(n16293), .B2(n12972), .ZN(
        n12875) );
  OAI211_X1 U16053 ( .C1(n13402), .C2(n16284), .A(n12876), .B(n12875), .ZN(
        P2_U3013) );
  INV_X1 U16054 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U16055 ( .A1(n13000), .A2(n19950), .ZN(n12877) );
  NAND2_X1 U16056 ( .A1(n12911), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U16057 ( .A1(n19267), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12880) );
  INV_X1 U16058 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16587) );
  OR2_X1 U16059 ( .A1(n19267), .A2(n16587), .ZN(n12879) );
  NAND2_X1 U16060 ( .A1(n12880), .A2(n12879), .ZN(n19286) );
  NAND2_X1 U16061 ( .A1(n19383), .A2(n19286), .ZN(n12882) );
  OAI211_X1 U16062 ( .C1(n12914), .C2(n14823), .A(n12881), .B(n12882), .ZN(
        P2_U2960) );
  INV_X1 U16063 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19350) );
  NAND2_X1 U16064 ( .A1(n12911), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12883) );
  OAI211_X1 U16065 ( .C1(n19350), .C2(n12914), .A(n12883), .B(n12882), .ZN(
        P2_U2975) );
  INV_X1 U16066 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U16067 ( .A1(n12911), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U16068 ( .A1(n19267), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12885) );
  INV_X1 U16069 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16581) );
  OR2_X1 U16070 ( .A1(n19267), .A2(n16581), .ZN(n12884) );
  NAND2_X1 U16071 ( .A1(n12885), .A2(n12884), .ZN(n19278) );
  NAND2_X1 U16072 ( .A1(n19383), .A2(n19278), .ZN(n12912) );
  OAI211_X1 U16073 ( .C1(n12904), .C2(n12914), .A(n12886), .B(n12912), .ZN(
        P2_U2963) );
  INV_X1 U16074 ( .A(n12887), .ZN(n15786) );
  OAI22_X1 U16075 ( .A1(n12909), .A2(n10153), .B1(n12888), .B2(n15789), .ZN(
        n15779) );
  NOR2_X1 U16076 ( .A1(n15779), .A2(n15829), .ZN(n12890) );
  INV_X1 U16077 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21102) );
  NAND3_X1 U16078 ( .A1(n16093), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20625), 
        .ZN(n12889) );
  OAI21_X1 U16079 ( .B1(n12890), .B2(n21102), .A(n12889), .ZN(P1_U2803) );
  INV_X1 U16080 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14817) );
  NAND2_X1 U16081 ( .A1(n16438), .A2(n13000), .ZN(n12977) );
  INV_X1 U16082 ( .A(n12891), .ZN(n12892) );
  OAI21_X1 U16083 ( .B1(n12977), .B2(n12892), .A(n12914), .ZN(n12893) );
  INV_X1 U16084 ( .A(n14670), .ZN(n19967) );
  NAND2_X1 U16085 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13203) );
  CLKBUF_X1 U16086 ( .A(n19335), .Z(n19366) );
  INV_X2 U16087 ( .A(n19333), .ZN(n19363) );
  AOI22_X1 U16088 ( .A1(n19366), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12894) );
  OAI21_X1 U16089 ( .B1(n14817), .B2(n19327), .A(n12894), .ZN(P2_U2926) );
  INV_X1 U16090 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14829) );
  AOI22_X1 U16091 ( .A1(n19335), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12895) );
  OAI21_X1 U16092 ( .B1(n14829), .B2(n19327), .A(n12895), .ZN(P2_U2929) );
  AOI22_X1 U16093 ( .A1(n19335), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U16094 ( .B1(n14823), .B2(n19327), .A(n12896), .ZN(P2_U2927) );
  INV_X1 U16095 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14844) );
  AOI22_X1 U16096 ( .A1(n19335), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12897) );
  OAI21_X1 U16097 ( .B1(n14844), .B2(n19327), .A(n12897), .ZN(P2_U2931) );
  AOI22_X1 U16098 ( .A1(n19335), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12898) );
  OAI21_X1 U16099 ( .B1(n14859), .B2(n19327), .A(n12898), .ZN(P2_U2933) );
  INV_X1 U16100 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U16101 ( .A1(n19366), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12899) );
  OAI21_X1 U16102 ( .B1(n14790), .B2(n19327), .A(n12899), .ZN(P2_U2923) );
  INV_X1 U16103 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16104 ( .A1(n19335), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12900) );
  OAI21_X1 U16105 ( .B1(n12901), .B2(n19327), .A(n12900), .ZN(P2_U2928) );
  INV_X1 U16106 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14851) );
  AOI22_X1 U16107 ( .A1(n19335), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12902) );
  OAI21_X1 U16108 ( .B1(n14851), .B2(n19327), .A(n12902), .ZN(P2_U2932) );
  AOI22_X1 U16109 ( .A1(n19366), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12903) );
  OAI21_X1 U16110 ( .B1(n12904), .B2(n19327), .A(n12903), .ZN(P2_U2924) );
  INV_X1 U16111 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U16112 ( .A1(n19366), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12905) );
  OAI21_X1 U16113 ( .B1(n14807), .B2(n19327), .A(n12905), .ZN(P2_U2925) );
  INV_X1 U16114 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U16115 ( .A1(n19335), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12906) );
  OAI21_X1 U16116 ( .B1(n14867), .B2(n19327), .A(n12906), .ZN(P2_U2934) );
  INV_X1 U16117 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16118 ( .A1(n19335), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12907) );
  OAI21_X1 U16119 ( .B1(n14835), .B2(n19327), .A(n12907), .ZN(P2_U2930) );
  AOI22_X1 U16120 ( .A1(n19335), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12908) );
  OAI21_X1 U16121 ( .B1(n13740), .B2(n19327), .A(n12908), .ZN(P2_U2935) );
  NAND2_X1 U16122 ( .A1(n12909), .A2(n20107), .ZN(n12915) );
  AND2_X1 U16123 ( .A1(n20848), .A2(n16101), .ZN(n13811) );
  AOI211_X1 U16124 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12915), .A(n13811), 
        .B(n10165), .ZN(n12910) );
  INV_X1 U16125 ( .A(n12910), .ZN(P1_U2801) );
  NAND2_X1 U16126 ( .A1(n19406), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12913) );
  OAI211_X1 U16127 ( .C1(n12564), .C2(n12914), .A(n12913), .B(n12912), .ZN(
        P2_U2978) );
  OAI21_X1 U16128 ( .B1(n13811), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n10163), 
        .ZN(n12916) );
  OAI21_X1 U16129 ( .B1(n12917), .B2(n10163), .A(n12916), .ZN(P1_U3487) );
  NAND2_X1 U16130 ( .A1(n12951), .A2(n12978), .ZN(n12929) );
  AOI21_X1 U16131 ( .B1(n12918), .B2(n16440), .A(n19452), .ZN(n12919) );
  NAND2_X1 U16132 ( .A1(n12977), .A2(n12919), .ZN(n12928) );
  INV_X1 U16133 ( .A(n12920), .ZN(n16432) );
  OAI211_X1 U16134 ( .C1(n16462), .C2(n12403), .A(n19950), .B(n12394), .ZN(
        n12924) );
  NAND2_X1 U16135 ( .A1(n12921), .A2(n12978), .ZN(n12922) );
  AND2_X1 U16136 ( .A1(n12923), .A2(n12922), .ZN(n12975) );
  OAI21_X1 U16137 ( .B1(n16432), .B2(n12924), .A(n12975), .ZN(n12926) );
  NOR2_X1 U16138 ( .A1(n12926), .A2(n12925), .ZN(n12927) );
  OAI211_X1 U16139 ( .C1(n12977), .C2(n12929), .A(n12928), .B(n12927), .ZN(
        n12930) );
  INV_X1 U16140 ( .A(n12931), .ZN(n12932) );
  OR2_X1 U16141 ( .A1(n16433), .A2(n12932), .ZN(n15515) );
  NAND2_X1 U16142 ( .A1(n15515), .A2(n12403), .ZN(n12934) );
  NAND2_X1 U16143 ( .A1(n12934), .A2(n12933), .ZN(n12935) );
  NOR2_X1 U16144 ( .A1(n12813), .A2(n12936), .ZN(n20091) );
  NAND2_X2 U16145 ( .A1(n12967), .A2(n20091), .ZN(n16402) );
  INV_X1 U16146 ( .A(n16402), .ZN(n16379) );
  INV_X1 U16147 ( .A(n12967), .ZN(n12937) );
  INV_X1 U16148 ( .A(n19412), .ZN(n16334) );
  NAND2_X1 U16149 ( .A1(n12937), .A2(n16334), .ZN(n16398) );
  OAI21_X1 U16150 ( .B1(n16398), .B2(n13765), .A(n12938), .ZN(n12971) );
  AND2_X1 U16151 ( .A1(n16433), .A2(n13000), .ZN(n12940) );
  OR2_X1 U16152 ( .A1(n16434), .A2(n12940), .ZN(n12941) );
  NAND2_X1 U16153 ( .A1(n12943), .A2(n12942), .ZN(n12944) );
  NAND2_X1 U16154 ( .A1(n12945), .A2(n12944), .ZN(n20076) );
  AOI22_X1 U16155 ( .A1(n16393), .A2(n12946), .B1(n16399), .B2(n20076), .ZN(
        n12969) );
  NAND2_X1 U16156 ( .A1(n12967), .A2(n16431), .ZN(n15414) );
  NAND2_X1 U16157 ( .A1(n12947), .A2(n13000), .ZN(n13793) );
  NAND2_X1 U16158 ( .A1(n13793), .A2(n12948), .ZN(n12950) );
  NAND2_X1 U16159 ( .A1(n12950), .A2(n12949), .ZN(n12964) );
  NAND2_X1 U16160 ( .A1(n12956), .A2(n19452), .ZN(n12953) );
  AOI22_X1 U16161 ( .A1(n12954), .A2(n12953), .B1(n12952), .B2(n12951), .ZN(
        n12961) );
  NOR2_X1 U16162 ( .A1(n12957), .A2(n12956), .ZN(n12958) );
  NAND2_X1 U16163 ( .A1(n12955), .A2(n12958), .ZN(n12960) );
  AND4_X1 U16164 ( .A1(n12962), .A2(n12961), .A3(n12960), .A4(n12959), .ZN(
        n12963) );
  NAND2_X1 U16165 ( .A1(n12964), .A2(n12963), .ZN(n15524) );
  OR2_X1 U16166 ( .A1(n15524), .A2(n12965), .ZN(n12966) );
  NAND2_X1 U16167 ( .A1(n12967), .A2(n12966), .ZN(n15418) );
  NAND2_X1 U16168 ( .A1(n15414), .A2(n15418), .ZN(n15419) );
  NAND2_X1 U16169 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13536) );
  OAI211_X1 U16170 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15419), .B(n13536), .ZN(n12968) );
  NAND2_X1 U16171 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  AOI211_X1 U16172 ( .C1(n16379), .C2(n12972), .A(n12971), .B(n12970), .ZN(
        n12973) );
  OAI21_X1 U16173 ( .B1(n13402), .B2(n16365), .A(n12973), .ZN(P2_U3045) );
  INV_X1 U16174 ( .A(n16438), .ZN(n12974) );
  NAND2_X1 U16175 ( .A1(n12974), .A2(n16434), .ZN(n12991) );
  AND3_X1 U16176 ( .A1(n12976), .A2(n12991), .A3(n12975), .ZN(n12981) );
  INV_X1 U16177 ( .A(n12977), .ZN(n12979) );
  INV_X1 U16178 ( .A(n16442), .ZN(n12984) );
  NAND3_X1 U16179 ( .A1(n12979), .A2(n12984), .A3(n12978), .ZN(n12980) );
  NOR2_X1 U16180 ( .A1(n19034), .A2(n13203), .ZN(n16457) );
  INV_X1 U16181 ( .A(n16457), .ZN(n16473) );
  OAI22_X1 U16182 ( .A1(n16430), .A2(n16471), .B1(n12982), .B2(n16473), .ZN(
        n12983) );
  NAND4_X1 U16183 ( .A1(n12984), .A2(n12403), .A3(n13836), .A4(n16439), .ZN(
        n12986) );
  NAND2_X1 U16184 ( .A1(n15527), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12985) );
  OAI21_X1 U16185 ( .B1(n15527), .B2(n12986), .A(n12985), .ZN(P2_U3595) );
  NAND2_X1 U16186 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  INV_X1 U16187 ( .A(n12965), .ZN(n13770) );
  NAND2_X1 U16188 ( .A1(n12991), .A2(n13770), .ZN(n12993) );
  OR2_X2 U16189 ( .A1(n14749), .A2(n11744), .ZN(n14779) );
  NOR2_X1 U16190 ( .A1(n14769), .A2(n11855), .ZN(n12994) );
  OAI21_X1 U16191 ( .B1(n20065), .B2(n14779), .A(n9960), .ZN(P2_U2885) );
  MUX2_X1 U16192 ( .A(n11823), .B(n13402), .S(n14769), .Z(n12999) );
  OAI21_X1 U16193 ( .B1(n13276), .B2(n14779), .A(n12999), .ZN(P2_U2886) );
  NAND2_X1 U16194 ( .A1(n13000), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13001) );
  NAND4_X1 U16195 ( .A1(n11868), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13001), 
        .A4(n20079), .ZN(n13002) );
  MUX2_X1 U16196 ( .A(n10090), .B(n11841), .S(n14749), .Z(n13004) );
  OAI21_X1 U16197 ( .B1(n20081), .B2(n14779), .A(n13004), .ZN(P2_U2887) );
  NOR2_X1 U16198 ( .A1(n13401), .A2(n14776), .ZN(n13009) );
  AOI21_X1 U16199 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n14776), .A(n13009), .ZN(
        n13010) );
  OAI21_X1 U16200 ( .B1(n15526), .B2(n14779), .A(n13010), .ZN(P2_U2884) );
  INV_X1 U16201 ( .A(n13011), .ZN(n13012) );
  NAND2_X1 U16202 ( .A1(n13013), .A2(n13012), .ZN(n13015) );
  OAI21_X1 U16203 ( .B1(n13016), .B2(n13015), .A(n13014), .ZN(n19236) );
  AOI21_X1 U16204 ( .B1(n13018), .B2(n13017), .A(n9952), .ZN(n19419) );
  NOR2_X1 U16205 ( .A1(n14769), .A2(n13019), .ZN(n13020) );
  AOI21_X1 U16206 ( .B1(n19419), .B2(n14769), .A(n13020), .ZN(n13021) );
  OAI21_X1 U16207 ( .B1(n19236), .B2(n14779), .A(n13021), .ZN(P2_U2883) );
  INV_X1 U16208 ( .A(n13536), .ZN(n13038) );
  INV_X1 U16209 ( .A(n15418), .ZN(n13539) );
  NAND2_X1 U16210 ( .A1(n13539), .A2(n13537), .ZN(n13543) );
  OAI21_X1 U16211 ( .B1(n15414), .B2(n13537), .A(n13543), .ZN(n13037) );
  NAND2_X1 U16212 ( .A1(n13022), .A2(n13454), .ZN(n13033) );
  OAI21_X1 U16213 ( .B1(n13025), .B2(n13024), .A(n13023), .ZN(n20067) );
  NAND2_X1 U16214 ( .A1(n13537), .A2(n13536), .ZN(n15248) );
  NOR2_X1 U16215 ( .A1(n15414), .A2(n15248), .ZN(n13026) );
  OR2_X1 U16216 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  AOI21_X1 U16217 ( .B1(n16399), .B2(n20067), .A(n13028), .ZN(n13032) );
  NAND3_X1 U16218 ( .A1(n13030), .A2(n16393), .A3(n13029), .ZN(n13031) );
  OAI211_X1 U16219 ( .C1(n16402), .C2(n13033), .A(n13032), .B(n13031), .ZN(
        n13036) );
  OR2_X1 U16220 ( .A1(n15418), .A2(n13038), .ZN(n13034) );
  AND2_X1 U16221 ( .A1(n13034), .A2(n16398), .ZN(n13544) );
  NOR2_X1 U16222 ( .A1(n13544), .A2(n13537), .ZN(n13035) );
  AOI211_X1 U16223 ( .C1(n13038), .C2(n13037), .A(n13036), .B(n13035), .ZN(
        n13039) );
  OAI21_X1 U16224 ( .B1(n13040), .B2(n16365), .A(n13039), .ZN(P2_U3044) );
  XOR2_X1 U16225 ( .A(n13014), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13043)
         );
  OAI21_X1 U16226 ( .B1(n9952), .B2(n10355), .A(n13054), .ZN(n19229) );
  MUX2_X1 U16227 ( .A(n12708), .B(n19229), .S(n14769), .Z(n13042) );
  OAI21_X1 U16228 ( .B1(n13043), .B2(n14779), .A(n13042), .ZN(P2_U2882) );
  XNOR2_X1 U16229 ( .A(n13044), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U16230 ( .B1(n9957), .B2(n13045), .A(n13101), .ZN(n19206) );
  MUX2_X1 U16231 ( .A(n12716), .B(n19206), .S(n14769), .Z(n13046) );
  OAI21_X1 U16232 ( .B1(n13047), .B2(n14779), .A(n13046), .ZN(P2_U2880) );
  INV_X1 U16233 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13077) );
  NAND3_X1 U16234 ( .A1(n15800), .A2(n20107), .A3(n15789), .ZN(n13048) );
  OAI21_X1 U16235 ( .B1(n13060), .B2(n13496), .A(n13048), .ZN(n13049) );
  NAND2_X1 U16236 ( .A1(n20212), .A2(n13599), .ZN(n13130) );
  NAND2_X1 U16237 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16102) );
  NOR2_X1 U16238 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16102), .ZN(n13128) );
  NOR2_X4 U16239 ( .A1(n20212), .A2(n20241), .ZN(n20224) );
  AOI22_X1 U16240 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20224), .B1(n20241), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13050) );
  OAI21_X1 U16241 ( .B1(n13077), .B2(n13130), .A(n13050), .ZN(P1_U2906) );
  NOR2_X1 U16242 ( .A1(n13014), .A2(n12103), .ZN(n13052) );
  INV_X1 U16243 ( .A(n13044), .ZN(n13051) );
  OAI211_X1 U16244 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13052), .A(
        n13051), .B(n14746), .ZN(n13057) );
  AND2_X1 U16245 ( .A1(n13054), .A2(n13053), .ZN(n13055) );
  OR2_X1 U16246 ( .A1(n13055), .A2(n9957), .ZN(n19216) );
  INV_X1 U16247 ( .A(n19216), .ZN(n16380) );
  NAND2_X1 U16248 ( .A1(n16380), .A2(n14769), .ZN(n13056) );
  OAI211_X1 U16249 ( .C1(n14769), .C2(n13058), .A(n13057), .B(n13056), .ZN(
        P2_U2881) );
  OAI21_X4 U16250 ( .B1(n21010), .B2(n16097), .A(n10165), .ZN(n20286) );
  INV_X1 U16251 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20228) );
  MUX2_X1 U16252 ( .A(BUF1_REG_8__SCAN_IN), .B(DATAI_8_), .S(n14369), .Z(
        n14332) );
  NAND2_X1 U16253 ( .A1(n20283), .A2(n14332), .ZN(n13062) );
  NAND2_X1 U16254 ( .A1(n20286), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13061) );
  OAI211_X1 U16255 ( .C1(n20245), .C2(n20228), .A(n13062), .B(n13061), .ZN(
        P1_U2960) );
  NAND2_X1 U16256 ( .A1(n20286), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13063) );
  OAI211_X1 U16257 ( .C1(n20245), .C2(n11268), .A(n13063), .B(n13062), .ZN(
        P1_U2945) );
  AOI22_X1 U16258 ( .A1(n20241), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13064) );
  OAI21_X1 U16259 ( .B1(n10660), .B2(n13130), .A(n13064), .ZN(P1_U2907) );
  INV_X1 U16260 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16261 ( .A1(n13128), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13065) );
  OAI21_X1 U16262 ( .B1(n13066), .B2(n13130), .A(n13065), .ZN(P1_U2913) );
  AOI22_X1 U16263 ( .A1(n13128), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13067) );
  OAI21_X1 U16264 ( .B1(n11268), .B2(n13130), .A(n13067), .ZN(P1_U2912) );
  AOI22_X1 U16265 ( .A1(n13128), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13068) );
  OAI21_X1 U16266 ( .B1(n11279), .B2(n13130), .A(n13068), .ZN(P1_U2911) );
  AOI22_X1 U16267 ( .A1(n20241), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13069) );
  OAI21_X1 U16268 ( .B1(n11294), .B2(n13130), .A(n13069), .ZN(P1_U2909) );
  INV_X1 U16269 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U16270 ( .A1(n20241), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13070) );
  OAI21_X1 U16271 ( .B1(n21053), .B2(n13130), .A(n13070), .ZN(P1_U2908) );
  MUX2_X1 U16272 ( .A(BUF1_REG_12__SCAN_IN), .B(DATAI_12_), .S(n14369), .Z(
        n20276) );
  AOI22_X1 U16273 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20276), .ZN(n13071) );
  OAI21_X1 U16274 ( .B1(n20245), .B2(n21053), .A(n13071), .ZN(P1_U2949) );
  MUX2_X1 U16275 ( .A(BUF1_REG_13__SCAN_IN), .B(DATAI_13_), .S(n14369), .Z(
        n20279) );
  AOI22_X1 U16276 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20279), .ZN(n13072) );
  OAI21_X1 U16277 ( .B1(n20245), .B2(n10660), .A(n13072), .ZN(P1_U2950) );
  MUX2_X1 U16278 ( .A(BUF1_REG_9__SCAN_IN), .B(DATAI_9_), .S(n14369), .Z(
        n20267) );
  AOI22_X1 U16279 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20267), .ZN(n13073) );
  OAI21_X1 U16280 ( .B1(n20245), .B2(n11279), .A(n13073), .ZN(P1_U2946) );
  MUX2_X1 U16281 ( .A(BUF1_REG_11__SCAN_IN), .B(DATAI_11_), .S(n14369), .Z(
        n20273) );
  AOI22_X1 U16282 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20273), .ZN(n13074) );
  OAI21_X1 U16283 ( .B1(n20245), .B2(n11294), .A(n13074), .ZN(P1_U2948) );
  INV_X1 U16284 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21171) );
  MUX2_X1 U16285 ( .A(BUF1_REG_10__SCAN_IN), .B(DATAI_10_), .S(n14369), .Z(
        n20270) );
  AOI22_X1 U16286 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20270), .ZN(n13075) );
  OAI21_X1 U16287 ( .B1(n20245), .B2(n21171), .A(n13075), .ZN(P1_U2947) );
  MUX2_X1 U16288 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n14369), .Z(
        n20282) );
  AOI22_X1 U16289 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20286), .B1(n20283), 
        .B2(n20282), .ZN(n13076) );
  OAI21_X1 U16290 ( .B1(n20245), .B2(n13077), .A(n13076), .ZN(P1_U2951) );
  INV_X1 U16291 ( .A(n13078), .ZN(n13081) );
  OAI21_X1 U16292 ( .B1(n13081), .B2(n13080), .A(n13079), .ZN(n14264) );
  NAND2_X1 U16293 ( .A1(n10743), .A2(n10695), .ZN(n13082) );
  INV_X1 U16294 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20244) );
  INV_X1 U16295 ( .A(n13082), .ZN(n13083) );
  OR2_X1 U16296 ( .A1(n14369), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13085) );
  INV_X1 U16297 ( .A(DATAI_0_), .ZN(n21405) );
  NAND2_X1 U16298 ( .A1(n14369), .A2(n21405), .ZN(n13084) );
  NAND2_X1 U16299 ( .A1(n13085), .A2(n13084), .ZN(n20255) );
  OAI222_X1 U16300 ( .A1(n14264), .A2(n14382), .B1(n14380), .B2(n20244), .C1(
        n14379), .C2(n20255), .ZN(P1_U2904) );
  OAI21_X1 U16301 ( .B1(n13087), .B2(n13086), .A(n13220), .ZN(n13512) );
  INV_X1 U16302 ( .A(n13088), .ZN(n13090) );
  NAND2_X1 U16303 ( .A1(n13090), .A2(n13089), .ZN(n13092) );
  AND2_X1 U16304 ( .A1(n13092), .A2(n13091), .ZN(n20343) );
  OAI222_X1 U16305 ( .A1(n14318), .A2(n13512), .B1(n20211), .B2(n10416), .C1(
        n14312), .C2(n20343), .ZN(P1_U2871) );
  OAI21_X1 U16306 ( .B1(n13094), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13093), .ZN(n13198) );
  INV_X1 U16307 ( .A(n13198), .ZN(n13098) );
  AND2_X1 U16308 ( .A1(n20317), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13195) );
  INV_X1 U16309 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13095) );
  AOI21_X1 U16310 ( .B1(n13821), .B2(n13096), .A(n13095), .ZN(n13097) );
  AOI211_X1 U16311 ( .C1(n13098), .C2(n20298), .A(n13195), .B(n13097), .ZN(
        n13099) );
  OAI21_X1 U16312 ( .B1(n13826), .B2(n14264), .A(n13099), .ZN(P1_U2999) );
  NAND2_X1 U16313 ( .A1(n13101), .A2(n13100), .ZN(n13102) );
  INV_X1 U16314 ( .A(n19193), .ZN(n13107) );
  OAI211_X1 U16315 ( .C1(n10513), .C2(n11927), .A(n14746), .B(n13104), .ZN(
        n13106) );
  NAND2_X1 U16316 ( .A1(n14749), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13105) );
  OAI211_X1 U16317 ( .C1(n13107), .C2(n14749), .A(n13106), .B(n13105), .ZN(
        P2_U2879) );
  XNOR2_X1 U16318 ( .A(n13104), .B(n13108), .ZN(n13112) );
  NAND2_X1 U16319 ( .A1(n9885), .A2(n13109), .ZN(n13110) );
  NAND2_X1 U16320 ( .A1(n13178), .A2(n13110), .ZN(n19182) );
  MUX2_X1 U16321 ( .A(n19182), .B(n12724), .S(n14749), .Z(n13111) );
  OAI21_X1 U16322 ( .B1(n13112), .B2(n14779), .A(n13111), .ZN(P2_U2878) );
  INV_X1 U16323 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20240) );
  INV_X1 U16324 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13113) );
  OR2_X1 U16325 ( .A1(n14369), .A2(n13113), .ZN(n13115) );
  NAND2_X1 U16326 ( .A1(n14369), .A2(DATAI_1_), .ZN(n13114) );
  OAI222_X1 U16327 ( .A1(n14382), .A2(n13512), .B1(n14380), .B2(n20240), .C1(
        n14379), .C2(n20357), .ZN(P1_U2903) );
  INV_X1 U16328 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16329 ( .A1(n20241), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16330 ( .B1(n13117), .B2(n13130), .A(n13116), .ZN(P1_U2920) );
  INV_X1 U16331 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16332 ( .A1(n13128), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13118) );
  OAI21_X1 U16333 ( .B1(n13119), .B2(n13130), .A(n13118), .ZN(P1_U2914) );
  AOI22_X1 U16334 ( .A1(n13128), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13120) );
  OAI21_X1 U16335 ( .B1(n21171), .B2(n13130), .A(n13120), .ZN(P1_U2910) );
  INV_X1 U16336 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16337 ( .A1(n13128), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16338 ( .B1(n13122), .B2(n13130), .A(n13121), .ZN(P1_U2917) );
  INV_X1 U16339 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16340 ( .A1(n13128), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13123) );
  OAI21_X1 U16341 ( .B1(n13124), .B2(n13130), .A(n13123), .ZN(P1_U2918) );
  INV_X1 U16342 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16343 ( .A1(n13128), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13125) );
  OAI21_X1 U16344 ( .B1(n13126), .B2(n13130), .A(n13125), .ZN(P1_U2919) );
  INV_X1 U16345 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U16346 ( .A1(n13128), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13127) );
  OAI21_X1 U16347 ( .B1(n21079), .B2(n13130), .A(n13127), .ZN(P1_U2916) );
  INV_X1 U16348 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16349 ( .A1(n13128), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13129) );
  OAI21_X1 U16350 ( .B1(n13131), .B2(n13130), .A(n13129), .ZN(P1_U2915) );
  NOR2_X1 U16351 ( .A1(n13132), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20341) );
  NOR2_X1 U16352 ( .A1(n20341), .A2(n20108), .ZN(n13135) );
  AOI22_X1 U16353 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13133) );
  OAI21_X1 U16354 ( .B1(n20302), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13133), .ZN(n13134) );
  AOI21_X1 U16355 ( .B1(n13135), .B2(n20346), .A(n13134), .ZN(n13136) );
  OAI21_X1 U16356 ( .B1(n13826), .B2(n13512), .A(n13136), .ZN(P1_U2998) );
  INV_X1 U16357 ( .A(n13138), .ZN(n13140) );
  NAND2_X1 U16358 ( .A1(n13140), .A2(n13139), .ZN(n13141) );
  NOR2_X1 U16359 ( .A1(n13155), .A2(n13141), .ZN(n13143) );
  AND3_X1 U16360 ( .A1(n11657), .A2(n13143), .A3(n13142), .ZN(n15798) );
  OR2_X1 U16361 ( .A1(n20720), .A2(n15798), .ZN(n13152) );
  NAND2_X1 U16362 ( .A1(n15800), .A2(n10521), .ZN(n14658) );
  NAND2_X1 U16363 ( .A1(n15800), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13144) );
  MUX2_X1 U16364 ( .A(n14658), .B(n13144), .S(n13320), .Z(n13150) );
  AND2_X1 U16365 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  NAND2_X1 U16366 ( .A1(n13148), .A2(n13147), .ZN(n13312) );
  NAND3_X1 U16367 ( .A1(n10751), .A2(n20355), .A3(n14656), .ZN(n13310) );
  XNOR2_X1 U16368 ( .A(n13305), .B(n13320), .ZN(n13153) );
  MUX2_X1 U16369 ( .A(n13312), .B(n13310), .S(n13153), .Z(n13149) );
  AND2_X1 U16370 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  NAND2_X1 U16371 ( .A1(n13152), .A2(n13151), .ZN(n13318) );
  AOI22_X1 U16372 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20350), .B2(n11616), .ZN(
        n14666) );
  NOR2_X1 U16373 ( .A1(n16101), .A2(n20324), .ZN(n20989) );
  AOI222_X1 U16374 ( .A1(n13318), .A2(n16093), .B1(n14666), .B2(n20989), .C1(
        n13153), .C2(n15825), .ZN(n13163) );
  INV_X1 U16375 ( .A(n13154), .ZN(n15778) );
  OAI211_X1 U16376 ( .C1(n15800), .C2(n13155), .A(n15778), .B(n15789), .ZN(
        n13156) );
  INV_X1 U16377 ( .A(n13156), .ZN(n13161) );
  AOI22_X1 U16378 ( .A1(n15788), .A2(n15783), .B1(n13157), .B2(n15776), .ZN(
        n13158) );
  NAND2_X1 U16379 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  INV_X1 U16380 ( .A(n16102), .ZN(n13329) );
  NAND2_X1 U16381 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13329), .ZN(n13330) );
  INV_X1 U16382 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21213) );
  OAI22_X1 U16383 ( .A1(n13327), .A2(n15829), .B1(n13330), .B2(n21213), .ZN(
        n16092) );
  AOI21_X1 U16384 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21012), .A(n16092), 
        .ZN(n20992) );
  MUX2_X1 U16385 ( .A(n13163), .B(n13320), .S(n20992), .Z(n13164) );
  INV_X1 U16386 ( .A(n13164), .ZN(P1_U3472) );
  OR2_X1 U16387 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13166) );
  NAND2_X1 U16388 ( .A1(n13167), .A2(n13166), .ZN(n14259) );
  INV_X1 U16389 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n21106) );
  OAI222_X1 U16390 ( .A1(n14259), .A2(n14312), .B1(n21106), .B2(n20211), .C1(
        n14264), .C2(n14318), .ZN(P1_U2872) );
  OAI21_X1 U16391 ( .B1(n13170), .B2(n13169), .A(n13168), .ZN(n13272) );
  OAI21_X1 U16392 ( .B1(n13224), .B2(n13171), .A(n13360), .ZN(n13172) );
  INV_X1 U16393 ( .A(n13172), .ZN(n20315) );
  AOI22_X1 U16394 ( .A1(n20315), .A2(n20206), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14316), .ZN(n13173) );
  OAI21_X1 U16395 ( .B1(n13272), .B2(n14318), .A(n13173), .ZN(P1_U2869) );
  OAI211_X1 U16396 ( .C1(n13176), .C2(n13175), .A(n13174), .B(n14746), .ZN(
        n13181) );
  AND2_X1 U16397 ( .A1(n13178), .A2(n13177), .ZN(n13179) );
  OR2_X1 U16398 ( .A1(n13179), .A2(n13184), .ZN(n15474) );
  NAND2_X1 U16399 ( .A1(n19170), .A2(n14769), .ZN(n13180) );
  OAI211_X1 U16400 ( .C1(n14769), .C2(n13182), .A(n13181), .B(n13180), .ZN(
        P2_U2877) );
  XNOR2_X1 U16401 ( .A(n13174), .B(n13294), .ZN(n13188) );
  OR2_X1 U16402 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  NAND2_X1 U16403 ( .A1(n13298), .A2(n13185), .ZN(n19162) );
  MUX2_X1 U16404 ( .A(n19162), .B(n13186), .S(n14776), .Z(n13187) );
  OAI21_X1 U16405 ( .B1(n13188), .B2(n14779), .A(n13187), .ZN(P2_U2876) );
  INV_X1 U16406 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20236) );
  INV_X1 U16407 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13189) );
  OR2_X1 U16408 ( .A1(n14369), .A2(n13189), .ZN(n13191) );
  NAND2_X1 U16409 ( .A1(n14369), .A2(DATAI_3_), .ZN(n13190) );
  AND2_X1 U16410 ( .A1(n13191), .A2(n13190), .ZN(n20260) );
  OAI222_X1 U16411 ( .A1(n14382), .A2(n13272), .B1(n14380), .B2(n20236), .C1(
        n14379), .C2(n20260), .ZN(P1_U2901) );
  INV_X1 U16412 ( .A(n14259), .ZN(n13196) );
  AOI21_X1 U16413 ( .B1(n13561), .B2(n20324), .A(n20325), .ZN(n20349) );
  INV_X1 U16414 ( .A(n14608), .ZN(n13192) );
  NOR3_X1 U16415 ( .A1(n13561), .A2(n13192), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13193) );
  AOI21_X1 U16416 ( .B1(n20349), .B2(n14614), .A(n13193), .ZN(n13194) );
  AOI211_X1 U16417 ( .C1(n20316), .C2(n13196), .A(n13195), .B(n13194), .ZN(
        n13197) );
  OAI21_X1 U16418 ( .B1(n13198), .B2(n20340), .A(n13197), .ZN(P1_U3031) );
  NAND2_X1 U16419 ( .A1(n15526), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19660) );
  OAI21_X1 U16420 ( .B1(n19660), .B2(n19789), .A(n20057), .ZN(n13212) );
  NAND3_X1 U16421 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20062), .A3(
        n20078), .ZN(n19577) );
  INV_X1 U16422 ( .A(n19577), .ZN(n13199) );
  OR2_X1 U16423 ( .A1(n13212), .A2(n13199), .ZN(n13209) );
  INV_X1 U16424 ( .A(n13277), .ZN(n13201) );
  NAND2_X1 U16425 ( .A1(n13201), .A2(n13200), .ZN(n13228) );
  INV_X1 U16426 ( .A(n13228), .ZN(n13202) );
  OR2_X1 U16427 ( .A1(n13387), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13207) );
  NOR2_X1 U16428 ( .A1(n20086), .A2(n19577), .ZN(n19629) );
  NOR2_X1 U16429 ( .A1(n20057), .A2(n19629), .ZN(n13206) );
  AOI21_X1 U16430 ( .B1(n19822), .B2(n13767), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n14672) );
  NAND2_X1 U16431 ( .A1(n14672), .A2(n13203), .ZN(n13204) );
  AOI21_X1 U16432 ( .B1(n13207), .B2(n13206), .A(n19826), .ZN(n13208) );
  NAND2_X1 U16433 ( .A1(n13209), .A2(n13208), .ZN(n19620) );
  INV_X1 U16434 ( .A(n19620), .ZN(n19608) );
  INV_X1 U16435 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U16436 ( .A1(n19268), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19267), .ZN(n19386) );
  OAI21_X1 U16437 ( .B1(n14881), .B2(n19629), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13211) );
  OAI21_X1 U16438 ( .B1(n13212), .B2(n19577), .A(n13211), .ZN(n19619) );
  INV_X1 U16439 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16559) );
  INV_X1 U16440 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18375) );
  OAI22_X2 U16441 ( .A1(n16559), .A2(n19468), .B1(n18375), .B2(n19466), .ZN(
        n19832) );
  AOI22_X1 U16442 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19464), .ZN(n19835) );
  INV_X1 U16443 ( .A(n19835), .ZN(n19857) );
  INV_X1 U16444 ( .A(n20081), .ZN(n19322) );
  NOR2_X2 U16445 ( .A1(n16440), .A2(n19470), .ZN(n19856) );
  AOI22_X1 U16446 ( .A1(n19857), .A2(n19649), .B1(n19856), .B2(n19629), .ZN(
        n13214) );
  OAI21_X1 U16447 ( .B1(n19871), .B2(n19611), .A(n13214), .ZN(n13215) );
  AOI21_X1 U16448 ( .B1(n13210), .B2(n19619), .A(n13215), .ZN(n13216) );
  OAI21_X1 U16449 ( .B1(n19608), .B2(n13217), .A(n13216), .ZN(P2_U3088) );
  INV_X1 U16450 ( .A(n13218), .ZN(n13219) );
  AOI21_X1 U16451 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n14069) );
  INV_X1 U16452 ( .A(n14318), .ZN(n20207) );
  AND2_X1 U16453 ( .A1(n13223), .A2(n13222), .ZN(n13225) );
  OR2_X1 U16454 ( .A1(n13225), .A2(n13224), .ZN(n20329) );
  OAI22_X1 U16455 ( .A1(n20329), .A2(n14312), .B1(n21243), .B2(n20211), .ZN(
        n13226) );
  AOI21_X1 U16456 ( .B1(n14069), .B2(n20207), .A(n13226), .ZN(n13227) );
  INV_X1 U16457 ( .A(n13227), .ZN(P1_U2870) );
  NAND2_X1 U16458 ( .A1(n20069), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19758) );
  NOR2_X1 U16459 ( .A1(n19479), .A2(n19758), .ZN(n19727) );
  AOI21_X1 U16460 ( .B1(n13434), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13230) );
  NOR2_X1 U16461 ( .A1(n15526), .A2(n19627), .ZN(n19829) );
  AOI21_X1 U16462 ( .B1(n19829), .B2(n19477), .A(n19861), .ZN(n13232) );
  OR2_X1 U16463 ( .A1(n19758), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19684) );
  NAND2_X1 U16464 ( .A1(n13232), .A2(n19684), .ZN(n13229) );
  OAI211_X1 U16465 ( .C1(n19727), .C2(n13230), .A(n13229), .B(n19863), .ZN(
        n19730) );
  INV_X1 U16466 ( .A(n19730), .ZN(n13242) );
  INV_X1 U16467 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16468 ( .A1(n19268), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19267), .ZN(n19388) );
  INV_X1 U16469 ( .A(n13232), .ZN(n13234) );
  INV_X1 U16470 ( .A(n13434), .ZN(n14876) );
  OAI21_X1 U16471 ( .B1(n14876), .B2(n19727), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13233) );
  OAI21_X1 U16472 ( .B1(n13234), .B2(n19684), .A(n13233), .ZN(n19729) );
  INV_X1 U16473 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20354) );
  INV_X1 U16474 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18378) );
  OAI22_X2 U16475 ( .A1(n20354), .A2(n19468), .B1(n18378), .B2(n19466), .ZN(
        n19900) );
  AOI22_X1 U16476 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19464), .ZN(n19903) );
  INV_X1 U16477 ( .A(n19903), .ZN(n19798) );
  NOR2_X2 U16478 ( .A1(n12403), .A2(n19470), .ZN(n19899) );
  AOI22_X1 U16479 ( .A1(n19798), .A2(n19751), .B1(n19899), .B2(n19727), .ZN(
        n13235) );
  OAI21_X1 U16480 ( .B1(n19801), .B2(n19724), .A(n13235), .ZN(n13236) );
  AOI21_X1 U16481 ( .B1(n13231), .B2(n19729), .A(n13236), .ZN(n13237) );
  OAI21_X1 U16482 ( .B1(n13242), .B2(n13376), .A(n13237), .ZN(P2_U3121) );
  INV_X1 U16483 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U16484 ( .A1(n19857), .A2(n19751), .B1(n19727), .B2(n19856), .ZN(
        n13238) );
  OAI21_X1 U16485 ( .B1(n19871), .B2(n19724), .A(n13238), .ZN(n13239) );
  AOI21_X1 U16486 ( .B1(n13210), .B2(n19729), .A(n13239), .ZN(n13240) );
  OAI21_X1 U16487 ( .B1(n13242), .B2(n13241), .A(n13240), .ZN(P2_U3120) );
  INV_X1 U16488 ( .A(n14069), .ZN(n13245) );
  INV_X1 U16489 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20238) );
  OR2_X1 U16490 ( .A1(n14369), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13244) );
  INV_X1 U16491 ( .A(DATAI_2_), .ZN(n21142) );
  NAND2_X1 U16492 ( .A1(n14369), .A2(n21142), .ZN(n13243) );
  NAND2_X1 U16493 ( .A1(n13244), .A2(n13243), .ZN(n20258) );
  OAI222_X1 U16494 ( .A1(n13245), .A2(n14382), .B1(n14380), .B2(n20238), .C1(
        n14379), .C2(n20258), .ZN(P1_U2902) );
  OAI21_X1 U16495 ( .B1(n13248), .B2(n13247), .A(n13246), .ZN(n20328) );
  AOI22_X1 U16496 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16497 ( .B1(n20302), .B2(n14071), .A(n13249), .ZN(n13250) );
  AOI21_X1 U16498 ( .B1(n14069), .B2(n15981), .A(n13250), .ZN(n13251) );
  OAI21_X1 U16499 ( .B1(n20108), .B2(n20328), .A(n13251), .ZN(P1_U2997) );
  NAND2_X1 U16500 ( .A1(n13253), .A2(n13252), .ZN(n13255) );
  INV_X1 U16501 ( .A(n13260), .ZN(n13254) );
  NAND2_X1 U16502 ( .A1(n13255), .A2(n13254), .ZN(n13693) );
  INV_X1 U16503 ( .A(n13693), .ZN(n20058) );
  XNOR2_X1 U16504 ( .A(n20059), .B(n13693), .ZN(n19302) );
  INV_X1 U16505 ( .A(n20065), .ZN(n13259) );
  XNOR2_X1 U16506 ( .A(n20065), .B(n20067), .ZN(n19308) );
  XNOR2_X1 U16507 ( .A(n13276), .B(n20076), .ZN(n19313) );
  OR2_X1 U16508 ( .A1(n13257), .A2(n13256), .ZN(n13258) );
  NAND2_X1 U16509 ( .A1(n12471), .A2(n13258), .ZN(n13709) );
  INV_X1 U16510 ( .A(n13709), .ZN(n19321) );
  NAND2_X1 U16511 ( .A1(n19322), .A2(n19321), .ZN(n19320) );
  NAND2_X1 U16512 ( .A1(n19313), .A2(n19320), .ZN(n19312) );
  OAI21_X1 U16513 ( .B1(n20076), .B2(n20072), .A(n19312), .ZN(n19307) );
  NAND2_X1 U16514 ( .A1(n19308), .A2(n19307), .ZN(n19306) );
  OAI21_X1 U16515 ( .B1(n13259), .B2(n20067), .A(n19306), .ZN(n19301) );
  NAND2_X1 U16516 ( .A1(n19302), .A2(n19301), .ZN(n19300) );
  OAI21_X1 U16517 ( .B1(n20059), .B2(n20058), .A(n19300), .ZN(n13262) );
  OAI21_X1 U16518 ( .B1(n13261), .B2(n13260), .A(n13719), .ZN(n19231) );
  NAND2_X1 U16519 ( .A1(n13262), .A2(n19231), .ZN(n19297) );
  XOR2_X1 U16520 ( .A(n19236), .B(n19297), .Z(n13268) );
  INV_X1 U16521 ( .A(n19231), .ZN(n13263) );
  AOI22_X1 U16522 ( .A1(n19318), .A2(n13263), .B1(n19317), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13267) );
  NAND2_X1 U16523 ( .A1(n14868), .A2(n13264), .ZN(n19285) );
  AOI22_X1 U16524 ( .A1(n19268), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19267), .ZN(n19453) );
  INV_X1 U16525 ( .A(n19453), .ZN(n13265) );
  NAND2_X1 U16526 ( .A1(n19285), .A2(n13265), .ZN(n13266) );
  OAI211_X1 U16527 ( .C1(n13268), .C2(n19269), .A(n13267), .B(n13266), .ZN(
        P2_U2915) );
  OAI21_X1 U16528 ( .B1(n13271), .B2(n13270), .A(n13269), .ZN(n20313) );
  INV_X1 U16529 ( .A(n13272), .ZN(n20198) );
  AOI22_X1 U16530 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13273) );
  OAI21_X1 U16531 ( .B1(n20302), .B2(n20189), .A(n13273), .ZN(n13274) );
  AOI21_X1 U16532 ( .B1(n20198), .B2(n15981), .A(n13274), .ZN(n13275) );
  OAI21_X1 U16533 ( .B1(n20108), .B2(n20313), .A(n13275), .ZN(P1_U2996) );
  NOR2_X1 U16534 ( .A1(n20062), .A2(n19855), .ZN(n13284) );
  AOI21_X1 U16535 ( .B1(n19829), .B2(n19655), .A(n13284), .ZN(n13282) );
  INV_X1 U16536 ( .A(n19427), .ZN(n19938) );
  NAND2_X1 U16537 ( .A1(n13200), .A2(n13277), .ZN(n13373) );
  INV_X1 U16538 ( .A(n13373), .ZN(n13278) );
  NAND2_X1 U16539 ( .A1(n13374), .A2(n13278), .ZN(n13367) );
  INV_X1 U16540 ( .A(n13367), .ZN(n13279) );
  NAND2_X1 U16541 ( .A1(n19427), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13280) );
  OAI211_X1 U16542 ( .C1(n19938), .C2(n20079), .A(n13283), .B(n19863), .ZN(
        n13281) );
  NOR2_X1 U16543 ( .A1(n13282), .A2(n13281), .ZN(n19936) );
  INV_X1 U16544 ( .A(n13283), .ZN(n13286) );
  AOI21_X1 U16545 ( .B1(n20079), .B2(n13284), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13285) );
  NOR2_X1 U16546 ( .A1(n13286), .A2(n13285), .ZN(n19939) );
  INV_X1 U16547 ( .A(n19856), .ZN(n13289) );
  AOI22_X1 U16548 ( .A1(n19931), .A2(n19832), .B1(n19942), .B2(n19857), .ZN(
        n13288) );
  OAI21_X1 U16549 ( .B1(n13289), .B2(n19427), .A(n13288), .ZN(n13290) );
  AOI21_X1 U16550 ( .B1(n19939), .B2(n13210), .A(n13290), .ZN(n13291) );
  OAI21_X1 U16551 ( .B1(n19936), .B2(n13292), .A(n13291), .ZN(P2_U3168) );
  OAI21_X1 U16552 ( .B1(n13174), .B2(n13294), .A(n13293), .ZN(n13296) );
  NAND3_X1 U16553 ( .A1(n13296), .A2(n14746), .A3(n13295), .ZN(n13301) );
  NAND2_X1 U16554 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U16555 ( .A1(n19150), .A2(n14769), .ZN(n13300) );
  OAI211_X1 U16556 ( .C1(n14769), .C2(n12733), .A(n13301), .B(n13300), .ZN(
        P2_U2875) );
  NOR2_X1 U16557 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n13327), .ZN(n13324) );
  INV_X1 U16558 ( .A(n15798), .ZN(n13317) );
  INV_X1 U16559 ( .A(n13303), .ZN(n13307) );
  NAND2_X1 U16560 ( .A1(n13307), .A2(n13302), .ZN(n13314) );
  MUX2_X1 U16561 ( .A(n13303), .B(n10519), .S(n13305), .Z(n13304) );
  INV_X1 U16562 ( .A(n13305), .ZN(n14661) );
  NAND2_X1 U16563 ( .A1(n14661), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13306) );
  NAND2_X1 U16564 ( .A1(n13307), .A2(n13306), .ZN(n13309) );
  NOR2_X1 U16565 ( .A1(n13309), .A2(n13308), .ZN(n14668) );
  OAI22_X1 U16566 ( .A1(n13312), .A2(n13311), .B1(n13310), .B2(n14668), .ZN(
        n13313) );
  AOI21_X1 U16567 ( .B1(n15800), .B2(n13314), .A(n13313), .ZN(n13315) );
  OAI21_X1 U16568 ( .B1(n14658), .B2(n10519), .A(n13315), .ZN(n13316) );
  AOI21_X1 U16569 ( .B1(n20594), .B2(n13317), .A(n13316), .ZN(n15793) );
  NAND2_X1 U16570 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21213), .ZN(n13321) );
  NAND3_X1 U16571 ( .A1(n15793), .A2(n13321), .A3(n15795), .ZN(n13323) );
  MUX2_X1 U16572 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13318), .S(
        n15795), .Z(n13319) );
  OAI22_X1 U16573 ( .A1(n15808), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13321), 
        .B2(n13320), .ZN(n13322) );
  OAI211_X1 U16574 ( .C1(n13324), .C2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13323), .B(n13322), .ZN(n15811) );
  INV_X1 U16575 ( .A(n20477), .ZN(n20719) );
  OR2_X1 U16576 ( .A1(n13325), .A2(n20719), .ZN(n13326) );
  XNOR2_X1 U16577 ( .A(n13326), .B(n16096), .ZN(n20173) );
  NOR2_X1 U16578 ( .A1(n20173), .A2(n11657), .ZN(n16094) );
  MUX2_X1 U16579 ( .A(n21213), .B(n13327), .S(n16101), .Z(n13328) );
  AOI22_X1 U16580 ( .A1(n16094), .A2(n16101), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13328), .ZN(n15812) );
  OAI21_X1 U16581 ( .B1(n15811), .B2(n14655), .A(n15812), .ZN(n13338) );
  NOR2_X1 U16582 ( .A1(n13338), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13331) );
  NAND2_X1 U16583 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20985), .ZN(n14651) );
  INV_X1 U16584 ( .A(n14651), .ZN(n14645) );
  INV_X1 U16585 ( .A(n13332), .ZN(n13333) );
  OAI21_X1 U16586 ( .B1(n13333), .B2(n21346), .A(n20848), .ZN(n20443) );
  NAND2_X1 U16587 ( .A1(n13332), .A2(n13334), .ZN(n20856) );
  OAI21_X1 U16588 ( .B1(n14645), .B2(n20720), .A(n13335), .ZN(n13336) );
  NAND2_X1 U16589 ( .A1(n20352), .A2(n13336), .ZN(n13337) );
  OAI21_X1 U16590 ( .B1(n20352), .B2(n11313), .A(n13337), .ZN(P1_U3476) );
  NOR2_X1 U16591 ( .A1(n13338), .A2(n16102), .ZN(n15827) );
  INV_X1 U16592 ( .A(n10883), .ZN(n15799) );
  OAI22_X1 U16593 ( .A1(n13339), .A2(n20804), .B1(n15799), .B2(n14645), .ZN(
        n13340) );
  OAI21_X1 U16594 ( .B1(n15827), .B2(n13340), .A(n20352), .ZN(n13341) );
  OAI21_X1 U16595 ( .B1(n20352), .B2(n20766), .A(n13341), .ZN(P1_U3478) );
  INV_X1 U16596 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13342) );
  OR2_X1 U16597 ( .A1(n14369), .A2(n13342), .ZN(n13344) );
  NAND2_X1 U16598 ( .A1(n14369), .A2(DATAI_4_), .ZN(n13343) );
  AND2_X1 U16599 ( .A1(n13344), .A2(n13343), .ZN(n20262) );
  XOR2_X1 U16600 ( .A(n13168), .B(n13345), .Z(n20297) );
  INV_X1 U16601 ( .A(n20297), .ZN(n13362) );
  INV_X1 U16602 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20234) );
  OAI222_X1 U16603 ( .A1(n14379), .A2(n20262), .B1(n14382), .B2(n13362), .C1(
        n20234), .C2(n14380), .ZN(P1_U2900) );
  INV_X1 U16604 ( .A(n13346), .ZN(n13471) );
  XNOR2_X1 U16605 ( .A(n13295), .B(n13471), .ZN(n13351) );
  AND2_X1 U16606 ( .A1(n13348), .A2(n13347), .ZN(n13349) );
  OR2_X1 U16607 ( .A1(n13349), .A2(n13467), .ZN(n16248) );
  MUX2_X1 U16608 ( .A(n16248), .B(n12737), .S(n14749), .Z(n13350) );
  OAI21_X1 U16609 ( .B1(n13351), .B2(n14779), .A(n13350), .ZN(P2_U2874) );
  OR2_X1 U16610 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  AND2_X1 U16611 ( .A1(n13352), .A2(n13355), .ZN(n20208) );
  INV_X1 U16612 ( .A(n20208), .ZN(n13358) );
  OR2_X1 U16613 ( .A1(n14369), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13357) );
  INV_X1 U16614 ( .A(DATAI_5_), .ZN(n21129) );
  NAND2_X1 U16615 ( .A1(n14369), .A2(n21129), .ZN(n13356) );
  NAND2_X1 U16616 ( .A1(n13357), .A2(n13356), .ZN(n20367) );
  OAI222_X1 U16617 ( .A1(n13358), .A2(n14382), .B1(n14380), .B2(n10962), .C1(
        n14379), .C2(n20367), .ZN(P1_U2899) );
  NAND2_X1 U16618 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  NAND2_X1 U16619 ( .A1(n16084), .A2(n13361), .ZN(n20306) );
  INV_X1 U16620 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21157) );
  OAI222_X1 U16621 ( .A1(n20306), .A2(n14312), .B1(n20211), .B2(n21157), .C1(
        n14318), .C2(n13362), .ZN(P1_U2868) );
  INV_X1 U16622 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U16623 ( .A1(n9850), .A2(n13390), .ZN(n13403) );
  INV_X1 U16624 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13365) );
  OAI22_X1 U16625 ( .A1(n13366), .A2(n19691), .B1(n19786), .B2(n13365), .ZN(
        n13381) );
  INV_X1 U16626 ( .A(n13368), .ZN(n13369) );
  NAND2_X1 U16627 ( .A1(n13369), .A2(n13364), .ZN(n13643) );
  INV_X1 U16628 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U16629 ( .A1(n13639), .A2(n13371), .B1(n13643), .B2(n13370), .ZN(
        n13372) );
  INV_X1 U16630 ( .A(n13372), .ZN(n13379) );
  INV_X1 U16631 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13375) );
  OAI22_X1 U16632 ( .A1(n13376), .A2(n13434), .B1(n13424), .B2(n13375), .ZN(
        n13377) );
  INV_X1 U16633 ( .A(n13377), .ZN(n13378) );
  NAND2_X1 U16634 ( .A1(n13379), .A2(n13378), .ZN(n13380) );
  NOR2_X1 U16635 ( .A1(n13381), .A2(n13380), .ZN(n13410) );
  INV_X1 U16636 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13521) );
  AOI21_X1 U16637 ( .B1(n14880), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n12403), .ZN(n13384) );
  NOR2_X1 U16638 ( .A1(n9851), .A2(n19250), .ZN(n13382) );
  NAND2_X1 U16639 ( .A1(n13382), .A2(n9854), .ZN(n13648) );
  OAI211_X1 U16640 ( .C1(n14893), .C2(n13521), .A(n13384), .B(n13383), .ZN(
        n13385) );
  INV_X1 U16641 ( .A(n13385), .ZN(n13409) );
  INV_X1 U16642 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13386) );
  INV_X1 U16643 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13393) );
  OAI22_X1 U16644 ( .A1(n13393), .A2(n19542), .B1(n19624), .B2(n13392), .ZN(
        n13394) );
  NOR2_X1 U16645 ( .A1(n9851), .A2(n13402), .ZN(n13397) );
  INV_X1 U16646 ( .A(n19507), .ZN(n13398) );
  NAND2_X1 U16647 ( .A1(n13398), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13406) );
  OR2_X2 U16648 ( .A1(n13403), .A2(n13402), .ZN(n13654) );
  NAND4_X1 U16649 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13414) );
  NAND2_X1 U16650 ( .A1(n13412), .A2(n13411), .ZN(n13413) );
  INV_X1 U16651 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13416) );
  OAI22_X1 U16652 ( .A1(n13416), .A2(n19576), .B1(n19624), .B2(n13415), .ZN(
        n13420) );
  OAI22_X1 U16653 ( .A1(n13418), .A2(n13648), .B1(n19507), .B2(n13417), .ZN(
        n13419) );
  NOR2_X1 U16654 ( .A1(n13420), .A2(n13419), .ZN(n13440) );
  INV_X1 U16655 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13422) );
  INV_X1 U16656 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13421) );
  OAI22_X1 U16657 ( .A1(n19478), .A2(n13422), .B1(n13643), .B2(n13421), .ZN(
        n13423) );
  INV_X1 U16658 ( .A(n13423), .ZN(n13426) );
  OAI22_X1 U16659 ( .A1(n13430), .A2(n19542), .B1(n13639), .B2(n13429), .ZN(
        n13438) );
  OAI22_X1 U16660 ( .A1(n13432), .A2(n19786), .B1(n13654), .B2(n13431), .ZN(
        n13437) );
  NAND4_X1 U16661 ( .A1(n13440), .A2(n10511), .A3(n9908), .A4(n13439), .ZN(
        n13441) );
  NAND2_X1 U16662 ( .A1(n13441), .A2(n13442), .ZN(n13445) );
  NAND2_X1 U16663 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  NAND2_X1 U16664 ( .A1(n9926), .A2(n13450), .ZN(n13692) );
  NAND2_X1 U16665 ( .A1(n13524), .A2(n13523), .ZN(n13455) );
  INV_X1 U16666 ( .A(n13631), .ZN(n13452) );
  NAND2_X1 U16667 ( .A1(n13452), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13453) );
  AND2_X1 U16668 ( .A1(n13454), .A2(n13453), .ZN(n13522) );
  XNOR2_X1 U16669 ( .A(n13455), .B(n13522), .ZN(n16397) );
  NOR2_X1 U16670 ( .A1(n13456), .A2(n13537), .ZN(n13458) );
  NOR2_X1 U16671 ( .A1(n13458), .A2(n13457), .ZN(n13530) );
  XNOR2_X1 U16672 ( .A(n13451), .B(n13530), .ZN(n13459) );
  AND2_X1 U16673 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NOR2_X1 U16674 ( .A1(n13533), .A2(n13461), .ZN(n16394) );
  INV_X1 U16675 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13694) );
  OAI22_X1 U16676 ( .A1(n13694), .A2(n19423), .B1(n16277), .B2(n13690), .ZN(
        n13462) );
  AOI21_X1 U16677 ( .B1(n19412), .B2(P2_REIP_REG_3__SCAN_IN), .A(n13462), .ZN(
        n13463) );
  OAI21_X1 U16678 ( .B1(n13401), .B2(n16284), .A(n13463), .ZN(n13464) );
  AOI21_X1 U16679 ( .B1(n16394), .B2(n16294), .A(n13464), .ZN(n13465) );
  OAI21_X1 U16680 ( .B1(n16397), .B2(n19415), .A(n13465), .ZN(P2_U3011) );
  NOR2_X1 U16681 ( .A1(n13467), .A2(n13466), .ZN(n13468) );
  OR2_X1 U16682 ( .A1(n13478), .A2(n13468), .ZN(n15436) );
  INV_X1 U16683 ( .A(n13469), .ZN(n13473) );
  OAI21_X1 U16684 ( .B1(n13295), .B2(n13471), .A(n13470), .ZN(n13472) );
  NAND3_X1 U16685 ( .A1(n13473), .A2(n14746), .A3(n13472), .ZN(n13475) );
  NAND2_X1 U16686 ( .A1(n14749), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13474) );
  OAI211_X1 U16687 ( .C1(n15436), .C2(n14749), .A(n13475), .B(n13474), .ZN(
        P2_U2873) );
  XNOR2_X1 U16688 ( .A(n13469), .B(n13476), .ZN(n13480) );
  OAI21_X1 U16689 ( .B1(n13478), .B2(n13477), .A(n13625), .ZN(n16229) );
  MUX2_X1 U16690 ( .A(n12744), .B(n16229), .S(n14769), .Z(n13479) );
  OAI21_X1 U16691 ( .B1(n13480), .B2(n14779), .A(n13479), .ZN(P2_U2872) );
  XOR2_X1 U16692 ( .A(n13352), .B(n13481), .Z(n20156) );
  OR2_X1 U16693 ( .A1(n16086), .A2(n13482), .ZN(n13483) );
  NAND2_X1 U16694 ( .A1(n13617), .A2(n13483), .ZN(n20151) );
  OAI22_X1 U16695 ( .A1(n20151), .A2(n14312), .B1(n21334), .B2(n20211), .ZN(
        n13484) );
  AOI21_X1 U16696 ( .B1(n20156), .B2(n20207), .A(n13484), .ZN(n13485) );
  INV_X1 U16697 ( .A(n13485), .ZN(P1_U2866) );
  NAND2_X1 U16698 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21018), .ZN(n15823) );
  NAND2_X1 U16699 ( .A1(n10916), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13486) );
  MUX2_X1 U16700 ( .A(n15823), .B(n13486), .S(n21012), .Z(n13487) );
  INV_X1 U16701 ( .A(n13487), .ZN(n13488) );
  INV_X1 U16702 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13490) );
  OAI21_X1 U16703 ( .B1(n13507), .B2(n13493), .A(n20133), .ZN(n20197) );
  INV_X1 U16704 ( .A(n20197), .ZN(n14263) );
  INV_X1 U16705 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21352) );
  NAND2_X1 U16706 ( .A1(n13496), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13498) );
  AND2_X1 U16707 ( .A1(n16097), .A2(n21346), .ZN(n15818) );
  NOR2_X1 U16708 ( .A1(n13498), .A2(n15818), .ZN(n13497) );
  INV_X1 U16709 ( .A(n13498), .ZN(n13499) );
  NOR2_X1 U16710 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  OAI22_X1 U16711 ( .A1(n20343), .A2(n20174), .B1(n10416), .B2(n20201), .ZN(
        n13504) );
  NOR2_X1 U16712 ( .A1(n20161), .A2(n21352), .ZN(n13503) );
  AOI211_X1 U16713 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13504), .B(n13503), .ZN(n13505) );
  OAI21_X1 U16714 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20184), .A(
        n13505), .ZN(n13510) );
  INV_X1 U16715 ( .A(n13507), .ZN(n13508) );
  NAND2_X1 U16716 ( .A1(n13508), .A2(n15776), .ZN(n20187) );
  NOR2_X1 U16717 ( .A1(n20595), .A2(n20187), .ZN(n13509) );
  AOI211_X1 U16718 ( .C1(n20179), .C2(n21352), .A(n13510), .B(n13509), .ZN(
        n13511) );
  OAI21_X1 U16719 ( .B1(n13512), .B2(n14263), .A(n13511), .ZN(P1_U2839) );
  INV_X1 U16720 ( .A(n14893), .ZN(n13517) );
  NOR2_X1 U16721 ( .A1(n19822), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13515) );
  NOR2_X1 U16722 ( .A1(n19508), .A2(n19758), .ZN(n19749) );
  AOI221_X1 U16723 ( .B1(n19751), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19781), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19727), .ZN(n13513) );
  NOR2_X1 U16724 ( .A1(n13513), .A2(n19861), .ZN(n13514) );
  AOI211_X1 U16725 ( .C1(n13517), .C2(n13515), .A(n19749), .B(n13514), .ZN(
        n13516) );
  AOI22_X1 U16726 ( .A1(n19751), .A2(n19900), .B1(n19781), .B2(n19798), .ZN(
        n13520) );
  OAI21_X1 U16727 ( .B1(n13517), .B2(n19749), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13518) );
  OAI21_X1 U16728 ( .B1(n19758), .B2(n19509), .A(n13518), .ZN(n19750) );
  AOI22_X1 U16729 ( .A1(n19750), .A2(n13231), .B1(n19899), .B2(n19749), .ZN(
        n13519) );
  OAI211_X1 U16730 ( .C1(n19755), .C2(n13521), .A(n13520), .B(n13519), .ZN(
        P2_U3129) );
  NAND2_X1 U16731 ( .A1(n13523), .A2(n13522), .ZN(n13525) );
  NAND2_X1 U16732 ( .A1(n13525), .A2(n13524), .ZN(n13674) );
  NAND2_X1 U16733 ( .A1(n9926), .A2(n10196), .ZN(n13527) );
  NAND2_X1 U16734 ( .A1(n9927), .A2(n13527), .ZN(n19234) );
  INV_X1 U16735 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13677) );
  XNOR2_X1 U16736 ( .A(n19234), .B(n13677), .ZN(n13673) );
  XNOR2_X1 U16737 ( .A(n13674), .B(n13673), .ZN(n19414) );
  NOR2_X1 U16738 ( .A1(n13530), .A2(n13451), .ZN(n13532) );
  OAI21_X1 U16739 ( .B1(n13533), .B2(n13532), .A(n13531), .ZN(n13676) );
  INV_X1 U16740 ( .A(n13676), .ZN(n13534) );
  NOR2_X1 U16741 ( .A1(n13675), .A2(n13534), .ZN(n13535) );
  XNOR2_X1 U16742 ( .A(n13535), .B(n13677), .ZN(n19413) );
  NOR2_X1 U16743 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  NAND2_X1 U16744 ( .A1(n13539), .A2(n13538), .ZN(n13542) );
  INV_X1 U16745 ( .A(n15248), .ZN(n13540) );
  OR2_X1 U16746 ( .A1(n15414), .A2(n13540), .ZN(n13541) );
  NOR2_X1 U16747 ( .A1(n16390), .A2(n13451), .ZN(n16383) );
  AND2_X1 U16748 ( .A1(n13544), .A2(n13543), .ZN(n15250) );
  OAI21_X1 U16749 ( .B1(n15414), .B2(n15248), .A(n15250), .ZN(n16392) );
  AOI21_X1 U16750 ( .B1(n13451), .B2(n15419), .A(n16392), .ZN(n16372) );
  INV_X1 U16751 ( .A(n16372), .ZN(n13546) );
  INV_X1 U16752 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19985) );
  NOR2_X1 U16753 ( .A1(n19985), .A2(n16334), .ZN(n13545) );
  AOI221_X1 U16754 ( .B1(n16383), .B2(n13677), .C1(n13546), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n13545), .ZN(n13548) );
  NAND2_X1 U16755 ( .A1(n19419), .A2(n16407), .ZN(n13547) );
  OAI211_X1 U16756 ( .C1(n16364), .C2(n19231), .A(n13548), .B(n13547), .ZN(
        n13549) );
  AOI21_X1 U16757 ( .B1(n19413), .B2(n16393), .A(n13549), .ZN(n13550) );
  OAI21_X1 U16758 ( .B1(n16402), .B2(n19414), .A(n13550), .ZN(P2_U3042) );
  INV_X1 U16759 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13551) );
  OR2_X1 U16760 ( .A1(n14369), .A2(n13551), .ZN(n13553) );
  NAND2_X1 U16761 ( .A1(n14369), .A2(DATAI_6_), .ZN(n13552) );
  AND2_X1 U16762 ( .A1(n13553), .A2(n13552), .ZN(n20376) );
  INV_X1 U16763 ( .A(n20156), .ZN(n13554) );
  OAI222_X1 U16764 ( .A1(n14379), .A2(n20376), .B1(n14382), .B2(n13554), .C1(
        n10981), .C2(n14380), .ZN(P1_U2898) );
  OAI21_X1 U16765 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(n15973) );
  NAND2_X1 U16766 ( .A1(n20307), .A2(n13559), .ZN(n16091) );
  AOI21_X1 U16767 ( .B1(n13561), .B2(n13560), .A(n20325), .ZN(n16052) );
  OAI21_X1 U16768 ( .B1(n16055), .B2(n13562), .A(n16052), .ZN(n16087) );
  INV_X1 U16769 ( .A(n16087), .ZN(n13563) );
  OAI211_X1 U16770 ( .C1(n13558), .C2(n16091), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13563), .ZN(n13749) );
  OAI21_X1 U16771 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16044), .A(
        n13749), .ZN(n13567) );
  INV_X1 U16772 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13564) );
  OAI22_X1 U16773 ( .A1(n20151), .A2(n20344), .B1(n20342), .B2(n13564), .ZN(
        n13565) );
  INV_X1 U16774 ( .A(n13565), .ZN(n13566) );
  OAI211_X1 U16775 ( .C1(n15973), .C2(n20340), .A(n13567), .B(n13566), .ZN(
        P1_U3025) );
  OAI21_X1 U16776 ( .B1(n20407), .B2(n20911), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13571) );
  NAND2_X1 U16777 ( .A1(n13571), .A2(n20848), .ZN(n13584) );
  INV_X1 U16778 ( .A(n13584), .ZN(n13576) );
  INV_X1 U16779 ( .A(n20720), .ZN(n13572) );
  OR2_X1 U16780 ( .A1(n20594), .A2(n13572), .ZN(n20446) );
  OR2_X1 U16781 ( .A1(n20446), .A2(n10856), .ZN(n13583) );
  NAND3_X1 U16782 ( .A1(n20653), .A2(n11313), .A3(n20723), .ZN(n20387) );
  NOR2_X1 U16783 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20387), .ZN(
        n20356) );
  INV_X1 U16784 ( .A(n13573), .ZN(n20597) );
  NAND2_X1 U16785 ( .A1(n20597), .A2(n20654), .ZN(n20479) );
  NAND2_X1 U16786 ( .A1(n20479), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13574) );
  NOR2_X1 U16787 ( .A1(n13581), .A2(n20625), .ZN(n20722) );
  NOR2_X1 U16788 ( .A1(n20483), .A2(n20722), .ZN(n20604) );
  OAI211_X1 U16789 ( .C1(n20356), .C2(n20985), .A(n13574), .B(n20604), .ZN(
        n13575) );
  INV_X1 U16790 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16569) );
  INV_X1 U16791 ( .A(DATAI_18_), .ZN(n21340) );
  OAI22_X1 U16792 ( .A1(n16569), .A2(n20377), .B1(n21340), .B2(n20379), .ZN(
        n20873) );
  INV_X1 U16793 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19438) );
  INV_X1 U16794 ( .A(DATAI_26_), .ZN(n21144) );
  OAI22_X1 U16795 ( .A1(n19438), .A2(n20377), .B1(n21144), .B2(n20379), .ZN(
        n20818) );
  INV_X1 U16796 ( .A(n20818), .ZN(n20876) );
  INV_X1 U16797 ( .A(n20356), .ZN(n20374) );
  NAND3_X1 U16798 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21012), .A3(n13578), 
        .ZN(n20365) );
  NAND2_X1 U16799 ( .A1(n20373), .A2(n13579), .ZN(n20871) );
  OAI22_X1 U16800 ( .A1(n20904), .A2(n20876), .B1(n20374), .B2(n20871), .ZN(
        n13580) );
  AOI21_X1 U16801 ( .B1(n20407), .B2(n20873), .A(n13580), .ZN(n13586) );
  INV_X1 U16802 ( .A(n13581), .ZN(n13582) );
  NOR2_X1 U16803 ( .A1(n13582), .A2(n20625), .ZN(n20656) );
  INV_X1 U16804 ( .A(n20656), .ZN(n20598) );
  NAND2_X1 U16805 ( .A1(n20380), .A2(n20816), .ZN(n13585) );
  OAI211_X1 U16806 ( .C1(n20384), .C2(n13587), .A(n13586), .B(n13585), .ZN(
        P1_U3035) );
  INV_X1 U16807 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13593) );
  INV_X1 U16808 ( .A(DATAI_19_), .ZN(n21051) );
  INV_X1 U16809 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16567) );
  OAI22_X2 U16810 ( .A1(n21051), .A2(n20379), .B1(n16567), .B2(n20377), .ZN(
        n20880) );
  INV_X1 U16811 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19444) );
  INV_X1 U16812 ( .A(DATAI_27_), .ZN(n13588) );
  OAI22_X1 U16813 ( .A1(n19444), .A2(n20377), .B1(n13588), .B2(n20379), .ZN(
        n20824) );
  INV_X1 U16814 ( .A(n20824), .ZN(n20883) );
  NAND2_X1 U16815 ( .A1(n20373), .A2(n13589), .ZN(n20878) );
  OAI22_X1 U16816 ( .A1(n20904), .A2(n20883), .B1(n20374), .B2(n20878), .ZN(
        n13590) );
  AOI21_X1 U16817 ( .B1(n20407), .B2(n20880), .A(n13590), .ZN(n13592) );
  NAND2_X1 U16818 ( .A1(n20380), .A2(n20822), .ZN(n13591) );
  OAI211_X1 U16819 ( .C1(n20384), .C2(n13593), .A(n13592), .B(n13591), .ZN(
        P1_U3036) );
  INV_X1 U16820 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13598) );
  INV_X1 U16821 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16565) );
  INV_X1 U16822 ( .A(DATAI_20_), .ZN(n21101) );
  INV_X1 U16823 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19451) );
  INV_X1 U16824 ( .A(DATAI_28_), .ZN(n21369) );
  NAND2_X1 U16825 ( .A1(n20373), .A2(n13594), .ZN(n20887) );
  OAI22_X1 U16826 ( .A1(n20904), .A2(n9980), .B1(n20374), .B2(n20887), .ZN(
        n13595) );
  AOI21_X1 U16827 ( .B1(n20407), .B2(n20889), .A(n13595), .ZN(n13597) );
  NAND2_X1 U16828 ( .A1(n20380), .A2(n20828), .ZN(n13596) );
  OAI211_X1 U16829 ( .C1(n20384), .C2(n13598), .A(n13597), .B(n13596), .ZN(
        P1_U3037) );
  INV_X1 U16830 ( .A(DATAI_16_), .ZN(n21332) );
  INV_X1 U16831 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16572) );
  OAI22_X1 U16832 ( .A1(n21332), .A2(n20379), .B1(n16572), .B2(n20377), .ZN(
        n20773) );
  INV_X1 U16833 ( .A(DATAI_24_), .ZN(n21337) );
  OAI22_X2 U16834 ( .A1(n21337), .A2(n20379), .B1(n16559), .B2(n20377), .ZN(
        n20860) );
  INV_X1 U16835 ( .A(n20860), .ZN(n20776) );
  NAND2_X1 U16836 ( .A1(n20373), .A2(n13599), .ZN(n20853) );
  OAI22_X1 U16837 ( .A1(n20904), .A2(n20776), .B1(n20374), .B2(n20853), .ZN(
        n13600) );
  AOI21_X1 U16838 ( .B1(n20407), .B2(n20773), .A(n13600), .ZN(n13602) );
  NAND2_X1 U16839 ( .A1(n20380), .A2(n20805), .ZN(n13601) );
  OAI211_X1 U16840 ( .C1(n20384), .C2(n13603), .A(n13602), .B(n13601), .ZN(
        P1_U3033) );
  INV_X1 U16841 ( .A(DATAI_23_), .ZN(n21194) );
  INV_X1 U16842 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16561) );
  OAI22_X2 U16843 ( .A1(n21194), .A2(n20379), .B1(n16561), .B2(n20377), .ZN(
        n20910) );
  INV_X1 U16844 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19469) );
  OAI22_X1 U16845 ( .A1(n19469), .A2(n20377), .B1(n11679), .B2(n20379), .ZN(
        n20841) );
  INV_X1 U16846 ( .A(n20841), .ZN(n20916) );
  NAND2_X1 U16847 ( .A1(n20373), .A2(n10695), .ZN(n20758) );
  OAI22_X1 U16848 ( .A1(n20904), .A2(n20916), .B1(n20374), .B2(n20758), .ZN(
        n13604) );
  AOI21_X1 U16849 ( .B1(n20407), .B2(n20910), .A(n13604), .ZN(n13608) );
  INV_X1 U16850 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16589) );
  OR2_X1 U16851 ( .A1(n14369), .A2(n16589), .ZN(n13606) );
  NAND2_X1 U16852 ( .A1(n14369), .A2(DATAI_7_), .ZN(n13605) );
  AND2_X1 U16853 ( .A1(n13606), .A2(n13605), .ZN(n20266) );
  NAND2_X1 U16854 ( .A1(n20380), .A2(n20907), .ZN(n13607) );
  OAI211_X1 U16855 ( .C1(n20384), .C2(n13609), .A(n13608), .B(n13607), .ZN(
        P1_U3040) );
  NAND2_X1 U16856 ( .A1(n13614), .A2(n13613), .ZN(n13615) );
  AND2_X1 U16857 ( .A1(n13611), .A2(n13615), .ZN(n20148) );
  INV_X1 U16858 ( .A(n20148), .ZN(n13620) );
  INV_X1 U16859 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21181) );
  NAND2_X1 U16860 ( .A1(n13617), .A2(n13616), .ZN(n13618) );
  AND2_X1 U16861 ( .A1(n13735), .A2(n13618), .ZN(n20144) );
  INV_X1 U16862 ( .A(n20144), .ZN(n13619) );
  OAI222_X1 U16863 ( .A1(n13620), .A2(n14318), .B1(n20211), .B2(n21181), .C1(
        n13619), .C2(n14312), .ZN(P1_U2865) );
  INV_X1 U16864 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20230) );
  OAI222_X1 U16865 ( .A1(n14382), .A2(n13620), .B1(n14380), .B2(n20230), .C1(
        n14379), .C2(n20266), .ZN(P1_U2897) );
  OAI21_X1 U16866 ( .B1(n13623), .B2(n13622), .A(n13621), .ZN(n13745) );
  INV_X1 U16867 ( .A(n13730), .ZN(n13624) );
  AOI21_X1 U16868 ( .B1(n13626), .B2(n13625), .A(n13624), .ZN(n19105) );
  NOR2_X1 U16869 ( .A1(n14769), .A2(n14973), .ZN(n13627) );
  AOI21_X1 U16870 ( .B1(n19105), .B2(n14769), .A(n13627), .ZN(n13628) );
  OAI21_X1 U16871 ( .B1(n13745), .B2(n14779), .A(n13628), .ZN(P2_U2871) );
  NAND2_X1 U16872 ( .A1(n9831), .A2(n13761), .ZN(n13629) );
  XNOR2_X1 U16873 ( .A(n13630), .B(n13629), .ZN(n13637) );
  OAI22_X1 U16874 ( .A1(n19982), .A2(n19183), .B1(n13631), .B2(n19233), .ZN(
        n13633) );
  OAI22_X1 U16875 ( .A1(n19110), .A2(n11855), .B1(n12668), .B2(n19185), .ZN(
        n13632) );
  AOI211_X1 U16876 ( .C1(n19251), .C2(n20067), .A(n13633), .B(n13632), .ZN(
        n13635) );
  OAI211_X1 U16877 ( .C1(n13710), .C2(n20065), .A(n13635), .B(n13634), .ZN(
        n13636) );
  AOI21_X1 U16878 ( .B1(n13637), .B2(n19226), .A(n13636), .ZN(n13638) );
  INV_X1 U16879 ( .A(n13638), .ZN(P2_U2853) );
  AOI22_X1 U16880 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n14876), .B1(
        n19757), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13647) );
  INV_X1 U16881 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13641) );
  OAI22_X1 U16882 ( .A1(n13641), .A2(n19478), .B1(n13639), .B2(n13640), .ZN(
        n13642) );
  INV_X1 U16883 ( .A(n13642), .ZN(n13646) );
  INV_X1 U16884 ( .A(n13643), .ZN(n19823) );
  AOI22_X1 U16885 ( .A1(n19546), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n19823), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U16886 ( .A1(n14881), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14880), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13644) );
  OAI22_X1 U16887 ( .A1(n12103), .A2(n13648), .B1(n19507), .B2(n13649), .ZN(
        n13653) );
  INV_X1 U16888 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13651) );
  OAI22_X1 U16889 ( .A1(n13651), .A2(n19576), .B1(n19624), .B2(n13650), .ZN(
        n13652) );
  NOR2_X1 U16890 ( .A1(n13653), .A2(n13652), .ZN(n13663) );
  INV_X1 U16891 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13656) );
  OAI22_X1 U16892 ( .A1(n13656), .A2(n19691), .B1(n13654), .B2(n13655), .ZN(
        n13657) );
  INV_X1 U16893 ( .A(n13657), .ZN(n13662) );
  INV_X1 U16894 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13659) );
  OAI22_X1 U16895 ( .A1(n13659), .A2(n14893), .B1(n19786), .B2(n13658), .ZN(
        n13660) );
  INV_X1 U16896 ( .A(n13660), .ZN(n13661) );
  NAND2_X1 U16897 ( .A1(n13665), .A2(n12403), .ZN(n13666) );
  NAND2_X1 U16898 ( .A1(n13678), .A2(n15043), .ZN(n13671) );
  INV_X1 U16899 ( .A(n14917), .ZN(n13670) );
  NAND2_X1 U16900 ( .A1(n9927), .A2(n10195), .ZN(n13669) );
  NAND2_X1 U16901 ( .A1(n13670), .A2(n13669), .ZN(n19219) );
  NAND2_X1 U16902 ( .A1(n13671), .A2(n19219), .ZN(n14875) );
  INV_X1 U16903 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13672) );
  XNOR2_X1 U16904 ( .A(n14874), .B(n14873), .ZN(n13728) );
  INV_X1 U16905 ( .A(n13678), .ZN(n13679) );
  NAND2_X1 U16906 ( .A1(n13679), .A2(n13672), .ZN(n13681) );
  NAND2_X1 U16907 ( .A1(n13680), .A2(n13681), .ZN(n15045) );
  INV_X1 U16908 ( .A(n15049), .ZN(n13683) );
  AOI21_X1 U16909 ( .B1(n13683), .B2(n13681), .A(n9817), .ZN(n13682) );
  AOI21_X1 U16910 ( .B1(n9814), .B2(n13683), .A(n13682), .ZN(n13726) );
  INV_X1 U16911 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13684) );
  OAI22_X1 U16912 ( .A1(n13684), .A2(n19423), .B1(n16277), .B2(n19223), .ZN(
        n13685) );
  AOI21_X1 U16913 ( .B1(n19412), .B2(P2_REIP_REG_5__SCAN_IN), .A(n13685), .ZN(
        n13686) );
  OAI21_X1 U16914 ( .B1(n16284), .B2(n19229), .A(n13686), .ZN(n13687) );
  AOI21_X1 U16915 ( .B1(n13726), .B2(n16294), .A(n13687), .ZN(n13688) );
  OAI21_X1 U16916 ( .B1(n19415), .B2(n13728), .A(n13688), .ZN(P2_U3009) );
  NOR2_X1 U16917 ( .A1(n9835), .A2(n13689), .ZN(n13691) );
  XNOR2_X1 U16918 ( .A(n13691), .B(n13690), .ZN(n13700) );
  OAI22_X1 U16919 ( .A1(n19984), .A2(n19183), .B1(n13692), .B2(n19233), .ZN(
        n13696) );
  OAI22_X1 U16920 ( .A1(n13694), .A2(n19185), .B1(n19232), .B2(n13693), .ZN(
        n13695) );
  AOI211_X1 U16921 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19189), .A(n13696), .B(
        n13695), .ZN(n13698) );
  NAND2_X1 U16922 ( .A1(n13396), .A2(n19249), .ZN(n13697) );
  OAI211_X1 U16923 ( .C1(n13710), .C2(n15526), .A(n13698), .B(n13697), .ZN(
        n13699) );
  AOI21_X1 U16924 ( .B1(n13700), .B2(n19226), .A(n13699), .ZN(n13701) );
  INV_X1 U16925 ( .A(n13701), .ZN(P2_U2852) );
  NAND2_X1 U16926 ( .A1(n13611), .A2(n13703), .ZN(n13704) );
  NAND2_X1 U16927 ( .A1(n13702), .A2(n13704), .ZN(n20134) );
  AOI22_X1 U16928 ( .A1(n14375), .A2(n14332), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14374), .ZN(n13705) );
  OAI21_X1 U16929 ( .B1(n20134), .B2(n14382), .A(n13705), .ZN(P1_U2896) );
  NOR2_X1 U16930 ( .A1(n9835), .A2(n13764), .ZN(n13766) );
  INV_X1 U16931 ( .A(n13766), .ZN(n13715) );
  NAND2_X1 U16932 ( .A1(n19226), .A2(n9835), .ZN(n19141) );
  INV_X1 U16933 ( .A(n19141), .ZN(n19256) );
  OAI21_X1 U16934 ( .B1(n19245), .B2(n19256), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U16935 ( .A1(n19248), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19247), 
        .B2(n13706), .ZN(n13708) );
  NAND2_X1 U16936 ( .A1(n19244), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n13707) );
  OAI211_X1 U16937 ( .C1(n13709), .C2(n19232), .A(n13708), .B(n13707), .ZN(
        n13712) );
  NOR2_X1 U16938 ( .A1(n20081), .A2(n13710), .ZN(n13711) );
  AOI211_X1 U16939 ( .C1(n19249), .C2(n13200), .A(n13712), .B(n13711), .ZN(
        n13713) );
  OAI211_X1 U16940 ( .C1(n13715), .C2(n19953), .A(n13714), .B(n13713), .ZN(
        P2_U2855) );
  NAND2_X1 U16941 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19412), .ZN(n13717) );
  NAND2_X1 U16942 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16371) );
  OAI211_X1 U16943 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16383), .B(n16371), .ZN(n13716) );
  OAI211_X1 U16944 ( .C1(n16372), .C2(n13672), .A(n13717), .B(n13716), .ZN(
        n13725) );
  INV_X1 U16945 ( .A(n13718), .ZN(n13720) );
  NAND2_X1 U16946 ( .A1(n13720), .A2(n13719), .ZN(n13722) );
  AND2_X1 U16947 ( .A1(n13722), .A2(n13721), .ZN(n19295) );
  INV_X1 U16948 ( .A(n19295), .ZN(n13723) );
  OAI22_X1 U16949 ( .A1(n19229), .A2(n16365), .B1(n16364), .B2(n13723), .ZN(
        n13724) );
  AOI211_X1 U16950 ( .C1(n13726), .C2(n16393), .A(n13725), .B(n13724), .ZN(
        n13727) );
  OAI21_X1 U16951 ( .B1(n16402), .B2(n13728), .A(n13727), .ZN(P2_U3041) );
  OAI21_X1 U16952 ( .B1(n10412), .B2(n10505), .A(n13756), .ZN(n14872) );
  NAND2_X1 U16953 ( .A1(n14749), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13733) );
  AND2_X1 U16954 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  OR2_X1 U16955 ( .A1(n13731), .A2(n9932), .ZN(n19095) );
  INV_X1 U16956 ( .A(n19095), .ZN(n15212) );
  NAND2_X1 U16957 ( .A1(n15212), .A2(n14769), .ZN(n13732) );
  OAI211_X1 U16958 ( .C1(n14872), .C2(n14779), .A(n13733), .B(n13732), .ZN(
        P2_U2870) );
  INV_X1 U16959 ( .A(n20134), .ZN(n13786) );
  NAND2_X1 U16960 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  NAND2_X1 U16961 ( .A1(n16066), .A2(n13736), .ZN(n20130) );
  OAI22_X1 U16962 ( .A1(n20130), .A2(n14312), .B1(n21250), .B2(n20211), .ZN(
        n13737) );
  AOI21_X1 U16963 ( .B1(n13786), .B2(n20207), .A(n13737), .ZN(n13738) );
  INV_X1 U16964 ( .A(n13738), .ZN(P1_U2864) );
  OAI21_X1 U16965 ( .B1(n13739), .B2(n16313), .A(n14865), .ZN(n19108) );
  INV_X1 U16966 ( .A(n19108), .ZN(n13742) );
  OAI22_X1 U16967 ( .A1(n14868), .A2(n19386), .B1(n19282), .B2(n13740), .ZN(
        n13741) );
  AOI21_X1 U16968 ( .B1(n19318), .B2(n13742), .A(n13741), .ZN(n13744) );
  AOI22_X1 U16969 ( .A1(n19262), .A2(BUF1_REG_16__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n13743) );
  OAI211_X1 U16970 ( .C1(n13745), .C2(n19269), .A(n13744), .B(n13743), .ZN(
        P2_U2903) );
  XNOR2_X1 U16971 ( .A(n13746), .B(n13751), .ZN(n13747) );
  XNOR2_X1 U16972 ( .A(n13748), .B(n13747), .ZN(n13788) );
  INV_X1 U16973 ( .A(n20130), .ZN(n13753) );
  AND2_X1 U16974 ( .A1(n20317), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13783) );
  NAND2_X1 U16975 ( .A1(n16057), .A2(n13749), .ZN(n16078) );
  NAND2_X1 U16976 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16044), .ZN(
        n16080) );
  OAI21_X1 U16977 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16061), .ZN(n13750) );
  OAI22_X1 U16978 ( .A1(n13751), .A2(n16078), .B1(n16080), .B2(n13750), .ZN(
        n13752) );
  AOI211_X1 U16979 ( .C1(n20316), .C2(n13753), .A(n13783), .B(n13752), .ZN(
        n13754) );
  OAI21_X1 U16980 ( .B1(n13788), .B2(n20340), .A(n13754), .ZN(P1_U3023) );
  AOI21_X1 U16981 ( .B1(n13757), .B2(n13756), .A(n13755), .ZN(n13758) );
  INV_X1 U16982 ( .A(n13758), .ZN(n14863) );
  OAI21_X1 U16983 ( .B1(n9932), .B2(n13759), .A(n14774), .ZN(n16308) );
  MUX2_X1 U16984 ( .A(n14955), .B(n16308), .S(n14769), .Z(n13760) );
  OAI21_X1 U16985 ( .B1(n14863), .B2(n14779), .A(n13760), .ZN(P2_U2869) );
  OAI211_X1 U16986 ( .C1(n13764), .C2(n13763), .A(n9831), .B(n13761), .ZN(
        n19261) );
  OAI21_X1 U16987 ( .B1(n9831), .B2(n13765), .A(n19261), .ZN(n13833) );
  AOI21_X1 U16988 ( .B1(n9835), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13766), .ZN(n13796) );
  NOR2_X1 U16989 ( .A1(n13796), .A2(n13767), .ZN(n13834) );
  INV_X1 U16990 ( .A(n16465), .ZN(n15525) );
  NOR2_X1 U16991 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13837), .ZN(
        n13778) );
  INV_X1 U16992 ( .A(n13768), .ZN(n13769) );
  NAND2_X1 U16993 ( .A1(n15515), .A2(n13769), .ZN(n15519) );
  OR2_X1 U16994 ( .A1(n16431), .A2(n16434), .ZN(n15516) );
  NAND2_X1 U16995 ( .A1(n13770), .A2(n12933), .ZN(n13771) );
  NAND2_X1 U16996 ( .A1(n13771), .A2(n13773), .ZN(n15518) );
  NOR2_X1 U16997 ( .A1(n13828), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13772) );
  NOR2_X1 U16998 ( .A1(n15518), .A2(n13772), .ZN(n13776) );
  INV_X1 U16999 ( .A(n15518), .ZN(n13775) );
  INV_X1 U17000 ( .A(n13772), .ZN(n15517) );
  NAND2_X1 U17001 ( .A1(n13773), .A2(n15517), .ZN(n13774) );
  OAI22_X1 U17002 ( .A1(n15516), .A2(n13776), .B1(n13775), .B2(n13774), .ZN(
        n13777) );
  OAI21_X1 U17003 ( .B1(n13778), .B2(n15519), .A(n13777), .ZN(n13779) );
  INV_X1 U17004 ( .A(n13836), .ZN(n20054) );
  OAI22_X1 U17005 ( .A1(n20065), .A2(n15525), .B1(n16414), .B2(n20054), .ZN(
        n13780) );
  AOI21_X1 U17006 ( .B1(n13833), .B2(n13834), .A(n13780), .ZN(n13782) );
  NAND2_X1 U17007 ( .A1(n15527), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13781) );
  OAI21_X1 U17008 ( .B1(n13782), .B2(n15527), .A(n13781), .ZN(P2_U3599) );
  AOI21_X1 U17009 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13783), .ZN(n13784) );
  OAI21_X1 U17010 ( .B1(n20302), .B2(n20132), .A(n13784), .ZN(n13785) );
  AOI21_X1 U17011 ( .B1(n13786), .B2(n15981), .A(n13785), .ZN(n13787) );
  OAI21_X1 U17012 ( .B1(n13788), .B2(n20108), .A(n13787), .ZN(P1_U2991) );
  AOI21_X1 U17013 ( .B1(n13790), .B2(n13702), .A(n13789), .ZN(n20204) );
  INV_X1 U17014 ( .A(n20204), .ZN(n13825) );
  AOI22_X1 U17015 ( .A1(n14375), .A2(n20267), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14374), .ZN(n13791) );
  OAI21_X1 U17016 ( .B1(n13825), .B2(n14382), .A(n13791), .ZN(P1_U2895) );
  INV_X1 U17017 ( .A(n15527), .ZN(n13802) );
  NOR2_X1 U17018 ( .A1(n13792), .A2(n15525), .ZN(n13799) );
  NAND2_X1 U17019 ( .A1(n13794), .A2(n13793), .ZN(n13830) );
  MUX2_X1 U17020 ( .A(n15515), .B(n13830), .S(n13801), .Z(n13795) );
  AOI21_X1 U17021 ( .B1(n13200), .B2(n15524), .A(n13795), .ZN(n16418) );
  INV_X1 U17022 ( .A(n13796), .ZN(n13797) );
  OAI22_X1 U17023 ( .A1(n16418), .A2(n20054), .B1(n13767), .B2(n13797), .ZN(
        n13798) );
  OAI21_X1 U17024 ( .B1(n13799), .B2(n13798), .A(n13802), .ZN(n13800) );
  OAI21_X1 U17025 ( .B1(n13802), .B2(n13801), .A(n13800), .ZN(P2_U3601) );
  XOR2_X1 U17026 ( .A(n13803), .B(n13789), .Z(n14524) );
  NOR2_X1 U17027 ( .A1(n16065), .A2(n13804), .ZN(n13805) );
  OR2_X1 U17028 ( .A1(n15916), .A2(n13805), .ZN(n16058) );
  OAI22_X1 U17029 ( .A1(n16058), .A2(n14312), .B1(n21347), .B2(n20211), .ZN(
        n13806) );
  AOI21_X1 U17030 ( .B1(n14524), .B2(n20207), .A(n13806), .ZN(n13807) );
  INV_X1 U17031 ( .A(n13807), .ZN(P1_U2862) );
  INV_X1 U17032 ( .A(n14524), .ZN(n13818) );
  INV_X1 U17033 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21219) );
  INV_X1 U17034 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20941) );
  INV_X1 U17035 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20935) );
  NOR2_X1 U17036 ( .A1(n20935), .A2(n21352), .ZN(n20178) );
  AND3_X1 U17037 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(n20178), .ZN(n20162) );
  NAND3_X1 U17038 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20162), .ZN(n13809) );
  INV_X1 U17039 ( .A(n13809), .ZN(n13808) );
  INV_X1 U17040 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21364) );
  OAI21_X1 U17041 ( .B1(n21219), .B2(n20129), .A(n21364), .ZN(n13815) );
  INV_X1 U17042 ( .A(n20161), .ZN(n13810) );
  NAND2_X1 U17043 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14050) );
  NOR2_X1 U17044 ( .A1(n13810), .A2(n13809), .ZN(n20140) );
  NAND3_X1 U17045 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n20140), .ZN(n20122) );
  NOR2_X1 U17046 ( .A1(n14050), .A2(n20122), .ZN(n14054) );
  NOR2_X1 U17047 ( .A1(n20160), .A2(n14054), .ZN(n15922) );
  OAI22_X1 U17048 ( .A1(n21347), .A2(n20201), .B1(n20174), .B2(n16058), .ZN(
        n13812) );
  NAND2_X1 U17049 ( .A1(n13811), .A2(n20161), .ZN(n20170) );
  AOI211_X1 U17050 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n13812), .B(n20153), .ZN(n13813) );
  OAI21_X1 U17051 ( .B1(n14522), .B2(n20184), .A(n13813), .ZN(n13814) );
  AOI21_X1 U17052 ( .B1(n13815), .B2(n15922), .A(n13814), .ZN(n13816) );
  OAI21_X1 U17053 ( .B1(n13818), .B2(n20133), .A(n13816), .ZN(P1_U2830) );
  AOI22_X1 U17054 ( .A1(n14375), .A2(n20270), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14374), .ZN(n13817) );
  OAI21_X1 U17055 ( .B1(n13818), .B2(n14382), .A(n13817), .ZN(P1_U2894) );
  XNOR2_X1 U17056 ( .A(n15938), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13819) );
  XNOR2_X1 U17057 ( .A(n13820), .B(n13819), .ZN(n16071) );
  NAND2_X1 U17058 ( .A1(n16071), .A2(n20298), .ZN(n13824) );
  INV_X1 U17059 ( .A(n20302), .ZN(n15956) );
  NAND2_X1 U17060 ( .A1(n20317), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16068) );
  OAI21_X1 U17061 ( .B1(n13821), .B2(n10664), .A(n16068), .ZN(n13822) );
  AOI21_X1 U17062 ( .B1(n15956), .B2(n20126), .A(n13822), .ZN(n13823) );
  OAI211_X1 U17063 ( .C1(n13826), .C2(n13825), .A(n13824), .B(n13823), .ZN(
        P1_U2990) );
  NAND2_X1 U17064 ( .A1(n19250), .A2(n15524), .ZN(n13832) );
  NOR2_X1 U17065 ( .A1(n13827), .A2(n13828), .ZN(n13829) );
  AOI22_X1 U17066 ( .A1(n10233), .A2(n15515), .B1(n13830), .B2(n13829), .ZN(
        n13831) );
  NAND2_X1 U17067 ( .A1(n13832), .A2(n13831), .ZN(n16419) );
  INV_X1 U17068 ( .A(n13833), .ZN(n13835) );
  AOI222_X1 U17069 ( .A1(n16419), .A2(n13836), .B1(n20072), .B2(n16465), .C1(
        n13835), .C2(n13834), .ZN(n13839) );
  NAND2_X1 U17070 ( .A1(n15527), .A2(n13837), .ZN(n13838) );
  OAI21_X1 U17071 ( .B1(n13839), .B2(n15527), .A(n13838), .ZN(P2_U3600) );
  INV_X1 U17072 ( .A(n13840), .ZN(n13843) );
  INV_X1 U17073 ( .A(n13841), .ZN(n13842) );
  NAND2_X1 U17074 ( .A1(n13843), .A2(n13842), .ZN(n13845) );
  INV_X1 U17075 ( .A(n15964), .ZN(n13847) );
  AOI22_X1 U17076 ( .A1(n14375), .A2(n20273), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14374), .ZN(n13846) );
  OAI21_X1 U17077 ( .B1(n13847), .B2(n14382), .A(n13846), .ZN(P1_U2893) );
  AND2_X1 U17078 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17060) );
  NAND3_X1 U17079 ( .A1(n13850), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13859) );
  INV_X1 U17080 ( .A(n13859), .ZN(n13849) );
  INV_X2 U17081 ( .A(n17293), .ZN(n15677) );
  OR3_X2 U17082 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18967), .A3(
        n18828), .ZN(n13966) );
  INV_X1 U17083 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17253) );
  INV_X4 U17084 ( .A(n9813), .ZN(n17328) );
  BUF_X2 U17085 ( .A(n15612), .Z(n17350) );
  AOI22_X1 U17086 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17087 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17351), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13853) );
  OAI211_X1 U17088 ( .C1(n17349), .C2(n17253), .A(n13854), .B(n13853), .ZN(
        n13865) );
  AOI22_X1 U17089 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n15618), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17323), .ZN(n13863) );
  AOI22_X1 U17090 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9810), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13862) );
  INV_X1 U17091 ( .A(n13870), .ZN(n13922) );
  INV_X2 U17092 ( .A(n13922), .ZN(n17242) );
  AOI22_X1 U17093 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17324), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17242), .ZN(n13861) );
  NAND2_X1 U17094 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13860) );
  NAND4_X1 U17095 ( .A1(n13863), .A2(n13862), .A3(n13861), .A4(n13860), .ZN(
        n13864) );
  INV_X1 U17096 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U17097 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13869) );
  OAI21_X1 U17098 ( .B1(n17144), .B2(n17206), .A(n13869), .ZN(n13877) );
  AOI22_X1 U17099 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17100 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13871) );
  OAI21_X1 U17101 ( .B1(n13901), .B2(n18415), .A(n13871), .ZN(n13875) );
  INV_X1 U17102 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17103 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17104 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17105 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13878) );
  OAI21_X1 U17106 ( .B1(n15538), .B2(n17221), .A(n13878), .ZN(n13888) );
  AOI22_X1 U17107 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13886) );
  INV_X1 U17108 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17348) );
  OAI22_X1 U17109 ( .A1(n13934), .A2(n17348), .B1(n13901), .B2(n18412), .ZN(
        n13884) );
  AOI22_X1 U17110 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17111 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17112 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13880) );
  NAND3_X1 U17113 ( .A1(n13882), .A2(n13881), .A3(n13880), .ZN(n13883) );
  AOI211_X1 U17114 ( .C1(n17352), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n13884), .B(n13883), .ZN(n13885) );
  OAI211_X1 U17115 ( .C1(n17293), .C2(n18689), .A(n13886), .B(n13885), .ZN(
        n13887) );
  AOI211_X4 U17116 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n13888), .B(n13887), .ZN(n16997) );
  INV_X1 U17117 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U17118 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13898) );
  INV_X1 U17119 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U17120 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U17121 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13889) );
  OAI211_X1 U17122 ( .C1(n17349), .C2(n13978), .A(n13890), .B(n13889), .ZN(
        n13896) );
  AOI22_X1 U17123 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17124 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17125 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U17126 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13891) );
  NAND4_X1 U17127 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n13895) );
  AOI211_X1 U17128 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13896), .B(n13895), .ZN(n13897) );
  OAI211_X1 U17129 ( .C1(n17293), .C2(n17175), .A(n13898), .B(n13897), .ZN(
        n18385) );
  AOI22_X1 U17130 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13899) );
  OAI21_X1 U17131 ( .B1(n17275), .B2(n14023), .A(n13899), .ZN(n13910) );
  AOI22_X1 U17132 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13908) );
  INV_X1 U17133 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13900) );
  INV_X1 U17134 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17317) );
  OAI22_X1 U17135 ( .A1(n17349), .A2(n13900), .B1(n13933), .B2(n17317), .ZN(
        n13906) );
  AOI22_X1 U17136 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17137 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17138 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13902) );
  NAND3_X1 U17139 ( .A1(n13904), .A2(n13903), .A3(n13902), .ZN(n13905) );
  AOI211_X1 U17140 ( .C1(n17352), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n13906), .B(n13905), .ZN(n13907) );
  OAI211_X1 U17141 ( .C1(n17339), .C2(n17389), .A(n13908), .B(n13907), .ZN(
        n13909) );
  AOI211_X4 U17142 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n13910), .B(n13909), .ZN(n15727) );
  INV_X1 U17143 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U17144 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13921) );
  INV_X1 U17145 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U17146 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17147 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U17148 ( .C1(n17349), .C2(n15531), .A(n13913), .B(n13912), .ZN(
        n13919) );
  AOI22_X1 U17149 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17150 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17151 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U17152 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13914) );
  NAND4_X1 U17153 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13918) );
  AOI211_X1 U17154 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13919), .B(n13918), .ZN(n13920) );
  NAND2_X1 U17155 ( .A1(n15727), .A2(n18393), .ZN(n15551) );
  AOI22_X1 U17156 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U17157 ( .B1(n9813), .B2(n17128), .A(n13923), .ZN(n13932) );
  INV_X1 U17158 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U17159 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13930) );
  INV_X1 U17160 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U17161 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U17162 ( .B1(n17339), .B2(n17370), .A(n13924), .ZN(n13928) );
  INV_X1 U17163 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U17164 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17165 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13925) );
  OAI211_X1 U17166 ( .C1(n17349), .C2(n17259), .A(n13926), .B(n13925), .ZN(
        n13927) );
  AOI211_X1 U17167 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n13928), .B(n13927), .ZN(n13929) );
  OAI211_X1 U17168 ( .C1(n17302), .C2(n17268), .A(n13930), .B(n13929), .ZN(
        n13931) );
  AOI211_X2 U17169 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n13932), .B(n13931), .ZN(n15719) );
  AOI22_X1 U17170 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13944) );
  INV_X1 U17171 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U17172 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17173 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13935) );
  OAI211_X1 U17174 ( .C1(n17349), .C2(n17274), .A(n13936), .B(n13935), .ZN(
        n13942) );
  AOI22_X1 U17175 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17176 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17177 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U17178 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13937) );
  NAND4_X1 U17179 ( .A1(n13940), .A2(n13939), .A3(n13938), .A4(n13937), .ZN(
        n13941) );
  AOI211_X1 U17180 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n13942), .B(n13941), .ZN(n13943) );
  OAI211_X1 U17181 ( .C1(n17302), .C2(n17284), .A(n13944), .B(n13943), .ZN(
        n18389) );
  NAND2_X1 U17182 ( .A1(n15719), .A2(n18389), .ZN(n18809) );
  OAI21_X1 U17183 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18822), .A(
        n15569), .ZN(n15722) );
  INV_X1 U17184 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U17185 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18373), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18974), .ZN(n13951) );
  INV_X1 U17186 ( .A(n15569), .ZN(n13945) );
  NAND2_X1 U17187 ( .A1(n15570), .A2(n13945), .ZN(n13946) );
  OAI21_X1 U17188 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n13850), .A(
        n13946), .ZN(n13950) );
  NAND2_X1 U17189 ( .A1(n13951), .A2(n13950), .ZN(n13947) );
  OAI21_X1 U17190 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18974), .A(
        n13947), .ZN(n13948) );
  OAI22_X1 U17191 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18369), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13948), .ZN(n13952) );
  NOR2_X1 U17192 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18369), .ZN(
        n13949) );
  NAND2_X1 U17193 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13948), .ZN(
        n13953) );
  AOI22_X1 U17194 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13952), .B1(
        n13949), .B2(n13953), .ZN(n13956) );
  NAND2_X1 U17195 ( .A1(n15570), .A2(n13956), .ZN(n13958) );
  XOR2_X1 U17196 ( .A(n13951), .B(n13950), .Z(n13957) );
  AOI21_X1 U17197 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13953), .A(
        n13952), .ZN(n13954) );
  INV_X1 U17198 ( .A(n15567), .ZN(n13955) );
  INV_X1 U17199 ( .A(n18803), .ZN(n15582) );
  INV_X1 U17200 ( .A(n18393), .ZN(n15550) );
  INV_X1 U17201 ( .A(n15719), .ZN(n18397) );
  NAND2_X1 U17202 ( .A1(n15550), .A2(n18397), .ZN(n15573) );
  NOR3_X1 U17203 ( .A1(n18400), .A2(n18389), .A3(n15562), .ZN(n13959) );
  NAND2_X1 U17204 ( .A1(n17445), .A2(n17399), .ZN(n17393) );
  INV_X2 U17205 ( .A(n17396), .ZN(n17390) );
  INV_X1 U17206 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16750) );
  INV_X1 U17207 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17061) );
  INV_X1 U17208 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16790) );
  INV_X1 U17209 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17202) );
  INV_X1 U17210 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n13961) );
  INV_X1 U17211 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17027) );
  NAND2_X1 U17212 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17385) );
  NOR2_X1 U17213 ( .A1(n17027), .A2(n17385), .ZN(n17376) );
  NAND3_X1 U17214 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17376), .ZN(n17371) );
  NAND4_X1 U17215 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n13960) );
  NOR4_X1 U17216 ( .A1(n13961), .A2(n16910), .A3(n17371), .A4(n13960), .ZN(
        n13962) );
  NAND4_X1 U17217 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n13962), .ZN(n17234) );
  NAND3_X1 U17218 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .ZN(n17201) );
  NOR2_X1 U17219 ( .A1(n17234), .A2(n17201), .ZN(n17217) );
  NAND3_X1 U17220 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17399), .A3(n17217), 
        .ZN(n17189) );
  NOR2_X1 U17221 ( .A1(n17202), .A2(n17189), .ZN(n17187) );
  NAND2_X1 U17222 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17187), .ZN(n17186) );
  NOR2_X1 U17223 ( .A1(n18400), .A2(n17186), .ZN(n17171) );
  NAND2_X1 U17224 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17171), .ZN(n17158) );
  NAND2_X1 U17225 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17126), .ZN(n17120) );
  NAND2_X1 U17226 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17125), .ZN(n17110) );
  NAND2_X1 U17227 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17114), .ZN(n17104) );
  NAND2_X1 U17228 ( .A1(n17390), .A2(n17104), .ZN(n13963) );
  OAI21_X1 U17229 ( .B1(n17060), .B2(n17393), .A(n13963), .ZN(n17099) );
  INV_X1 U17230 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U17231 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13964) );
  OAI21_X1 U17232 ( .B1(n13879), .B2(n17145), .A(n13964), .ZN(n13975) );
  INV_X1 U17233 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U17234 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13973) );
  INV_X1 U17235 ( .A(n13965), .ZN(n17222) );
  INV_X1 U17236 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17143) );
  OAI22_X1 U17237 ( .A1(n17222), .A2(n15531), .B1(n13966), .B2(n17143), .ZN(
        n13971) );
  AOI22_X1 U17238 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13969) );
  AOI22_X1 U17239 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13968) );
  AOI22_X1 U17240 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13967) );
  NAND3_X1 U17241 ( .A1(n13969), .A2(n13968), .A3(n13967), .ZN(n13970) );
  AOI211_X1 U17242 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n13971), .B(n13970), .ZN(n13972) );
  OAI211_X1 U17243 ( .C1(n13933), .C2(n17373), .A(n13973), .B(n13972), .ZN(
        n13974) );
  AOI211_X1 U17244 ( .C1(n17350), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13975), .B(n13974), .ZN(n14038) );
  INV_X1 U17245 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U17246 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13976) );
  OAI21_X1 U17247 ( .B1(n17302), .B2(n17174), .A(n13976), .ZN(n13986) );
  AOI22_X1 U17248 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U17249 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17241), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13977) );
  OAI21_X1 U17250 ( .B1(n17222), .B2(n13978), .A(n13977), .ZN(n13982) );
  AOI22_X1 U17251 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U17252 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13979) );
  OAI211_X1 U17253 ( .C1(n17349), .C2(n17175), .A(n13980), .B(n13979), .ZN(
        n13981) );
  AOI211_X1 U17254 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n13982), .B(n13981), .ZN(n13983) );
  OAI211_X1 U17255 ( .C1(n13933), .C2(n17383), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI211_X1 U17256 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n13986), .B(n13985), .ZN(n17106) );
  INV_X1 U17257 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15610) );
  AOI22_X1 U17258 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13987) );
  OAI21_X1 U17259 ( .B1(n9813), .B2(n15610), .A(n13987), .ZN(n13996) );
  AOI22_X1 U17260 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13994) );
  INV_X1 U17261 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U17262 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17241), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13988) );
  OAI21_X1 U17263 ( .B1(n17144), .B2(n17332), .A(n13988), .ZN(n13992) );
  INV_X1 U17264 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18693) );
  AOI22_X1 U17265 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17351), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17266 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13989) );
  OAI211_X1 U17267 ( .C1(n17349), .C2(n18693), .A(n13990), .B(n13989), .ZN(
        n13991) );
  AOI211_X1 U17268 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n13992), .B(n13991), .ZN(n13993) );
  OAI211_X1 U17269 ( .C1(n17293), .C2(n18415), .A(n13994), .B(n13993), .ZN(
        n13995) );
  AOI211_X1 U17270 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n13996), .B(n13995), .ZN(n17116) );
  INV_X1 U17271 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U17272 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17273 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13997) );
  OAI21_X1 U17274 ( .B1(n13879), .B2(n17221), .A(n13997), .ZN(n14004) );
  INV_X1 U17275 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15676) );
  OAI22_X1 U17276 ( .A1(n17302), .A2(n15676), .B1(n17293), .B2(n18412), .ZN(
        n13998) );
  AOI21_X1 U17277 ( .B1(n17335), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n13998), .ZN(n14002) );
  AOI22_X1 U17278 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17279 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U17280 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13999) );
  NAND4_X1 U17281 ( .A1(n14002), .A2(n14001), .A3(n14000), .A4(n13999), .ZN(
        n14003) );
  AOI211_X1 U17282 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n14004), .B(n14003), .ZN(n14005) );
  OAI211_X1 U17283 ( .C1(n13933), .C2(n17361), .A(n14006), .B(n14005), .ZN(
        n17122) );
  AOI22_X1 U17284 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14016) );
  INV_X1 U17285 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U17286 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n9810), .ZN(n14007) );
  OAI21_X1 U17287 ( .B1(n13934), .B2(n17240), .A(n14007), .ZN(n14014) );
  AOI22_X1 U17288 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17241), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14012) );
  INV_X1 U17289 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U17290 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17324), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n15633), .ZN(n14009) );
  AOI22_X1 U17291 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17323), .ZN(n14008) );
  OAI211_X1 U17292 ( .C1(n17090), .C2(n13966), .A(n14009), .B(n14008), .ZN(
        n14010) );
  AOI21_X1 U17293 ( .B1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17335), .A(
        n14010), .ZN(n14011) );
  OAI211_X1 U17294 ( .C1(n17367), .C2(n17293), .A(n14012), .B(n14011), .ZN(
        n14013) );
  AOI211_X1 U17295 ( .C1(n17328), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n14014), .B(n14013), .ZN(n14015) );
  OAI211_X1 U17296 ( .C1(n17302), .C2(n17253), .A(n14016), .B(n14015), .ZN(
        n17123) );
  NAND2_X1 U17297 ( .A1(n17122), .A2(n17123), .ZN(n17121) );
  NOR2_X1 U17298 ( .A1(n17116), .A2(n17121), .ZN(n17115) );
  AOI22_X1 U17299 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U17300 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14017) );
  OAI21_X1 U17301 ( .B1(n13933), .B2(n17389), .A(n14017), .ZN(n14025) );
  AOI22_X1 U17302 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14022) );
  INV_X1 U17303 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U17304 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17305 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14018) );
  OAI211_X1 U17306 ( .C1(n13901), .C2(n17191), .A(n14019), .B(n14018), .ZN(
        n14020) );
  AOI21_X1 U17307 ( .B1(n17335), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n14020), .ZN(n14021) );
  OAI211_X1 U17308 ( .C1(n13868), .C2(n14023), .A(n14022), .B(n14021), .ZN(
        n14024) );
  AOI211_X1 U17309 ( .C1(n17351), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n14025), .B(n14024), .ZN(n14026) );
  OAI211_X1 U17310 ( .C1(n15538), .C2(n17317), .A(n14027), .B(n14026), .ZN(
        n17112) );
  NAND2_X1 U17311 ( .A1(n17115), .A2(n17112), .ZN(n17111) );
  NOR2_X1 U17312 ( .A1(n17106), .A2(n17111), .ZN(n17105) );
  AOI22_X1 U17313 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14037) );
  INV_X1 U17314 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U17315 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17351), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17316 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14028) );
  OAI211_X1 U17317 ( .C1(n17349), .C2(n15598), .A(n14029), .B(n14028), .ZN(
        n14035) );
  AOI22_X1 U17318 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17319 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17320 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U17321 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14030) );
  NAND4_X1 U17322 ( .A1(n14033), .A2(n14032), .A3(n14031), .A4(n14030), .ZN(
        n14034) );
  AOI211_X1 U17323 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n14035), .B(n14034), .ZN(n14036) );
  OAI211_X1 U17324 ( .C1(n13933), .C2(n17381), .A(n14037), .B(n14036), .ZN(
        n17102) );
  NAND2_X1 U17325 ( .A1(n17105), .A2(n17102), .ZN(n17101) );
  NOR2_X1 U17326 ( .A1(n14038), .A2(n17101), .ZN(n17096) );
  AOI21_X1 U17327 ( .B1(n14038), .B2(n17101), .A(n17096), .ZN(n17415) );
  AOI22_X1 U17328 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17099), .B1(n17415), 
        .B2(n17396), .ZN(n14041) );
  INV_X1 U17329 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14039) );
  INV_X1 U17330 ( .A(n17104), .ZN(n17109) );
  NAND3_X1 U17331 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14039), .A3(n17109), 
        .ZN(n14040) );
  NAND2_X1 U17332 ( .A1(n14041), .A2(n14040), .ZN(P3_U2675) );
  AOI22_X1 U17333 ( .A1(n14361), .A2(DATAI_30_), .B1(n14374), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14046) );
  AND2_X1 U17334 ( .A1(n9845), .A2(n10695), .ZN(n14044) );
  AOI22_X1 U17335 ( .A1(n14364), .A2(n20282), .B1(n14362), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14045) );
  OAI211_X1 U17336 ( .C1(n14062), .C2(n14382), .A(n14046), .B(n14045), .ZN(
        P1_U2874) );
  OAI22_X1 U17337 ( .A1(n14048), .A2(n20172), .B1(n20184), .B2(n14047), .ZN(
        n14049) );
  INV_X1 U17338 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21128) );
  INV_X1 U17339 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21376) );
  NAND2_X1 U17340 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15921), .ZN(n14252) );
  NAND3_X1 U17341 ( .A1(n15906), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_13__SCAN_IN), .ZN(n15905) );
  NAND2_X1 U17342 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15886) );
  NAND2_X1 U17343 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15882), .ZN(n14226) );
  NAND3_X1 U17344 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n14171) );
  INV_X1 U17345 ( .A(n14171), .ZN(n14051) );
  AND2_X1 U17346 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U17347 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14057) );
  AND2_X1 U17348 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14053) );
  NAND2_X1 U17349 ( .A1(n14151), .A2(n14053), .ZN(n14122) );
  INV_X1 U17350 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21249) );
  NAND2_X1 U17351 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14109) );
  INV_X1 U17352 ( .A(n14109), .ZN(n14059) );
  NAND2_X1 U17353 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14056) );
  NAND2_X1 U17354 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14055) );
  NAND3_X1 U17355 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n14054), .ZN(n14238) );
  NOR2_X1 U17356 ( .A1(n14055), .A2(n14238), .ZN(n15887) );
  NAND4_X1 U17357 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n15887), .ZN(n14225) );
  NOR3_X1 U17358 ( .A1(n21128), .A2(n14056), .A3(n14225), .ZN(n14202) );
  AND2_X1 U17359 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14187) );
  NAND3_X1 U17360 ( .A1(n14202), .A2(P1_REIP_REG_23__SCAN_IN), .A3(n14187), 
        .ZN(n14172) );
  INV_X1 U17361 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20962) );
  NOR3_X1 U17362 ( .A1(n14172), .A2(n14057), .A3(n20962), .ZN(n14144) );
  NAND3_X1 U17363 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14144), .ZN(n14115) );
  INV_X1 U17364 ( .A(n14115), .ZN(n14058) );
  NAND2_X1 U17365 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  NAND2_X1 U17366 ( .A1(n20123), .A2(n14060), .ZN(n14108) );
  INV_X1 U17367 ( .A(n14108), .ZN(n14061) );
  AOI21_X1 U17368 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14063), .ZN(n14064) );
  OAI21_X1 U17369 ( .B1(n20302), .B2(n14065), .A(n14064), .ZN(n14066) );
  OAI21_X1 U17370 ( .B1(n14068), .B2(n20108), .A(n14067), .ZN(P1_U2968) );
  NAND2_X1 U17371 ( .A1(n14069), .A2(n20197), .ZN(n14078) );
  AOI21_X1 U17372 ( .B1(n20178), .B2(n20161), .A(n20160), .ZN(n20185) );
  INV_X1 U17373 ( .A(n20179), .ZN(n14070) );
  OAI21_X1 U17374 ( .B1(n14070), .B2(n21352), .A(n20935), .ZN(n14076) );
  NOR2_X1 U17375 ( .A1(n20174), .A2(n20329), .ZN(n14075) );
  INV_X1 U17376 ( .A(n14071), .ZN(n14072) );
  AOI22_X1 U17377 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20190), .B1(
        n20191), .B2(n14072), .ZN(n14073) );
  OAI21_X1 U17378 ( .B1(n20201), .B2(n21243), .A(n14073), .ZN(n14074) );
  AOI211_X1 U17379 ( .C1(n20185), .C2(n14076), .A(n14075), .B(n14074), .ZN(
        n14077) );
  OAI211_X1 U17380 ( .C1(n20187), .C2(n20720), .A(n14078), .B(n14077), .ZN(
        P1_U2838) );
  INV_X1 U17381 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14998) );
  NAND2_X1 U17382 ( .A1(n14680), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U17383 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14079) );
  AOI21_X1 U17384 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14081), .ZN(n14741) );
  INV_X1 U17385 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15004) );
  NAND2_X1 U17386 ( .A1(n14680), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n14083) );
  NAND2_X1 U17387 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14082) );
  AOI21_X1 U17388 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14084), .ZN(n14735) );
  INV_X1 U17389 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14728) );
  NAND2_X1 U17390 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14086) );
  AOI22_X1 U17391 ( .A1(n14680), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n14085) );
  INV_X1 U17392 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n14089) );
  NAND2_X1 U17393 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14088) );
  AOI22_X1 U17394 ( .A1(n14680), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n14087) );
  INV_X1 U17395 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U17396 ( .A1(n14680), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14091) );
  NAND2_X1 U17397 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14090) );
  AOI21_X1 U17398 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14093), .ZN(n14709) );
  INV_X1 U17399 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U17400 ( .A1(n14680), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U17401 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14094) );
  AOI21_X1 U17402 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14096), .ZN(n14701) );
  INV_X1 U17403 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U17404 ( .A1(n14685), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14098) );
  AOI22_X1 U17405 ( .A1(n14680), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n14097) );
  INV_X1 U17406 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U17407 ( .A1(n14680), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14101) );
  NAND2_X1 U17408 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14100) );
  AOI21_X1 U17409 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14102), .ZN(n14679) );
  NOR2_X1 U17410 ( .A1(n16120), .A2(n14776), .ZN(n14103) );
  AOI21_X1 U17411 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14776), .A(n14103), .ZN(
        n14104) );
  OAI21_X1 U17412 ( .B1(n14105), .B2(n14779), .A(n14104), .ZN(P2_U2857) );
  INV_X1 U17413 ( .A(n14106), .ZN(n14113) );
  INV_X1 U17414 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U17415 ( .A1(n20177), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20190), .ZN(n14107) );
  OAI21_X1 U17416 ( .B1(n14108), .B2(n20971), .A(n14107), .ZN(n14111) );
  NOR3_X1 U17417 ( .A1(n14122), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14109), 
        .ZN(n14110) );
  AOI211_X1 U17418 ( .C1(n14265), .C2(n20186), .A(n14111), .B(n14110), .ZN(
        n14112) );
  OAI21_X1 U17419 ( .B1(n14113), .B2(n20133), .A(n14112), .ZN(P1_U2809) );
  NAND2_X1 U17420 ( .A1(n14390), .A2(n20155), .ZN(n14121) );
  INV_X1 U17421 ( .A(n14114), .ZN(n14540) );
  NAND2_X1 U17422 ( .A1(n20123), .A2(n14115), .ZN(n14132) );
  OAI22_X1 U17423 ( .A1(n14116), .A2(n20172), .B1(n21191), .B2(n20201), .ZN(
        n14117) );
  AOI21_X1 U17424 ( .B1(n20191), .B2(n14386), .A(n14117), .ZN(n14118) );
  OAI21_X1 U17425 ( .B1(n14132), .B2(n21249), .A(n14118), .ZN(n14119) );
  AOI21_X1 U17426 ( .B1(n14540), .B2(n20186), .A(n14119), .ZN(n14120) );
  OAI211_X1 U17427 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14122), .A(n14121), 
        .B(n14120), .ZN(P1_U2811) );
  OAI21_X2 U17428 ( .B1(n14123), .B2(n14125), .A(n14124), .ZN(n14398) );
  OR2_X1 U17429 ( .A1(n14143), .A2(n14126), .ZN(n14127) );
  NAND2_X1 U17430 ( .A1(n14128), .A2(n14127), .ZN(n14551) );
  INV_X1 U17431 ( .A(n14551), .ZN(n14134) );
  INV_X1 U17432 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21220) );
  OAI22_X1 U17433 ( .A1(n14129), .A2(n20172), .B1(n20184), .B2(n14400), .ZN(
        n14130) );
  AOI21_X1 U17434 ( .B1(n20177), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14130), .ZN(
        n14131) );
  OAI21_X1 U17435 ( .B1(n14132), .B2(n21220), .A(n14131), .ZN(n14133) );
  AOI21_X1 U17436 ( .B1(n14134), .B2(n20186), .A(n14133), .ZN(n14136) );
  NAND3_X1 U17437 ( .A1(n14151), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n21220), 
        .ZN(n14135) );
  OAI211_X1 U17438 ( .C1(n14398), .C2(n20133), .A(n14136), .B(n14135), .ZN(
        P1_U2812) );
  INV_X1 U17439 ( .A(n14123), .ZN(n14138) );
  INV_X1 U17440 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21384) );
  INV_X1 U17441 ( .A(n14139), .ZN(n14156) );
  INV_X1 U17442 ( .A(n14140), .ZN(n14141) );
  AOI21_X1 U17443 ( .B1(n14166), .B2(n14156), .A(n14141), .ZN(n14142) );
  OR2_X1 U17444 ( .A1(n14143), .A2(n14142), .ZN(n14559) );
  NOR2_X1 U17445 ( .A1(n14144), .A2(n20160), .ZN(n14162) );
  NAND2_X1 U17446 ( .A1(n14162), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14149) );
  INV_X1 U17447 ( .A(n14145), .ZN(n14410) );
  OAI22_X1 U17448 ( .A1(n14146), .A2(n20172), .B1(n20184), .B2(n14410), .ZN(
        n14147) );
  AOI21_X1 U17449 ( .B1(n20177), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14147), .ZN(
        n14148) );
  OAI211_X1 U17450 ( .C1(n14559), .C2(n20174), .A(n14149), .B(n14148), .ZN(
        n14150) );
  AOI21_X1 U17451 ( .B1(n14151), .B2(n21384), .A(n14150), .ZN(n14152) );
  OAI21_X1 U17452 ( .B1(n14408), .B2(n20133), .A(n14152), .ZN(P1_U2813) );
  INV_X1 U17453 ( .A(n14154), .ZN(n14155) );
  AOI21_X1 U17454 ( .B1(n10133), .B2(n14155), .A(n10488), .ZN(n14420) );
  INV_X1 U17455 ( .A(n14420), .ZN(n14328) );
  XNOR2_X1 U17456 ( .A(n14166), .B(n14156), .ZN(n14570) );
  OAI22_X1 U17457 ( .A1(n14157), .A2(n20172), .B1(n20184), .B2(n14418), .ZN(
        n14158) );
  AOI21_X1 U17458 ( .B1(n20177), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14158), .ZN(
        n14159) );
  OAI21_X1 U17459 ( .B1(n14570), .B2(n20174), .A(n14159), .ZN(n14161) );
  INV_X1 U17460 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21120) );
  NOR3_X1 U17461 ( .A1(n9937), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n21120), .ZN(
        n14160) );
  AOI211_X1 U17462 ( .C1(n14162), .C2(P1_REIP_REG_26__SCAN_IN), .A(n14161), 
        .B(n14160), .ZN(n14163) );
  OAI21_X1 U17463 ( .B1(n14328), .B2(n20133), .A(n14163), .ZN(P1_U2814) );
  AOI21_X1 U17464 ( .B1(n14165), .B2(n14164), .A(n14154), .ZN(n14431) );
  INV_X1 U17465 ( .A(n14431), .ZN(n14331) );
  AOI21_X1 U17466 ( .B1(n14167), .B2(n9882), .A(n14166), .ZN(n14577) );
  AOI22_X1 U17467 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20190), .B1(
        n20191), .B2(n14427), .ZN(n14168) );
  OAI21_X1 U17468 ( .B1(n20201), .B2(n21159), .A(n14168), .ZN(n14170) );
  NOR2_X1 U17469 ( .A1(n9937), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14169) );
  AOI211_X1 U17470 ( .C1(n14577), .C2(n20186), .A(n14170), .B(n14169), .ZN(
        n14174) );
  INV_X1 U17471 ( .A(n14222), .ZN(n14209) );
  NOR3_X1 U17472 ( .A1(n14209), .A2(n14171), .A3(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14184) );
  AND2_X1 U17473 ( .A1(n14172), .A2(n20123), .ZN(n14188) );
  OAI21_X1 U17474 ( .B1(n14184), .B2(n14188), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14173) );
  OAI211_X1 U17475 ( .C1(n14331), .C2(n20133), .A(n14174), .B(n14173), .ZN(
        P1_U2815) );
  INV_X1 U17476 ( .A(n14164), .ZN(n14176) );
  AOI21_X1 U17477 ( .B1(n14177), .B2(n14175), .A(n14176), .ZN(n14441) );
  INV_X1 U17478 ( .A(n14441), .ZN(n14335) );
  NAND2_X1 U17479 ( .A1(n9893), .A2(n14178), .ZN(n14179) );
  NAND2_X1 U17480 ( .A1(n9882), .A2(n14179), .ZN(n14582) );
  INV_X1 U17481 ( .A(n14180), .ZN(n14439) );
  OAI22_X1 U17482 ( .A1(n14181), .A2(n20172), .B1(n20184), .B2(n14439), .ZN(
        n14182) );
  AOI21_X1 U17483 ( .B1(n20177), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14182), .ZN(
        n14183) );
  OAI21_X1 U17484 ( .B1(n14582), .B2(n20174), .A(n14183), .ZN(n14185) );
  AOI211_X1 U17485 ( .C1(n14188), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14185), 
        .B(n14184), .ZN(n14186) );
  OAI21_X1 U17486 ( .B1(n14335), .B2(n20133), .A(n14186), .ZN(P1_U2816) );
  AOI21_X1 U17487 ( .B1(n14222), .B2(n14187), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14198) );
  INV_X1 U17488 ( .A(n14188), .ZN(n14197) );
  INV_X1 U17489 ( .A(n14189), .ZN(n14200) );
  OAI21_X1 U17490 ( .B1(n14200), .B2(n9956), .A(n14175), .ZN(n14339) );
  INV_X1 U17491 ( .A(n14339), .ZN(n14447) );
  NAND2_X1 U17492 ( .A1(n14447), .A2(n20155), .ZN(n14196) );
  INV_X1 U17493 ( .A(n14190), .ZN(n14445) );
  OAI22_X1 U17494 ( .A1(n14191), .A2(n20172), .B1(n20184), .B2(n14445), .ZN(
        n14194) );
  OAI21_X1 U17495 ( .B1(n14203), .B2(n14192), .A(n9893), .ZN(n14593) );
  NOR2_X1 U17496 ( .A1(n14593), .A2(n20174), .ZN(n14193) );
  AOI211_X1 U17497 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20177), .A(n14194), .B(
        n14193), .ZN(n14195) );
  OAI211_X1 U17498 ( .C1(n14198), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        P1_U2817) );
  INV_X1 U17499 ( .A(n14199), .ZN(n14201) );
  AOI21_X1 U17500 ( .B1(n14201), .B2(n9860), .A(n14200), .ZN(n14456) );
  INV_X1 U17501 ( .A(n14456), .ZN(n14343) );
  OR2_X1 U17502 ( .A1(n14202), .A2(n20160), .ZN(n15864) );
  INV_X1 U17503 ( .A(n15864), .ZN(n14212) );
  INV_X1 U17504 ( .A(n14203), .ZN(n14204) );
  OAI21_X1 U17505 ( .B1(n14217), .B2(n14205), .A(n14204), .ZN(n15987) );
  AOI22_X1 U17506 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20190), .B1(
        n20191), .B2(n14452), .ZN(n14207) );
  NAND2_X1 U17507 ( .A1(n20177), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14206) );
  OAI211_X1 U17508 ( .C1(n15987), .C2(n20174), .A(n14207), .B(n14206), .ZN(
        n14211) );
  XNOR2_X1 U17509 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14208) );
  NOR2_X1 U17510 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  AOI211_X1 U17511 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14212), .A(n14211), 
        .B(n14210), .ZN(n14213) );
  OAI21_X1 U17512 ( .B1(n14343), .B2(n20133), .A(n14213), .ZN(P1_U2818) );
  OAI21_X1 U17513 ( .B1(n9891), .B2(n14214), .A(n9860), .ZN(n14464) );
  INV_X1 U17514 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21273) );
  INV_X1 U17515 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14215) );
  OAI22_X1 U17516 ( .A1(n14466), .A2(n20184), .B1(n20172), .B2(n14215), .ZN(
        n14216) );
  AOI21_X1 U17517 ( .B1(n20177), .B2(P1_EBX_REG_21__SCAN_IN), .A(n14216), .ZN(
        n14220) );
  AOI21_X1 U17518 ( .B1(n14218), .B2(n14276), .A(n14217), .ZN(n15833) );
  NAND2_X1 U17519 ( .A1(n15833), .A2(n20186), .ZN(n14219) );
  OAI211_X1 U17520 ( .C1(n15864), .C2(n21273), .A(n14220), .B(n14219), .ZN(
        n14221) );
  AOI21_X1 U17521 ( .B1(n14222), .B2(n21273), .A(n14221), .ZN(n14223) );
  OAI21_X1 U17522 ( .B1(n14464), .B2(n20133), .A(n14223), .ZN(P1_U2819) );
  OAI21_X1 U17523 ( .B1(n11194), .B2(n9955), .A(n14224), .ZN(n14473) );
  INV_X1 U17524 ( .A(n15861), .ZN(n14228) );
  AND2_X1 U17525 ( .A1(n20123), .A2(n14225), .ZN(n15881) );
  NOR2_X1 U17526 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14226), .ZN(n15873) );
  NOR2_X1 U17527 ( .A1(n15881), .A2(n15873), .ZN(n14227) );
  MUX2_X1 U17528 ( .A(n14228), .B(n14227), .S(P1_REIP_REG_19__SCAN_IN), .Z(
        n14235) );
  NAND2_X1 U17529 ( .A1(n14285), .A2(n14229), .ZN(n14230) );
  NAND2_X1 U17530 ( .A1(n14274), .A2(n14230), .ZN(n14279) );
  INV_X1 U17531 ( .A(n14279), .ZN(n15996) );
  AOI22_X1 U17532 ( .A1(n14474), .A2(n20191), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n20177), .ZN(n14231) );
  OAI211_X1 U17533 ( .C1(n20172), .C2(n14232), .A(n14231), .B(n20170), .ZN(
        n14233) );
  AOI21_X1 U17534 ( .B1(n15996), .B2(n20186), .A(n14233), .ZN(n14234) );
  OAI211_X1 U17535 ( .C1(n14473), .C2(n20133), .A(n14235), .B(n14234), .ZN(
        P1_U2821) );
  AOI21_X1 U17536 ( .B1(n14237), .B2(n14236), .A(n9859), .ZN(n14512) );
  INV_X1 U17537 ( .A(n14512), .ZN(n14377) );
  INV_X1 U17538 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21363) );
  NAND2_X1 U17539 ( .A1(n20123), .A2(n14238), .ZN(n14251) );
  AOI21_X1 U17540 ( .B1(n10425), .B2(n14248), .A(n14239), .ZN(n14240) );
  NOR2_X1 U17541 ( .A1(n14240), .A2(n10428), .ZN(n16027) );
  AOI22_X1 U17542 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20177), .B1(n20186), 
        .B2(n16027), .ZN(n14241) );
  OAI21_X1 U17543 ( .B1(n21363), .B2(n14251), .A(n14241), .ZN(n14244) );
  AOI21_X1 U17544 ( .B1(n20190), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20153), .ZN(n14242) );
  OAI21_X1 U17545 ( .B1(n20184), .B2(n14510), .A(n14242), .ZN(n14243) );
  AOI211_X1 U17546 ( .C1(n15906), .C2(n21363), .A(n14244), .B(n14243), .ZN(
        n14245) );
  OAI21_X1 U17547 ( .B1(n14377), .B2(n20133), .A(n14245), .ZN(P1_U2827) );
  OAI21_X1 U17548 ( .B1(n14246), .B2(n14247), .A(n14236), .ZN(n15954) );
  XNOR2_X1 U17549 ( .A(n15918), .B(n14248), .ZN(n16036) );
  AOI22_X1 U17550 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(n20177), .B1(n20186), 
        .B2(n16036), .ZN(n14249) );
  OAI211_X1 U17551 ( .C1(n20172), .C2(n14250), .A(n14249), .B(n20170), .ZN(
        n14254) );
  AOI21_X1 U17552 ( .B1(n21376), .B2(n14252), .A(n14251), .ZN(n14253) );
  AOI211_X1 U17553 ( .C1(n15955), .C2(n20191), .A(n14254), .B(n14253), .ZN(
        n14255) );
  OAI21_X1 U17554 ( .B1(n15954), .B2(n20133), .A(n14255), .ZN(P1_U2828) );
  INV_X1 U17555 ( .A(n20187), .ZN(n14261) );
  NAND2_X1 U17556 ( .A1(n20123), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U17557 ( .A1(n20172), .A2(n20184), .ZN(n14256) );
  AOI22_X1 U17558 ( .A1(n20177), .A2(P1_EBX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14256), .ZN(n14257) );
  OAI211_X1 U17559 ( .C1(n20174), .C2(n14259), .A(n14258), .B(n14257), .ZN(
        n14260) );
  AOI21_X1 U17560 ( .B1(n10883), .B2(n14261), .A(n14260), .ZN(n14262) );
  OAI21_X1 U17561 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(P1_U2840) );
  INV_X1 U17562 ( .A(n14265), .ZN(n14267) );
  INV_X1 U17563 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14266) );
  OAI22_X1 U17564 ( .A1(n14267), .A2(n14312), .B1(n20211), .B2(n14266), .ZN(
        P1_U2841) );
  INV_X1 U17565 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14268) );
  OAI222_X1 U17566 ( .A1(n14398), .A2(n14318), .B1(n14268), .B2(n20211), .C1(
        n14551), .C2(n14312), .ZN(P1_U2844) );
  INV_X1 U17567 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21349) );
  OAI222_X1 U17568 ( .A1(n14408), .A2(n14318), .B1(n21349), .B2(n20211), .C1(
        n14559), .C2(n14312), .ZN(P1_U2845) );
  OAI222_X1 U17569 ( .A1(n14328), .A2(n14318), .B1(n21132), .B2(n20211), .C1(
        n14312), .C2(n14570), .ZN(P1_U2846) );
  INV_X1 U17570 ( .A(n14577), .ZN(n14269) );
  OAI222_X1 U17571 ( .A1(n14318), .A2(n14331), .B1(n21159), .B2(n20211), .C1(
        n14269), .C2(n14312), .ZN(P1_U2847) );
  INV_X1 U17572 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21228) );
  OAI222_X1 U17573 ( .A1(n14318), .A2(n14335), .B1(n21228), .B2(n20211), .C1(
        n14582), .C2(n14312), .ZN(P1_U2848) );
  OAI222_X1 U17574 ( .A1(n14339), .A2(n14318), .B1(n21229), .B2(n20211), .C1(
        n14593), .C2(n14312), .ZN(P1_U2849) );
  INV_X1 U17575 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21339) );
  OAI222_X1 U17576 ( .A1(n15987), .A2(n14312), .B1(n21339), .B2(n20211), .C1(
        n14343), .C2(n14318), .ZN(P1_U2850) );
  AOI22_X1 U17577 ( .A1(n15833), .A2(n20206), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14316), .ZN(n14270) );
  OAI21_X1 U17578 ( .B1(n14464), .B2(n14318), .A(n14270), .ZN(P1_U2851) );
  AND2_X1 U17579 ( .A1(n14224), .A2(n14271), .ZN(n14272) );
  OR2_X1 U17580 ( .A1(n14272), .A2(n9891), .ZN(n15860) );
  NAND2_X1 U17581 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  NAND2_X1 U17582 ( .A1(n14276), .A2(n14275), .ZN(n15862) );
  OAI22_X1 U17583 ( .A1(n15862), .A2(n14312), .B1(n21353), .B2(n20211), .ZN(
        n14277) );
  INV_X1 U17584 ( .A(n14277), .ZN(n14278) );
  OAI21_X1 U17585 ( .B1(n15860), .B2(n14318), .A(n14278), .ZN(P1_U2852) );
  INV_X1 U17586 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14280) );
  OAI222_X1 U17587 ( .A1(n14473), .A2(n14318), .B1(n14280), .B2(n20211), .C1(
        n14312), .C2(n14279), .ZN(P1_U2853) );
  OR2_X1 U17588 ( .A1(n9890), .A2(n14281), .ZN(n14282) );
  AND2_X1 U17589 ( .A1(n10127), .A2(n14282), .ZN(n15875) );
  INV_X1 U17590 ( .A(n15875), .ZN(n14356) );
  OR2_X1 U17591 ( .A1(n9931), .A2(n14283), .ZN(n14284) );
  NAND2_X1 U17592 ( .A1(n14285), .A2(n14284), .ZN(n16003) );
  OAI22_X1 U17593 ( .A1(n16003), .A2(n14312), .B1(n21379), .B2(n20211), .ZN(
        n14286) );
  INV_X1 U17594 ( .A(n14286), .ZN(n14287) );
  OAI21_X1 U17595 ( .B1(n14356), .B2(n14318), .A(n14287), .ZN(P1_U2854) );
  AND2_X1 U17596 ( .A1(n14288), .A2(n14289), .ZN(n14290) );
  NOR2_X1 U17597 ( .A1(n9890), .A2(n14290), .ZN(n15880) );
  INV_X1 U17598 ( .A(n15880), .ZN(n14360) );
  INV_X1 U17599 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14293) );
  AOI21_X1 U17600 ( .B1(n14291), .B2(n14296), .A(n9931), .ZN(n14292) );
  INV_X1 U17601 ( .A(n14292), .ZN(n15885) );
  OAI222_X1 U17602 ( .A1(n14360), .A2(n14318), .B1(n20211), .B2(n14293), .C1(
        n15885), .C2(n14312), .ZN(P1_U2855) );
  NAND2_X1 U17603 ( .A1(n14304), .A2(n14294), .ZN(n14295) );
  NAND2_X1 U17604 ( .A1(n14296), .A2(n14295), .ZN(n15893) );
  INV_X1 U17605 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21188) );
  INV_X1 U17606 ( .A(n14288), .ZN(n14299) );
  AOI21_X1 U17607 ( .B1(n14300), .B2(n14298), .A(n14299), .ZN(n15934) );
  INV_X1 U17608 ( .A(n15934), .ZN(n14367) );
  OAI222_X1 U17609 ( .A1(n15893), .A2(n14312), .B1(n20211), .B2(n21188), .C1(
        n14367), .C2(n14318), .ZN(P1_U2856) );
  NAND2_X1 U17610 ( .A1(n14301), .A2(n14302), .ZN(n14303) );
  AND2_X1 U17611 ( .A1(n14298), .A2(n14303), .ZN(n15902) );
  INV_X1 U17612 ( .A(n15902), .ZN(n14372) );
  INV_X1 U17613 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14306) );
  OAI21_X1 U17614 ( .B1(n14310), .B2(n14305), .A(n14304), .ZN(n15898) );
  OAI222_X1 U17615 ( .A1(n14372), .A2(n14318), .B1(n14306), .B2(n20211), .C1(
        n14312), .C2(n15898), .ZN(P1_U2857) );
  OAI21_X1 U17616 ( .B1(n9859), .B2(n14307), .A(n14301), .ZN(n15910) );
  AND2_X1 U17617 ( .A1(n14309), .A2(n14308), .ZN(n14311) );
  OR2_X1 U17618 ( .A1(n14311), .A2(n14310), .ZN(n16018) );
  OAI22_X1 U17619 ( .A1(n16018), .A2(n14312), .B1(n15908), .B2(n20211), .ZN(
        n14313) );
  INV_X1 U17620 ( .A(n14313), .ZN(n14314) );
  OAI21_X1 U17621 ( .B1(n15910), .B2(n14318), .A(n14314), .ZN(P1_U2858) );
  AOI22_X1 U17622 ( .A1(n16027), .A2(n20206), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14316), .ZN(n14315) );
  OAI21_X1 U17623 ( .B1(n14377), .B2(n14318), .A(n14315), .ZN(P1_U2859) );
  AOI22_X1 U17624 ( .A1(n16036), .A2(n20206), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14316), .ZN(n14317) );
  OAI21_X1 U17625 ( .B1(n15954), .B2(n14318), .A(n14317), .ZN(P1_U2860) );
  AOI22_X1 U17626 ( .A1(n14361), .A2(DATAI_29_), .B1(n14374), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17627 ( .A1(n14364), .A2(n20279), .B1(n14362), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14319) );
  OAI211_X1 U17628 ( .C1(n14321), .C2(n14382), .A(n14320), .B(n14319), .ZN(
        P1_U2875) );
  AOI22_X1 U17629 ( .A1(n14361), .A2(DATAI_28_), .B1(n14374), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17630 ( .A1(n14364), .A2(n20276), .B1(n14362), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14322) );
  OAI211_X1 U17631 ( .C1(n14398), .C2(n14382), .A(n14323), .B(n14322), .ZN(
        P1_U2876) );
  AOI22_X1 U17632 ( .A1(n14361), .A2(DATAI_27_), .B1(n14374), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14325) );
  AOI22_X1 U17633 ( .A1(n14364), .A2(n20273), .B1(n14362), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14324) );
  OAI211_X1 U17634 ( .C1(n14408), .C2(n14382), .A(n14325), .B(n14324), .ZN(
        P1_U2877) );
  AOI22_X1 U17635 ( .A1(n14361), .A2(DATAI_26_), .B1(n14374), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U17636 ( .A1(n14364), .A2(n20270), .B1(n14362), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14326) );
  OAI211_X1 U17637 ( .C1(n14328), .C2(n14382), .A(n14327), .B(n14326), .ZN(
        P1_U2878) );
  AOI22_X1 U17638 ( .A1(n14361), .A2(DATAI_25_), .B1(n14374), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17639 ( .A1(n14364), .A2(n20267), .B1(n14362), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14329) );
  OAI211_X1 U17640 ( .C1(n14331), .C2(n14382), .A(n14330), .B(n14329), .ZN(
        P1_U2879) );
  AOI22_X1 U17641 ( .A1(n14361), .A2(DATAI_24_), .B1(n14374), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17642 ( .A1(n14364), .A2(n14332), .B1(n14362), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14333) );
  OAI211_X1 U17643 ( .C1(n14335), .C2(n14382), .A(n14334), .B(n14333), .ZN(
        P1_U2880) );
  AOI22_X1 U17644 ( .A1(n14361), .A2(DATAI_23_), .B1(n14374), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14338) );
  INV_X1 U17645 ( .A(n20266), .ZN(n14336) );
  AOI22_X1 U17646 ( .A1(n14364), .A2(n14336), .B1(n14362), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14337) );
  OAI211_X1 U17647 ( .C1(n14339), .C2(n14382), .A(n14338), .B(n14337), .ZN(
        P1_U2881) );
  AOI22_X1 U17648 ( .A1(n14361), .A2(DATAI_22_), .B1(n14374), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14342) );
  INV_X1 U17649 ( .A(n20376), .ZN(n14340) );
  AOI22_X1 U17650 ( .A1(n14364), .A2(n14340), .B1(n14362), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14341) );
  OAI211_X1 U17651 ( .C1(n14343), .C2(n14382), .A(n14342), .B(n14341), .ZN(
        P1_U2882) );
  AOI22_X1 U17652 ( .A1(n14361), .A2(DATAI_21_), .B1(n14374), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14346) );
  INV_X1 U17653 ( .A(n20367), .ZN(n14344) );
  AOI22_X1 U17654 ( .A1(n14364), .A2(n14344), .B1(n14362), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14345) );
  OAI211_X1 U17655 ( .C1(n14464), .C2(n14382), .A(n14346), .B(n14345), .ZN(
        P1_U2883) );
  AOI22_X1 U17656 ( .A1(n14361), .A2(DATAI_20_), .B1(n14374), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14349) );
  INV_X1 U17657 ( .A(n20262), .ZN(n14347) );
  AOI22_X1 U17658 ( .A1(n14364), .A2(n14347), .B1(n14362), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14348) );
  OAI211_X1 U17659 ( .C1(n15860), .C2(n14382), .A(n14349), .B(n14348), .ZN(
        P1_U2884) );
  AOI22_X1 U17660 ( .A1(n14361), .A2(DATAI_19_), .B1(n14374), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14352) );
  INV_X1 U17661 ( .A(n20260), .ZN(n14350) );
  AOI22_X1 U17662 ( .A1(n14364), .A2(n14350), .B1(n14362), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14351) );
  OAI211_X1 U17663 ( .C1(n14473), .C2(n14382), .A(n14352), .B(n14351), .ZN(
        P1_U2885) );
  AOI22_X1 U17664 ( .A1(n14361), .A2(DATAI_18_), .B1(n14374), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14355) );
  INV_X1 U17665 ( .A(n20258), .ZN(n14353) );
  AOI22_X1 U17666 ( .A1(n14364), .A2(n14353), .B1(n14362), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U17667 ( .C1(n14356), .C2(n14382), .A(n14355), .B(n14354), .ZN(
        P1_U2886) );
  AOI22_X1 U17668 ( .A1(n14361), .A2(DATAI_17_), .B1(n14374), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14359) );
  INV_X1 U17669 ( .A(n20357), .ZN(n14357) );
  AOI22_X1 U17670 ( .A1(n14364), .A2(n14357), .B1(n14362), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14358) );
  OAI211_X1 U17671 ( .C1(n14360), .C2(n14382), .A(n14359), .B(n14358), .ZN(
        P1_U2887) );
  AOI22_X1 U17672 ( .A1(n14361), .A2(DATAI_16_), .B1(n14374), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14366) );
  INV_X1 U17673 ( .A(n20255), .ZN(n14363) );
  AOI22_X1 U17674 ( .A1(n14364), .A2(n14363), .B1(n14362), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14365) );
  OAI211_X1 U17675 ( .C1(n14367), .C2(n14382), .A(n14366), .B(n14365), .ZN(
        P1_U2888) );
  INV_X1 U17676 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20214) );
  INV_X1 U17677 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14368) );
  OR2_X1 U17678 ( .A1(n14369), .A2(n14368), .ZN(n14371) );
  NAND2_X1 U17679 ( .A1(n14369), .A2(DATAI_15_), .ZN(n14370) );
  AND2_X1 U17680 ( .A1(n14371), .A2(n14370), .ZN(n20290) );
  OAI222_X1 U17681 ( .A1(n14382), .A2(n14372), .B1(n14380), .B2(n20214), .C1(
        n14379), .C2(n20290), .ZN(P1_U2889) );
  AOI22_X1 U17682 ( .A1(n14375), .A2(n20282), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14374), .ZN(n14373) );
  OAI21_X1 U17683 ( .B1(n15910), .B2(n14382), .A(n14373), .ZN(P1_U2890) );
  AOI22_X1 U17684 ( .A1(n14375), .A2(n20279), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14374), .ZN(n14376) );
  OAI21_X1 U17685 ( .B1(n14377), .B2(n14382), .A(n14376), .ZN(P1_U2891) );
  INV_X1 U17686 ( .A(n20276), .ZN(n14378) );
  OAI222_X1 U17687 ( .A1(n15954), .A2(n14382), .B1(n14381), .B2(n14380), .C1(
        n14379), .C2(n14378), .ZN(P1_U2892) );
  MUX2_X1 U17688 ( .A(n14384), .B(n9825), .S(n11531), .Z(n14385) );
  XNOR2_X1 U17689 ( .A(n14385), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14544) );
  INV_X1 U17690 ( .A(n14386), .ZN(n14388) );
  AND2_X1 U17691 ( .A1(n20317), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14539) );
  AOI21_X1 U17692 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14539), .ZN(n14387) );
  OAI21_X1 U17693 ( .B1(n20302), .B2(n14388), .A(n14387), .ZN(n14389) );
  AOI21_X1 U17694 ( .B1(n14390), .B2(n15981), .A(n14389), .ZN(n14391) );
  OAI21_X1 U17695 ( .B1(n20108), .B2(n14544), .A(n14391), .ZN(P1_U2970) );
  NAND2_X1 U17696 ( .A1(n15938), .A2(n14566), .ZN(n14413) );
  NAND3_X1 U17697 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14413), .ZN(n14393) );
  OAI21_X1 U17698 ( .B1(n9838), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14393), .ZN(n14395) );
  MUX2_X1 U17699 ( .A(n14556), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15938), .Z(n14394) );
  NAND2_X1 U17700 ( .A1(n14395), .A2(n14394), .ZN(n14397) );
  XNOR2_X1 U17701 ( .A(n14397), .B(n14396), .ZN(n14554) );
  INV_X1 U17702 ( .A(n14398), .ZN(n14402) );
  AND2_X1 U17703 ( .A1(n20317), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14546) );
  AOI21_X1 U17704 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14546), .ZN(n14399) );
  OAI21_X1 U17705 ( .B1(n20302), .B2(n14400), .A(n14399), .ZN(n14401) );
  OAI21_X1 U17706 ( .B1(n20108), .B2(n14554), .A(n14403), .ZN(P1_U2971) );
  NOR3_X1 U17707 ( .A1(n14412), .A2(n14404), .A3(n15938), .ZN(n14405) );
  NOR2_X1 U17708 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  AND2_X1 U17709 ( .A1(n20317), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14555) );
  AOI21_X1 U17710 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14555), .ZN(n14409) );
  OAI21_X1 U17711 ( .B1(n20302), .B2(n14410), .A(n14409), .ZN(n14411) );
  INV_X1 U17712 ( .A(n14392), .ZN(n14433) );
  OAI21_X1 U17713 ( .B1(n14433), .B2(n11531), .A(n9838), .ZN(n14414) );
  NAND2_X1 U17714 ( .A1(n14414), .A2(n14413), .ZN(n14416) );
  XNOR2_X1 U17715 ( .A(n14416), .B(n14415), .ZN(n14574) );
  AND2_X1 U17716 ( .A1(n20317), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14568) );
  AOI21_X1 U17717 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14568), .ZN(n14417) );
  OAI21_X1 U17718 ( .B1(n20302), .B2(n14418), .A(n14417), .ZN(n14419) );
  AOI21_X1 U17719 ( .B1(n14420), .B2(n20296), .A(n14419), .ZN(n14421) );
  OAI21_X1 U17720 ( .B1(n20108), .B2(n14574), .A(n14421), .ZN(P1_U2973) );
  NOR2_X1 U17721 ( .A1(n14392), .A2(n14422), .ZN(n14425) );
  NAND2_X1 U17722 ( .A1(n14423), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14435) );
  NOR2_X1 U17723 ( .A1(n14435), .A2(n14436), .ZN(n14424) );
  MUX2_X1 U17724 ( .A(n14425), .B(n14424), .S(n15938), .Z(n14426) );
  XNOR2_X1 U17725 ( .A(n14426), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14581) );
  INV_X1 U17726 ( .A(n14427), .ZN(n14429) );
  AND2_X1 U17727 ( .A1(n20317), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14576) );
  AOI21_X1 U17728 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14576), .ZN(n14428) );
  OAI21_X1 U17729 ( .B1(n20302), .B2(n14429), .A(n14428), .ZN(n14430) );
  AOI21_X1 U17730 ( .B1(n14431), .B2(n15981), .A(n14430), .ZN(n14432) );
  OAI21_X1 U17731 ( .B1(n20108), .B2(n14581), .A(n14432), .ZN(P1_U2974) );
  NAND2_X1 U17732 ( .A1(n14433), .A2(n14435), .ZN(n14434) );
  MUX2_X1 U17733 ( .A(n14435), .B(n14434), .S(n11531), .Z(n14437) );
  XNOR2_X1 U17734 ( .A(n14437), .B(n14436), .ZN(n14591) );
  AND2_X1 U17735 ( .A1(n20317), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14584) );
  AOI21_X1 U17736 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14584), .ZN(n14438) );
  OAI21_X1 U17737 ( .B1(n20302), .B2(n14439), .A(n14438), .ZN(n14440) );
  AOI21_X1 U17738 ( .B1(n14441), .B2(n15981), .A(n14440), .ZN(n14442) );
  OAI21_X1 U17739 ( .B1(n20108), .B2(n14591), .A(n14442), .ZN(P1_U2975) );
  XNOR2_X1 U17740 ( .A(n11533), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14443) );
  XNOR2_X1 U17741 ( .A(n14392), .B(n14443), .ZN(n14601) );
  AND2_X1 U17742 ( .A1(n20317), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14595) );
  AOI21_X1 U17743 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14595), .ZN(n14444) );
  OAI21_X1 U17744 ( .B1(n20302), .B2(n14445), .A(n14444), .ZN(n14446) );
  AOI21_X1 U17745 ( .B1(n14447), .B2(n20296), .A(n14446), .ZN(n14448) );
  OAI21_X1 U17746 ( .B1(n14601), .B2(n20108), .A(n14448), .ZN(P1_U2976) );
  NAND2_X1 U17747 ( .A1(n9820), .A2(n14449), .ZN(n14451) );
  XNOR2_X1 U17748 ( .A(n14451), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15989) );
  INV_X1 U17749 ( .A(n15989), .ZN(n14458) );
  INV_X1 U17750 ( .A(n14452), .ZN(n14454) );
  AOI22_X1 U17751 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14453) );
  OAI21_X1 U17752 ( .B1(n20302), .B2(n14454), .A(n14453), .ZN(n14455) );
  AOI21_X1 U17753 ( .B1(n14456), .B2(n20296), .A(n14455), .ZN(n14457) );
  OAI21_X1 U17754 ( .B1(n20108), .B2(n14458), .A(n14457), .ZN(P1_U2977) );
  OR2_X1 U17755 ( .A1(n14515), .A2(n16001), .ZN(n14459) );
  NAND2_X1 U17756 ( .A1(n14603), .A2(n14459), .ZN(n14470) );
  INV_X1 U17757 ( .A(n14605), .ZN(n14462) );
  NAND2_X1 U17758 ( .A1(n15938), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14602) );
  NOR2_X1 U17759 ( .A1(n14602), .A2(n14461), .ZN(n14460) );
  AOI22_X1 U17760 ( .A1(n14462), .A2(n14461), .B1(n14460), .B2(n14470), .ZN(
        n14463) );
  XNOR2_X1 U17761 ( .A(n14463), .B(n11545), .ZN(n15832) );
  INV_X1 U17762 ( .A(n14464), .ZN(n14468) );
  AOI22_X1 U17763 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U17764 ( .B1(n20302), .B2(n14466), .A(n14465), .ZN(n14467) );
  AOI21_X1 U17765 ( .B1(n14468), .B2(n15981), .A(n14467), .ZN(n14469) );
  OAI21_X1 U17766 ( .B1(n20108), .B2(n15832), .A(n14469), .ZN(P1_U2978) );
  INV_X1 U17767 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14613) );
  MUX2_X1 U17768 ( .A(n14613), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n15938), .Z(n14471) );
  MUX2_X1 U17769 ( .A(n14602), .B(n14471), .S(n14470), .Z(n14472) );
  AND2_X1 U17770 ( .A1(n14472), .A2(n14605), .ZN(n15995) );
  INV_X1 U17771 ( .A(n14473), .ZN(n14478) );
  INV_X1 U17772 ( .A(n14474), .ZN(n14476) );
  AOI22_X1 U17773 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14475) );
  OAI21_X1 U17774 ( .B1(n20302), .B2(n14476), .A(n14475), .ZN(n14477) );
  AOI21_X1 U17775 ( .B1(n14478), .B2(n20296), .A(n14477), .ZN(n14479) );
  OAI21_X1 U17776 ( .B1(n15995), .B2(n20108), .A(n14479), .ZN(P1_U2980) );
  OAI21_X1 U17777 ( .B1(n14481), .B2(n14480), .A(n14603), .ZN(n16004) );
  AOI22_X1 U17778 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14482) );
  OAI21_X1 U17779 ( .B1(n20302), .B2(n14483), .A(n14482), .ZN(n14484) );
  AOI21_X1 U17780 ( .B1(n15875), .B2(n15981), .A(n14484), .ZN(n14485) );
  OAI21_X1 U17781 ( .B1(n20108), .B2(n16004), .A(n14485), .ZN(P1_U2981) );
  NOR2_X1 U17782 ( .A1(n15938), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14490) );
  INV_X1 U17783 ( .A(n15960), .ZN(n14486) );
  NOR2_X1 U17784 ( .A1(n14486), .A2(n14506), .ZN(n15940) );
  AOI21_X1 U17785 ( .B1(n15940), .B2(n14488), .A(n14487), .ZN(n14489) );
  MUX2_X1 U17786 ( .A(n14490), .B(n14515), .S(n14489), .Z(n14491) );
  XNOR2_X1 U17787 ( .A(n14491), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14629) );
  INV_X1 U17788 ( .A(n15877), .ZN(n14493) );
  AND2_X1 U17789 ( .A1(n20317), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14626) );
  AOI21_X1 U17790 ( .B1(n20291), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14626), .ZN(n14492) );
  OAI21_X1 U17791 ( .B1(n20302), .B2(n14493), .A(n14492), .ZN(n14494) );
  AOI21_X1 U17792 ( .B1(n15880), .B2(n20296), .A(n14494), .ZN(n14495) );
  OAI21_X1 U17793 ( .B1(n14629), .B2(n20108), .A(n14495), .ZN(P1_U2982) );
  INV_X1 U17794 ( .A(n14496), .ZN(n14498) );
  NOR2_X1 U17795 ( .A1(n15940), .A2(n14497), .ZN(n14633) );
  AOI21_X1 U17796 ( .B1(n11531), .B2(n14498), .A(n14633), .ZN(n14500) );
  OAI21_X1 U17797 ( .B1(n14515), .B2(n14636), .A(n14631), .ZN(n14499) );
  XNOR2_X1 U17798 ( .A(n14500), .B(n14499), .ZN(n16012) );
  AOI22_X1 U17799 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14501) );
  OAI21_X1 U17800 ( .B1(n20302), .B2(n14502), .A(n14501), .ZN(n14503) );
  AOI21_X1 U17801 ( .B1(n15902), .B2(n20296), .A(n14503), .ZN(n14504) );
  OAI21_X1 U17802 ( .B1(n16012), .B2(n20108), .A(n14504), .ZN(P1_U2984) );
  NOR2_X1 U17803 ( .A1(n15960), .A2(n14505), .ZN(n15949) );
  OAI21_X1 U17804 ( .B1(n15949), .B2(n14506), .A(n15951), .ZN(n14507) );
  XOR2_X1 U17805 ( .A(n14508), .B(n14507), .Z(n16028) );
  INV_X1 U17806 ( .A(n16028), .ZN(n14514) );
  AOI22_X1 U17807 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14509) );
  OAI21_X1 U17808 ( .B1(n20302), .B2(n14510), .A(n14509), .ZN(n14511) );
  AOI21_X1 U17809 ( .B1(n14512), .B2(n15981), .A(n14511), .ZN(n14513) );
  OAI21_X1 U17810 ( .B1(n14514), .B2(n20108), .A(n14513), .ZN(P1_U2986) );
  NAND2_X1 U17811 ( .A1(n9819), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14517) );
  XNOR2_X1 U17812 ( .A(n15960), .B(n16064), .ZN(n14516) );
  MUX2_X1 U17813 ( .A(n14517), .B(n14516), .S(n14515), .Z(n14520) );
  NOR3_X1 U17814 ( .A1(n9819), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15938), .ZN(n15961) );
  INV_X1 U17815 ( .A(n15961), .ZN(n14519) );
  NAND2_X1 U17816 ( .A1(n14520), .A2(n14519), .ZN(n16060) );
  INV_X1 U17817 ( .A(n16060), .ZN(n14526) );
  AOI22_X1 U17818 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U17819 ( .B1(n20302), .B2(n14522), .A(n14521), .ZN(n14523) );
  AOI21_X1 U17820 ( .B1(n14524), .B2(n15981), .A(n14523), .ZN(n14525) );
  OAI21_X1 U17821 ( .B1(n14526), .B2(n20108), .A(n14525), .ZN(P1_U2989) );
  INV_X1 U17822 ( .A(n14527), .ZN(n14534) );
  NAND3_X1 U17823 ( .A1(n14557), .A2(n14528), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14530) );
  AOI21_X1 U17824 ( .B1(n14531), .B2(n14530), .A(n14529), .ZN(n14532) );
  AOI211_X1 U17825 ( .C1(n14534), .C2(n20316), .A(n14533), .B(n14532), .ZN(
        n14535) );
  OAI21_X1 U17826 ( .B1(n14536), .B2(n20340), .A(n14535), .ZN(P1_U3001) );
  INV_X1 U17827 ( .A(n14557), .ZN(n14537) );
  NOR3_X1 U17828 ( .A1(n14537), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14548), .ZN(n14538) );
  AOI211_X1 U17829 ( .C1(n14540), .C2(n20316), .A(n14539), .B(n14538), .ZN(
        n14543) );
  NAND2_X1 U17830 ( .A1(n14541), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14542) );
  OAI211_X1 U17831 ( .C1(n14544), .C2(n20340), .A(n14543), .B(n14542), .ZN(
        P1_U3002) );
  INV_X1 U17832 ( .A(n14545), .ZN(n14562) );
  INV_X1 U17833 ( .A(n14546), .ZN(n14550) );
  NAND3_X1 U17834 ( .A1(n14557), .A2(n14548), .A3(n14547), .ZN(n14549) );
  OAI211_X1 U17835 ( .C1(n14551), .C2(n20344), .A(n14550), .B(n14549), .ZN(
        n14552) );
  AOI21_X1 U17836 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14562), .A(
        n14552), .ZN(n14553) );
  OAI21_X1 U17837 ( .B1(n14554), .B2(n20340), .A(n14553), .ZN(P1_U3003) );
  AOI21_X1 U17838 ( .B1(n14557), .B2(n14556), .A(n14555), .ZN(n14558) );
  OAI21_X1 U17839 ( .B1(n14559), .B2(n20344), .A(n14558), .ZN(n14561) );
  NAND2_X1 U17840 ( .A1(n14564), .A2(n14563), .ZN(n14565) );
  NOR2_X1 U17841 ( .A1(n14592), .A2(n14565), .ZN(n14575) );
  OR2_X1 U17842 ( .A1(n14578), .A2(n14575), .ZN(n14569) );
  NOR3_X1 U17843 ( .A1(n14592), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14566), .ZN(n14567) );
  AOI211_X1 U17844 ( .C1(n14569), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14568), .B(n14567), .ZN(n14573) );
  INV_X1 U17845 ( .A(n14570), .ZN(n14571) );
  NAND2_X1 U17846 ( .A1(n14571), .A2(n20316), .ZN(n14572) );
  OAI211_X1 U17847 ( .C1(n14574), .C2(n20340), .A(n14573), .B(n14572), .ZN(
        P1_U3005) );
  AOI211_X1 U17848 ( .C1(n14577), .C2(n20316), .A(n14576), .B(n14575), .ZN(
        n14580) );
  NAND2_X1 U17849 ( .A1(n14578), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14579) );
  OAI211_X1 U17850 ( .C1(n14581), .C2(n20340), .A(n14580), .B(n14579), .ZN(
        P1_U3006) );
  INV_X1 U17851 ( .A(n14582), .ZN(n14585) );
  NOR3_X1 U17852 ( .A1(n14592), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14596), .ZN(n14583) );
  AOI211_X1 U17853 ( .C1(n14585), .C2(n20316), .A(n14584), .B(n14583), .ZN(
        n14590) );
  INV_X1 U17854 ( .A(n14586), .ZN(n14587) );
  AOI21_X1 U17855 ( .B1(n14587), .B2(n20323), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14588) );
  OAI21_X1 U17856 ( .B1(n14598), .B2(n14588), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14589) );
  OAI211_X1 U17857 ( .C1(n14591), .C2(n20340), .A(n14590), .B(n14589), .ZN(
        P1_U3007) );
  INV_X1 U17858 ( .A(n14592), .ZN(n14597) );
  NOR2_X1 U17859 ( .A1(n14593), .A2(n20344), .ZN(n14594) );
  AOI211_X1 U17860 ( .C1(n14597), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        n14600) );
  NAND2_X1 U17861 ( .A1(n14598), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14599) );
  OAI211_X1 U17862 ( .C1(n14601), .C2(n20340), .A(n14600), .B(n14599), .ZN(
        P1_U3008) );
  OR2_X1 U17863 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  NAND2_X1 U17864 ( .A1(n14605), .A2(n14604), .ZN(n14606) );
  XNOR2_X1 U17865 ( .A(n14606), .B(n14461), .ZN(n15928) );
  INV_X1 U17866 ( .A(n14607), .ZN(n14612) );
  NOR3_X1 U17867 ( .A1(n14608), .A2(n20324), .A3(n14611), .ZN(n14610) );
  NOR2_X1 U17868 ( .A1(n14610), .A2(n14609), .ZN(n14615) );
  OAI21_X1 U17869 ( .B1(n14614), .B2(n14611), .A(n14615), .ZN(n16026) );
  NAND2_X1 U17870 ( .A1(n14612), .A2(n16026), .ZN(n16000) );
  NOR3_X1 U17871 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14613), .A3(
        n16000), .ZN(n14620) );
  AOI21_X1 U17872 ( .B1(n14615), .B2(n14614), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14616) );
  OAI21_X1 U17873 ( .B1(n14616), .B2(n15994), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14618) );
  INV_X1 U17874 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21246) );
  NOR2_X1 U17875 ( .A1(n20342), .A2(n21246), .ZN(n15927) );
  INV_X1 U17876 ( .A(n15927), .ZN(n14617) );
  OAI211_X1 U17877 ( .C1(n20344), .C2(n15862), .A(n14618), .B(n14617), .ZN(
        n14619) );
  AOI211_X1 U17878 ( .C1(n15928), .C2(n20332), .A(n14620), .B(n14619), .ZN(
        n14621) );
  INV_X1 U17879 ( .A(n14621), .ZN(P1_U3011) );
  OR2_X1 U17880 ( .A1(n16025), .A2(n16010), .ZN(n16017) );
  OAI21_X1 U17881 ( .B1(n14639), .B2(n16017), .A(n14622), .ZN(n14627) );
  NOR2_X1 U17882 ( .A1(n16021), .A2(n20323), .ZN(n14623) );
  AOI211_X1 U17883 ( .C1(n20327), .C2(n14624), .A(n14623), .B(n20325), .ZN(
        n16032) );
  OAI21_X1 U17884 ( .B1(n14630), .B2(n16002), .A(n16032), .ZN(n16006) );
  NOR2_X1 U17885 ( .A1(n15885), .A2(n20344), .ZN(n14625) );
  AOI211_X1 U17886 ( .C1(n14627), .C2(n16006), .A(n14626), .B(n14625), .ZN(
        n14628) );
  OAI21_X1 U17887 ( .B1(n14629), .B2(n20340), .A(n14628), .ZN(P1_U3014) );
  OAI21_X1 U17888 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14630), .A(
        n16032), .ZN(n16011) );
  INV_X1 U17889 ( .A(n16011), .ZN(n14644) );
  OAI21_X1 U17890 ( .B1(n14633), .B2(n14632), .A(n14631), .ZN(n14635) );
  XNOR2_X1 U17891 ( .A(n14635), .B(n14634), .ZN(n15933) );
  NAND2_X1 U17892 ( .A1(n15933), .A2(n20332), .ZN(n14642) );
  AOI21_X1 U17893 ( .B1(n14636), .B2(n14643), .A(n16017), .ZN(n14640) );
  INV_X1 U17894 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14637) );
  OAI22_X1 U17895 ( .A1(n15893), .A2(n20344), .B1(n20342), .B2(n14637), .ZN(
        n14638) );
  AOI21_X1 U17896 ( .B1(n14640), .B2(n14639), .A(n14638), .ZN(n14641) );
  OAI211_X1 U17897 ( .C1(n14644), .C2(n14643), .A(n14642), .B(n14641), .ZN(
        P1_U3015) );
  NOR2_X1 U17898 ( .A1(n13332), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14646) );
  OAI22_X1 U17899 ( .A1(n20443), .A2(n14646), .B1(n20595), .B2(n14645), .ZN(
        n14647) );
  MUX2_X1 U17900 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14647), .S(
        n20352), .Z(P1_U3477) );
  NOR2_X1 U17901 ( .A1(n20857), .A2(n13332), .ZN(n20716) );
  NOR2_X1 U17902 ( .A1(n20532), .A2(n20856), .ZN(n20566) );
  AOI21_X1 U17903 ( .B1(n14651), .B2(n20594), .A(n20566), .ZN(n14652) );
  OAI21_X1 U17904 ( .B1(n14653), .B2(n20804), .A(n14652), .ZN(n14654) );
  MUX2_X1 U17905 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14654), .S(
        n20352), .Z(P1_U3475) );
  INV_X1 U17906 ( .A(n20989), .ZN(n14665) );
  OR2_X1 U17907 ( .A1(n20595), .A2(n15798), .ZN(n14660) );
  INV_X1 U17908 ( .A(n14655), .ZN(n14662) );
  NAND3_X1 U17909 ( .A1(n14656), .A2(n14661), .A3(n14662), .ZN(n14657) );
  AND2_X1 U17910 ( .A1(n14658), .A2(n14657), .ZN(n14659) );
  NAND2_X1 U17911 ( .A1(n14660), .A2(n14659), .ZN(n15796) );
  NAND2_X1 U17912 ( .A1(n15796), .A2(n16093), .ZN(n14664) );
  NAND3_X1 U17913 ( .A1(n14662), .A2(n15825), .A3(n14661), .ZN(n14663) );
  OAI211_X1 U17914 ( .C1(n14666), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14667) );
  MUX2_X1 U17915 ( .A(n14667), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20992), .Z(P1_U3473) );
  OAI22_X1 U17916 ( .A1(n15793), .A2(n20995), .B1(n14668), .B2(n20987), .ZN(
        n14669) );
  MUX2_X1 U17917 ( .A(n14669), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20992), .Z(P1_U3469) );
  AOI22_X1 U17918 ( .A1(n14671), .A2(n19627), .B1(n14670), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14675) );
  INV_X1 U17919 ( .A(n14672), .ZN(n16466) );
  OAI21_X1 U17920 ( .B1(n19958), .B2(n19822), .A(n16466), .ZN(n14673) );
  OAI21_X1 U17921 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14678) );
  AOI21_X1 U17922 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16459), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14676) );
  AOI211_X1 U17923 ( .C1(n19950), .C2(n19366), .A(n14676), .B(n19032), .ZN(
        n14677) );
  MUX2_X1 U17924 ( .A(n14678), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14677), 
        .Z(P2_U3610) );
  NAND2_X1 U17925 ( .A1(n14680), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U17926 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14681) );
  AOI21_X1 U17927 ( .B1(n14685), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14684), .ZN(n14686) );
  INV_X1 U17928 ( .A(n16115), .ZN(n14688) );
  NAND2_X1 U17929 ( .A1(n14688), .A2(n14769), .ZN(n14689) );
  OAI21_X1 U17930 ( .B1(n14769), .B2(n14683), .A(n14689), .ZN(P2_U2856) );
  OR2_X1 U17931 ( .A1(n14702), .A2(n14690), .ZN(n14691) );
  NAND2_X1 U17932 ( .A1(n14692), .A2(n14691), .ZN(n16131) );
  OR2_X1 U17933 ( .A1(n14694), .A2(n14693), .ZN(n14780) );
  NAND3_X1 U17934 ( .A1(n14780), .A2(n14695), .A3(n14746), .ZN(n14697) );
  NAND2_X1 U17935 ( .A1(n14749), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14696) );
  OAI211_X1 U17936 ( .C1(n14749), .C2(n16131), .A(n14697), .B(n14696), .ZN(
        P2_U2858) );
  NOR2_X1 U17937 ( .A1(n12258), .A2(n14698), .ZN(n14700) );
  XNOR2_X1 U17938 ( .A(n14700), .B(n14699), .ZN(n14794) );
  AND2_X1 U17939 ( .A1(n14711), .A2(n14701), .ZN(n14703) );
  OR2_X1 U17940 ( .A1(n14703), .A2(n14702), .ZN(n16140) );
  NOR2_X1 U17941 ( .A1(n16140), .A2(n14776), .ZN(n14704) );
  AOI21_X1 U17942 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14776), .A(n14704), .ZN(
        n14705) );
  OAI21_X1 U17943 ( .B1(n14794), .B2(n14779), .A(n14705), .ZN(P2_U2859) );
  OAI21_X1 U17944 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14802) );
  NAND2_X1 U17945 ( .A1(n14749), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14713) );
  NAND2_X1 U17946 ( .A1(n14718), .A2(n14709), .ZN(n14710) );
  NAND2_X1 U17947 ( .A1(n14711), .A2(n14710), .ZN(n16158) );
  OR2_X1 U17948 ( .A1(n16158), .A2(n14749), .ZN(n14712) );
  OAI211_X1 U17949 ( .C1(n14802), .C2(n14779), .A(n14713), .B(n14712), .ZN(
        P2_U2860) );
  AOI21_X1 U17950 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14717) );
  INV_X1 U17951 ( .A(n14717), .ZN(n14811) );
  OAI21_X1 U17952 ( .B1(n14727), .B2(n14719), .A(n14718), .ZN(n15114) );
  NOR2_X1 U17953 ( .A1(n15114), .A2(n14776), .ZN(n14720) );
  AOI21_X1 U17954 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14749), .A(n14720), .ZN(
        n14721) );
  OAI21_X1 U17955 ( .B1(n14811), .B2(n14779), .A(n14721), .ZN(P2_U2861) );
  OAI21_X1 U17956 ( .B1(n14722), .B2(n14724), .A(n14723), .ZN(n14821) );
  NOR2_X1 U17957 ( .A1(n14734), .A2(n14725), .ZN(n14726) );
  OR2_X1 U17958 ( .A1(n14727), .A2(n14726), .ZN(n16177) );
  MUX2_X1 U17959 ( .A(n16177), .B(n14728), .S(n14749), .Z(n14729) );
  OAI21_X1 U17960 ( .B1(n14821), .B2(n14779), .A(n14729), .ZN(P2_U2862) );
  AOI21_X1 U17961 ( .B1(n14731), .B2(n14730), .A(n9938), .ZN(n14732) );
  XOR2_X1 U17962 ( .A(n14733), .B(n14732), .Z(n14828) );
  AOI21_X1 U17963 ( .B1(n14735), .B2(n14738), .A(n14734), .ZN(n16187) );
  INV_X1 U17964 ( .A(n16187), .ZN(n15344) );
  NOR2_X1 U17965 ( .A1(n15344), .A2(n14776), .ZN(n14736) );
  AOI21_X1 U17966 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14749), .A(n14736), .ZN(
        n14737) );
  OAI21_X1 U17967 ( .B1(n14828), .B2(n14779), .A(n14737), .ZN(P2_U2863) );
  INV_X1 U17968 ( .A(n14738), .ZN(n14739) );
  AOI21_X1 U17969 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n16196) );
  INV_X1 U17970 ( .A(n16196), .ZN(n15151) );
  NOR2_X1 U17971 ( .A1(n14742), .A2(n14743), .ZN(n14745) );
  NOR2_X1 U17972 ( .A1(n14745), .A2(n14744), .ZN(n16209) );
  NAND2_X1 U17973 ( .A1(n16209), .A2(n14746), .ZN(n14748) );
  NAND2_X1 U17974 ( .A1(n14749), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14747) );
  OAI211_X1 U17975 ( .C1(n15151), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        P2_U2864) );
  OR2_X1 U17976 ( .A1(n14763), .A2(n14757), .ZN(n14758) );
  INV_X1 U17977 ( .A(n14758), .ZN(n14753) );
  INV_X1 U17978 ( .A(n14751), .ZN(n14752) );
  OAI21_X1 U17979 ( .B1(n14753), .B2(n14752), .A(n12162), .ZN(n14834) );
  MUX2_X1 U17980 ( .A(n14755), .B(n14754), .S(n14749), .Z(n14756) );
  OAI21_X1 U17981 ( .B1(n14834), .B2(n14779), .A(n14756), .ZN(P2_U2865) );
  INV_X1 U17982 ( .A(n14757), .ZN(n14759) );
  OAI21_X1 U17983 ( .B1(n12127), .B2(n14759), .A(n14758), .ZN(n14840) );
  MUX2_X1 U17984 ( .A(n15385), .B(n14760), .S(n14749), .Z(n14761) );
  OAI21_X1 U17985 ( .B1(n14840), .B2(n14779), .A(n14761), .ZN(P2_U2866) );
  OAI21_X1 U17986 ( .B1(n14762), .B2(n14764), .A(n14763), .ZN(n14849) );
  INV_X1 U17987 ( .A(n14765), .ZN(n14766) );
  AOI21_X1 U17988 ( .B1(n14767), .B2(n14773), .A(n14766), .ZN(n19062) );
  NOR2_X1 U17989 ( .A1(n14769), .A2(n14952), .ZN(n14768) );
  AOI21_X1 U17990 ( .B1(n19062), .B2(n14769), .A(n14768), .ZN(n14770) );
  OAI21_X1 U17991 ( .B1(n14849), .B2(n14779), .A(n14770), .ZN(P2_U2867) );
  INV_X1 U17992 ( .A(n14762), .ZN(n14771) );
  OAI21_X1 U17993 ( .B1(n13755), .B2(n14772), .A(n14771), .ZN(n14856) );
  AOI21_X1 U17994 ( .B1(n14775), .B2(n14774), .A(n12757), .ZN(n19072) );
  INV_X1 U17995 ( .A(n19072), .ZN(n15192) );
  NOR2_X1 U17996 ( .A1(n15192), .A2(n14776), .ZN(n14777) );
  AOI21_X1 U17997 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14749), .A(n14777), .ZN(
        n14778) );
  OAI21_X1 U17998 ( .B1(n14779), .B2(n14856), .A(n14778), .ZN(P2_U2868) );
  NAND3_X1 U17999 ( .A1(n14780), .A2(n14695), .A3(n19319), .ZN(n14786) );
  INV_X1 U18000 ( .A(n14868), .ZN(n16207) );
  MUX2_X1 U18001 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n19267), .Z(n19380) );
  AOI22_X1 U18002 ( .A1(n16207), .A2(n19380), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19317), .ZN(n14785) );
  AOI22_X1 U18003 ( .A1(n19262), .A2(BUF1_REG_29__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14784) );
  OR2_X1 U18004 ( .A1(n14789), .A2(n14781), .ZN(n14782) );
  NAND2_X1 U18005 ( .A1(n16133), .A2(n19318), .ZN(n14783) );
  NAND4_X1 U18006 ( .A1(n14786), .A2(n14785), .A3(n14784), .A4(n14783), .ZN(
        P2_U2890) );
  NOR2_X1 U18007 ( .A1(n14797), .A2(n14787), .ZN(n14788) );
  INV_X1 U18008 ( .A(n15294), .ZN(n16141) );
  AOI22_X1 U18009 ( .A1(n19268), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19267), .ZN(n19400) );
  OAI22_X1 U18010 ( .A1(n14868), .A2(n19400), .B1(n19282), .B2(n14790), .ZN(
        n14791) );
  AOI21_X1 U18011 ( .B1(n16141), .B2(n19318), .A(n14791), .ZN(n14793) );
  AOI22_X1 U18012 ( .A1(n19262), .A2(BUF1_REG_28__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14792) );
  OAI211_X1 U18013 ( .C1(n14794), .C2(n19269), .A(n14793), .B(n14792), .ZN(
        P2_U2891) );
  NOR2_X1 U18014 ( .A1(n14804), .A2(n14795), .ZN(n14796) );
  OR2_X1 U18015 ( .A1(n14797), .A2(n14796), .ZN(n15306) );
  INV_X1 U18016 ( .A(n15306), .ZN(n16161) );
  INV_X1 U18017 ( .A(n19278), .ZN(n14798) );
  OAI22_X1 U18018 ( .A1(n14868), .A2(n14798), .B1(n19282), .B2(n12904), .ZN(
        n14799) );
  AOI21_X1 U18019 ( .B1(n16161), .B2(n19318), .A(n14799), .ZN(n14801) );
  AOI22_X1 U18020 ( .A1(n19262), .A2(BUF1_REG_27__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U18021 ( .C1(n14802), .C2(n19269), .A(n14801), .B(n14800), .ZN(
        P2_U2892) );
  AND2_X1 U18022 ( .A1(n14815), .A2(n14803), .ZN(n14805) );
  OR2_X1 U18023 ( .A1(n14805), .A2(n14804), .ZN(n16169) );
  INV_X1 U18024 ( .A(n16169), .ZN(n15317) );
  INV_X1 U18025 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16583) );
  NOR2_X1 U18026 ( .A1(n19267), .A2(n16583), .ZN(n14806) );
  AOI21_X1 U18027 ( .B1(n19267), .B2(BUF2_REG_10__SCAN_IN), .A(n14806), .ZN(
        n19398) );
  OAI22_X1 U18028 ( .A1(n14868), .A2(n19398), .B1(n19282), .B2(n14807), .ZN(
        n14808) );
  AOI21_X1 U18029 ( .B1(n19318), .B2(n15317), .A(n14808), .ZN(n14810) );
  AOI22_X1 U18030 ( .A1(n19262), .A2(BUF1_REG_26__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14809) );
  OAI211_X1 U18031 ( .C1(n14811), .C2(n19269), .A(n14810), .B(n14809), .ZN(
        P2_U2893) );
  NAND2_X1 U18032 ( .A1(n14813), .A2(n14812), .ZN(n14814) );
  NAND2_X1 U18033 ( .A1(n14815), .A2(n14814), .ZN(n16184) );
  INV_X1 U18034 ( .A(n16184), .ZN(n15329) );
  INV_X1 U18035 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16585) );
  NOR2_X1 U18036 ( .A1(n19267), .A2(n16585), .ZN(n14816) );
  AOI21_X1 U18037 ( .B1(n19267), .B2(BUF2_REG_9__SCAN_IN), .A(n14816), .ZN(
        n19396) );
  OAI22_X1 U18038 ( .A1(n14868), .A2(n19396), .B1(n19282), .B2(n14817), .ZN(
        n14818) );
  AOI21_X1 U18039 ( .B1(n19318), .B2(n15329), .A(n14818), .ZN(n14820) );
  AOI22_X1 U18040 ( .A1(n19262), .A2(BUF1_REG_25__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14819) );
  OAI211_X1 U18041 ( .C1(n14821), .C2(n19269), .A(n14820), .B(n14819), .ZN(
        P2_U2894) );
  INV_X1 U18042 ( .A(n19318), .ZN(n19270) );
  XOR2_X1 U18043 ( .A(n14822), .B(n15356), .Z(n16186) );
  INV_X1 U18044 ( .A(n16186), .ZN(n14824) );
  OAI22_X1 U18045 ( .A1(n19270), .A2(n14824), .B1(n19282), .B2(n14823), .ZN(
        n14825) );
  AOI21_X1 U18046 ( .B1(n16207), .B2(n19286), .A(n14825), .ZN(n14827) );
  AOI22_X1 U18047 ( .A1(n19262), .A2(BUF1_REG_24__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14826) );
  OAI211_X1 U18048 ( .C1(n14828), .C2(n19269), .A(n14827), .B(n14826), .ZN(
        P2_U2895) );
  INV_X1 U18049 ( .A(n15373), .ZN(n14831) );
  AOI22_X1 U18050 ( .A1(n19268), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19267), .ZN(n19461) );
  OAI22_X1 U18051 ( .A1(n14868), .A2(n19461), .B1(n19282), .B2(n14829), .ZN(
        n14830) );
  AOI21_X1 U18052 ( .B1(n19318), .B2(n14831), .A(n14830), .ZN(n14833) );
  AOI22_X1 U18053 ( .A1(n19262), .A2(BUF1_REG_22__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n14832) );
  OAI211_X1 U18054 ( .C1(n14834), .C2(n19269), .A(n14833), .B(n14832), .ZN(
        P2_U2897) );
  AOI22_X1 U18055 ( .A1(n19268), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19267), .ZN(n19457) );
  OAI22_X1 U18056 ( .A1(n14868), .A2(n19457), .B1(n19282), .B2(n14835), .ZN(
        n14836) );
  AOI21_X1 U18057 ( .B1(n19318), .B2(n14837), .A(n14836), .ZN(n14839) );
  AOI22_X1 U18058 ( .A1(n19262), .A2(BUF1_REG_21__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14838) );
  OAI211_X1 U18059 ( .C1(n14840), .C2(n19269), .A(n14839), .B(n14838), .ZN(
        P2_U2898) );
  OAI21_X1 U18060 ( .B1(n14843), .B2(n14842), .A(n14841), .ZN(n19059) );
  INV_X1 U18061 ( .A(n19059), .ZN(n14846) );
  OAI22_X1 U18062 ( .A1(n14868), .A2(n19453), .B1(n19282), .B2(n14844), .ZN(
        n14845) );
  AOI21_X1 U18063 ( .B1(n19318), .B2(n14846), .A(n14845), .ZN(n14848) );
  AOI22_X1 U18064 ( .A1(n19262), .A2(BUF1_REG_20__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n14847) );
  OAI211_X1 U18065 ( .C1(n14849), .C2(n19269), .A(n14848), .B(n14847), .ZN(
        P2_U2899) );
  XNOR2_X1 U18066 ( .A(n14850), .B(n14857), .ZN(n19074) );
  INV_X1 U18067 ( .A(n19074), .ZN(n14853) );
  AOI22_X1 U18068 ( .A1(n19268), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19267), .ZN(n19446) );
  OAI22_X1 U18069 ( .A1(n14868), .A2(n19446), .B1(n19282), .B2(n14851), .ZN(
        n14852) );
  AOI21_X1 U18070 ( .B1(n19318), .B2(n14853), .A(n14852), .ZN(n14855) );
  AOI22_X1 U18071 ( .A1(n19262), .A2(BUF1_REG_19__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U18072 ( .C1(n14856), .C2(n19269), .A(n14855), .B(n14854), .ZN(
        P2_U2900) );
  OAI21_X1 U18073 ( .B1(n14858), .B2(n14864), .A(n14857), .ZN(n19084) );
  INV_X1 U18074 ( .A(n19084), .ZN(n16303) );
  AOI22_X1 U18075 ( .A1(n19268), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19267), .ZN(n19440) );
  OAI22_X1 U18076 ( .A1(n14868), .A2(n19440), .B1(n19282), .B2(n14859), .ZN(
        n14860) );
  AOI21_X1 U18077 ( .B1(n19318), .B2(n16303), .A(n14860), .ZN(n14862) );
  AOI22_X1 U18078 ( .A1(n19262), .A2(BUF1_REG_18__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n14861) );
  OAI211_X1 U18079 ( .C1(n14863), .C2(n19269), .A(n14862), .B(n14861), .ZN(
        P2_U2901) );
  AOI21_X1 U18080 ( .B1(n14866), .B2(n14865), .A(n14864), .ZN(n19089) );
  OAI22_X1 U18081 ( .A1(n14868), .A2(n19388), .B1(n19282), .B2(n14867), .ZN(
        n14869) );
  AOI21_X1 U18082 ( .B1(n19318), .B2(n19089), .A(n14869), .ZN(n14871) );
  AOI22_X1 U18083 ( .A1(n19262), .A2(BUF1_REG_17__SCAN_IN), .B1(n19264), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14870) );
  OAI211_X1 U18084 ( .C1(n14872), .C2(n19269), .A(n14871), .B(n14870), .ZN(
        P2_U2902) );
  INV_X1 U18085 ( .A(n14908), .ZN(n14906) );
  AOI22_X1 U18086 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n14876), .B1(
        n19757), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14885) );
  INV_X1 U18087 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14878) );
  OAI22_X1 U18088 ( .A1(n14878), .A2(n19478), .B1(n13639), .B2(n14877), .ZN(
        n14879) );
  INV_X1 U18089 ( .A(n14879), .ZN(n14884) );
  AOI22_X1 U18090 ( .A1(n19546), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14880), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U18091 ( .A1(n14881), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n19823), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14882) );
  INV_X1 U18092 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14887) );
  INV_X1 U18093 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14886) );
  OAI22_X1 U18094 ( .A1(n14887), .A2(n13648), .B1(n19576), .B2(n14886), .ZN(
        n14891) );
  INV_X1 U18095 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14889) );
  OAI22_X1 U18096 ( .A1(n14889), .A2(n19507), .B1(n19624), .B2(n14888), .ZN(
        n14890) );
  NOR2_X1 U18097 ( .A1(n14891), .A2(n14890), .ZN(n14901) );
  INV_X1 U18098 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14894) );
  OAI22_X1 U18099 ( .A1(n14894), .A2(n14893), .B1(n19691), .B2(n14892), .ZN(
        n14895) );
  INV_X1 U18100 ( .A(n14895), .ZN(n14900) );
  INV_X1 U18101 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14897) );
  OAI22_X1 U18102 ( .A1(n14897), .A2(n19786), .B1(n13654), .B2(n14896), .ZN(
        n14898) );
  INV_X1 U18103 ( .A(n14898), .ZN(n14899) );
  NAND4_X1 U18104 ( .A1(n14902), .A2(n14901), .A3(n14900), .A4(n14899), .ZN(
        n14905) );
  NAND2_X1 U18105 ( .A1(n14903), .A2(n12403), .ZN(n14904) );
  INV_X1 U18106 ( .A(n14907), .ZN(n15048) );
  NAND2_X1 U18107 ( .A1(n14908), .A2(n15048), .ZN(n14909) );
  INV_X1 U18108 ( .A(n14910), .ZN(n14916) );
  XNOR2_X1 U18109 ( .A(n14917), .B(n14916), .ZN(n19208) );
  INV_X1 U18110 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16382) );
  XNOR2_X1 U18111 ( .A(n14911), .B(n16382), .ZN(n16292) );
  NAND2_X1 U18112 ( .A1(n14911), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14912) );
  OAI21_X1 U18113 ( .B1(n14915), .B2(n14913), .A(n14925), .ZN(n19184) );
  OR2_X1 U18114 ( .A1(n19184), .A2(n15043), .ZN(n14923) );
  INV_X1 U18115 ( .A(n14923), .ZN(n14914) );
  NAND2_X1 U18116 ( .A1(n14914), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15501) );
  INV_X1 U18117 ( .A(n14915), .ZN(n14921) );
  NAND2_X1 U18118 ( .A1(n14917), .A2(n14916), .ZN(n14919) );
  NAND2_X1 U18119 ( .A1(n14919), .A2(n14918), .ZN(n14920) );
  NAND2_X1 U18120 ( .A1(n14921), .A2(n14920), .ZN(n19198) );
  INV_X1 U18121 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16358) );
  OR2_X1 U18122 ( .A1(n19198), .A2(n16358), .ZN(n15498) );
  INV_X1 U18123 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U18124 ( .A1(n14923), .A2(n14922), .ZN(n15500) );
  NAND2_X1 U18125 ( .A1(n19198), .A2(n16358), .ZN(n15497) );
  AND2_X1 U18126 ( .A1(n15500), .A2(n15497), .ZN(n14924) );
  INV_X1 U18127 ( .A(n14929), .ZN(n14928) );
  NAND2_X1 U18128 ( .A1(n12683), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14926) );
  MUX2_X1 U18129 ( .A(n9853), .B(n14926), .S(n14925), .Z(n14927) );
  NAND2_X1 U18130 ( .A1(n14928), .A2(n14927), .ZN(n19174) );
  INV_X1 U18131 ( .A(n19174), .ZN(n14941) );
  AOI21_X1 U18132 ( .B1(n14941), .B2(n15087), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15482) );
  NAND2_X1 U18133 ( .A1(n9853), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14930) );
  MUX2_X1 U18134 ( .A(n14930), .B(P2_EBX_REG_10__SCAN_IN), .S(n14929), .Z(
        n14931) );
  AND2_X1 U18135 ( .A1(n14931), .A2(n15012), .ZN(n19163) );
  NAND2_X1 U18136 ( .A1(n19163), .A2(n15087), .ZN(n14938) );
  INV_X1 U18137 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15471) );
  NAND2_X1 U18138 ( .A1(n14938), .A2(n15471), .ZN(n15466) );
  INV_X1 U18139 ( .A(n14932), .ZN(n14936) );
  INV_X1 U18140 ( .A(n14933), .ZN(n14934) );
  NAND3_X1 U18141 ( .A1(n12683), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n14934), 
        .ZN(n14935) );
  NAND2_X1 U18142 ( .A1(n14936), .A2(n14935), .ZN(n19154) );
  OR2_X1 U18143 ( .A1(n19154), .A2(n15043), .ZN(n14937) );
  OR2_X1 U18144 ( .A1(n14938), .A2(n15471), .ZN(n15467) );
  INV_X1 U18145 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14939) );
  NOR2_X1 U18146 ( .A1(n15043), .A2(n14939), .ZN(n14940) );
  NAND2_X1 U18147 ( .A1(n14941), .A2(n14940), .ZN(n15465) );
  NAND2_X1 U18148 ( .A1(n15467), .A2(n15465), .ZN(n16258) );
  OR2_X1 U18149 ( .A1(n15043), .A2(n16265), .ZN(n14942) );
  NOR2_X1 U18150 ( .A1(n19154), .A2(n14942), .ZN(n16259) );
  NOR2_X1 U18151 ( .A1(n16258), .A2(n16259), .ZN(n14943) );
  NAND3_X1 U18152 ( .A1(n9853), .A2(n14944), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n14945) );
  AND2_X1 U18153 ( .A1(n14947), .A2(n14945), .ZN(n19143) );
  NAND2_X1 U18154 ( .A1(n19143), .A2(n15087), .ZN(n14949) );
  INV_X1 U18155 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16326) );
  NOR2_X1 U18156 ( .A1(n14949), .A2(n16326), .ZN(n15454) );
  NAND2_X1 U18157 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  NAND2_X1 U18158 ( .A1(n14964), .A2(n14948), .ZN(n19136) );
  INV_X1 U18159 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14988) );
  OAI21_X1 U18160 ( .B1(n19136), .B2(n15043), .A(n14988), .ZN(n16245) );
  NAND2_X1 U18161 ( .A1(n14949), .A2(n16326), .ZN(n16242) );
  AND2_X1 U18162 ( .A1(n16245), .A2(n16242), .ZN(n14950) );
  NOR2_X1 U18163 ( .A1(n14951), .A2(n15043), .ZN(n14991) );
  NOR2_X1 U18164 ( .A1(n14991), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15161) );
  NOR2_X1 U18165 ( .A1(n12404), .A2(n14952), .ZN(n14953) );
  XNOR2_X1 U18166 ( .A(n14954), .B(n14953), .ZN(n19056) );
  AOI21_X1 U18167 ( .B1(n19056), .B2(n15087), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15177) );
  INV_X1 U18168 ( .A(n14969), .ZN(n14956) );
  NAND2_X1 U18169 ( .A1(n14956), .A2(n14955), .ZN(n14971) );
  NAND3_X1 U18170 ( .A1(n14971), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n12683), 
        .ZN(n14957) );
  NAND2_X1 U18171 ( .A1(n10199), .A2(n14957), .ZN(n19069) );
  OR2_X1 U18172 ( .A1(n19069), .A2(n15043), .ZN(n14958) );
  INV_X1 U18173 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15189) );
  NAND2_X1 U18174 ( .A1(n14958), .A2(n15189), .ZN(n15185) );
  NOR2_X1 U18175 ( .A1(n12404), .A2(n14959), .ZN(n14960) );
  NAND2_X1 U18176 ( .A1(n14976), .A2(n14960), .ZN(n14961) );
  NAND2_X1 U18177 ( .A1(n14961), .A2(n14969), .ZN(n19086) );
  INV_X1 U18178 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15211) );
  INV_X1 U18179 ( .A(n14962), .ZN(n14963) );
  XNOR2_X1 U18180 ( .A(n14964), .B(n14963), .ZN(n19122) );
  NAND2_X1 U18181 ( .A1(n19122), .A2(n15087), .ZN(n14965) );
  INV_X1 U18182 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U18183 ( .A1(n14965), .A2(n15443), .ZN(n15447) );
  OR2_X1 U18184 ( .A1(n14967), .A2(n14966), .ZN(n14968) );
  AND2_X1 U18185 ( .A1(n14968), .A2(n14975), .ZN(n19113) );
  NAND2_X1 U18186 ( .A1(n19113), .A2(n15087), .ZN(n14983) );
  INV_X1 U18187 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16318) );
  NAND2_X1 U18188 ( .A1(n14983), .A2(n16318), .ZN(n16220) );
  NAND4_X1 U18189 ( .A1(n15185), .A2(n15158), .A3(n15447), .A4(n16220), .ZN(
        n14979) );
  NAND2_X1 U18190 ( .A1(n9853), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14970) );
  MUX2_X1 U18191 ( .A(n12683), .B(n14970), .S(n14969), .Z(n14972) );
  NAND2_X1 U18192 ( .A1(n14972), .A2(n14971), .ZN(n19079) );
  INV_X1 U18193 ( .A(n19079), .ZN(n14993) );
  AOI21_X1 U18194 ( .B1(n14993), .B2(n15087), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15198) );
  NOR2_X1 U18195 ( .A1(n12404), .A2(n14973), .ZN(n14974) );
  INV_X1 U18196 ( .A(n15012), .ZN(n15005) );
  AOI21_X1 U18197 ( .B1(n14975), .B2(n14974), .A(n15005), .ZN(n14977) );
  NAND2_X1 U18198 ( .A1(n19096), .A2(n15087), .ZN(n14978) );
  XNOR2_X1 U18199 ( .A(n14978), .B(n15430), .ZN(n15214) );
  INV_X1 U18200 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14981) );
  NOR2_X1 U18201 ( .A1(n15043), .A2(n14981), .ZN(n14982) );
  INV_X1 U18202 ( .A(n14983), .ZN(n14984) );
  NAND2_X1 U18203 ( .A1(n14984), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16221) );
  NOR2_X1 U18204 ( .A1(n15043), .A2(n15443), .ZN(n14985) );
  NAND2_X1 U18205 ( .A1(n19122), .A2(n14985), .ZN(n16223) );
  AND2_X1 U18206 ( .A1(n16221), .A2(n16223), .ZN(n15154) );
  NOR2_X1 U18207 ( .A1(n15043), .A2(n15430), .ZN(n14986) );
  NAND2_X1 U18208 ( .A1(n19096), .A2(n14986), .ZN(n15156) );
  OR2_X1 U18209 ( .A1(n15043), .A2(n15211), .ZN(n14987) );
  OR2_X1 U18210 ( .A1(n19086), .A2(n14987), .ZN(n15157) );
  INV_X1 U18211 ( .A(n19136), .ZN(n14990) );
  NOR2_X1 U18212 ( .A1(n15043), .A2(n14988), .ZN(n14989) );
  NAND2_X1 U18213 ( .A1(n14990), .A2(n14989), .ZN(n16244) );
  NAND4_X1 U18214 ( .A1(n15154), .A2(n15156), .A3(n15157), .A4(n16244), .ZN(
        n14995) );
  NAND2_X1 U18215 ( .A1(n14991), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15162) );
  NOR2_X1 U18216 ( .A1(n15043), .A2(n16300), .ZN(n14992) );
  NAND2_X1 U18217 ( .A1(n14993), .A2(n14992), .ZN(n15199) );
  OR2_X1 U18218 ( .A1(n15043), .A2(n15189), .ZN(n14994) );
  OR2_X1 U18219 ( .A1(n19069), .A2(n14994), .ZN(n15184) );
  AND2_X1 U18220 ( .A1(n15199), .A2(n15184), .ZN(n15159) );
  INV_X1 U18221 ( .A(n14996), .ZN(n14997) );
  AOI21_X1 U18222 ( .B1(n14997), .B2(n15087), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15363) );
  NAND3_X1 U18223 ( .A1(n14997), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15087), .ZN(n15364) );
  NOR2_X1 U18224 ( .A1(n12404), .A2(n14998), .ZN(n14999) );
  NAND2_X1 U18225 ( .A1(n15000), .A2(n14999), .ZN(n15001) );
  NAND2_X1 U18226 ( .A1(n15006), .A2(n15001), .ZN(n16201) );
  NOR2_X1 U18227 ( .A1(n16201), .A2(n15043), .ZN(n15002) );
  INV_X1 U18228 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15352) );
  XNOR2_X1 U18229 ( .A(n15002), .B(n15352), .ZN(n15144) );
  NOR2_X1 U18230 ( .A1(n12404), .A2(n15004), .ZN(n15007) );
  AOI211_X1 U18231 ( .C1(n15007), .C2(n15006), .A(n15005), .B(n15010), .ZN(
        n16185) );
  INV_X1 U18232 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15255) );
  NAND2_X1 U18233 ( .A1(n12683), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U18234 ( .A1(n15010), .A2(n14728), .ZN(n15013) );
  INV_X1 U18235 ( .A(n15083), .ZN(n15011) );
  NAND2_X1 U18236 ( .A1(n15012), .A2(n15011), .ZN(n15035) );
  NAND2_X1 U18237 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n15013), .ZN(n15014) );
  NOR2_X1 U18238 ( .A1(n12404), .A2(n15014), .ZN(n15015) );
  NOR2_X1 U18239 ( .A1(n15035), .A2(n15015), .ZN(n16166) );
  NAND2_X1 U18240 ( .A1(n16166), .A2(n15087), .ZN(n15022) );
  XNOR2_X1 U18241 ( .A(n15022), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15113) );
  INV_X1 U18242 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15302) );
  NAND2_X1 U18243 ( .A1(n9853), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15084) );
  NAND2_X1 U18244 ( .A1(n15035), .A2(n15084), .ZN(n15086) );
  NOR2_X1 U18245 ( .A1(n12404), .A2(n15016), .ZN(n15017) );
  AND2_X1 U18246 ( .A1(n15086), .A2(n15017), .ZN(n15018) );
  NOR2_X2 U18247 ( .A1(n15086), .A2(n15017), .ZN(n15029) );
  OR2_X1 U18248 ( .A1(n15018), .A2(n15029), .ZN(n16147) );
  INV_X1 U18249 ( .A(n16147), .ZN(n15019) );
  NAND2_X1 U18250 ( .A1(n15019), .A2(n15087), .ZN(n15092) );
  AOI21_X1 U18251 ( .B1(n15081), .B2(n15302), .A(n15092), .ZN(n15024) );
  INV_X1 U18252 ( .A(n15020), .ZN(n15021) );
  INV_X1 U18253 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15331) );
  INV_X1 U18254 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15315) );
  OR2_X1 U18255 ( .A1(n15022), .A2(n15315), .ZN(n15023) );
  NAND2_X1 U18256 ( .A1(n15111), .A2(n15023), .ZN(n15082) );
  NAND2_X1 U18257 ( .A1(n15025), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15026) );
  NAND2_X1 U18258 ( .A1(n12683), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15028) );
  XOR2_X1 U18259 ( .A(n15028), .B(n15029), .Z(n16128) );
  AOI21_X1 U18260 ( .B1(n16128), .B2(n15087), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15069) );
  INV_X1 U18261 ( .A(n15069), .ZN(n15027) );
  NAND2_X1 U18262 ( .A1(n15029), .A2(n15028), .ZN(n15036) );
  NOR2_X1 U18263 ( .A1(n12404), .A2(n15030), .ZN(n15031) );
  XNOR2_X1 U18264 ( .A(n15036), .B(n15031), .ZN(n16118) );
  OR2_X1 U18265 ( .A1(n16118), .A2(n15043), .ZN(n15032) );
  INV_X1 U18266 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U18267 ( .A1(n15032), .A2(n15269), .ZN(n15060) );
  INV_X1 U18268 ( .A(n15068), .ZN(n15033) );
  INV_X1 U18269 ( .A(n15035), .ZN(n15038) );
  NOR2_X1 U18270 ( .A1(n15036), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15037) );
  MUX2_X1 U18271 ( .A(n15038), .B(n15037), .S(n9853), .Z(n16103) );
  NAND2_X1 U18272 ( .A1(n16103), .A2(n15087), .ZN(n15039) );
  XOR2_X1 U18273 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15039), .Z(
        n15040) );
  XNOR2_X1 U18274 ( .A(n15041), .B(n15040), .ZN(n15267) );
  NAND2_X1 U18275 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15050), .ZN(
        n15051) );
  NOR2_X1 U18277 ( .A1(n15049), .A2(n15044), .ZN(n15046) );
  MUX2_X1 U18278 ( .A(n15044), .B(n15046), .S(n15045), .Z(n15047) );
  XNOR2_X1 U18279 ( .A(n14922), .B(n15050), .ZN(n15495) );
  NAND2_X1 U18280 ( .A1(n9836), .A2(n10178), .ZN(n15494) );
  INV_X1 U18281 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15378) );
  NAND2_X1 U18282 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16349) );
  NOR2_X1 U18283 ( .A1(n14939), .A2(n16349), .ZN(n15440) );
  NAND2_X1 U18284 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15442) );
  NOR2_X1 U18285 ( .A1(n15443), .A2(n15442), .ZN(n15441) );
  NAND2_X1 U18286 ( .A1(n15440), .A2(n15441), .ZN(n15413) );
  NAND2_X1 U18287 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15411) );
  NOR2_X1 U18288 ( .A1(n15211), .A2(n15411), .ZN(n16302) );
  NAND2_X1 U18289 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16302), .ZN(
        n15391) );
  NOR2_X1 U18290 ( .A1(n15413), .A2(n15391), .ZN(n15392) );
  NAND3_X1 U18291 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n15392), .ZN(n15166) );
  NOR2_X1 U18292 ( .A1(n15378), .A2(n15166), .ZN(n15252) );
  NAND2_X1 U18293 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15350) );
  NAND3_X1 U18294 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U18295 ( .A1(n15072), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15052) );
  XNOR2_X1 U18296 ( .A(n15052), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15265) );
  INV_X1 U18297 ( .A(n15053), .ZN(n15056) );
  NAND2_X1 U18298 ( .A1(n19412), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15243) );
  OAI21_X1 U18299 ( .B1(n19423), .B2(n15054), .A(n15243), .ZN(n15055) );
  AOI21_X1 U18300 ( .B1(n19411), .B2(n15056), .A(n15055), .ZN(n15057) );
  OAI21_X1 U18301 ( .B1(n16115), .B2(n16284), .A(n15057), .ZN(n15058) );
  AOI21_X1 U18302 ( .B1(n15265), .B2(n16294), .A(n15058), .ZN(n15059) );
  OAI21_X1 U18303 ( .B1(n15267), .B2(n19415), .A(n15059), .ZN(P2_U2983) );
  NAND2_X1 U18304 ( .A1(n9887), .A2(n15060), .ZN(n15061) );
  XNOR2_X1 U18305 ( .A(n15062), .B(n15061), .ZN(n15278) );
  XNOR2_X1 U18306 ( .A(n15072), .B(n15269), .ZN(n15276) );
  XNOR2_X1 U18307 ( .A(n9970), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16116) );
  INV_X1 U18308 ( .A(n16116), .ZN(n15064) );
  NAND2_X1 U18309 ( .A1(n19412), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15270) );
  OAI21_X1 U18310 ( .B1(n19423), .B2(n10336), .A(n15270), .ZN(n15063) );
  AOI21_X1 U18311 ( .B1(n19411), .B2(n15064), .A(n15063), .ZN(n15065) );
  OAI21_X1 U18312 ( .B1(n16120), .B2(n16284), .A(n15065), .ZN(n15066) );
  AOI21_X1 U18313 ( .B1(n15276), .B2(n16294), .A(n15066), .ZN(n15067) );
  OAI21_X1 U18314 ( .B1(n15278), .B2(n19415), .A(n15067), .ZN(P2_U2984) );
  NOR2_X1 U18315 ( .A1(n15069), .A2(n15068), .ZN(n15071) );
  AOI21_X1 U18316 ( .B1(n15102), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15073) );
  NOR2_X1 U18317 ( .A1(n15073), .A2(n15072), .ZN(n15288) );
  AND2_X1 U18318 ( .A1(n15074), .A2(n15076), .ZN(n15075) );
  NOR2_X1 U18319 ( .A1(n9970), .A2(n15075), .ZN(n16125) );
  NAND2_X1 U18320 ( .A1(n19412), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15281) );
  OAI21_X1 U18321 ( .B1(n19423), .B2(n15076), .A(n15281), .ZN(n15077) );
  AOI21_X1 U18322 ( .B1(n19411), .B2(n16125), .A(n15077), .ZN(n15078) );
  OAI21_X1 U18323 ( .B1(n16131), .B2(n16284), .A(n15078), .ZN(n15079) );
  AOI21_X1 U18324 ( .B1(n15288), .B2(n16294), .A(n15079), .ZN(n15080) );
  OAI21_X1 U18325 ( .B1(n15290), .B2(n19415), .A(n15080), .ZN(P2_U2985) );
  OR2_X1 U18326 ( .A1(n15084), .A2(n15083), .ZN(n15085) );
  AND2_X1 U18327 ( .A1(n15086), .A2(n15085), .ZN(n16155) );
  NAND2_X1 U18328 ( .A1(n16155), .A2(n15087), .ZN(n15089) );
  XNOR2_X1 U18329 ( .A(n15090), .B(n15088), .ZN(n15101) );
  NAND2_X1 U18330 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15100) );
  OR2_X1 U18331 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  NAND2_X1 U18332 ( .A1(n15100), .A2(n15091), .ZN(n15094) );
  XNOR2_X1 U18333 ( .A(n15092), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15093) );
  XNOR2_X1 U18334 ( .A(n15094), .B(n15093), .ZN(n15300) );
  XOR2_X1 U18335 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15102), .Z(
        n15298) );
  INV_X1 U18336 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20033) );
  NOR2_X1 U18337 ( .A1(n16334), .A2(n20033), .ZN(n15291) );
  OAI21_X1 U18338 ( .B1(n15095), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15074), .ZN(n16109) );
  NOR2_X1 U18339 ( .A1(n16277), .A2(n16109), .ZN(n15096) );
  AOI211_X1 U18340 ( .C1(n16270), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15291), .B(n15096), .ZN(n15097) );
  OAI21_X1 U18341 ( .B1(n16140), .B2(n16284), .A(n15097), .ZN(n15098) );
  AOI21_X1 U18342 ( .B1(n15298), .B2(n16294), .A(n15098), .ZN(n15099) );
  OAI21_X1 U18343 ( .B1(n15300), .B2(n19415), .A(n15099), .ZN(P2_U2986) );
  OR2_X1 U18344 ( .A1(n15101), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15301) );
  NAND3_X1 U18345 ( .A1(n15100), .A2(n16293), .A3(n15301), .ZN(n15110) );
  AOI21_X1 U18346 ( .B1(n15302), .B2(n15118), .A(n15102), .ZN(n15311) );
  NOR2_X1 U18347 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n15103), .ZN(
        n15104) );
  NOR2_X1 U18348 ( .A1(n15095), .A2(n15104), .ZN(n16154) );
  INV_X1 U18349 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U18350 ( .A1(n19412), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15305) );
  OAI21_X1 U18351 ( .B1(n19423), .B2(n15105), .A(n15305), .ZN(n15106) );
  AOI21_X1 U18352 ( .B1(n19411), .B2(n16154), .A(n15106), .ZN(n15107) );
  OAI21_X1 U18353 ( .B1(n16158), .B2(n16284), .A(n15107), .ZN(n15108) );
  AOI21_X1 U18354 ( .B1(n15311), .B2(n16294), .A(n15108), .ZN(n15109) );
  NAND2_X1 U18355 ( .A1(n15110), .A2(n15109), .ZN(P2_U2987) );
  NOR2_X1 U18356 ( .A1(n15122), .A2(n15126), .ZN(n15112) );
  XOR2_X1 U18357 ( .A(n15113), .B(n15112), .Z(n15314) );
  INV_X1 U18358 ( .A(n15114), .ZN(n16172) );
  OAI21_X1 U18359 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n15115), .A(
        n15116), .ZN(n16110) );
  NAND2_X1 U18360 ( .A1(n19412), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15318) );
  NAND2_X1 U18361 ( .A1(n16270), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15117) );
  OAI211_X1 U18362 ( .C1(n16277), .C2(n16110), .A(n15318), .B(n15117), .ZN(
        n15120) );
  OAI21_X1 U18363 ( .B1(n15128), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15118), .ZN(n15325) );
  NOR2_X1 U18364 ( .A1(n15325), .A2(n19416), .ZN(n15119) );
  AOI211_X1 U18365 ( .C1(n16172), .C2(n19420), .A(n15120), .B(n15119), .ZN(
        n15121) );
  OAI21_X1 U18366 ( .B1(n15314), .B2(n19415), .A(n15121), .ZN(P2_U2988) );
  INV_X1 U18367 ( .A(n15122), .ZN(n15127) );
  OAI21_X1 U18368 ( .B1(n15124), .B2(n15126), .A(n15123), .ZN(n15125) );
  OAI21_X1 U18369 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15337) );
  AOI21_X1 U18370 ( .B1(n15331), .B2(n15140), .A(n15128), .ZN(n15335) );
  AOI21_X1 U18371 ( .B1(n15131), .B2(n15130), .A(n15115), .ZN(n16180) );
  NAND2_X1 U18372 ( .A1(n19412), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15326) );
  OAI21_X1 U18373 ( .B1(n19423), .B2(n15131), .A(n15326), .ZN(n15132) );
  AOI21_X1 U18374 ( .B1(n19411), .B2(n16180), .A(n15132), .ZN(n15133) );
  OAI21_X1 U18375 ( .B1(n16177), .B2(n16284), .A(n15133), .ZN(n15134) );
  AOI21_X1 U18376 ( .B1(n15335), .B2(n16294), .A(n15134), .ZN(n15135) );
  OAI21_X1 U18377 ( .B1(n19415), .B2(n15337), .A(n15135), .ZN(P2_U2989) );
  XNOR2_X1 U18378 ( .A(n10507), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15137) );
  XNOR2_X1 U18379 ( .A(n10072), .B(n15137), .ZN(n15348) );
  OAI21_X1 U18380 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15138), .A(
        n15130), .ZN(n16111) );
  INV_X1 U18381 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20025) );
  NOR2_X1 U18382 ( .A1(n16334), .A2(n20025), .ZN(n15339) );
  AOI21_X1 U18383 ( .B1(n16270), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15339), .ZN(n15139) );
  OAI21_X1 U18384 ( .B1(n16277), .B2(n16111), .A(n15139), .ZN(n15142) );
  OAI21_X1 U18385 ( .B1(n15146), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15140), .ZN(n15338) );
  NOR2_X1 U18386 ( .A1(n15338), .A2(n19416), .ZN(n15141) );
  AOI211_X1 U18387 ( .C1(n19420), .C2(n16187), .A(n15142), .B(n15141), .ZN(
        n15143) );
  OAI21_X1 U18388 ( .B1(n15348), .B2(n19415), .A(n15143), .ZN(P2_U2990) );
  XNOR2_X1 U18389 ( .A(n15145), .B(n15144), .ZN(n15362) );
  AOI21_X1 U18390 ( .B1(n9883), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15147) );
  NOR2_X1 U18391 ( .A1(n15147), .A2(n15146), .ZN(n15349) );
  AOI22_X1 U18392 ( .A1(n16270), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19412), .ZN(n15150) );
  AOI21_X1 U18393 ( .B1(n15148), .B2(n12778), .A(n15138), .ZN(n16199) );
  NAND2_X1 U18394 ( .A1(n19411), .A2(n16199), .ZN(n15149) );
  OAI211_X1 U18395 ( .C1(n15151), .C2(n16284), .A(n15150), .B(n15149), .ZN(
        n15152) );
  AOI21_X1 U18396 ( .B1(n15349), .B2(n16294), .A(n15152), .ZN(n15153) );
  OAI21_X1 U18397 ( .B1(n15362), .B2(n19415), .A(n15153), .ZN(P2_U2991) );
  INV_X1 U18398 ( .A(n15447), .ZN(n16222) );
  OAI21_X1 U18399 ( .B1(n16224), .B2(n16222), .A(n15154), .ZN(n15155) );
  NAND2_X1 U18400 ( .A1(n15155), .A2(n16220), .ZN(n15215) );
  OAI21_X1 U18401 ( .B1(n15215), .B2(n15214), .A(n15156), .ZN(n15209) );
  NAND2_X1 U18402 ( .A1(n15158), .A2(n15157), .ZN(n15208) );
  OR2_X1 U18403 ( .A1(n15174), .A2(n15175), .ZN(n15178) );
  INV_X1 U18404 ( .A(n15177), .ZN(n15160) );
  NAND2_X1 U18405 ( .A1(n15178), .A2(n15160), .ZN(n15165) );
  INV_X1 U18406 ( .A(n15161), .ZN(n15163) );
  NAND2_X1 U18407 ( .A1(n15163), .A2(n15162), .ZN(n15164) );
  XNOR2_X1 U18408 ( .A(n15165), .B(n15164), .ZN(n15389) );
  INV_X1 U18409 ( .A(n15166), .ZN(n15377) );
  NAND2_X1 U18410 ( .A1(n15195), .A2(n15377), .ZN(n15173) );
  AOI21_X1 U18411 ( .B1(n15378), .B2(n15173), .A(n9883), .ZN(n15387) );
  NAND2_X1 U18412 ( .A1(n19412), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15379) );
  OAI21_X1 U18413 ( .B1(n19423), .B2(n15167), .A(n15379), .ZN(n15168) );
  AOI21_X1 U18414 ( .B1(n19411), .B2(n15169), .A(n15168), .ZN(n15170) );
  OAI21_X1 U18415 ( .B1(n15385), .B2(n16284), .A(n15170), .ZN(n15171) );
  AOI21_X1 U18416 ( .B1(n15387), .B2(n16294), .A(n15171), .ZN(n15172) );
  OAI21_X1 U18417 ( .B1(n15389), .B2(n19415), .A(n15172), .ZN(P2_U2993) );
  NAND2_X1 U18418 ( .A1(n15195), .A2(n15392), .ZN(n15197) );
  NOR2_X1 U18419 ( .A1(n15197), .A2(n15189), .ZN(n15188) );
  OAI21_X1 U18420 ( .B1(n15188), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15173), .ZN(n15400) );
  OAI21_X1 U18421 ( .B1(n15177), .B2(n15175), .A(n15174), .ZN(n15176) );
  OAI21_X1 U18422 ( .B1(n15178), .B2(n15177), .A(n15176), .ZN(n15390) );
  NAND2_X1 U18423 ( .A1(n15390), .A2(n16293), .ZN(n15183) );
  INV_X1 U18424 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20017) );
  NOR2_X1 U18425 ( .A1(n16334), .A2(n20017), .ZN(n15394) );
  AOI21_X1 U18426 ( .B1(n16270), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15394), .ZN(n15179) );
  OAI21_X1 U18427 ( .B1(n16277), .B2(n15180), .A(n15179), .ZN(n15181) );
  AOI21_X1 U18428 ( .B1(n19062), .B2(n19420), .A(n15181), .ZN(n15182) );
  OAI211_X1 U18429 ( .C1(n19416), .C2(n15400), .A(n15183), .B(n15182), .ZN(
        P2_U2994) );
  NAND2_X1 U18430 ( .A1(n15185), .A2(n15184), .ZN(n15187) );
  OAI21_X1 U18431 ( .B1(n15200), .B2(n15198), .A(n15199), .ZN(n15186) );
  XOR2_X1 U18432 ( .A(n15187), .B(n15186), .Z(n15410) );
  AOI21_X1 U18433 ( .B1(n15189), .B2(n15197), .A(n15188), .ZN(n15408) );
  AOI22_X1 U18434 ( .A1(n16270), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19412), .ZN(n15191) );
  NAND2_X1 U18435 ( .A1(n19411), .A2(n19066), .ZN(n15190) );
  OAI211_X1 U18436 ( .C1(n15192), .C2(n16284), .A(n15191), .B(n15190), .ZN(
        n15193) );
  AOI21_X1 U18437 ( .B1(n15408), .B2(n16294), .A(n15193), .ZN(n15194) );
  OAI21_X1 U18438 ( .B1(n15410), .B2(n19415), .A(n15194), .ZN(P2_U2995) );
  INV_X1 U18439 ( .A(n15411), .ZN(n15196) );
  NOR2_X1 U18440 ( .A1(n15211), .A2(n15415), .ZN(n15210) );
  OAI21_X1 U18441 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15210), .A(
        n15197), .ZN(n16312) );
  NAND2_X1 U18442 ( .A1(n10240), .A2(n15199), .ZN(n15201) );
  XOR2_X1 U18443 ( .A(n15201), .B(n15200), .Z(n16309) );
  NAND2_X1 U18444 ( .A1(n16309), .A2(n16293), .ZN(n15206) );
  OAI22_X1 U18445 ( .A1(n20013), .A2(n16334), .B1(n16277), .B2(n15202), .ZN(
        n15204) );
  NOR2_X1 U18446 ( .A1(n16308), .A2(n16284), .ZN(n15203) );
  AOI211_X1 U18447 ( .C1(n16270), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15204), .B(n15203), .ZN(n15205) );
  OAI211_X1 U18448 ( .C1(n19416), .C2(n16312), .A(n15206), .B(n15205), .ZN(
        P2_U2996) );
  AOI21_X1 U18449 ( .B1(n15209), .B2(n15208), .A(n15207), .ZN(n15426) );
  AND2_X1 U18450 ( .A1(n19412), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15423) );
  OAI21_X1 U18451 ( .B1(n15426), .B2(n19415), .A(n15213), .ZN(P2_U2997) );
  XNOR2_X1 U18452 ( .A(n15215), .B(n15214), .ZN(n15434) );
  INV_X1 U18453 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15216) );
  OAI22_X1 U18454 ( .A1(n15216), .A2(n19423), .B1(n16277), .B2(n19104), .ZN(
        n15221) );
  NOR2_X1 U18455 ( .A1(n20009), .A2(n16334), .ZN(n15220) );
  INV_X1 U18456 ( .A(n9892), .ZN(n16228) );
  NOR2_X1 U18457 ( .A1(n16318), .A2(n16228), .ZN(n16227) );
  INV_X1 U18458 ( .A(n16227), .ZN(n15218) );
  INV_X1 U18459 ( .A(n15415), .ZN(n15217) );
  AOI211_X1 U18460 ( .C1(n15430), .C2(n15218), .A(n15217), .B(n19416), .ZN(
        n15219) );
  NOR3_X1 U18461 ( .A1(n15221), .A2(n15220), .A3(n15219), .ZN(n15223) );
  NAND2_X1 U18462 ( .A1(n19105), .A2(n19420), .ZN(n15222) );
  OAI211_X1 U18463 ( .C1(n15434), .C2(n19415), .A(n15223), .B(n15222), .ZN(
        P2_U2998) );
  XNOR2_X1 U18464 ( .A(n15226), .B(n16358), .ZN(n16370) );
  NAND2_X1 U18465 ( .A1(n15498), .A2(n15497), .ZN(n15228) );
  XNOR2_X1 U18466 ( .A(n15227), .B(n15228), .ZN(n16368) );
  INV_X1 U18467 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15229) );
  OAI22_X1 U18468 ( .A1(n15229), .A2(n19423), .B1(n16277), .B2(n19201), .ZN(
        n15230) );
  AOI21_X1 U18469 ( .B1(n19412), .B2(P2_REIP_REG_7__SCAN_IN), .A(n15230), .ZN(
        n15231) );
  OAI21_X1 U18470 ( .B1(n19206), .B2(n16284), .A(n15231), .ZN(n15232) );
  AOI21_X1 U18471 ( .B1(n16368), .B2(n16293), .A(n15232), .ZN(n15233) );
  OAI21_X1 U18472 ( .B1(n16370), .B2(n19416), .A(n15233), .ZN(P2_U3007) );
  INV_X1 U18473 ( .A(n15234), .ZN(n15236) );
  AOI22_X1 U18474 ( .A1(n12510), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12453), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U18475 ( .A1(n12567), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U18476 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  XNOR2_X1 U18477 ( .A(n15240), .B(n15239), .ZN(n19263) );
  NAND2_X1 U18478 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15257) );
  INV_X1 U18479 ( .A(n15257), .ZN(n15241) );
  NOR2_X1 U18480 ( .A1(n16382), .A2(n16371), .ZN(n15504) );
  NAND4_X1 U18481 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n15504), .ZN(n15246) );
  NAND2_X1 U18482 ( .A1(n15252), .A2(n15439), .ZN(n15367) );
  NOR2_X1 U18483 ( .A1(n15350), .A2(n15367), .ZN(n15341) );
  AND2_X1 U18484 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15341), .ZN(
        n15316) );
  NAND2_X1 U18485 ( .A1(n15241), .A2(n15316), .ZN(n15284) );
  INV_X1 U18486 ( .A(n15279), .ZN(n15268) );
  NAND3_X1 U18487 ( .A1(n15242), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15268), .ZN(n15244) );
  OAI21_X1 U18488 ( .B1(n15284), .B2(n15244), .A(n15243), .ZN(n15245) );
  AOI21_X1 U18489 ( .B1(n19263), .B2(n16399), .A(n15245), .ZN(n15263) );
  INV_X1 U18490 ( .A(n15246), .ZN(n15247) );
  NAND2_X1 U18491 ( .A1(n15248), .A2(n15247), .ZN(n15249) );
  NAND2_X1 U18492 ( .A1(n15419), .A2(n15249), .ZN(n15251) );
  INV_X1 U18493 ( .A(n15252), .ZN(n15253) );
  NAND2_X1 U18494 ( .A1(n15419), .A2(n15253), .ZN(n15254) );
  AND2_X1 U18495 ( .A1(n15486), .A2(n15254), .ZN(n15368) );
  AOI21_X1 U18496 ( .B1(n15419), .B2(n15350), .A(n15255), .ZN(n15256) );
  NAND2_X1 U18497 ( .A1(n15368), .A2(n15256), .ZN(n15340) );
  INV_X1 U18498 ( .A(n15419), .ZN(n16410) );
  NAND2_X1 U18499 ( .A1(n15486), .A2(n16410), .ZN(n15258) );
  NAND2_X1 U18500 ( .A1(n15340), .A2(n15258), .ZN(n15332) );
  NAND2_X1 U18501 ( .A1(n15258), .A2(n15257), .ZN(n15259) );
  NAND2_X1 U18502 ( .A1(n15332), .A2(n15259), .ZN(n15308) );
  AND2_X1 U18503 ( .A1(n15419), .A2(n15279), .ZN(n15260) );
  OR2_X1 U18504 ( .A1(n15308), .A2(n15260), .ZN(n15273) );
  AND2_X1 U18505 ( .A1(n15419), .A2(n15269), .ZN(n15261) );
  OAI21_X1 U18506 ( .B1(n15273), .B2(n15261), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15262) );
  OAI211_X1 U18507 ( .C1(n16115), .C2(n16365), .A(n15263), .B(n15262), .ZN(
        n15264) );
  AOI21_X1 U18508 ( .B1(n15265), .B2(n16393), .A(n15264), .ZN(n15266) );
  OAI21_X1 U18509 ( .B1(n15267), .B2(n16402), .A(n15266), .ZN(P2_U3015) );
  INV_X1 U18510 ( .A(n15284), .ZN(n15303) );
  NAND3_X1 U18511 ( .A1(n15303), .A2(n15269), .A3(n15268), .ZN(n15271) );
  OAI211_X1 U18512 ( .C1(n16119), .C2(n16364), .A(n15271), .B(n15270), .ZN(
        n15272) );
  OAI21_X1 U18513 ( .B1(n16120), .B2(n16365), .A(n15274), .ZN(n15275) );
  AOI21_X1 U18514 ( .B1(n15276), .B2(n16393), .A(n15275), .ZN(n15277) );
  OAI21_X1 U18515 ( .B1(n15278), .B2(n16402), .A(n15277), .ZN(P2_U3016) );
  AND2_X1 U18516 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U18517 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15280), .A(
        n15279), .ZN(n15283) );
  NAND2_X1 U18518 ( .A1(n16133), .A2(n16399), .ZN(n15282) );
  OAI211_X1 U18519 ( .C1(n15284), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        n15285) );
  OAI21_X1 U18520 ( .B1(n16131), .B2(n16365), .A(n15286), .ZN(n15287) );
  AOI21_X1 U18521 ( .B1(n15288), .B2(n16393), .A(n15287), .ZN(n15289) );
  OAI21_X1 U18522 ( .B1(n15290), .B2(n16402), .A(n15289), .ZN(P2_U3017) );
  XNOR2_X1 U18523 ( .A(n15302), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15292) );
  AOI21_X1 U18524 ( .B1(n15303), .B2(n15292), .A(n15291), .ZN(n15293) );
  OAI21_X1 U18525 ( .B1(n15294), .B2(n16364), .A(n15293), .ZN(n15295) );
  AOI21_X1 U18526 ( .B1(n15308), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15295), .ZN(n15296) );
  OAI21_X1 U18527 ( .B1(n16140), .B2(n16365), .A(n15296), .ZN(n15297) );
  AOI21_X1 U18528 ( .B1(n15298), .B2(n16393), .A(n15297), .ZN(n15299) );
  OAI21_X1 U18529 ( .B1(n15300), .B2(n16402), .A(n15299), .ZN(P2_U3018) );
  NAND3_X1 U18530 ( .A1(n15100), .A2(n16379), .A3(n15301), .ZN(n15313) );
  NAND2_X1 U18531 ( .A1(n15303), .A2(n15302), .ZN(n15304) );
  OAI211_X1 U18532 ( .C1(n16364), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15307) );
  AOI21_X1 U18533 ( .B1(n15308), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15307), .ZN(n15309) );
  OAI21_X1 U18534 ( .B1(n16158), .B2(n16365), .A(n15309), .ZN(n15310) );
  AOI21_X1 U18535 ( .B1(n15311), .B2(n16393), .A(n15310), .ZN(n15312) );
  NAND2_X1 U18536 ( .A1(n15313), .A2(n15312), .ZN(P2_U3019) );
  NOR2_X1 U18537 ( .A1(n15332), .A2(n15315), .ZN(n15322) );
  INV_X1 U18538 ( .A(n15316), .ZN(n15327) );
  XNOR2_X1 U18539 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U18540 ( .A1(n15317), .A2(n16399), .ZN(n15319) );
  OAI211_X1 U18541 ( .C1(n15327), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        n15321) );
  AOI211_X1 U18542 ( .C1(n16172), .C2(n16407), .A(n15322), .B(n15321), .ZN(
        n15323) );
  OAI211_X1 U18543 ( .C1(n15325), .C2(n16404), .A(n15324), .B(n15323), .ZN(
        P2_U3020) );
  NOR2_X1 U18544 ( .A1(n16177), .A2(n16365), .ZN(n15334) );
  OAI21_X1 U18545 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15327), .A(
        n15326), .ZN(n15328) );
  AOI21_X1 U18546 ( .B1(n16399), .B2(n15329), .A(n15328), .ZN(n15330) );
  OAI21_X1 U18547 ( .B1(n15332), .B2(n15331), .A(n15330), .ZN(n15333) );
  AOI211_X1 U18548 ( .C1(n15335), .C2(n16393), .A(n15334), .B(n15333), .ZN(
        n15336) );
  OAI21_X1 U18549 ( .B1(n16402), .B2(n15337), .A(n15336), .ZN(P2_U3021) );
  INV_X1 U18550 ( .A(n15338), .ZN(n15346) );
  AOI21_X1 U18551 ( .B1(n16399), .B2(n16186), .A(n15339), .ZN(n15343) );
  OAI21_X1 U18552 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15341), .A(
        n15340), .ZN(n15342) );
  OAI211_X1 U18553 ( .C1(n15344), .C2(n16365), .A(n15343), .B(n15342), .ZN(
        n15345) );
  AOI21_X1 U18554 ( .B1(n15346), .B2(n16393), .A(n15345), .ZN(n15347) );
  OAI21_X1 U18555 ( .B1(n15348), .B2(n16402), .A(n15347), .ZN(P2_U3022) );
  NAND2_X1 U18556 ( .A1(n15349), .A2(n16393), .ZN(n15361) );
  OAI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15350), .ZN(n15351) );
  OAI22_X1 U18558 ( .A1(n15368), .A2(n15352), .B1(n15367), .B2(n15351), .ZN(
        n15359) );
  OR2_X1 U18559 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  AND2_X1 U18560 ( .A1(n15356), .A2(n15355), .ZN(n16208) );
  INV_X1 U18561 ( .A(n16208), .ZN(n15357) );
  INV_X1 U18562 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20023) );
  OAI22_X1 U18563 ( .A1(n16364), .A2(n15357), .B1(n20023), .B2(n16334), .ZN(
        n15358) );
  AOI211_X1 U18564 ( .C1(n16196), .C2(n16407), .A(n15359), .B(n15358), .ZN(
        n15360) );
  OAI211_X1 U18565 ( .C1(n15362), .C2(n16402), .A(n15361), .B(n15360), .ZN(
        P2_U3023) );
  NAND2_X1 U18566 ( .A1(n10064), .A2(n15364), .ZN(n15365) );
  XNOR2_X1 U18567 ( .A(n15366), .B(n15365), .ZN(n16213) );
  INV_X1 U18568 ( .A(n15367), .ZN(n15371) );
  INV_X1 U18569 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15370) );
  INV_X1 U18570 ( .A(n15368), .ZN(n15383) );
  NOR2_X1 U18571 ( .A1(n20021), .A2(n16334), .ZN(n15369) );
  AOI221_X1 U18572 ( .B1(n15371), .B2(n15370), .C1(n15383), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15369), .ZN(n15372) );
  OAI21_X1 U18573 ( .B1(n16364), .B2(n15373), .A(n15372), .ZN(n15375) );
  XNOR2_X1 U18574 ( .A(n9883), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16214) );
  NOR2_X1 U18575 ( .A1(n16214), .A2(n16404), .ZN(n15374) );
  AOI211_X1 U18576 ( .C1(n16407), .C2(n16216), .A(n15375), .B(n15374), .ZN(
        n15376) );
  OAI21_X1 U18577 ( .B1(n16213), .B2(n16402), .A(n15376), .ZN(P2_U3024) );
  NAND3_X1 U18578 ( .A1(n15439), .A2(n15378), .A3(n15377), .ZN(n15380) );
  OAI211_X1 U18579 ( .C1(n16364), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        n15382) );
  AOI21_X1 U18580 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15383), .A(
        n15382), .ZN(n15384) );
  OAI21_X1 U18581 ( .B1(n15385), .B2(n16365), .A(n15384), .ZN(n15386) );
  AOI21_X1 U18582 ( .B1(n15387), .B2(n16393), .A(n15386), .ZN(n15388) );
  OAI21_X1 U18583 ( .B1(n15389), .B2(n16402), .A(n15388), .ZN(P2_U3025) );
  NAND2_X1 U18584 ( .A1(n15390), .A2(n16379), .ZN(n15399) );
  INV_X1 U18585 ( .A(n15439), .ZN(n15487) );
  NOR2_X1 U18586 ( .A1(n15413), .A2(n15487), .ZN(n16301) );
  INV_X1 U18587 ( .A(n16301), .ZN(n16319) );
  OR2_X1 U18588 ( .A1(n15391), .A2(n16319), .ZN(n15406) );
  XNOR2_X1 U18589 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15396) );
  OAI21_X1 U18590 ( .B1(n16410), .B2(n15392), .A(n15486), .ZN(n15403) );
  NOR2_X1 U18591 ( .A1(n16364), .A2(n19059), .ZN(n15393) );
  AOI211_X1 U18592 ( .C1(n15403), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15394), .B(n15393), .ZN(n15395) );
  OAI21_X1 U18593 ( .B1(n15406), .B2(n15396), .A(n15395), .ZN(n15397) );
  AOI21_X1 U18594 ( .B1(n19062), .B2(n16407), .A(n15397), .ZN(n15398) );
  OAI211_X1 U18595 ( .C1(n15400), .C2(n16404), .A(n15399), .B(n15398), .ZN(
        P2_U3026) );
  NAND2_X1 U18596 ( .A1(n19072), .A2(n16407), .ZN(n15405) );
  INV_X1 U18597 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20015) );
  NOR2_X1 U18598 ( .A1(n20015), .A2(n16334), .ZN(n15402) );
  NOR2_X1 U18599 ( .A1(n16364), .A2(n19074), .ZN(n15401) );
  AOI211_X1 U18600 ( .C1(n15403), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15402), .B(n15401), .ZN(n15404) );
  OAI211_X1 U18601 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15406), .A(
        n15405), .B(n15404), .ZN(n15407) );
  AOI21_X1 U18602 ( .B1(n15408), .B2(n16393), .A(n15407), .ZN(n15409) );
  OAI21_X1 U18603 ( .B1(n15410), .B2(n16402), .A(n15409), .ZN(P2_U3027) );
  AOI21_X1 U18604 ( .B1(n16393), .B2(n9892), .A(n16301), .ZN(n15427) );
  NOR2_X1 U18605 ( .A1(n15427), .A2(n15411), .ZN(n15420) );
  INV_X1 U18606 ( .A(n15486), .ZN(n15412) );
  AOI21_X1 U18607 ( .B1(n15413), .B2(n15419), .A(n15412), .ZN(n16317) );
  INV_X1 U18608 ( .A(n15414), .ZN(n15416) );
  OAI21_X1 U18609 ( .B1(n15416), .B2(n16393), .A(n15415), .ZN(n15417) );
  OAI211_X1 U18610 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15418), .A(
        n16317), .B(n15417), .ZN(n15429) );
  INV_X1 U18611 ( .A(n15421), .ZN(n15425) );
  NOR2_X1 U18612 ( .A1(n19095), .A2(n16365), .ZN(n15422) );
  AOI211_X1 U18613 ( .C1(n16399), .C2(n19089), .A(n15423), .B(n15422), .ZN(
        n15424) );
  OAI211_X1 U18614 ( .C1(n15426), .C2(n16402), .A(n15425), .B(n15424), .ZN(
        P2_U3029) );
  OAI21_X1 U18615 ( .B1(n16318), .B2(n15427), .A(n15430), .ZN(n15428) );
  OAI21_X1 U18616 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15433) );
  OAI22_X1 U18617 ( .A1(n16364), .A2(n19108), .B1(n20009), .B2(n16334), .ZN(
        n15431) );
  AOI21_X1 U18618 ( .B1(n19105), .B2(n16407), .A(n15431), .ZN(n15432) );
  OAI211_X1 U18619 ( .C1(n15434), .C2(n16402), .A(n15433), .B(n15432), .ZN(
        P2_U3030) );
  INV_X1 U18620 ( .A(n16349), .ZN(n15435) );
  NOR2_X1 U18621 ( .A1(n15442), .A2(n15452), .ZN(n16240) );
  OAI21_X1 U18622 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16240), .A(
        n16228), .ZN(n16234) );
  OR2_X1 U18623 ( .A1(n15437), .A2(n9933), .ZN(n15438) );
  NAND2_X1 U18624 ( .A1(n15438), .A2(n16314), .ZN(n19274) );
  OAI21_X1 U18625 ( .B1(n15440), .B2(n16410), .A(n15486), .ZN(n16327) );
  INV_X1 U18626 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20005) );
  NOR2_X1 U18627 ( .A1(n20005), .A2(n16334), .ZN(n15445) );
  NAND2_X1 U18628 ( .A1(n15440), .A2(n15439), .ZN(n16325) );
  AOI211_X1 U18629 ( .C1(n15443), .C2(n15442), .A(n15441), .B(n16325), .ZN(
        n15444) );
  AOI211_X1 U18630 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16327), .A(
        n15445), .B(n15444), .ZN(n15446) );
  OAI21_X1 U18631 ( .B1(n16364), .B2(n19274), .A(n15446), .ZN(n15450) );
  NAND2_X1 U18632 ( .A1(n15447), .A2(n16223), .ZN(n15448) );
  XNOR2_X1 U18633 ( .A(n16224), .B(n15448), .ZN(n16233) );
  NOR2_X1 U18634 ( .A1(n16233), .A2(n16402), .ZN(n15449) );
  AOI211_X1 U18635 ( .C1(n16407), .C2(n19128), .A(n15450), .B(n15449), .ZN(
        n15451) );
  OAI21_X1 U18636 ( .B1(n16234), .B2(n16404), .A(n15451), .ZN(P2_U3032) );
  NAND2_X1 U18637 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16263), .ZN(
        n16241) );
  INV_X1 U18638 ( .A(n16242), .ZN(n15453) );
  NOR2_X1 U18639 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  XNOR2_X1 U18640 ( .A(n15456), .B(n15455), .ZN(n16253) );
  NOR2_X1 U18641 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16325), .ZN(
        n16328) );
  INV_X1 U18642 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20001) );
  NOR2_X1 U18643 ( .A1(n20001), .A2(n16334), .ZN(n15457) );
  AOI211_X1 U18644 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16327), .A(
        n16328), .B(n15457), .ZN(n15462) );
  OR2_X1 U18645 ( .A1(n15458), .A2(n16341), .ZN(n15459) );
  NAND2_X1 U18646 ( .A1(n15459), .A2(n16331), .ZN(n19277) );
  INV_X1 U18647 ( .A(n19277), .ZN(n15460) );
  AOI22_X1 U18648 ( .A1(n19150), .A2(n16407), .B1(n16399), .B2(n15460), .ZN(
        n15461) );
  OAI211_X1 U18649 ( .C1(n16253), .C2(n16402), .A(n15462), .B(n15461), .ZN(
        n15463) );
  INV_X1 U18650 ( .A(n15463), .ZN(n15464) );
  OAI21_X1 U18651 ( .B1(n16254), .B2(n16404), .A(n15464), .ZN(P2_U3034) );
  NAND2_X1 U18652 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15480), .ZN(
        n16264) );
  OAI21_X1 U18653 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15480), .A(
        n16264), .ZN(n16272) );
  INV_X1 U18654 ( .A(n15465), .ZN(n15481) );
  OR2_X1 U18655 ( .A1(n9919), .A2(n15481), .ZN(n15469) );
  AND2_X1 U18656 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  XNOR2_X1 U18657 ( .A(n15469), .B(n15468), .ZN(n16271) );
  NOR2_X1 U18658 ( .A1(n14939), .A2(n15487), .ZN(n16350) );
  OAI21_X1 U18659 ( .B1(n16410), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15486), .ZN(n16344) );
  INV_X1 U18660 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19997) );
  NOR2_X1 U18661 ( .A1(n19997), .A2(n16334), .ZN(n15470) );
  AOI221_X1 U18662 ( .B1(n16350), .B2(n15471), .C1(n16344), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15470), .ZN(n15477) );
  OR2_X1 U18663 ( .A1(n15472), .A2(n15488), .ZN(n15473) );
  NAND2_X1 U18664 ( .A1(n15473), .A2(n16342), .ZN(n19281) );
  OAI22_X1 U18665 ( .A1(n15474), .A2(n16365), .B1(n16364), .B2(n19281), .ZN(
        n15475) );
  INV_X1 U18666 ( .A(n15475), .ZN(n15476) );
  OAI211_X1 U18667 ( .C1(n16271), .C2(n16402), .A(n15477), .B(n15476), .ZN(
        n15478) );
  INV_X1 U18668 ( .A(n15478), .ZN(n15479) );
  OAI21_X1 U18669 ( .B1(n16272), .B2(n16404), .A(n15479), .ZN(P2_U3036) );
  NOR2_X1 U18670 ( .A1(n15482), .A2(n15481), .ZN(n15483) );
  XNOR2_X1 U18671 ( .A(n15484), .B(n15483), .ZN(n16280) );
  NAND2_X1 U18672 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19412), .ZN(n15485) );
  OAI221_X1 U18673 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15487), .C1(
        n14939), .C2(n15486), .A(n15485), .ZN(n15492) );
  AOI21_X1 U18674 ( .B1(n15489), .B2(n15508), .A(n15488), .ZN(n19283) );
  INV_X1 U18675 ( .A(n19283), .ZN(n15490) );
  OAI22_X1 U18676 ( .A1(n19182), .A2(n16365), .B1(n16364), .B2(n15490), .ZN(
        n15491) );
  AOI211_X1 U18677 ( .C1(n16280), .C2(n16379), .A(n15492), .B(n15491), .ZN(
        n15493) );
  OAI21_X1 U18678 ( .B1(n10269), .B2(n16404), .A(n15493), .ZN(P2_U3037) );
  OAI21_X1 U18679 ( .B1(n15496), .B2(n15495), .A(n15494), .ZN(n16286) );
  NAND2_X1 U18680 ( .A1(n15227), .A2(n15497), .ZN(n15499) );
  NAND2_X1 U18681 ( .A1(n15499), .A2(n15498), .ZN(n15503) );
  AND2_X1 U18682 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  XNOR2_X1 U18683 ( .A(n15503), .B(n15502), .ZN(n16285) );
  OAI21_X1 U18684 ( .B1(n16410), .B2(n15504), .A(n16372), .ZN(n16355) );
  INV_X1 U18685 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19993) );
  NOR2_X1 U18686 ( .A1(n19993), .A2(n16334), .ZN(n15506) );
  NAND2_X1 U18687 ( .A1(n15504), .A2(n16383), .ZN(n16359) );
  AOI221_X1 U18688 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n16358), .C2(n14922), .A(
        n16359), .ZN(n15505) );
  AOI211_X1 U18689 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16355), .A(
        n15506), .B(n15505), .ZN(n15512) );
  OR2_X1 U18690 ( .A1(n15507), .A2(n16360), .ZN(n15509) );
  NAND2_X1 U18691 ( .A1(n15509), .A2(n15508), .ZN(n19288) );
  INV_X1 U18692 ( .A(n19288), .ZN(n15510) );
  AOI22_X1 U18693 ( .A1(n19193), .A2(n16407), .B1(n16399), .B2(n15510), .ZN(
        n15511) );
  OAI211_X1 U18694 ( .C1(n16285), .C2(n16402), .A(n15512), .B(n15511), .ZN(
        n15513) );
  INV_X1 U18695 ( .A(n15513), .ZN(n15514) );
  OAI21_X1 U18696 ( .B1(n16286), .B2(n16404), .A(n15514), .ZN(P2_U3038) );
  AOI22_X1 U18697 ( .A1(n15516), .A2(n15517), .B1(n13768), .B2(n15515), .ZN(
        n15521) );
  AND3_X1 U18698 ( .A1(n15519), .A2(n15518), .A3(n15517), .ZN(n15520) );
  MUX2_X1 U18699 ( .A(n15521), .B(n15520), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15522) );
  NAND2_X1 U18700 ( .A1(n15522), .A2(n10501), .ZN(n15523) );
  AOI21_X1 U18701 ( .B1(n13396), .B2(n15524), .A(n15523), .ZN(n16411) );
  OAI22_X1 U18702 ( .A1(n15526), .A2(n15525), .B1(n16411), .B2(n20054), .ZN(
        n15528) );
  MUX2_X1 U18703 ( .A(n15528), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15527), .Z(P2_U3596) );
  AOI22_X1 U18704 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15529) );
  OAI21_X1 U18705 ( .B1(n17339), .B2(n17143), .A(n15529), .ZN(n15540) );
  AOI22_X1 U18706 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15537) );
  AOI22_X1 U18707 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15530) );
  OAI21_X1 U18708 ( .B1(n17275), .B2(n15531), .A(n15530), .ZN(n15535) );
  AOI22_X1 U18709 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18710 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17351), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15532) );
  OAI211_X1 U18711 ( .C1(n13966), .C2(n17373), .A(n15533), .B(n15532), .ZN(
        n15534) );
  AOI211_X1 U18712 ( .C1(n17335), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15535), .B(n15534), .ZN(n15536) );
  OAI211_X1 U18713 ( .C1(n15538), .C2(n15653), .A(n15537), .B(n15536), .ZN(
        n15539) );
  AOI211_X1 U18714 ( .C1(n17328), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n15540), .B(n15539), .ZN(n17491) );
  INV_X1 U18715 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16940) );
  INV_X1 U18716 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16960) );
  INV_X1 U18717 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16989) );
  INV_X1 U18718 ( .A(n17399), .ZN(n17384) );
  NAND2_X1 U18719 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17375), .ZN(n17368) );
  NAND2_X1 U18720 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17344), .ZN(n17321) );
  NAND2_X1 U18721 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17343), .ZN(n17318) );
  NAND2_X1 U18722 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17306), .ZN(n15541) );
  NOR2_X1 U18723 ( .A1(n18400), .A2(n15541), .ZN(n17288) );
  INV_X1 U18724 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16882) );
  NOR2_X1 U18725 ( .A1(n17396), .A2(n16882), .ZN(n15542) );
  OAI22_X1 U18726 ( .A1(n17288), .A2(n15542), .B1(n15541), .B2(n16882), .ZN(
        n15543) );
  OAI21_X1 U18727 ( .B1(n17491), .B2(n17390), .A(n15543), .ZN(P3_U2690) );
  NOR2_X1 U18728 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18960), .ZN(
        n18408) );
  INV_X1 U18729 ( .A(n18408), .ZN(n15544) );
  NAND3_X1 U18730 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18959)
         );
  INV_X1 U18731 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16999) );
  OAI21_X1 U18732 ( .B1(n18828), .B2(n18967), .A(n16999), .ZN(n15584) );
  NOR2_X1 U18733 ( .A1(n15677), .A2(n15584), .ZN(n18362) );
  INV_X1 U18734 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16651) );
  OR2_X1 U18735 ( .A1(n16651), .A2(n18959), .ZN(n15583) );
  OAI211_X1 U18736 ( .C1(n18959), .C2(n18362), .A(n18455), .B(n15583), .ZN(
        n18368) );
  NAND2_X1 U18737 ( .A1(n15544), .A2(n18368), .ZN(n15547) );
  INV_X1 U18738 ( .A(n15547), .ZN(n15546) );
  NOR3_X1 U18739 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19011), .ZN(n16476) );
  INV_X1 U18740 ( .A(n16476), .ZN(n18712) );
  NOR2_X1 U18741 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18984) );
  INV_X1 U18742 ( .A(n18984), .ZN(n19022) );
  NAND2_X1 U18743 ( .A1(n18856), .A2(n18960), .ZN(n16644) );
  NAND2_X1 U18744 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17989) );
  INV_X1 U18745 ( .A(n17989), .ZN(n17923) );
  OAI22_X1 U18746 ( .A1(n19004), .A2(n17923), .B1(n18822), .B2(n18960), .ZN(
        n15549) );
  NAND3_X1 U18747 ( .A1(n18823), .A2(n18368), .A3(n15549), .ZN(n15545) );
  OAI221_X1 U18748 ( .B1(n18823), .B2(n15546), .C1(n18823), .C2(n18712), .A(
        n15545), .ZN(P3_U2864) );
  NAND2_X1 U18749 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18522) );
  NOR2_X1 U18750 ( .A1(n19004), .A2(n17923), .ZN(n15548) );
  AOI221_X1 U18751 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18522), .C1(n15548), 
        .C2(n18522), .A(n15547), .ZN(n18367) );
  OAI221_X1 U18752 ( .B1(n16476), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n16476), .C2(n15549), .A(n18368), .ZN(n18365) );
  AOI22_X1 U18753 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18367), .B1(
        n18365), .B2(n18373), .ZN(P3_U2865) );
  NAND3_X1 U18754 ( .A1(n15727), .A2(n15719), .A3(n15725), .ZN(n15552) );
  NAND2_X1 U18755 ( .A1(n10113), .A2(n17590), .ZN(n15571) );
  NOR2_X1 U18756 ( .A1(n15550), .A2(n15719), .ZN(n15554) );
  NAND4_X1 U18757 ( .A1(n15559), .A2(n15725), .A3(n15564), .A4(n15554), .ZN(
        n15560) );
  NAND2_X1 U18758 ( .A1(n15719), .A2(n18393), .ZN(n18817) );
  AND2_X1 U18759 ( .A1(n18400), .A2(n18817), .ZN(n15857) );
  NOR3_X1 U18760 ( .A1(n16997), .A2(n15857), .A3(n10113), .ZN(n15579) );
  AOI21_X1 U18761 ( .B1(n15551), .B2(n15552), .A(n15579), .ZN(n15558) );
  INV_X1 U18762 ( .A(n15551), .ZN(n15730) );
  NAND2_X1 U18763 ( .A1(n15730), .A2(n18397), .ZN(n15724) );
  AOI21_X1 U18764 ( .B1(n15552), .B2(n15724), .A(n18372), .ZN(n15557) );
  OAI22_X1 U18765 ( .A1(n15564), .A2(n18385), .B1(n18389), .B2(n18817), .ZN(
        n15556) );
  INV_X1 U18766 ( .A(n15727), .ZN(n18381) );
  AOI21_X1 U18767 ( .B1(n16997), .B2(n10113), .A(n18381), .ZN(n15574) );
  OAI21_X1 U18768 ( .B1(n15554), .B2(n17445), .A(n18389), .ZN(n15553) );
  OAI21_X1 U18769 ( .B1(n15554), .B2(n15574), .A(n15553), .ZN(n15555) );
  INV_X1 U18770 ( .A(n15571), .ZN(n15561) );
  INV_X1 U18771 ( .A(n15562), .ZN(n15563) );
  NAND3_X1 U18772 ( .A1(n15564), .A2(n19012), .A3(n15563), .ZN(n15565) );
  NAND2_X1 U18773 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19013) );
  OAI21_X1 U18774 ( .B1(n15570), .B2(n15569), .A(n15567), .ZN(n15568) );
  NAND2_X1 U18775 ( .A1(n18799), .A2(n19013), .ZN(n15580) );
  NAND2_X2 U18776 ( .A1(n18999), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18945) );
  INV_X1 U18777 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n16640) );
  NAND2_X1 U18778 ( .A1(n16640), .A2(n18883), .ZN(n18869) );
  NAND3_X1 U18779 ( .A1(n18880), .A2(n18945), .A3(n18869), .ZN(n19010) );
  INV_X1 U18780 ( .A(n19010), .ZN(n15729) );
  NAND2_X1 U18781 ( .A1(n15574), .A2(n15573), .ZN(n15575) );
  AOI21_X1 U18782 ( .B1(n15720), .B2(n15577), .A(n15576), .ZN(n15578) );
  OAI21_X1 U18783 ( .B1(n15580), .B2(n17551), .A(n15735), .ZN(n15581) );
  INV_X1 U18784 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U18785 ( .A1(n18957), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18370) );
  INV_X1 U18786 ( .A(n15584), .ZN(n15585) );
  NOR2_X1 U18787 ( .A1(n15585), .A2(n16666), .ZN(n18806) );
  NAND3_X1 U18788 ( .A1(n18986), .A2(n18984), .A3(n18806), .ZN(n15586) );
  OAI21_X1 U18789 ( .B1(n18986), .B2(n16999), .A(n15586), .ZN(P3_U3284) );
  INV_X1 U18790 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U18791 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15596) );
  INV_X1 U18792 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U18793 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18794 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15587) );
  OAI211_X1 U18795 ( .C1(n13966), .C2(n17261), .A(n15588), .B(n15587), .ZN(
        n15594) );
  AOI22_X1 U18796 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U18797 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15591) );
  AOI22_X1 U18798 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15590) );
  NAND2_X1 U18799 ( .A1(n17335), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n15589) );
  NAND4_X1 U18800 ( .A1(n15592), .A2(n15591), .A3(n15590), .A4(n15589), .ZN(
        n15593) );
  AOI211_X1 U18801 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n15594), .B(n15593), .ZN(n15595) );
  OAI211_X1 U18802 ( .C1(n13933), .C2(n17069), .A(n15596), .B(n15595), .ZN(
        n17954) );
  AOI22_X1 U18803 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15597) );
  OAI21_X1 U18804 ( .B1(n17144), .B2(n17381), .A(n15597), .ZN(n15608) );
  AOI22_X1 U18805 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15606) );
  AOI22_X1 U18806 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U18807 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15604) );
  INV_X1 U18808 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17277) );
  OAI22_X1 U18809 ( .A1(n17293), .A2(n17277), .B1(n13933), .B2(n15598), .ZN(
        n15602) );
  INV_X1 U18810 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U18811 ( .A1(n13911), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15599) );
  OAI21_X1 U18812 ( .B1(n17349), .B2(n15600), .A(n15599), .ZN(n15601) );
  NAND4_X1 U18813 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15607) );
  INV_X1 U18814 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U18815 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15620) );
  OAI22_X1 U18816 ( .A1(n17293), .A2(n15610), .B1(n13922), .B2(n17332), .ZN(
        n15617) );
  AOI22_X1 U18817 ( .A1(n15611), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U18818 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15614) );
  NAND3_X1 U18819 ( .A1(n15615), .A2(n15614), .A3(n15613), .ZN(n15616) );
  AOI211_X1 U18820 ( .C1(n15618), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n15617), .B(n15616), .ZN(n15619) );
  AOI22_X1 U18821 ( .A1(n13911), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15621) );
  OAI21_X1 U18822 ( .B1(n13933), .B2(n18693), .A(n15621), .ZN(n15623) );
  AOI22_X1 U18823 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15626) );
  OAI21_X1 U18824 ( .B1(n17144), .B2(n17389), .A(n15626), .ZN(n15629) );
  AOI22_X1 U18825 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15627) );
  OAI21_X1 U18826 ( .B1(n13879), .B2(n17191), .A(n15627), .ZN(n15628) );
  AOI211_X1 U18827 ( .C1(n13852), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n15629), .B(n15628), .ZN(n15639) );
  AOI22_X1 U18828 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15632) );
  INV_X1 U18829 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15630) );
  INV_X1 U18830 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U18831 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U18832 ( .A1(n13911), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15634) );
  OAI211_X1 U18833 ( .C1(n17349), .C2(n15636), .A(n15635), .B(n15634), .ZN(
        n15637) );
  INV_X1 U18834 ( .A(n15637), .ZN(n15638) );
  NAND3_X1 U18835 ( .A1(n15639), .A2(n10500), .A3(n15638), .ZN(n15640) );
  AOI22_X1 U18836 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15650) );
  INV_X1 U18837 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U18838 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18839 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15641) );
  OAI211_X1 U18840 ( .C1(n13966), .C2(n17292), .A(n15642), .B(n15641), .ZN(
        n15648) );
  AOI22_X1 U18841 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18842 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15645) );
  AOI22_X1 U18843 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15644) );
  NAND2_X1 U18844 ( .A1(n17335), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n15643) );
  NAND4_X1 U18845 ( .A1(n15646), .A2(n15645), .A3(n15644), .A4(n15643), .ZN(
        n15647) );
  AOI211_X1 U18846 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15648), .B(n15647), .ZN(n15649) );
  OAI211_X1 U18847 ( .C1(n17144), .C2(n17383), .A(n15650), .B(n15649), .ZN(
        n15687) );
  NAND2_X1 U18848 ( .A1(n15746), .A2(n15687), .ZN(n15691) );
  AOI22_X1 U18849 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18850 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18851 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15651) );
  OAI211_X1 U18852 ( .C1(n17349), .C2(n15653), .A(n15652), .B(n15651), .ZN(
        n15659) );
  AOI22_X1 U18853 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18854 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18855 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U18856 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n15654) );
  NAND4_X1 U18857 ( .A1(n15657), .A2(n15656), .A3(n15655), .A4(n15654), .ZN(
        n15658) );
  AOI211_X1 U18858 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n15659), .B(n15658), .ZN(n15660) );
  NAND2_X1 U18859 ( .A1(n15694), .A2(n15740), .ZN(n15698) );
  AOI22_X1 U18860 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15662) );
  OAI21_X1 U18861 ( .B1(n17339), .B2(n17090), .A(n15662), .ZN(n15672) );
  AOI22_X1 U18862 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18863 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U18864 ( .B1(n17293), .B2(n17240), .A(n15663), .ZN(n15668) );
  INV_X1 U18865 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18866 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18867 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15664) );
  OAI211_X1 U18868 ( .C1(n17349), .C2(n15666), .A(n15665), .B(n15664), .ZN(
        n15667) );
  AOI211_X1 U18869 ( .C1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .C2(n17176), .A(
        n15668), .B(n15667), .ZN(n15669) );
  OAI211_X1 U18870 ( .C1(n17144), .C2(n17367), .A(n15670), .B(n15669), .ZN(
        n15671) );
  INV_X1 U18871 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17661) );
  INV_X1 U18872 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U18873 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18874 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15611), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18875 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15674) );
  OAI211_X1 U18876 ( .C1(n17349), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        n15681) );
  AOI22_X1 U18877 ( .A1(n13852), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18878 ( .A1(n13870), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U18879 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15678) );
  INV_X1 U18880 ( .A(n18027), .ZN(n15683) );
  INV_X1 U18881 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18328) );
  NOR2_X1 U18882 ( .A1(n18328), .A2(n15685), .ZN(n15686) );
  INV_X1 U18883 ( .A(n15687), .ZN(n17533) );
  XOR2_X1 U18884 ( .A(n15746), .B(n17533), .Z(n15688) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18317) );
  NOR2_X1 U18886 ( .A1(n15689), .A2(n15688), .ZN(n15690) );
  INV_X1 U18887 ( .A(n15736), .ZN(n17527) );
  XNOR2_X1 U18888 ( .A(n15691), .B(n17527), .ZN(n15692) );
  XNOR2_X1 U18889 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15692), .ZN(
        n17988) );
  NOR2_X2 U18890 ( .A1(n17987), .A2(n15693), .ZN(n15696) );
  INV_X1 U18891 ( .A(n15740), .ZN(n17524) );
  XOR2_X1 U18892 ( .A(n15694), .B(n17524), .Z(n15695) );
  XNOR2_X1 U18893 ( .A(n15696), .B(n15695), .ZN(n17974) );
  INV_X1 U18894 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17973) );
  NOR2_X1 U18895 ( .A1(n15696), .A2(n15695), .ZN(n15697) );
  XNOR2_X1 U18896 ( .A(n15699), .B(n18285), .ZN(n17964) );
  OAI21_X1 U18897 ( .B1(n16538), .B2(n15738), .A(n17811), .ZN(n15700) );
  XNOR2_X1 U18898 ( .A(n17812), .B(n15700), .ZN(n17944) );
  NOR2_X1 U18899 ( .A1(n17945), .A2(n17944), .ZN(n17943) );
  NOR2_X1 U18900 ( .A1(n17812), .A2(n15700), .ZN(n15701) );
  NOR2_X1 U18901 ( .A1(n17943), .A2(n15701), .ZN(n15702) );
  NAND2_X1 U18902 ( .A1(n15702), .A2(n17930), .ZN(n17826) );
  NOR2_X1 U18903 ( .A1(n18248), .A2(n18237), .ZN(n18230) );
  NAND2_X1 U18904 ( .A1(n18230), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18207) );
  NAND2_X1 U18905 ( .A1(n18183), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18189) );
  NOR2_X1 U18906 ( .A1(n18198), .A2(n18189), .ZN(n17830) );
  NAND2_X1 U18907 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17830), .ZN(
        n16534) );
  INV_X1 U18908 ( .A(n17826), .ZN(n15704) );
  NOR2_X1 U18909 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17904) );
  NOR4_X1 U18910 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15703) );
  NAND4_X1 U18911 ( .A1(n15704), .A2(n17904), .A3(n15703), .A4(n18173), .ZN(
        n15705) );
  NAND2_X1 U18912 ( .A1(n17811), .A2(n15705), .ZN(n15706) );
  INV_X1 U18913 ( .A(n15706), .ZN(n15708) );
  INV_X1 U18914 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18152) );
  NOR2_X1 U18915 ( .A1(n18164), .A2(n18152), .ZN(n18142) );
  INV_X1 U18916 ( .A(n18142), .ZN(n18140) );
  INV_X1 U18917 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17795) );
  INV_X1 U18918 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17783) );
  INV_X1 U18919 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17771) );
  NOR2_X1 U18920 ( .A1(n17783), .A2(n17771), .ZN(n18115) );
  AND2_X1 U18921 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18115), .ZN(
        n18101) );
  NAND2_X1 U18922 ( .A1(n18101), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18080) );
  INV_X1 U18923 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18079) );
  NAND2_X1 U18924 ( .A1(n18142), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18082) );
  INV_X1 U18925 ( .A(n18082), .ZN(n18113) );
  NAND2_X1 U18926 ( .A1(n18113), .A2(n18101), .ZN(n18095) );
  NAND2_X1 U18927 ( .A1(n18100), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18088) );
  NOR2_X1 U18928 ( .A1(n18079), .A2(n18088), .ZN(n17713) );
  INV_X1 U18929 ( .A(n17713), .ZN(n17722) );
  NAND2_X1 U18930 ( .A1(n17811), .A2(n17795), .ZN(n17794) );
  NOR2_X1 U18931 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17794), .ZN(
        n15709) );
  NAND2_X1 U18932 ( .A1(n15709), .A2(n17771), .ZN(n17758) );
  INV_X1 U18933 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18096) );
  NAND3_X1 U18934 ( .A1(n17740), .A2(n18079), .A3(n18096), .ZN(n15710) );
  INV_X1 U18935 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U18936 ( .A1(n17721), .A2(n17725), .ZN(n17720) );
  NAND2_X1 U18937 ( .A1(n15716), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15715) );
  INV_X1 U18938 ( .A(n17720), .ZN(n17708) );
  NAND2_X1 U18939 ( .A1(n17720), .A2(n17811), .ZN(n15714) );
  INV_X1 U18940 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18058) );
  AND3_X2 U18941 ( .A1(n15715), .A2(n15714), .A3(n15713), .ZN(n17695) );
  INV_X1 U18942 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18048) );
  NAND2_X1 U18943 ( .A1(n17933), .A2(n15716), .ZN(n17707) );
  NOR2_X1 U18944 ( .A1(n18058), .A2(n18048), .ZN(n15762) );
  NAND2_X2 U18945 ( .A1(n17694), .A2(n15717), .ZN(n16546) );
  NOR2_X4 U18946 ( .A1(n17686), .A2(n16546), .ZN(n17675) );
  NAND2_X1 U18947 ( .A1(n15841), .A2(n15840), .ZN(n15718) );
  XNOR2_X1 U18948 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15718), .ZN(
        n16520) );
  NAND2_X1 U18949 ( .A1(n15727), .A2(n10113), .ZN(n15726) );
  NOR2_X1 U18950 ( .A1(n15719), .A2(n15726), .ZN(n15733) );
  AOI21_X1 U18951 ( .B1(n15723), .B2(n15722), .A(n15721), .ZN(n16474) );
  INV_X1 U18952 ( .A(n16474), .ZN(n18798) );
  AOI21_X1 U18953 ( .B1(n15725), .B2(n15724), .A(n18803), .ZN(n15732) );
  OAI21_X1 U18954 ( .B1(n15727), .B2(n10113), .A(n15726), .ZN(n15728) );
  OAI21_X1 U18955 ( .B1(n15729), .B2(n15728), .A(n19013), .ZN(n16646) );
  NOR3_X1 U18956 ( .A1(n15730), .A2(n16648), .A3(n16646), .ZN(n15731) );
  AOI211_X1 U18957 ( .C1(n15733), .C2(n18798), .A(n15732), .B(n15731), .ZN(
        n15734) );
  INV_X1 U18958 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17866) );
  NAND2_X1 U18959 ( .A1(n18172), .A2(n17713), .ZN(n18076) );
  INV_X1 U18960 ( .A(n18041), .ZN(n17660) );
  NOR2_X1 U18961 ( .A1(n15738), .A2(n18797), .ZN(n18201) );
  NAND2_X1 U18962 ( .A1(n18334), .A2(n18201), .ZN(n18272) );
  INV_X1 U18963 ( .A(n18272), .ZN(n15770) );
  INV_X1 U18964 ( .A(n15858), .ZN(n15747) );
  NOR2_X1 U18965 ( .A1(n17550), .A2(n15747), .ZN(n15748) );
  NOR2_X1 U18966 ( .A1(n15736), .A2(n15742), .ZN(n15739) );
  NAND2_X1 U18967 ( .A1(n15739), .A2(n15740), .ZN(n17956) );
  INV_X1 U18968 ( .A(n17956), .ZN(n17958) );
  NAND2_X1 U18969 ( .A1(n17954), .A2(n17958), .ZN(n15737) );
  NOR2_X1 U18970 ( .A1(n15737), .A2(n17518), .ZN(n15760) );
  INV_X1 U18971 ( .A(n15760), .ZN(n15756) );
  XOR2_X1 U18972 ( .A(n15738), .B(n15737), .Z(n17947) );
  XNOR2_X1 U18973 ( .A(n17954), .B(n17956), .ZN(n15755) );
  XOR2_X1 U18974 ( .A(n15740), .B(n15739), .Z(n15741) );
  NAND2_X1 U18975 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15741), .ZN(
        n15754) );
  XNOR2_X1 U18976 ( .A(n17973), .B(n15741), .ZN(n17971) );
  XNOR2_X1 U18977 ( .A(n17527), .B(n15742), .ZN(n15743) );
  NAND2_X1 U18978 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15743), .ZN(
        n15753) );
  INV_X1 U18979 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18305) );
  XNOR2_X1 U18980 ( .A(n18305), .B(n15743), .ZN(n17984) );
  XOR2_X1 U18981 ( .A(n15745), .B(n17533), .Z(n15744) );
  NAND2_X1 U18982 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15744), .ZN(
        n15752) );
  XNOR2_X1 U18983 ( .A(n18317), .B(n15744), .ZN(n18313) );
  AOI21_X1 U18984 ( .B1(n15858), .B2(n15746), .A(n15745), .ZN(n15750) );
  OR2_X1 U18985 ( .A1(n18328), .A2(n15750), .ZN(n15751) );
  AND2_X1 U18986 ( .A1(n15673), .A2(n17550), .ZN(n15749) );
  INV_X1 U18987 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18985) );
  NAND2_X1 U18988 ( .A1(n15747), .A2(n18985), .ZN(n18026) );
  NOR2_X1 U18989 ( .A1(n18019), .A2(n18026), .ZN(n18018) );
  NOR3_X1 U18990 ( .A1(n15749), .A2(n15748), .A3(n18018), .ZN(n18011) );
  XNOR2_X1 U18991 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15750), .ZN(
        n18010) );
  NAND2_X1 U18992 ( .A1(n18011), .A2(n18010), .ZN(n18009) );
  NAND2_X1 U18993 ( .A1(n15751), .A2(n18009), .ZN(n18312) );
  NAND2_X1 U18994 ( .A1(n18313), .A2(n18312), .ZN(n18311) );
  NAND2_X1 U18995 ( .A1(n15752), .A2(n18311), .ZN(n17983) );
  NAND2_X1 U18996 ( .A1(n17984), .A2(n17983), .ZN(n17982) );
  NAND2_X1 U18997 ( .A1(n15753), .A2(n17982), .ZN(n17970) );
  NAND2_X1 U18998 ( .A1(n17971), .A2(n17970), .ZN(n17969) );
  NAND2_X1 U18999 ( .A1(n15754), .A2(n17969), .ZN(n17957) );
  AOI222_X1 U19000 ( .A1(n15755), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n15755), .B2(n17957), .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(
        n17957), .ZN(n17948) );
  NAND2_X1 U19001 ( .A1(n17947), .A2(n17948), .ZN(n17946) );
  NAND2_X1 U19002 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17946), .ZN(
        n15759) );
  NOR2_X1 U19003 ( .A1(n15756), .A2(n15759), .ZN(n15761) );
  NOR2_X1 U19004 ( .A1(n17947), .A2(n17948), .ZN(n15758) );
  NOR2_X1 U19005 ( .A1(n15760), .A2(n15759), .ZN(n15757) );
  AOI211_X1 U19006 ( .C1(n15760), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        n17931) );
  NOR2_X1 U19007 ( .A1(n17931), .A2(n17930), .ZN(n17929) );
  INV_X1 U19008 ( .A(n15762), .ZN(n18036) );
  INV_X1 U19009 ( .A(n18088), .ZN(n17726) );
  NAND3_X1 U19010 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17726), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18059) );
  NOR2_X1 U19011 ( .A1(n18036), .A2(n18059), .ZN(n16537) );
  NAND2_X1 U19012 ( .A1(n18169), .A2(n16537), .ZN(n17659) );
  AND2_X1 U19013 ( .A1(n15765), .A2(n16665), .ZN(n15767) );
  AOI21_X1 U19014 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18327) );
  NAND3_X1 U19015 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18135) );
  NOR2_X1 U19016 ( .A1(n18327), .A2(n18135), .ZN(n18259) );
  NOR3_X1 U19017 ( .A1(n17930), .A2(n18285), .A3(n17945), .ZN(n18136) );
  NAND2_X1 U19018 ( .A1(n18259), .A2(n18136), .ZN(n18184) );
  NOR2_X1 U19019 ( .A1(n16534), .A2(n18184), .ZN(n18081) );
  NAND2_X1 U19020 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18134) );
  NOR2_X1 U19021 ( .A1(n18135), .A2(n18134), .ZN(n18258) );
  NAND2_X1 U19022 ( .A1(n18136), .A2(n18258), .ZN(n18160) );
  NOR2_X1 U19023 ( .A1(n16534), .A2(n18160), .ZN(n18138) );
  OAI21_X1 U19024 ( .B1(n18985), .B2(n18818), .A(n18353), .ZN(n18329) );
  AOI22_X1 U19025 ( .A1(n18804), .A2(n18081), .B1(n18138), .B2(n18329), .ZN(
        n18060) );
  INV_X1 U19026 ( .A(n18060), .ZN(n16535) );
  NAND2_X1 U19027 ( .A1(n16537), .A2(n16535), .ZN(n16522) );
  OAI21_X1 U19028 ( .B1(n17659), .B2(n18332), .A(n16522), .ZN(n15769) );
  AOI22_X1 U19029 ( .A1(n17660), .A2(n15770), .B1(n18334), .B2(n15769), .ZN(
        n15848) );
  NAND2_X1 U19030 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16507) );
  INV_X1 U19031 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15839) );
  NOR2_X1 U19032 ( .A1(n16507), .A2(n15839), .ZN(n15838) );
  INV_X1 U19033 ( .A(n15838), .ZN(n16524) );
  OAI22_X1 U19034 ( .A1(n16508), .A2(n18349), .B1(n16506), .B2(n18272), .ZN(
        n15844) );
  NAND3_X2 U19035 ( .A1(n18984), .A2(n18957), .A3(n18856), .ZN(n18339) );
  INV_X2 U19036 ( .A(n18339), .ZN(n18357) );
  OR2_X1 U19037 ( .A1(n18985), .A2(n18160), .ZN(n18246) );
  NOR2_X1 U19038 ( .A1(n16534), .A2(n18246), .ZN(n18159) );
  NAND3_X1 U19039 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16537), .A3(
        n18159), .ZN(n15771) );
  AOI21_X1 U19040 ( .B1(n16537), .B2(n18081), .A(n18833), .ZN(n18035) );
  NOR2_X2 U19041 ( .A1(n18357), .A2(n18334), .ZN(n18346) );
  AOI211_X1 U19042 ( .C1(n18813), .C2(n15771), .A(n18035), .B(n18346), .ZN(
        n15772) );
  OAI221_X1 U19043 ( .B1(n18353), .B2(n16537), .C1(n18353), .C2(n18138), .A(
        n15772), .ZN(n15843) );
  AOI21_X1 U19044 ( .B1(n18204), .B2(n17686), .A(n15843), .ZN(n16542) );
  INV_X1 U19045 ( .A(n18261), .ZN(n18085) );
  NAND2_X1 U19046 ( .A1(n18334), .A2(n18085), .ZN(n18340) );
  OAI22_X1 U19047 ( .A1(n18357), .A2(n16542), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18340), .ZN(n15773) );
  NOR2_X1 U19048 ( .A1(n15844), .A2(n15773), .ZN(n15774) );
  MUX2_X1 U19049 ( .A(n10503), .B(n15774), .S(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n15775) );
  NAND2_X1 U19050 ( .A1(n18357), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16516) );
  OAI211_X1 U19051 ( .C1(n16520), .C2(n18270), .A(n15775), .B(n16516), .ZN(
        P3_U2833) );
  INV_X1 U19052 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21222) );
  NOR3_X1 U19053 ( .A1(n21010), .A2(n15776), .A3(n21005), .ZN(n15777) );
  OR3_X1 U19054 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n20106) );
  AOI21_X1 U19055 ( .B1(n21213), .B2(n21222), .A(n20106), .ZN(n15816) );
  INV_X1 U19056 ( .A(n15780), .ZN(n15781) );
  OR2_X1 U19057 ( .A1(n15782), .A2(n15781), .ZN(n15784) );
  OAI21_X1 U19058 ( .B1(n15784), .B2(n10153), .A(n15783), .ZN(n15792) );
  INV_X1 U19059 ( .A(n15785), .ZN(n15787) );
  NAND2_X1 U19060 ( .A1(n15787), .A2(n15786), .ZN(n15791) );
  NAND2_X1 U19061 ( .A1(n15789), .A2(n15788), .ZN(n15790) );
  AND3_X1 U19062 ( .A1(n15792), .A2(n15791), .A3(n15790), .ZN(n21003) );
  INV_X1 U19063 ( .A(n21003), .ZN(n15815) );
  INV_X1 U19064 ( .A(n15793), .ZN(n15794) );
  AND2_X1 U19065 ( .A1(n15795), .A2(n15794), .ZN(n15810) );
  AND2_X1 U19066 ( .A1(n15796), .A2(n15795), .ZN(n15806) );
  OAI22_X1 U19067 ( .A1(n15799), .A2(n15798), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15797), .ZN(n20986) );
  NAND2_X1 U19068 ( .A1(n15800), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n20994) );
  INV_X1 U19069 ( .A(n20994), .ZN(n15801) );
  NOR2_X1 U19070 ( .A1(n20986), .A2(n15801), .ZN(n15803) );
  NAND2_X1 U19071 ( .A1(n20723), .A2(n15806), .ZN(n15802) );
  NAND3_X1 U19072 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15803), .A3(
        n15802), .ZN(n15805) );
  NAND2_X1 U19073 ( .A1(n15808), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15804) );
  OAI211_X1 U19074 ( .C1(n15806), .C2(n20723), .A(n15805), .B(n15804), .ZN(
        n15807) );
  OAI21_X1 U19075 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15808), .A(
        n15807), .ZN(n15809) );
  AOI222_X1 U19076 ( .A1(n20653), .A2(n15810), .B1(n20653), .B2(n15809), .C1(
        n15810), .C2(n15809), .ZN(n15813) );
  OAI211_X1 U19077 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15813), .A(
        n15812), .B(n15811), .ZN(n15814) );
  NOR4_X1 U19078 ( .A1(n15817), .A2(n15816), .A3(n15815), .A4(n15814), .ZN(
        n15830) );
  INV_X1 U19079 ( .A(n15830), .ZN(n15822) );
  NAND4_X1 U19080 ( .A1(n11580), .A2(n20355), .A3(n15849), .A4(n15818), .ZN(
        n15821) );
  OAI21_X1 U19081 ( .B1(n15819), .B2(n16097), .A(n20917), .ZN(n15820) );
  NAND2_X1 U19082 ( .A1(n15821), .A2(n15820), .ZN(n16099) );
  AOI221_X1 U19083 ( .B1(n21012), .B2(n16101), .C1(n15822), .C2(n16101), .A(
        n16099), .ZN(n15824) );
  NOR2_X1 U19084 ( .A1(n15824), .A2(n21012), .ZN(n20918) );
  OAI211_X1 U19085 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n16097), .A(n20918), 
        .B(n15823), .ZN(n16100) );
  AOI21_X1 U19086 ( .B1(n21018), .B2(n15825), .A(n15824), .ZN(n15826) );
  OAI22_X1 U19087 ( .A1(n15827), .A2(n16100), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15826), .ZN(n15828) );
  OAI21_X1 U19088 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(P1_U3161) );
  NOR2_X1 U19089 ( .A1(n15831), .A2(n16000), .ZN(n15984) );
  AOI22_X1 U19090 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20317), .B1(n15984), 
        .B2(n11545), .ZN(n15836) );
  INV_X1 U19091 ( .A(n15832), .ZN(n15834) );
  AOI22_X1 U19092 ( .A1(n15834), .A2(n20332), .B1(n20316), .B2(n15833), .ZN(
        n15835) );
  OAI211_X1 U19093 ( .C1(n11545), .C2(n15985), .A(n15836), .B(n15835), .ZN(
        P1_U3010) );
  INV_X1 U19094 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15837) );
  NAND2_X1 U19095 ( .A1(n15838), .A2(n15837), .ZN(n16505) );
  NOR2_X1 U19096 ( .A1(n16486), .A2(n9914), .ZN(n15842) );
  XNOR2_X1 U19097 ( .A(n15842), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16501) );
  AOI22_X1 U19098 ( .A1(n18357), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n18253), 
        .B2(n16501), .ZN(n15847) );
  INV_X1 U19099 ( .A(n18340), .ZN(n18262) );
  AOI22_X1 U19100 ( .A1(n18262), .A2(n16524), .B1(n18339), .B2(n15843), .ZN(
        n16521) );
  INV_X1 U19101 ( .A(n16521), .ZN(n15845) );
  OAI21_X1 U19102 ( .B1(n15845), .B2(n15844), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15846) );
  OAI211_X1 U19103 ( .C1(n15848), .C2(n16505), .A(n15847), .B(n15846), .ZN(
        P3_U2832) );
  INV_X1 U19104 ( .A(HOLD), .ZN(n21254) );
  INV_X1 U19105 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20932) );
  NAND2_X1 U19106 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20932), .ZN(n20924) );
  INV_X1 U19107 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20920) );
  INV_X1 U19108 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21022) );
  NOR2_X1 U19109 ( .A1(n20920), .A2(n21022), .ZN(n20927) );
  AOI221_X1 U19110 ( .B1(n20932), .B2(n20927), .C1(n21254), .C2(n20927), .A(
        n15849), .ZN(n15851) );
  NAND2_X1 U19111 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21005), .ZN(n15850) );
  OAI211_X1 U19112 ( .C1(n21254), .C2(n20924), .A(n15851), .B(n15850), .ZN(
        P1_U3195) );
  AND2_X1 U19113 ( .A1(n20224), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19114 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15852) );
  NOR3_X1 U19115 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19034), .A3(n19950), 
        .ZN(n19951) );
  NOR4_X1 U19116 ( .A1(n15853), .A2(n15852), .A3(n19951), .A4(n16457), .ZN(
        P2_U3178) );
  AOI221_X1 U19117 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16457), .C1(n20092), .C2(
        n16457), .A(n19863), .ZN(n20087) );
  INV_X1 U19118 ( .A(n20087), .ZN(n20084) );
  NOR2_X1 U19119 ( .A1(n16427), .A2(n20084), .ZN(P2_U3047) );
  NAND2_X1 U19120 ( .A1(n17445), .A2(n17401), .ZN(n17544) );
  INV_X1 U19121 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17621) );
  NAND2_X1 U19122 ( .A1(n15857), .A2(n17401), .ZN(n17541) );
  AOI22_X1 U19123 ( .A1(n17543), .A2(BUF2_REG_0__SCAN_IN), .B1(n17528), .B2(
        n15858), .ZN(n15859) );
  OAI221_X1 U19124 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17544), .C1(n17621), 
        .C2(n17401), .A(n15859), .ZN(P3_U2735) );
  AOI22_X1 U19125 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20190), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n20177), .ZN(n15867) );
  INV_X1 U19126 ( .A(n15860), .ZN(n15929) );
  AOI21_X1 U19127 ( .B1(n15861), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15863) );
  OAI22_X1 U19128 ( .A1(n15864), .A2(n15863), .B1(n20174), .B2(n15862), .ZN(
        n15865) );
  AOI21_X1 U19129 ( .B1(n15929), .B2(n20155), .A(n15865), .ZN(n15866) );
  OAI211_X1 U19130 ( .C1(n15932), .C2(n20184), .A(n15867), .B(n15866), .ZN(
        P1_U2820) );
  AOI22_X1 U19131 ( .A1(n15868), .A2(n20191), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15881), .ZN(n15871) );
  AOI21_X1 U19132 ( .B1(n20190), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20153), .ZN(n15870) );
  NAND2_X1 U19133 ( .A1(n20177), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n15869) );
  NAND3_X1 U19134 ( .A1(n15871), .A2(n15870), .A3(n15869), .ZN(n15872) );
  OR2_X1 U19135 ( .A1(n15873), .A2(n15872), .ZN(n15874) );
  AOI21_X1 U19136 ( .B1(n15875), .B2(n20155), .A(n15874), .ZN(n15876) );
  OAI21_X1 U19137 ( .B1(n20174), .B2(n16003), .A(n15876), .ZN(P1_U2822) );
  AOI22_X1 U19138 ( .A1(n15877), .A2(n20191), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n20177), .ZN(n15878) );
  OAI211_X1 U19139 ( .C1(n20172), .C2(n11156), .A(n20170), .B(n15878), .ZN(
        n15879) );
  AOI21_X1 U19140 ( .B1(n15880), .B2(n20155), .A(n15879), .ZN(n15884) );
  OAI21_X1 U19141 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15882), .A(n15881), 
        .ZN(n15883) );
  OAI211_X1 U19142 ( .C1(n15885), .C2(n20174), .A(n15884), .B(n15883), .ZN(
        P1_U2823) );
  OAI21_X1 U19143 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), 
        .A(n15886), .ZN(n15896) );
  NOR2_X1 U19144 ( .A1(n20160), .A2(n15887), .ZN(n15907) );
  AOI22_X1 U19145 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20177), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n15907), .ZN(n15892) );
  INV_X1 U19146 ( .A(n15937), .ZN(n15890) );
  INV_X1 U19147 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15888) );
  NOR2_X1 U19148 ( .A1(n20172), .A2(n15888), .ZN(n15889) );
  AOI211_X1 U19149 ( .C1(n20191), .C2(n15890), .A(n20153), .B(n15889), .ZN(
        n15891) );
  OAI211_X1 U19150 ( .C1(n20174), .C2(n15893), .A(n15892), .B(n15891), .ZN(
        n15894) );
  AOI21_X1 U19151 ( .B1(n15934), .B2(n20155), .A(n15894), .ZN(n15895) );
  OAI21_X1 U19152 ( .B1(n15905), .B2(n15896), .A(n15895), .ZN(P1_U2824) );
  AOI22_X1 U19153 ( .A1(n15897), .A2(n20191), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15907), .ZN(n15904) );
  INV_X1 U19154 ( .A(n15898), .ZN(n16013) );
  AOI22_X1 U19155 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n20177), .B1(n20186), 
        .B2(n16013), .ZN(n15899) );
  OAI211_X1 U19156 ( .C1(n20172), .C2(n15900), .A(n20170), .B(n15899), .ZN(
        n15901) );
  AOI21_X1 U19157 ( .B1(n15902), .B2(n20155), .A(n15901), .ZN(n15903) );
  OAI211_X1 U19158 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15905), .A(n15904), 
        .B(n15903), .ZN(P1_U2825) );
  AOI21_X1 U19159 ( .B1(n15906), .B2(P1_REIP_REG_13__SCAN_IN), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15914) );
  INV_X1 U19160 ( .A(n15907), .ZN(n15913) );
  OAI22_X1 U19161 ( .A1(n15908), .A2(n20201), .B1(n20174), .B2(n16018), .ZN(
        n15909) );
  AOI211_X1 U19162 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20153), .B(n15909), .ZN(n15912) );
  INV_X1 U19163 ( .A(n15910), .ZN(n15944) );
  AOI22_X1 U19164 ( .A1(n15944), .A2(n20155), .B1(n20191), .B2(n15943), .ZN(
        n15911) );
  OAI211_X1 U19165 ( .C1(n15914), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        P1_U2826) );
  INV_X1 U19166 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20946) );
  OR2_X1 U19167 ( .A1(n15916), .A2(n15915), .ZN(n15917) );
  AND2_X1 U19168 ( .A1(n15918), .A2(n15917), .ZN(n16045) );
  AOI22_X1 U19169 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20177), .B1(n20186), 
        .B2(n16045), .ZN(n15919) );
  OAI211_X1 U19170 ( .C1(n20172), .C2(n11047), .A(n15919), .B(n20170), .ZN(
        n15920) );
  AOI221_X1 U19171 ( .B1(n15922), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15921), 
        .C2(n20946), .A(n15920), .ZN(n15924) );
  NAND2_X1 U19172 ( .A1(n15964), .A2(n20155), .ZN(n15923) );
  OAI211_X1 U19173 ( .C1(n20184), .C2(n15967), .A(n15924), .B(n15923), .ZN(
        P1_U2829) );
  INV_X1 U19174 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15926) );
  AOI22_X1 U19175 ( .A1(n15964), .A2(n20207), .B1(n20206), .B2(n16045), .ZN(
        n15925) );
  OAI21_X1 U19176 ( .B1(n20211), .B2(n15926), .A(n15925), .ZN(P1_U2861) );
  AOI21_X1 U19177 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20291), .A(
        n15927), .ZN(n15931) );
  AOI22_X1 U19178 ( .A1(n15929), .A2(n15981), .B1(n20298), .B2(n15928), .ZN(
        n15930) );
  OAI211_X1 U19179 ( .C1(n20302), .C2(n15932), .A(n15931), .B(n15930), .ZN(
        P1_U2979) );
  AOI22_X1 U19180 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15936) );
  AOI22_X1 U19181 ( .A1(n15934), .A2(n15981), .B1(n20298), .B2(n15933), .ZN(
        n15935) );
  OAI211_X1 U19182 ( .C1(n20302), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        P1_U2983) );
  OAI22_X1 U19183 ( .A1(n15940), .A2(n15939), .B1(n15938), .B2(n16031), .ZN(
        n15942) );
  XNOR2_X1 U19184 ( .A(n15938), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15941) );
  XNOR2_X1 U19185 ( .A(n15942), .B(n15941), .ZN(n16019) );
  AOI22_X1 U19186 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15946) );
  AOI22_X1 U19187 ( .A1(n15944), .A2(n15981), .B1(n15956), .B2(n15943), .ZN(
        n15945) );
  OAI211_X1 U19188 ( .C1(n16019), .C2(n20108), .A(n15946), .B(n15945), .ZN(
        P1_U2985) );
  INV_X1 U19189 ( .A(n15947), .ZN(n15948) );
  NOR2_X1 U19190 ( .A1(n15949), .A2(n15948), .ZN(n15953) );
  NAND2_X1 U19191 ( .A1(n15951), .A2(n15950), .ZN(n15952) );
  XNOR2_X1 U19192 ( .A(n15953), .B(n15952), .ZN(n16042) );
  AOI22_X1 U19193 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15959) );
  INV_X1 U19194 ( .A(n15954), .ZN(n15957) );
  AOI22_X1 U19195 ( .A1(n15957), .A2(n15981), .B1(n15956), .B2(n15955), .ZN(
        n15958) );
  OAI211_X1 U19196 ( .C1(n16042), .C2(n20108), .A(n15959), .B(n15958), .ZN(
        P1_U2987) );
  AOI22_X1 U19197 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15966) );
  NOR3_X1 U19198 ( .A1(n15960), .A2(n11531), .A3(n16064), .ZN(n15962) );
  NOR2_X1 U19199 ( .A1(n15962), .A2(n15961), .ZN(n15963) );
  XNOR2_X1 U19200 ( .A(n15963), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16046) );
  AOI22_X1 U19201 ( .A1(n16046), .A2(n20298), .B1(n20296), .B2(n15964), .ZN(
        n15965) );
  OAI211_X1 U19202 ( .C1(n20302), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        P1_U2988) );
  AOI22_X1 U19203 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15972) );
  XNOR2_X1 U19204 ( .A(n15968), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15969) );
  XNOR2_X1 U19205 ( .A(n15970), .B(n15969), .ZN(n16076) );
  AOI22_X1 U19206 ( .A1(n16076), .A2(n20298), .B1(n15981), .B2(n20148), .ZN(
        n15971) );
  OAI211_X1 U19207 ( .C1(n20302), .C2(n20150), .A(n15972), .B(n15971), .ZN(
        P1_U2992) );
  AOI22_X1 U19208 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15976) );
  INV_X1 U19209 ( .A(n15973), .ZN(n15974) );
  AOI22_X1 U19210 ( .A1(n15974), .A2(n20298), .B1(n15981), .B2(n20156), .ZN(
        n15975) );
  OAI211_X1 U19211 ( .C1(n20302), .C2(n20159), .A(n15976), .B(n15975), .ZN(
        P1_U2993) );
  AOI22_X1 U19212 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15983) );
  OAI21_X1 U19213 ( .B1(n15979), .B2(n15978), .A(n15977), .ZN(n15980) );
  INV_X1 U19214 ( .A(n15980), .ZN(n16088) );
  AOI22_X1 U19215 ( .A1(n16088), .A2(n20298), .B1(n15981), .B2(n20208), .ZN(
        n15982) );
  OAI211_X1 U19216 ( .C1(n20302), .C2(n20169), .A(n15983), .B(n15982), .ZN(
        P1_U2994) );
  OAI21_X1 U19217 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15984), .ZN(n15992) );
  OAI22_X1 U19218 ( .A1(n15987), .A2(n20344), .B1(n15986), .B2(n15985), .ZN(
        n15988) );
  AOI21_X1 U19219 ( .B1(n20332), .B2(n15989), .A(n15988), .ZN(n15991) );
  NAND2_X1 U19220 ( .A1(n20317), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15990) );
  OAI211_X1 U19221 ( .C1(n15993), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        P1_U3009) );
  AOI22_X1 U19222 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15994), .B1(
        n20317), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15999) );
  INV_X1 U19223 ( .A(n15995), .ZN(n15997) );
  AOI22_X1 U19224 ( .A1(n15997), .A2(n20332), .B1(n20316), .B2(n15996), .ZN(
        n15998) );
  OAI211_X1 U19225 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16000), .A(
        n15999), .B(n15998), .ZN(P1_U3012) );
  NAND2_X1 U19226 ( .A1(n16002), .A2(n16001), .ZN(n16009) );
  OAI22_X1 U19227 ( .A1(n16004), .A2(n20340), .B1(n20344), .B2(n16003), .ZN(
        n16005) );
  AOI21_X1 U19228 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16006), .A(
        n16005), .ZN(n16008) );
  NAND2_X1 U19229 ( .A1(n20317), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16007) );
  OAI211_X1 U19230 ( .C1(n16010), .C2(n16009), .A(n16008), .B(n16007), .ZN(
        P1_U3013) );
  AOI22_X1 U19231 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16011), .B1(
        n20317), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16016) );
  INV_X1 U19232 ( .A(n16012), .ZN(n16014) );
  AOI22_X1 U19233 ( .A1(n16014), .A2(n20332), .B1(n20316), .B2(n16013), .ZN(
        n16015) );
  OAI211_X1 U19234 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16017), .A(
        n16016), .B(n16015), .ZN(P1_U3016) );
  NOR2_X1 U19235 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16081), .ZN(
        n16022) );
  OAI22_X1 U19236 ( .A1(n16019), .A2(n20340), .B1(n20344), .B2(n16018), .ZN(
        n16020) );
  AOI21_X1 U19237 ( .B1(n16022), .B2(n16021), .A(n16020), .ZN(n16024) );
  NAND2_X1 U19238 ( .A1(n20317), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16023) );
  OAI211_X1 U19239 ( .C1(n16032), .C2(n16025), .A(n16024), .B(n16023), .ZN(
        P1_U3017) );
  INV_X1 U19240 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U19241 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n20317), .B1(n16031), 
        .B2(n16026), .ZN(n16030) );
  AOI22_X1 U19242 ( .A1(n16028), .A2(n20332), .B1(n20316), .B2(n16027), .ZN(
        n16029) );
  OAI211_X1 U19243 ( .C1(n16032), .C2(n16031), .A(n16030), .B(n16029), .ZN(
        P1_U3018) );
  NOR2_X1 U19244 ( .A1(n20342), .A2(n21376), .ZN(n16035) );
  AND3_X1 U19245 ( .A1(n16033), .A2(n16039), .A3(n16044), .ZN(n16034) );
  AOI211_X1 U19246 ( .C1(n20316), .C2(n16036), .A(n16035), .B(n16034), .ZN(
        n16041) );
  OAI21_X1 U19247 ( .B1(n16037), .B2(n16051), .A(n20327), .ZN(n16038) );
  OAI211_X1 U19248 ( .C1(n16039), .C2(n20323), .A(n16052), .B(n16038), .ZN(
        n16047) );
  OAI221_X1 U19249 ( .B1(n16047), .B2(n20322), .C1(n16047), .C2(n16043), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16040) );
  OAI211_X1 U19250 ( .C1(n16042), .C2(n20340), .A(n16041), .B(n16040), .ZN(
        P1_U3019) );
  NAND2_X1 U19251 ( .A1(n16044), .A2(n16043), .ZN(n16050) );
  AOI22_X1 U19252 ( .A1(n16045), .A2(n20316), .B1(n20317), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16049) );
  AOI22_X1 U19253 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16047), .B1(
        n20332), .B2(n16046), .ZN(n16048) );
  OAI211_X1 U19254 ( .C1(n16051), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        P1_U3020) );
  OAI211_X1 U19255 ( .C1(n16055), .C2(n16054), .A(n16053), .B(n16052), .ZN(
        n16056) );
  NAND2_X1 U19256 ( .A1(n16057), .A2(n16056), .ZN(n16074) );
  OAI22_X1 U19257 ( .A1(n16058), .A2(n20344), .B1(n21364), .B2(n20342), .ZN(
        n16059) );
  AOI21_X1 U19258 ( .B1(n20332), .B2(n16060), .A(n16059), .ZN(n16063) );
  NOR2_X1 U19259 ( .A1(n16061), .A2(n16080), .ZN(n16070) );
  OAI221_X1 U19260 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16064), .C2(n16075), .A(
        n16070), .ZN(n16062) );
  OAI211_X1 U19261 ( .C1(n16064), .C2(n16074), .A(n16063), .B(n16062), .ZN(
        P1_U3021) );
  AOI21_X1 U19262 ( .B1(n16067), .B2(n16066), .A(n16065), .ZN(n20203) );
  INV_X1 U19263 ( .A(n16068), .ZN(n16069) );
  AOI21_X1 U19264 ( .B1(n20203), .B2(n20316), .A(n16069), .ZN(n16073) );
  AOI22_X1 U19265 ( .A1(n16071), .A2(n20332), .B1(n16070), .B2(n16075), .ZN(
        n16072) );
  OAI211_X1 U19266 ( .C1(n16075), .C2(n16074), .A(n16073), .B(n16072), .ZN(
        P1_U3022) );
  INV_X1 U19267 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16079) );
  AOI222_X1 U19268 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20317), .B1(n20316), 
        .B2(n20144), .C1(n20332), .C2(n16076), .ZN(n16077) );
  OAI221_X1 U19269 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16080), .C1(
        n16079), .C2(n16078), .A(n16077), .ZN(P1_U3024) );
  INV_X1 U19270 ( .A(n16081), .ZN(n16082) );
  NAND2_X1 U19271 ( .A1(n20304), .A2(n16082), .ZN(n20321) );
  AND2_X1 U19272 ( .A1(n16084), .A2(n16083), .ZN(n16085) );
  AOI22_X1 U19273 ( .A1(n9951), .A2(n20316), .B1(n20317), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19274 ( .A1(n16088), .A2(n20332), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16087), .ZN(n16089) );
  OAI211_X1 U19275 ( .C1(n16091), .C2(n20321), .A(n16090), .B(n16089), .ZN(
        P1_U3026) );
  INV_X1 U19276 ( .A(n20992), .ZN(n20990) );
  NAND3_X1 U19277 ( .A1(n16094), .A2(n16093), .A3(n16092), .ZN(n16095) );
  OAI21_X1 U19278 ( .B1(n20990), .B2(n16096), .A(n16095), .ZN(P1_U3468) );
  OAI221_X1 U19279 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21012), .C2(n16097), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20919) );
  NAND2_X1 U19280 ( .A1(n16102), .A2(n20919), .ZN(n16098) );
  AOI22_X1 U19281 ( .A1(n16101), .A2(n16100), .B1(n16099), .B2(n16098), .ZN(
        P1_U3162) );
  OAI22_X1 U19282 ( .A1(n20918), .A2(n20985), .B1(n21012), .B2(n16102), .ZN(
        P1_U3466) );
  INV_X1 U19283 ( .A(n16103), .ZN(n16105) );
  OAI22_X1 U19284 ( .A1(n16105), .A2(n19233), .B1(n14683), .B2(n16104), .ZN(
        n16108) );
  AOI22_X1 U19285 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19217), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19248), .ZN(n16106) );
  INV_X1 U19286 ( .A(n16106), .ZN(n16107) );
  AOI211_X1 U19287 ( .C1(n19251), .C2(n19263), .A(n16108), .B(n16107), .ZN(
        n16114) );
  INV_X1 U19288 ( .A(n16109), .ZN(n16145) );
  INV_X1 U19289 ( .A(n16110), .ZN(n16165) );
  INV_X1 U19290 ( .A(n16111), .ZN(n16190) );
  NOR2_X1 U19291 ( .A1(n9835), .A2(n16112), .ZN(n16198) );
  NOR2_X1 U19292 ( .A1(n9835), .A2(n16188), .ZN(n16179) );
  NOR2_X1 U19293 ( .A1(n16180), .A2(n16179), .ZN(n16178) );
  NOR2_X1 U19294 ( .A1(n9835), .A2(n16178), .ZN(n16164) );
  NOR2_X1 U19295 ( .A1(n9835), .A2(n16163), .ZN(n16153) );
  NOR2_X1 U19296 ( .A1(n9835), .A2(n16152), .ZN(n16144) );
  NOR2_X1 U19297 ( .A1(n16145), .A2(n16144), .ZN(n16143) );
  NAND4_X1 U19298 ( .A1(n19226), .A2(n16127), .A3(n16116), .A4(n9831), .ZN(
        n16113) );
  OAI211_X1 U19299 ( .C1(n16115), .C2(n19230), .A(n16114), .B(n16113), .ZN(
        P2_U2824) );
  AOI22_X1 U19300 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19248), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19245), .ZN(n16117) );
  OAI21_X1 U19301 ( .B1(n16118), .B2(n19233), .A(n16117), .ZN(n16122) );
  OAI22_X1 U19302 ( .A1(n16120), .A2(n19230), .B1(n16119), .B2(n19232), .ZN(
        n16121) );
  OAI21_X1 U19303 ( .B1(n19953), .B2(n16124), .A(n16123), .ZN(P2_U2825) );
  AOI21_X1 U19304 ( .B1(n16126), .B2(n16125), .A(n19953), .ZN(n16138) );
  INV_X1 U19305 ( .A(n16127), .ZN(n16137) );
  AOI22_X1 U19306 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19244), .B1(n16128), 
        .B2(n19247), .ZN(n16130) );
  AOI22_X1 U19307 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19248), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19217), .ZN(n16129) );
  OAI211_X1 U19308 ( .C1(n16131), .C2(n19230), .A(n16130), .B(n16129), .ZN(
        n16132) );
  AOI21_X1 U19309 ( .B1(n16138), .B2(n16137), .A(n16136), .ZN(n16139) );
  INV_X1 U19310 ( .A(n16139), .ZN(P2_U2826) );
  INV_X1 U19311 ( .A(n16140), .ZN(n16142) );
  AOI22_X1 U19312 ( .A1(n16142), .A2(n19249), .B1(n16141), .B2(n19251), .ZN(
        n16151) );
  AOI211_X1 U19313 ( .C1(n16145), .C2(n16144), .A(n16143), .B(n19953), .ZN(
        n16149) );
  AOI22_X1 U19314 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19245), .ZN(n16146) );
  OAI21_X1 U19315 ( .B1(n16147), .B2(n19233), .A(n16146), .ZN(n16148) );
  AOI211_X1 U19316 ( .C1(n19248), .C2(P2_REIP_REG_28__SCAN_IN), .A(n16149), 
        .B(n16148), .ZN(n16150) );
  NAND2_X1 U19317 ( .A1(n16151), .A2(n16150), .ZN(P2_U2827) );
  AOI211_X1 U19318 ( .C1(n16154), .C2(n16153), .A(n16152), .B(n19953), .ZN(
        n16160) );
  AOI22_X1 U19319 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19248), .B1(n16155), 
        .B2(n19247), .ZN(n16157) );
  AOI22_X1 U19320 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19245), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19189), .ZN(n16156) );
  OAI211_X1 U19321 ( .C1(n16158), .C2(n19230), .A(n16157), .B(n16156), .ZN(
        n16159) );
  AOI211_X1 U19322 ( .C1(n19251), .C2(n16161), .A(n16160), .B(n16159), .ZN(
        n16162) );
  INV_X1 U19323 ( .A(n16162), .ZN(P2_U2828) );
  AOI211_X1 U19324 ( .C1(n16165), .C2(n16164), .A(n16163), .B(n19953), .ZN(
        n16171) );
  AOI22_X1 U19325 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19248), .B1(n16166), 
        .B2(n19247), .ZN(n16168) );
  AOI22_X1 U19326 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19245), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19189), .ZN(n16167) );
  OAI211_X1 U19327 ( .C1(n16169), .C2(n19232), .A(n16168), .B(n16167), .ZN(
        n16170) );
  AOI211_X1 U19328 ( .C1(n19249), .C2(n16172), .A(n16171), .B(n16170), .ZN(
        n16173) );
  INV_X1 U19329 ( .A(n16173), .ZN(P2_U2829) );
  AOI22_X1 U19330 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19248), .B1(n16174), 
        .B2(n19247), .ZN(n16176) );
  AOI22_X1 U19331 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19245), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19244), .ZN(n16175) );
  OAI211_X1 U19332 ( .C1(n16177), .C2(n19230), .A(n16176), .B(n16175), .ZN(
        n16182) );
  AOI211_X1 U19333 ( .C1(n16180), .C2(n16179), .A(n16178), .B(n19953), .ZN(
        n16181) );
  NOR2_X1 U19334 ( .A1(n16182), .A2(n16181), .ZN(n16183) );
  OAI21_X1 U19335 ( .B1(n16184), .B2(n19232), .A(n16183), .ZN(P2_U2830) );
  AOI22_X1 U19336 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19244), .B1(n16185), 
        .B2(n19247), .ZN(n16195) );
  AOI22_X1 U19337 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19248), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19245), .ZN(n16194) );
  AOI22_X1 U19338 ( .A1(n16187), .A2(n19249), .B1(n16186), .B2(n19251), .ZN(
        n16193) );
  AOI21_X1 U19339 ( .B1(n16190), .B2(n16189), .A(n16188), .ZN(n16191) );
  NAND2_X1 U19340 ( .A1(n19226), .A2(n16191), .ZN(n16192) );
  NAND4_X1 U19341 ( .A1(n16195), .A2(n16194), .A3(n16193), .A4(n16192), .ZN(
        P2_U2831) );
  AOI22_X1 U19342 ( .A1(n16196), .A2(n19249), .B1(n16208), .B2(n19251), .ZN(
        n16205) );
  AOI211_X1 U19343 ( .C1(n16199), .C2(n16198), .A(n16197), .B(n19953), .ZN(
        n16203) );
  AOI22_X1 U19344 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19245), .ZN(n16200) );
  OAI21_X1 U19345 ( .B1(n16201), .B2(n19233), .A(n16200), .ZN(n16202) );
  AOI211_X1 U19346 ( .C1(n19248), .C2(P2_REIP_REG_23__SCAN_IN), .A(n16203), 
        .B(n16202), .ZN(n16204) );
  NAND2_X1 U19347 ( .A1(n16205), .A2(n16204), .ZN(P2_U2832) );
  OAI22_X1 U19348 ( .A1(n19267), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19268), .ZN(n19472) );
  INV_X1 U19349 ( .A(n19472), .ZN(n16206) );
  AOI22_X1 U19350 ( .A1(n16207), .A2(n16206), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19317), .ZN(n16212) );
  AOI22_X1 U19351 ( .A1(n19264), .A2(BUF2_REG_23__SCAN_IN), .B1(n19262), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16211) );
  AOI22_X1 U19352 ( .A1(n16209), .A2(n19319), .B1(n19318), .B2(n16208), .ZN(
        n16210) );
  NAND3_X1 U19353 ( .A1(n16212), .A2(n16211), .A3(n16210), .ZN(P2_U2896) );
  AOI22_X1 U19354 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19412), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16270), .ZN(n16218) );
  OAI22_X1 U19355 ( .A1(n16214), .A2(n19416), .B1(n16213), .B2(n19415), .ZN(
        n16215) );
  AOI21_X1 U19356 ( .B1(n19420), .B2(n16216), .A(n16215), .ZN(n16217) );
  OAI211_X1 U19357 ( .C1(n16277), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        P2_U2992) );
  AOI22_X1 U19358 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n19112), .ZN(n16232) );
  NAND2_X1 U19359 ( .A1(n16221), .A2(n16220), .ZN(n16226) );
  AOI21_X1 U19360 ( .B1(n16224), .B2(n16223), .A(n16222), .ZN(n16225) );
  XOR2_X1 U19361 ( .A(n16226), .B(n16225), .Z(n16324) );
  INV_X1 U19362 ( .A(n16324), .ZN(n16230) );
  AOI21_X1 U19363 ( .B1(n16318), .B2(n16228), .A(n16227), .ZN(n16321) );
  INV_X1 U19364 ( .A(n16229), .ZN(n19114) );
  AOI222_X1 U19365 ( .A1(n16230), .A2(n16293), .B1(n16294), .B2(n16321), .C1(
        n19420), .C2(n19114), .ZN(n16231) );
  OAI211_X1 U19366 ( .C1(n19109), .C2(n19423), .A(n16232), .B(n16231), .ZN(
        P2_U2999) );
  AOI22_X1 U19367 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19412), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16270), .ZN(n16237) );
  OAI22_X1 U19368 ( .A1(n16234), .A2(n19416), .B1(n16233), .B2(n19415), .ZN(
        n16235) );
  AOI21_X1 U19369 ( .B1(n19420), .B2(n19128), .A(n16235), .ZN(n16236) );
  OAI211_X1 U19370 ( .C1(n16277), .C2(n16238), .A(n16237), .B(n16236), .ZN(
        P2_U3000) );
  AOI22_X1 U19371 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n16239), .ZN(n16251) );
  AOI21_X1 U19372 ( .B1(n14988), .B2(n16241), .A(n16240), .ZN(n16337) );
  NAND2_X1 U19373 ( .A1(n16243), .A2(n16242), .ZN(n16247) );
  NAND2_X1 U19374 ( .A1(n16245), .A2(n16244), .ZN(n16246) );
  XNOR2_X1 U19375 ( .A(n16247), .B(n16246), .ZN(n16340) );
  INV_X1 U19376 ( .A(n16340), .ZN(n16249) );
  INV_X1 U19377 ( .A(n16248), .ZN(n19138) );
  AOI222_X1 U19378 ( .A1(n16337), .A2(n16294), .B1(n16293), .B2(n16249), .C1(
        n19420), .C2(n19138), .ZN(n16250) );
  OAI211_X1 U19379 ( .C1(n16252), .C2(n19423), .A(n16251), .B(n16250), .ZN(
        P2_U3001) );
  AOI22_X1 U19380 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19412), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16270), .ZN(n16255) );
  AOI22_X1 U19381 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n16257), .ZN(n16268) );
  NOR2_X1 U19382 ( .A1(n9896), .A2(n16258), .ZN(n16262) );
  NOR2_X1 U19383 ( .A1(n16260), .A2(n16259), .ZN(n16261) );
  XNOR2_X1 U19384 ( .A(n16262), .B(n16261), .ZN(n16345) );
  INV_X1 U19385 ( .A(n19162), .ZN(n16266) );
  AOI21_X1 U19386 ( .B1(n16265), .B2(n16264), .A(n16263), .ZN(n16348) );
  AOI222_X1 U19387 ( .A1(n16345), .A2(n16293), .B1(n19420), .B2(n16266), .C1(
        n16294), .C2(n16348), .ZN(n16267) );
  OAI211_X1 U19388 ( .C1(n16269), .C2(n19423), .A(n16268), .B(n16267), .ZN(
        P2_U3003) );
  AOI22_X1 U19389 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19412), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16270), .ZN(n16275) );
  OAI22_X1 U19390 ( .A1(n16272), .A2(n19416), .B1(n16271), .B2(n19415), .ZN(
        n16273) );
  AOI21_X1 U19391 ( .B1(n19420), .B2(n19170), .A(n16273), .ZN(n16274) );
  OAI211_X1 U19392 ( .C1(n16277), .C2(n16276), .A(n16275), .B(n16274), .ZN(
        P2_U3004) );
  INV_X1 U19393 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16278) );
  OAI22_X1 U19394 ( .A1(n16278), .A2(n19423), .B1(n16277), .B2(n19177), .ZN(
        n16279) );
  AOI21_X1 U19395 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n19412), .A(n16279), .ZN(
        n16283) );
  AOI22_X1 U19396 ( .A1(n16281), .A2(n16294), .B1(n16293), .B2(n16280), .ZN(
        n16282) );
  OAI211_X1 U19397 ( .C1(n16284), .C2(n19182), .A(n16283), .B(n16282), .ZN(
        P2_U3005) );
  AOI22_X1 U19398 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n19192), .ZN(n16289) );
  OAI22_X1 U19399 ( .A1(n16286), .A2(n19416), .B1(n16285), .B2(n19415), .ZN(
        n16287) );
  AOI21_X1 U19400 ( .B1(n19420), .B2(n19193), .A(n16287), .ZN(n16288) );
  OAI211_X1 U19401 ( .C1(n19186), .C2(n19423), .A(n16289), .B(n16288), .ZN(
        P2_U3006) );
  AOI22_X1 U19402 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n19212), .ZN(n16298) );
  XNOR2_X1 U19403 ( .A(n16290), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16381) );
  XOR2_X1 U19404 ( .A(n16291), .B(n16292), .Z(n16378) );
  AOI22_X1 U19405 ( .A1(n16381), .A2(n16294), .B1(n16293), .B2(n16378), .ZN(
        n16295) );
  INV_X1 U19406 ( .A(n16295), .ZN(n16296) );
  AOI21_X1 U19407 ( .B1(n19420), .B2(n16380), .A(n16296), .ZN(n16297) );
  OAI211_X1 U19408 ( .C1(n16299), .C2(n19423), .A(n16298), .B(n16297), .ZN(
        P2_U3008) );
  OAI21_X1 U19409 ( .B1(n16302), .B2(n16410), .A(n16317), .ZN(n16307) );
  NAND3_X1 U19410 ( .A1(n16302), .A2(n16301), .A3(n16300), .ZN(n16305) );
  AOI22_X1 U19411 ( .A1(n16399), .A2(n16303), .B1(P2_REIP_REG_18__SCAN_IN), 
        .B2(n19412), .ZN(n16304) );
  NAND2_X1 U19412 ( .A1(n16305), .A2(n16304), .ZN(n16306) );
  AOI21_X1 U19413 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16307), .A(
        n16306), .ZN(n16311) );
  INV_X1 U19414 ( .A(n16308), .ZN(n19082) );
  AOI22_X1 U19415 ( .A1(n16309), .A2(n16379), .B1(n16407), .B2(n19082), .ZN(
        n16310) );
  OAI211_X1 U19416 ( .C1(n16404), .C2(n16312), .A(n16311), .B(n16310), .ZN(
        P2_U3028) );
  AOI21_X1 U19417 ( .B1(n16315), .B2(n16314), .A(n16313), .ZN(n19271) );
  NAND2_X1 U19418 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19412), .ZN(n16316) );
  OAI221_X1 U19419 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16319), 
        .C1(n16318), .C2(n16317), .A(n16316), .ZN(n16320) );
  AOI21_X1 U19420 ( .B1(n16399), .B2(n19271), .A(n16320), .ZN(n16323) );
  AOI22_X1 U19421 ( .A1(n19114), .A2(n16407), .B1(n16393), .B2(n16321), .ZN(
        n16322) );
  OAI211_X1 U19422 ( .C1(n16402), .C2(n16324), .A(n16323), .B(n16322), .ZN(
        P2_U3031) );
  NOR2_X1 U19423 ( .A1(n16326), .A2(n16325), .ZN(n16330) );
  OR2_X1 U19424 ( .A1(n16328), .A2(n16327), .ZN(n16329) );
  MUX2_X1 U19425 ( .A(n16330), .B(n16329), .S(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(n16336) );
  INV_X1 U19426 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20003) );
  AOI21_X1 U19427 ( .B1(n16332), .B2(n16331), .A(n9933), .ZN(n19275) );
  NAND2_X1 U19428 ( .A1(n16399), .A2(n19275), .ZN(n16333) );
  OAI21_X1 U19429 ( .B1(n20003), .B2(n16334), .A(n16333), .ZN(n16335) );
  NOR2_X1 U19430 ( .A1(n16336), .A2(n16335), .ZN(n16339) );
  AOI22_X1 U19431 ( .A1(n16337), .A2(n16393), .B1(n16407), .B2(n19138), .ZN(
        n16338) );
  OAI211_X1 U19432 ( .C1(n16402), .C2(n16340), .A(n16339), .B(n16338), .ZN(
        P2_U3033) );
  AOI21_X1 U19433 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n19279) );
  AOI22_X1 U19434 ( .A1(n16344), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16399), .B2(n19279), .ZN(n16354) );
  INV_X1 U19435 ( .A(n16345), .ZN(n16346) );
  OAI22_X1 U19436 ( .A1(n16346), .A2(n16402), .B1(n16365), .B2(n19162), .ZN(
        n16347) );
  AOI21_X1 U19437 ( .B1(n16393), .B2(n16348), .A(n16347), .ZN(n16353) );
  NAND2_X1 U19438 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19412), .ZN(n16352) );
  OAI211_X1 U19439 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16350), .B(n16349), .ZN(
        n16351) );
  NAND4_X1 U19440 ( .A1(n16354), .A2(n16353), .A3(n16352), .A4(n16351), .ZN(
        P2_U3035) );
  INV_X1 U19441 ( .A(n16355), .ZN(n16357) );
  NAND2_X1 U19442 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19412), .ZN(n16356) );
  OAI221_X1 U19443 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16359), .C1(
        n16358), .C2(n16357), .A(n16356), .ZN(n16367) );
  AOI21_X1 U19444 ( .B1(n16362), .B2(n16361), .A(n16360), .ZN(n19290) );
  INV_X1 U19445 ( .A(n19290), .ZN(n16363) );
  OAI22_X1 U19446 ( .A1(n19206), .A2(n16365), .B1(n16364), .B2(n16363), .ZN(
        n16366) );
  AOI211_X1 U19447 ( .C1(n16368), .C2(n16379), .A(n16367), .B(n16366), .ZN(
        n16369) );
  OAI21_X1 U19448 ( .B1(n16404), .B2(n16370), .A(n16369), .ZN(P2_U3039) );
  INV_X1 U19449 ( .A(n16371), .ZN(n16384) );
  OAI21_X1 U19450 ( .B1(n16410), .B2(n16384), .A(n16372), .ZN(n16377) );
  OAI21_X1 U19451 ( .B1(n16375), .B2(n16374), .A(n16373), .ZN(n16376) );
  INV_X1 U19452 ( .A(n16376), .ZN(n19292) );
  AOI22_X1 U19453 ( .A1(n16377), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16399), .B2(n19292), .ZN(n16388) );
  AOI222_X1 U19454 ( .A1(n16381), .A2(n16393), .B1(n16407), .B2(n16380), .C1(
        n16379), .C2(n16378), .ZN(n16387) );
  NAND2_X1 U19455 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19412), .ZN(n16386) );
  NAND3_X1 U19456 ( .A1(n16384), .A2(n16383), .A3(n16382), .ZN(n16385) );
  NAND4_X1 U19457 ( .A1(n16388), .A2(n16387), .A3(n16386), .A4(n16385), .ZN(
        P2_U3040) );
  AOI22_X1 U19458 ( .A1(n16399), .A2(n20058), .B1(n19412), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n16389) );
  OAI21_X1 U19459 ( .B1(n16390), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16389), .ZN(n16391) );
  AOI21_X1 U19460 ( .B1(n13396), .B2(n16407), .A(n16391), .ZN(n16396) );
  AOI22_X1 U19461 ( .A1(n16394), .A2(n16393), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16392), .ZN(n16395) );
  OAI211_X1 U19462 ( .C1(n16397), .C2(n16402), .A(n16396), .B(n16395), .ZN(
        P2_U3043) );
  INV_X1 U19463 ( .A(n16398), .ZN(n16400) );
  AOI22_X1 U19464 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16399), .B2(n19321), .ZN(n16409) );
  OAI22_X1 U19465 ( .A1(n16404), .A2(n16403), .B1(n16402), .B2(n16401), .ZN(
        n16405) );
  AOI211_X1 U19466 ( .C1(n16407), .C2(n13200), .A(n16406), .B(n16405), .ZN(
        n16408) );
  OAI211_X1 U19467 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16410), .A(
        n16409), .B(n16408), .ZN(P2_U3046) );
  INV_X1 U19468 ( .A(n16430), .ZN(n16413) );
  MUX2_X1 U19469 ( .A(n16412), .B(n16411), .S(n16413), .Z(n16429) );
  NAND2_X1 U19470 ( .A1(n16414), .A2(n16413), .ZN(n16417) );
  NAND2_X1 U19471 ( .A1(n16430), .A2(n16415), .ZN(n16416) );
  NAND2_X1 U19472 ( .A1(n16417), .A2(n16416), .ZN(n16423) );
  INV_X1 U19473 ( .A(n16423), .ZN(n16451) );
  NOR2_X1 U19474 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19538) );
  INV_X1 U19475 ( .A(n19538), .ZN(n19540) );
  OR2_X1 U19476 ( .A1(n16419), .A2(n20078), .ZN(n16421) );
  NAND2_X1 U19477 ( .A1(n16418), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16420) );
  AOI22_X1 U19478 ( .A1(n16421), .A2(n16420), .B1(n16419), .B2(n20078), .ZN(
        n16422) );
  OAI22_X1 U19479 ( .A1(n16423), .A2(n19540), .B1(n16430), .B2(n16422), .ZN(
        n16424) );
  OAI21_X1 U19480 ( .B1(n16451), .B2(n20069), .A(n16424), .ZN(n16425) );
  OAI21_X1 U19481 ( .B1(n16429), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16425), .ZN(n16428) );
  NAND2_X1 U19482 ( .A1(n16429), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16426) );
  NAND3_X1 U19483 ( .A1(n16428), .A2(n16427), .A3(n16426), .ZN(n16454) );
  INV_X1 U19484 ( .A(n16429), .ZN(n16452) );
  NAND2_X1 U19485 ( .A1(n16430), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16449) );
  INV_X1 U19486 ( .A(n16431), .ZN(n16437) );
  NAND2_X1 U19487 ( .A1(n16433), .A2(n16432), .ZN(n16436) );
  NAND2_X1 U19488 ( .A1(n16438), .A2(n16434), .ZN(n16435) );
  OAI211_X1 U19489 ( .C1(n16438), .C2(n16437), .A(n16436), .B(n16435), .ZN(
        n20095) );
  NOR2_X1 U19490 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16445) );
  NAND2_X1 U19491 ( .A1(n12403), .A2(n16439), .ZN(n16441) );
  OAI22_X1 U19492 ( .A1(n16442), .A2(n16441), .B1(n16440), .B2(n12813), .ZN(
        n16443) );
  INV_X1 U19493 ( .A(n16443), .ZN(n16444) );
  OAI21_X1 U19494 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(n16447) );
  NOR2_X1 U19495 ( .A1(n20095), .A2(n16447), .ZN(n16448) );
  NAND2_X1 U19496 ( .A1(n16449), .A2(n16448), .ZN(n16450) );
  AOI21_X1 U19497 ( .B1(n16452), .B2(n16451), .A(n16450), .ZN(n16453) );
  AND2_X1 U19498 ( .A1(n16454), .A2(n16453), .ZN(n16472) );
  INV_X1 U19499 ( .A(n20092), .ZN(n16456) );
  AOI211_X1 U19500 ( .C1(n16457), .C2(n16456), .A(n19951), .B(n16455), .ZN(
        n16470) );
  NAND2_X1 U19501 ( .A1(n16472), .A2(n13767), .ZN(n16458) );
  NAND2_X1 U19502 ( .A1(n16458), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16464) );
  NAND2_X1 U19503 ( .A1(n16459), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16460) );
  AOI21_X1 U19504 ( .B1(n16462), .B2(n16461), .A(n16460), .ZN(n16463) );
  AND2_X1 U19505 ( .A1(n16464), .A2(n16463), .ZN(n16468) );
  NOR2_X1 U19506 ( .A1(n19950), .A2(n19949), .ZN(n19952) );
  AOI211_X1 U19507 ( .C1(n16466), .C2(n16465), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n19952), .ZN(n16467) );
  AOI21_X1 U19508 ( .B1(n16468), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16467), 
        .ZN(n16469) );
  OAI211_X1 U19509 ( .C1(n16472), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        P2_U3176) );
  OAI221_X1 U19510 ( .B1(n20079), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n20079), 
        .C2(n19949), .A(n16473), .ZN(P2_U3593) );
  NAND2_X1 U19511 ( .A1(n16506), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16475) );
  XOR2_X1 U19512 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16475), .Z(
        n16533) );
  NAND4_X1 U19513 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16867) );
  NAND3_X1 U19514 ( .A1(n17854), .A2(n17852), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17815) );
  NAND2_X1 U19515 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17817) );
  NAND2_X1 U19516 ( .A1(n17803), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17776) );
  NAND2_X1 U19517 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17778) );
  NAND2_X1 U19518 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17746) );
  NAND2_X1 U19519 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U19520 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17663) );
  INV_X1 U19521 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18942) );
  NOR2_X1 U19522 ( .A1(n18942), .A2(n18339), .ZN(n16526) );
  NAND2_X1 U19523 ( .A1(n18957), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18029) );
  OAI21_X1 U19524 ( .B1(n18024), .B2(n17802), .A(n18685), .ZN(n17851) );
  INV_X1 U19525 ( .A(n17851), .ZN(n17777) );
  OR2_X1 U19526 ( .A1(n16477), .A2(n17777), .ZN(n16499) );
  XOR2_X1 U19527 ( .A(n10299), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16480) );
  NOR2_X1 U19528 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17802), .ZN(
        n16510) );
  NAND2_X1 U19529 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16512), .ZN(
        n16673) );
  INV_X1 U19530 ( .A(n16673), .ZN(n16479) );
  NAND2_X1 U19531 ( .A1(n18745), .A2(n16477), .ZN(n16478) );
  OAI211_X1 U19532 ( .C1(n16479), .C2(n18029), .A(n18028), .B(n16478), .ZN(
        n16511) );
  NOR2_X1 U19533 ( .A1(n16510), .A2(n16511), .ZN(n16498) );
  OAI22_X1 U19534 ( .A1(n16499), .A2(n16480), .B1(n16498), .B2(n10299), .ZN(
        n16481) );
  AOI211_X1 U19535 ( .C1(n17872), .C2(n17006), .A(n16526), .B(n16481), .ZN(
        n16496) );
  INV_X1 U19536 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16482) );
  AOI21_X1 U19537 ( .B1(n16486), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16483), .ZN(n16484) );
  NAND2_X1 U19538 ( .A1(n16482), .A2(n17811), .ZN(n16487) );
  NAND2_X1 U19539 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16482), .ZN(
        n16523) );
  NAND3_X1 U19540 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17933), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16488) );
  NAND2_X1 U19541 ( .A1(n16488), .A2(n16487), .ZN(n16489) );
  AND2_X2 U19542 ( .A1(n16492), .A2(n16491), .ZN(n16530) );
  NAND2_X1 U19543 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16508), .ZN(
        n16493) );
  XNOR2_X1 U19544 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16493), .ZN(
        n16528) );
  NOR2_X2 U19545 ( .A1(n10113), .A2(n16650), .ZN(n18000) );
  OAI211_X1 U19546 ( .C1(n17938), .C2(n16533), .A(n16496), .B(n16495), .ZN(
        P3_U2799) );
  INV_X2 U19547 ( .A(n17938), .ZN(n17889) );
  NAND2_X1 U19548 ( .A1(n16537), .A2(n9847), .ZN(n17685) );
  XOR2_X1 U19549 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9964), .Z(n16693) );
  NAND2_X1 U19550 ( .A1(n18357), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16497) );
  OAI221_X1 U19551 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16499), .C1(
        n10300), .C2(n16498), .A(n16497), .ZN(n16500) );
  AOI21_X1 U19552 ( .B1(n17872), .B2(n16693), .A(n16500), .ZN(n16504) );
  OAI22_X1 U19553 ( .A1(n16506), .A2(n17938), .B1(n16508), .B2(n18033), .ZN(
        n16502) );
  AOI22_X1 U19554 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16502), .B1(
        n17934), .B2(n16501), .ZN(n16503) );
  OAI211_X1 U19555 ( .C1(n17685), .C2(n16505), .A(n16504), .B(n16503), .ZN(
        P3_U2800) );
  NOR2_X1 U19556 ( .A1(n16506), .A2(n17938), .ZN(n16518) );
  NOR2_X1 U19557 ( .A1(n18041), .A2(n16507), .ZN(n16540) );
  NOR2_X1 U19558 ( .A1(n16507), .A2(n17659), .ZN(n16541) );
  NOR2_X1 U19559 ( .A1(n16508), .A2(n18033), .ZN(n16509) );
  OAI21_X1 U19560 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16541), .A(
        n16509), .ZN(n16515) );
  AOI21_X1 U19561 ( .B1(n10298), .B2(n16673), .A(n9964), .ZN(n16702) );
  OAI21_X1 U19562 ( .B1(n16510), .B2(n17872), .A(n16702), .ZN(n16514) );
  OAI221_X1 U19563 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16512), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18745), .A(n16511), .ZN(
        n16513) );
  NAND4_X1 U19564 ( .A1(n16516), .A2(n16515), .A3(n16514), .A4(n16513), .ZN(
        n16517) );
  AOI221_X1 U19565 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16518), 
        .C1(n16540), .C2(n16518), .A(n16517), .ZN(n16519) );
  OAI21_X1 U19566 ( .B1(n16520), .B2(n17893), .A(n16519), .ZN(P3_U2801) );
  OAI21_X1 U19567 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18340), .A(
        n16521), .ZN(n16527) );
  NOR4_X1 U19568 ( .A1(n16524), .A2(n16523), .A3(n18351), .A4(n16522), .ZN(
        n16525) );
  AOI211_X1 U19569 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16527), .A(
        n16526), .B(n16525), .ZN(n16532) );
  OAI211_X1 U19570 ( .C1(n16533), .C2(n18272), .A(n16532), .B(n16531), .ZN(
        P3_U2831) );
  INV_X1 U19571 ( .A(n18332), .ZN(n18802) );
  AOI22_X1 U19572 ( .A1(n18224), .A2(n18802), .B1(n18226), .B2(n18201), .ZN(
        n18137) );
  INV_X1 U19573 ( .A(n18137), .ZN(n16536) );
  NAND2_X1 U19574 ( .A1(n16537), .A2(n18110), .ZN(n18043) );
  NAND2_X1 U19575 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17661), .ZN(
        n17674) );
  AOI211_X1 U19576 ( .C1(n16538), .C2(n17675), .A(n17518), .B(n18797), .ZN(
        n16539) );
  AOI22_X1 U19577 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17661), .B2(n17811), .ZN(n17671) );
  NAND2_X1 U19578 ( .A1(n17671), .A2(n17670), .ZN(n17669) );
  INV_X1 U19579 ( .A(n18201), .ZN(n18225) );
  OAI22_X1 U19580 ( .A1(n16541), .A2(n18332), .B1(n16540), .B2(n18225), .ZN(
        n16544) );
  INV_X1 U19581 ( .A(n16542), .ZN(n16543) );
  NOR2_X1 U19582 ( .A1(n16544), .A2(n16543), .ZN(n16545) );
  NOR4_X1 U19583 ( .A1(n17811), .A2(n17686), .A3(n16546), .A4(n18361), .ZN(
        n16548) );
  NAND2_X1 U19584 ( .A1(n18357), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17664) );
  NOR3_X1 U19585 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16550) );
  NOR4_X1 U19586 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16549) );
  NAND4_X1 U19587 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16550), .A3(n16549), .A4(
        U215), .ZN(U213) );
  INV_X2 U19588 ( .A(U214), .ZN(n16598) );
  INV_X1 U19589 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16636) );
  OAI222_X1 U19590 ( .A1(U212), .A2(n19326), .B1(n16601), .B2(n19469), .C1(
        U214), .C2(n16636), .ZN(U216) );
  INV_X1 U19591 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16552) );
  INV_X1 U19592 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20372) );
  INV_X1 U19593 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19329) );
  OAI222_X1 U19594 ( .A1(U214), .A2(n16552), .B1(n16601), .B2(n20372), .C1(
        U212), .C2(n19329), .ZN(U217) );
  INV_X1 U19595 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n16553) );
  INV_X1 U19596 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20364) );
  INV_X1 U19597 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19332) );
  OAI222_X1 U19598 ( .A1(U214), .A2(n16553), .B1(n16601), .B2(n20364), .C1(
        U212), .C2(n19332), .ZN(U218) );
  INV_X2 U19599 ( .A(U212), .ZN(n16599) );
  AOI22_X1 U19600 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16598), .ZN(n16554) );
  OAI21_X1 U19601 ( .B1(n19451), .B2(n16601), .A(n16554), .ZN(U219) );
  AOI22_X1 U19602 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16598), .ZN(n16555) );
  OAI21_X1 U19603 ( .B1(n19444), .B2(n16601), .A(n16555), .ZN(U220) );
  AOI22_X1 U19604 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16598), .ZN(n16556) );
  OAI21_X1 U19605 ( .B1(n19438), .B2(n16601), .A(n16556), .ZN(U221) );
  AOI22_X1 U19606 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16598), .ZN(n16557) );
  OAI21_X1 U19607 ( .B1(n20354), .B2(n16601), .A(n16557), .ZN(U222) );
  AOI22_X1 U19608 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16598), .ZN(n16558) );
  OAI21_X1 U19609 ( .B1(n16559), .B2(n16601), .A(n16558), .ZN(U223) );
  AOI22_X1 U19610 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16598), .ZN(n16560) );
  OAI21_X1 U19611 ( .B1(n16561), .B2(n16601), .A(n16560), .ZN(U224) );
  INV_X1 U19612 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20378) );
  AOI22_X1 U19613 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16598), .ZN(n16562) );
  OAI21_X1 U19614 ( .B1(n20378), .B2(n16601), .A(n16562), .ZN(U225) );
  INV_X1 U19615 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20368) );
  AOI22_X1 U19616 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16598), .ZN(n16563) );
  OAI21_X1 U19617 ( .B1(n20368), .B2(n16601), .A(n16563), .ZN(U226) );
  AOI22_X1 U19618 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16598), .ZN(n16564) );
  OAI21_X1 U19619 ( .B1(n16565), .B2(n16601), .A(n16564), .ZN(U227) );
  AOI22_X1 U19620 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16598), .ZN(n16566) );
  OAI21_X1 U19621 ( .B1(n16567), .B2(n16601), .A(n16566), .ZN(U228) );
  AOI22_X1 U19622 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16598), .ZN(n16568) );
  OAI21_X1 U19623 ( .B1(n16569), .B2(n16601), .A(n16568), .ZN(U229) );
  INV_X1 U19624 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20359) );
  AOI22_X1 U19625 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16598), .ZN(n16570) );
  OAI21_X1 U19626 ( .B1(n20359), .B2(n16601), .A(n16570), .ZN(U230) );
  AOI22_X1 U19627 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16598), .ZN(n16571) );
  OAI21_X1 U19628 ( .B1(n16572), .B2(n16601), .A(n16571), .ZN(U231) );
  AOI22_X1 U19629 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16598), .ZN(n16573) );
  OAI21_X1 U19630 ( .B1(n14368), .B2(n16601), .A(n16573), .ZN(U232) );
  AOI22_X1 U19631 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16598), .ZN(n16574) );
  OAI21_X1 U19632 ( .B1(n16575), .B2(n16601), .A(n16574), .ZN(U233) );
  INV_X1 U19633 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16577) );
  AOI22_X1 U19634 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16598), .ZN(n16576) );
  OAI21_X1 U19635 ( .B1(n16577), .B2(n16601), .A(n16576), .ZN(U234) );
  INV_X1 U19636 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16579) );
  AOI22_X1 U19637 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16598), .ZN(n16578) );
  OAI21_X1 U19638 ( .B1(n16579), .B2(n16601), .A(n16578), .ZN(U235) );
  AOI22_X1 U19639 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16598), .ZN(n16580) );
  OAI21_X1 U19640 ( .B1(n16581), .B2(n16601), .A(n16580), .ZN(U236) );
  AOI22_X1 U19641 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16598), .ZN(n16582) );
  OAI21_X1 U19642 ( .B1(n16583), .B2(n16601), .A(n16582), .ZN(U237) );
  AOI22_X1 U19643 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16598), .ZN(n16584) );
  OAI21_X1 U19644 ( .B1(n16585), .B2(n16601), .A(n16584), .ZN(U238) );
  AOI22_X1 U19645 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16598), .ZN(n16586) );
  OAI21_X1 U19646 ( .B1(n16587), .B2(n16601), .A(n16586), .ZN(U239) );
  AOI22_X1 U19647 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16598), .ZN(n16588) );
  OAI21_X1 U19648 ( .B1(n16589), .B2(n16601), .A(n16588), .ZN(U240) );
  AOI22_X1 U19649 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16598), .ZN(n16590) );
  OAI21_X1 U19650 ( .B1(n13551), .B2(n16601), .A(n16590), .ZN(U241) );
  INV_X1 U19651 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16592) );
  AOI22_X1 U19652 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16598), .ZN(n16591) );
  OAI21_X1 U19653 ( .B1(n16592), .B2(n16601), .A(n16591), .ZN(U242) );
  AOI22_X1 U19654 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16598), .ZN(n16593) );
  OAI21_X1 U19655 ( .B1(n13342), .B2(n16601), .A(n16593), .ZN(U243) );
  AOI22_X1 U19656 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16598), .ZN(n16594) );
  OAI21_X1 U19657 ( .B1(n13189), .B2(n16601), .A(n16594), .ZN(U244) );
  INV_X1 U19658 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16596) );
  AOI22_X1 U19659 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16598), .ZN(n16595) );
  OAI21_X1 U19660 ( .B1(n16596), .B2(n16601), .A(n16595), .ZN(U245) );
  AOI22_X1 U19661 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16598), .ZN(n16597) );
  OAI21_X1 U19662 ( .B1(n13113), .B2(n16601), .A(n16597), .ZN(U246) );
  INV_X1 U19663 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16602) );
  AOI22_X1 U19664 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16599), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16598), .ZN(n16600) );
  OAI21_X1 U19665 ( .B1(n16602), .B2(n16601), .A(n16600), .ZN(U247) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16634), .ZN(n16603) );
  INV_X1 U19667 ( .A(n16603), .ZN(U251) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16631), .ZN(n16604) );
  INV_X1 U19669 ( .A(n16604), .ZN(U252) );
  INV_X1 U19670 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16605) );
  INV_X1 U19671 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U19672 ( .A1(n16634), .A2(n16605), .B1(n18382), .B2(U215), .ZN(U253) );
  INV_X1 U19673 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16606) );
  INV_X1 U19674 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18386) );
  AOI22_X1 U19675 ( .A1(n16634), .A2(n16606), .B1(n18386), .B2(U215), .ZN(U254) );
  OAI22_X1 U19676 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16631), .ZN(n16607) );
  INV_X1 U19677 ( .A(n16607), .ZN(U255) );
  INV_X1 U19678 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16608) );
  INV_X1 U19679 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U19680 ( .A1(n16634), .A2(n16608), .B1(n18394), .B2(U215), .ZN(U256) );
  OAI22_X1 U19681 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16631), .ZN(n16609) );
  INV_X1 U19682 ( .A(n16609), .ZN(U257) );
  INV_X1 U19683 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16610) );
  INV_X1 U19684 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18402) );
  AOI22_X1 U19685 ( .A1(n16634), .A2(n16610), .B1(n18402), .B2(U215), .ZN(U258) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16634), .ZN(n16611) );
  INV_X1 U19687 ( .A(n16611), .ZN(U259) );
  INV_X1 U19688 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16612) );
  INV_X1 U19689 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U19690 ( .A1(n16634), .A2(n16612), .B1(n17511), .B2(U215), .ZN(U260) );
  OAI22_X1 U19691 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16634), .ZN(n16613) );
  INV_X1 U19692 ( .A(n16613), .ZN(U261) );
  INV_X1 U19693 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16615) );
  INV_X1 U19694 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n16614) );
  AOI22_X1 U19695 ( .A1(n16631), .A2(n16615), .B1(n16614), .B2(U215), .ZN(U262) );
  INV_X1 U19696 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16616) );
  INV_X1 U19697 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U19698 ( .A1(n16631), .A2(n16616), .B1(n17499), .B2(U215), .ZN(U263) );
  INV_X1 U19699 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16617) );
  INV_X1 U19700 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U19701 ( .A1(n16634), .A2(n16617), .B1(n17494), .B2(U215), .ZN(U264) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16634), .ZN(n16618) );
  INV_X1 U19703 ( .A(n16618), .ZN(U265) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16634), .ZN(n16619) );
  INV_X1 U19705 ( .A(n16619), .ZN(U266) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16634), .ZN(n16620) );
  INV_X1 U19707 ( .A(n16620), .ZN(U267) );
  OAI22_X1 U19708 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16634), .ZN(n16621) );
  INV_X1 U19709 ( .A(n16621), .ZN(U268) );
  OAI22_X1 U19710 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16634), .ZN(n16622) );
  INV_X1 U19711 ( .A(n16622), .ZN(U269) );
  OAI22_X1 U19712 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16634), .ZN(n16623) );
  INV_X1 U19713 ( .A(n16623), .ZN(U270) );
  INV_X1 U19714 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16624) );
  INV_X1 U19715 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18390) );
  AOI22_X1 U19716 ( .A1(n16631), .A2(n16624), .B1(n18390), .B2(U215), .ZN(U271) );
  OAI22_X1 U19717 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16631), .ZN(n16625) );
  INV_X1 U19718 ( .A(n16625), .ZN(U272) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16631), .ZN(n16626) );
  INV_X1 U19720 ( .A(n16626), .ZN(U273) );
  OAI22_X1 U19721 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16631), .ZN(n16627) );
  INV_X1 U19722 ( .A(n16627), .ZN(U274) );
  INV_X1 U19723 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16628) );
  AOI22_X1 U19724 ( .A1(n16634), .A2(n16628), .B1(n18375), .B2(U215), .ZN(U275) );
  INV_X1 U19725 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19726 ( .A1(n16634), .A2(n16629), .B1(n18378), .B2(U215), .ZN(U276) );
  INV_X1 U19727 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16630) );
  INV_X1 U19728 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19437) );
  AOI22_X1 U19729 ( .A1(n16631), .A2(n16630), .B1(n19437), .B2(U215), .ZN(U277) );
  INV_X1 U19730 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16632) );
  INV_X1 U19731 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19445) );
  AOI22_X1 U19732 ( .A1(n16634), .A2(n16632), .B1(n19445), .B2(U215), .ZN(U278) );
  INV_X1 U19733 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16633) );
  INV_X1 U19734 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19450) );
  AOI22_X1 U19735 ( .A1(n16634), .A2(n16633), .B1(n19450), .B2(U215), .ZN(U279) );
  INV_X1 U19736 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19456) );
  AOI22_X1 U19737 ( .A1(n16634), .A2(n19332), .B1(n19456), .B2(U215), .ZN(U280) );
  INV_X1 U19738 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19460) );
  AOI22_X1 U19739 ( .A1(n16634), .A2(n19329), .B1(n19460), .B2(U215), .ZN(U281) );
  INV_X1 U19740 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19467) );
  AOI22_X1 U19741 ( .A1(n16634), .A2(n19326), .B1(n19467), .B2(U215), .ZN(U282) );
  INV_X1 U19742 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16635) );
  AOI222_X1 U19743 ( .A1(n19326), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16636), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16635), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16637) );
  INV_X2 U19744 ( .A(n16639), .ZN(n16638) );
  INV_X1 U19745 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18902) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19998) );
  AOI22_X1 U19747 ( .A1(n16638), .A2(n18902), .B1(n19998), .B2(n16639), .ZN(
        U347) );
  INV_X1 U19748 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18900) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19996) );
  AOI22_X1 U19750 ( .A1(n16638), .A2(n18900), .B1(n19996), .B2(n16639), .ZN(
        U348) );
  INV_X1 U19751 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18897) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19994) );
  AOI22_X1 U19753 ( .A1(n16638), .A2(n18897), .B1(n19994), .B2(n16639), .ZN(
        U349) );
  INV_X1 U19754 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18896) );
  INV_X1 U19755 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19992) );
  AOI22_X1 U19756 ( .A1(n16638), .A2(n18896), .B1(n19992), .B2(n16639), .ZN(
        U350) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18894) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19990) );
  AOI22_X1 U19759 ( .A1(n16638), .A2(n18894), .B1(n19990), .B2(n16639), .ZN(
        U351) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18892) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19988) );
  AOI22_X1 U19762 ( .A1(n16638), .A2(n18892), .B1(n19988), .B2(n16639), .ZN(
        U352) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18890) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U19765 ( .A1(n16638), .A2(n18890), .B1(n19986), .B2(n16639), .ZN(
        U353) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18888) );
  AOI22_X1 U19767 ( .A1(n16638), .A2(n18888), .B1(n19983), .B2(n16639), .ZN(
        U354) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18941) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20037) );
  AOI22_X1 U19770 ( .A1(n16638), .A2(n18941), .B1(n20037), .B2(n16639), .ZN(
        U356) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18938) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20034) );
  AOI22_X1 U19773 ( .A1(n16638), .A2(n18938), .B1(n20034), .B2(n16639), .ZN(
        U357) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18937) );
  INV_X1 U19775 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20031) );
  AOI22_X1 U19776 ( .A1(n16638), .A2(n18937), .B1(n20031), .B2(n16639), .ZN(
        U358) );
  INV_X1 U19777 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18934) );
  INV_X1 U19778 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20030) );
  AOI22_X1 U19779 ( .A1(n16638), .A2(n18934), .B1(n20030), .B2(n16639), .ZN(
        U359) );
  INV_X1 U19780 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18932) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U19782 ( .A1(n16638), .A2(n18932), .B1(n20028), .B2(n16639), .ZN(
        U360) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18930) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20026) );
  AOI22_X1 U19785 ( .A1(n16638), .A2(n18930), .B1(n20026), .B2(n16639), .ZN(
        U361) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18927) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U19788 ( .A1(n16638), .A2(n18927), .B1(n20024), .B2(n16639), .ZN(
        U362) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18926) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U19791 ( .A1(n16638), .A2(n18926), .B1(n20022), .B2(n16639), .ZN(
        U363) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18923) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20020) );
  AOI22_X1 U19794 ( .A1(n16638), .A2(n18923), .B1(n20020), .B2(n16639), .ZN(
        U364) );
  INV_X1 U19795 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18886) );
  INV_X1 U19796 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U19797 ( .A1(n16638), .A2(n18886), .B1(n19981), .B2(n16639), .ZN(
        U365) );
  INV_X1 U19798 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18922) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U19800 ( .A1(n16638), .A2(n18922), .B1(n20018), .B2(n16639), .ZN(
        U366) );
  INV_X1 U19801 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18919) );
  INV_X1 U19802 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U19803 ( .A1(n16638), .A2(n18919), .B1(n20016), .B2(n16639), .ZN(
        U367) );
  INV_X1 U19804 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18918) );
  INV_X1 U19805 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20014) );
  AOI22_X1 U19806 ( .A1(n16638), .A2(n18918), .B1(n20014), .B2(n16639), .ZN(
        U368) );
  INV_X1 U19807 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18916) );
  INV_X1 U19808 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U19809 ( .A1(n16638), .A2(n18916), .B1(n20012), .B2(n16639), .ZN(
        U369) );
  INV_X1 U19810 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18914) );
  INV_X1 U19811 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U19812 ( .A1(n16638), .A2(n18914), .B1(n20010), .B2(n16639), .ZN(
        U370) );
  INV_X1 U19813 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18912) );
  INV_X1 U19814 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U19815 ( .A1(n16638), .A2(n18912), .B1(n20008), .B2(n16639), .ZN(
        U371) );
  INV_X1 U19816 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18910) );
  INV_X1 U19817 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U19818 ( .A1(n16638), .A2(n18910), .B1(n20006), .B2(n16639), .ZN(
        U372) );
  INV_X1 U19819 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18908) );
  INV_X1 U19820 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U19821 ( .A1(n16638), .A2(n18908), .B1(n20004), .B2(n16639), .ZN(
        U373) );
  INV_X1 U19822 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18906) );
  INV_X1 U19823 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U19824 ( .A1(n16638), .A2(n18906), .B1(n20002), .B2(n16639), .ZN(
        U374) );
  INV_X1 U19825 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18904) );
  INV_X1 U19826 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U19827 ( .A1(n16638), .A2(n18904), .B1(n20000), .B2(n16639), .ZN(
        U375) );
  INV_X1 U19828 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18884) );
  INV_X1 U19829 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U19830 ( .A1(n16638), .A2(n18884), .B1(n19980), .B2(n16639), .ZN(
        U376) );
  INV_X1 U19831 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16642) );
  NAND2_X1 U19832 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18883), .ZN(n16641) );
  NAND2_X1 U19833 ( .A1(n18880), .A2(n16640), .ZN(n18870) );
  OAI21_X1 U19834 ( .B1(n16641), .B2(n18880), .A(n18870), .ZN(n18956) );
  OAI21_X1 U19835 ( .B1(n18880), .B2(n16642), .A(n9797), .ZN(P3_U2633) );
  OAI21_X1 U19836 ( .B1(n16649), .B2(n17588), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16643) );
  OAI21_X1 U19837 ( .B1(n16644), .B2(n18857), .A(n16643), .ZN(P3_U2634) );
  AOI21_X1 U19838 ( .B1(n18880), .B2(n18883), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16645) );
  AOI22_X1 U19839 ( .A1(n18999), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16645), 
        .B2(n19020), .ZN(P3_U2635) );
  INV_X1 U19840 ( .A(BS16), .ZN(n21108) );
  AOI21_X1 U19841 ( .B1(n18869), .B2(n21108), .A(n9797), .ZN(n18952) );
  INV_X1 U19842 ( .A(n18952), .ZN(n18954) );
  OAI21_X1 U19843 ( .B1(n18956), .B2(n19011), .A(n18954), .ZN(P3_U2636) );
  INV_X1 U19844 ( .A(n16646), .ZN(n16647) );
  NOR3_X1 U19845 ( .A1(n16649), .A2(n16648), .A3(n16647), .ZN(n18843) );
  NOR2_X1 U19846 ( .A1(n18843), .A2(n18847), .ZN(n19000) );
  OAI21_X1 U19847 ( .B1(n19000), .B2(n16651), .A(n16650), .ZN(P3_U2637) );
  NOR4_X1 U19848 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16655) );
  NOR4_X1 U19849 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16654) );
  NOR4_X1 U19850 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16653) );
  NOR4_X1 U19851 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16652) );
  NAND4_X1 U19852 ( .A1(n16655), .A2(n16654), .A3(n16653), .A4(n16652), .ZN(
        n16661) );
  NOR4_X1 U19853 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16659) );
  AOI211_X1 U19854 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16658) );
  NOR4_X1 U19855 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16657) );
  NOR4_X1 U19856 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16656) );
  NAND4_X1 U19857 ( .A1(n16659), .A2(n16658), .A3(n16657), .A4(n16656), .ZN(
        n16660) );
  NOR2_X1 U19858 ( .A1(n16661), .A2(n16660), .ZN(n18997) );
  INV_X1 U19859 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18950) );
  NOR3_X1 U19860 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16663) );
  OAI21_X1 U19861 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16663), .A(n18997), .ZN(
        n16662) );
  OAI21_X1 U19862 ( .B1(n18997), .B2(n18950), .A(n16662), .ZN(P3_U2638) );
  INV_X1 U19863 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18990) );
  INV_X1 U19864 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18955) );
  AOI21_X1 U19865 ( .B1(n18990), .B2(n18955), .A(n16663), .ZN(n16664) );
  INV_X1 U19866 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18947) );
  INV_X1 U19867 ( .A(n18997), .ZN(n18992) );
  AOI22_X1 U19868 ( .A1(n18997), .A2(n16664), .B1(n18947), .B2(n18992), .ZN(
        P3_U2639) );
  NAND2_X1 U19869 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18856), .ZN(n18858) );
  NAND3_X1 U19870 ( .A1(n18957), .A2(n18856), .A3(n19011), .ZN(n18865) );
  NOR2_X1 U19871 ( .A1(n18297), .A2(n17014), .ZN(n16667) );
  INV_X1 U19872 ( .A(n19009), .ZN(n19023) );
  AOI211_X1 U19873 ( .C1(n19012), .C2(n19010), .A(n19007), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18849) );
  NAND2_X1 U19874 ( .A1(n19009), .A2(n18372), .ZN(n16671) );
  AOI211_X4 U19875 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n10113), .A(n18849), .B(
        n16671), .ZN(n17052) );
  INV_X1 U19876 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18944) );
  INV_X1 U19877 ( .A(n16671), .ZN(n16668) );
  INV_X1 U19878 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18931) );
  INV_X1 U19879 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18928) );
  INV_X1 U19880 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18921) );
  INV_X1 U19881 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18917) );
  INV_X1 U19882 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18913) );
  INV_X1 U19883 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18911) );
  INV_X1 U19884 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18903) );
  INV_X1 U19885 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18898) );
  INV_X1 U19886 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18893) );
  INV_X1 U19887 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18889) );
  NAND3_X1 U19888 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16990) );
  NOR2_X1 U19889 ( .A1(n18889), .A2(n16990), .ZN(n16986) );
  NAND2_X1 U19890 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16986), .ZN(n16985) );
  NOR2_X1 U19891 ( .A1(n18893), .A2(n16985), .ZN(n16951) );
  NAND2_X1 U19892 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16951), .ZN(n16946) );
  OR2_X1 U19893 ( .A1(n18898), .A2(n16946), .ZN(n16913) );
  INV_X1 U19894 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18901) );
  INV_X1 U19895 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18899) );
  NOR4_X1 U19896 ( .A1(n18903), .A2(n16913), .A3(n18901), .A4(n18899), .ZN(
        n16893) );
  AND2_X1 U19897 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16893), .ZN(n16869) );
  NAND3_X1 U19898 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16869), .ZN(n16854) );
  NOR3_X1 U19899 ( .A1(n18913), .A2(n18911), .A3(n16854), .ZN(n16833) );
  NAND2_X1 U19900 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16833), .ZN(n16805) );
  NOR2_X1 U19901 ( .A1(n18917), .A2(n16805), .ZN(n16810) );
  NAND2_X1 U19902 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16810), .ZN(n16799) );
  NAND3_X1 U19903 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n16800), .ZN(n16768) );
  NOR2_X1 U19904 ( .A1(n18928), .A2(n16768), .ZN(n16766) );
  NAND2_X1 U19905 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16766), .ZN(n16746) );
  NOR2_X1 U19906 ( .A1(n18931), .A2(n16746), .ZN(n16732) );
  NAND2_X1 U19907 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16732), .ZN(n16684) );
  NOR2_X1 U19908 ( .A1(n17045), .A2(n16684), .ZN(n16727) );
  NAND4_X1 U19909 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16727), .ZN(n16683) );
  NOR3_X1 U19910 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18944), .A3(n16683), 
        .ZN(n16669) );
  AOI21_X1 U19911 ( .B1(n17052), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16669), .ZN(
        n16690) );
  NAND2_X1 U19912 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n10113), .ZN(n16670) );
  AOI211_X4 U19913 ( .C1(n19011), .C2(n19013), .A(n16671), .B(n16670), .ZN(
        n17051) );
  NOR3_X1 U19914 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17020) );
  INV_X1 U19915 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17377) );
  NAND2_X1 U19916 ( .A1(n17020), .A2(n17377), .ZN(n17015) );
  NOR2_X1 U19917 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17015), .ZN(n16991) );
  NAND2_X1 U19918 ( .A1(n16991), .A2(n16989), .ZN(n16981) );
  NAND2_X1 U19919 ( .A1(n16965), .A2(n16960), .ZN(n16959) );
  NAND2_X1 U19920 ( .A1(n16927), .A2(n16940), .ZN(n16915) );
  NAND2_X1 U19921 ( .A1(n16914), .A2(n16910), .ZN(n16909) );
  NAND2_X1 U19922 ( .A1(n16890), .A2(n16882), .ZN(n16881) );
  INV_X1 U19923 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17236) );
  NAND2_X1 U19924 ( .A1(n16868), .A2(n17236), .ZN(n16858) );
  INV_X1 U19925 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16841) );
  NAND2_X1 U19926 ( .A1(n16844), .A2(n16841), .ZN(n16838) );
  INV_X1 U19927 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16817) );
  NAND2_X1 U19928 ( .A1(n16818), .A2(n16817), .ZN(n16814) );
  NAND2_X1 U19929 ( .A1(n16796), .A2(n16790), .ZN(n16789) );
  NAND2_X1 U19930 ( .A1(n16775), .A2(n17061), .ZN(n16771) );
  NAND2_X1 U19931 ( .A1(n16755), .A2(n16750), .ZN(n16749) );
  NOR2_X1 U19932 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16749), .ZN(n16733) );
  INV_X1 U19933 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U19934 ( .A1(n16733), .A2(n16729), .ZN(n16728) );
  NOR2_X1 U19935 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16728), .ZN(n16712) );
  INV_X1 U19936 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17062) );
  NAND2_X1 U19937 ( .A1(n16712), .A2(n17062), .ZN(n16691) );
  NOR2_X1 U19938 ( .A1(n17044), .A2(n16691), .ZN(n16697) );
  INV_X1 U19939 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17067) );
  INV_X1 U19940 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17682) );
  INV_X1 U19941 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16680) );
  INV_X1 U19942 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16830) );
  NAND2_X1 U19943 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17803), .ZN(
        n16843) );
  INV_X1 U19944 ( .A(n17775), .ZN(n16672) );
  NOR2_X1 U19945 ( .A1(n17778), .A2(n16672), .ZN(n17742) );
  INV_X1 U19946 ( .A(n17742), .ZN(n16807) );
  NAND2_X1 U19947 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16682), .ZN(
        n16681) );
  NAND2_X1 U19948 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17700), .ZN(
        n16679) );
  NAND2_X1 U19949 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17657), .ZN(
        n16675) );
  NOR2_X1 U19950 ( .A1(n17682), .A2(n16675), .ZN(n16674) );
  OAI21_X1 U19951 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16674), .A(
        n16673), .ZN(n17666) );
  INV_X1 U19952 ( .A(n17666), .ZN(n16715) );
  AOI21_X1 U19953 ( .B1(n17682), .B2(n16675), .A(n16674), .ZN(n17678) );
  OAI21_X1 U19954 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17657), .A(
        n16675), .ZN(n16676) );
  INV_X1 U19955 ( .A(n16676), .ZN(n17693) );
  INV_X1 U19956 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17718) );
  NOR2_X1 U19957 ( .A1(n17718), .A2(n16679), .ZN(n16678) );
  INV_X1 U19958 ( .A(n17657), .ZN(n16677) );
  OAI21_X1 U19959 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16678), .A(
        n16677), .ZN(n17705) );
  INV_X1 U19960 ( .A(n17705), .ZN(n16744) );
  AOI21_X1 U19961 ( .B1(n17718), .B2(n16679), .A(n16678), .ZN(n17714) );
  OAI21_X1 U19962 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17700), .A(
        n16679), .ZN(n17732) );
  INV_X1 U19963 ( .A(n17732), .ZN(n16765) );
  AOI21_X1 U19964 ( .B1(n16680), .B2(n16681), .A(n17700), .ZN(n17744) );
  OAI21_X1 U19965 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16682), .A(
        n16681), .ZN(n17752) );
  INV_X1 U19966 ( .A(n17752), .ZN(n16785) );
  AOI21_X1 U19967 ( .B1(n10286), .B2(n16807), .A(n16682), .ZN(n17768) );
  NAND2_X1 U19968 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17775), .ZN(
        n16820) );
  INV_X1 U19969 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16861) );
  NOR2_X1 U19970 ( .A1(n18024), .A2(n17815), .ZN(n17816) );
  INV_X1 U19971 ( .A(n17816), .ZN(n16853) );
  NOR2_X1 U19972 ( .A1(n16861), .A2(n16853), .ZN(n16852) );
  INV_X1 U19973 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16978) );
  NAND2_X1 U19974 ( .A1(n16852), .A2(n16978), .ZN(n16845) );
  NOR2_X1 U19975 ( .A1(n16820), .A2(n16845), .ZN(n16806) );
  AOI21_X1 U19976 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16806), .A(
        n16977), .ZN(n16795) );
  NOR2_X1 U19977 ( .A1(n17768), .A2(n16795), .ZN(n16794) );
  NOR2_X1 U19978 ( .A1(n16794), .A2(n16977), .ZN(n16784) );
  NOR2_X1 U19979 ( .A1(n16785), .A2(n16784), .ZN(n16783) );
  NOR2_X1 U19980 ( .A1(n16783), .A2(n16977), .ZN(n16777) );
  NOR2_X1 U19981 ( .A1(n17744), .A2(n16777), .ZN(n16776) );
  NOR2_X1 U19982 ( .A1(n16776), .A2(n16977), .ZN(n16764) );
  NOR2_X1 U19983 ( .A1(n16765), .A2(n16764), .ZN(n16763) );
  NOR2_X1 U19984 ( .A1(n16763), .A2(n16977), .ZN(n16757) );
  NOR2_X1 U19985 ( .A1(n17714), .A2(n16757), .ZN(n16756) );
  NOR2_X1 U19986 ( .A1(n16756), .A2(n16977), .ZN(n16743) );
  NOR2_X1 U19987 ( .A1(n16744), .A2(n16743), .ZN(n16742) );
  NOR2_X1 U19988 ( .A1(n16742), .A2(n16977), .ZN(n16735) );
  NOR2_X1 U19989 ( .A1(n17693), .A2(n16735), .ZN(n16734) );
  NOR2_X1 U19990 ( .A1(n16734), .A2(n16977), .ZN(n16724) );
  NOR2_X1 U19991 ( .A1(n17678), .A2(n16724), .ZN(n16723) );
  NOR2_X1 U19992 ( .A1(n16723), .A2(n16977), .ZN(n16714) );
  NOR2_X1 U19993 ( .A1(n16715), .A2(n16714), .ZN(n16713) );
  NOR2_X1 U19994 ( .A1(n16713), .A2(n16977), .ZN(n16701) );
  NOR2_X1 U19995 ( .A1(n16702), .A2(n16701), .ZN(n16700) );
  NOR2_X1 U19996 ( .A1(n16700), .A2(n16977), .ZN(n16692) );
  NAND2_X1 U19997 ( .A1(n17006), .A2(n17014), .ZN(n16842) );
  NOR3_X1 U19998 ( .A1(n16693), .A2(n16692), .A3(n16842), .ZN(n16688) );
  NOR2_X1 U19999 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16683), .ZN(n16695) );
  INV_X1 U20000 ( .A(n16695), .ZN(n16686) );
  NAND3_X1 U20001 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16685) );
  INV_X1 U20002 ( .A(n17055), .ZN(n17043) );
  OR2_X1 U20003 ( .A1(n16684), .A2(n17043), .ZN(n16711) );
  NAND2_X1 U20004 ( .A1(n17045), .A2(n17055), .ZN(n17054) );
  OAI21_X1 U20005 ( .B1(n16685), .B2(n16711), .A(n17054), .ZN(n16710) );
  AOI21_X1 U20006 ( .B1(n16686), .B2(n16710), .A(n18942), .ZN(n16687) );
  AOI211_X1 U20007 ( .C1(n16697), .C2(n17067), .A(n16688), .B(n16687), .ZN(
        n16689) );
  OAI211_X1 U20008 ( .C1(n10299), .C2(n17019), .A(n16690), .B(n16689), .ZN(
        P3_U2640) );
  NAND2_X1 U20009 ( .A1(n17051), .A2(n16691), .ZN(n16706) );
  XOR2_X1 U20010 ( .A(n16693), .B(n16692), .Z(n16696) );
  OAI22_X1 U20011 ( .A1(n10300), .A2(n17019), .B1(n18944), .B2(n16710), .ZN(
        n16694) );
  AOI211_X1 U20012 ( .C1(n16696), .C2(n17014), .A(n16695), .B(n16694), .ZN(
        n16699) );
  OAI21_X1 U20013 ( .B1(n17052), .B2(n16697), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16698) );
  OAI211_X1 U20014 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16706), .A(n16699), .B(
        n16698), .ZN(P3_U2641) );
  INV_X1 U20015 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18940) );
  AOI211_X1 U20016 ( .C1(n16702), .C2(n16701), .A(n16700), .B(n18863), .ZN(
        n16705) );
  NAND3_X1 U20017 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16727), .ZN(n16703) );
  OAI22_X1 U20018 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16703), .B1(n10298), 
        .B2(n17019), .ZN(n16704) );
  AOI211_X1 U20019 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17052), .A(n16705), .B(
        n16704), .ZN(n16709) );
  INV_X1 U20020 ( .A(n16706), .ZN(n16707) );
  OAI21_X1 U20021 ( .B1(n16712), .B2(n17062), .A(n16707), .ZN(n16708) );
  OAI211_X1 U20022 ( .C1(n16710), .C2(n18940), .A(n16709), .B(n16708), .ZN(
        P3_U2642) );
  AOI22_X1 U20023 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17037), .B1(
        n17052), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16722) );
  NAND2_X1 U20024 ( .A1(n17054), .A2(n16711), .ZN(n16740) );
  INV_X1 U20025 ( .A(n16740), .ZN(n16718) );
  AOI211_X1 U20026 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16728), .A(n16712), .B(
        n17044), .ZN(n16717) );
  AOI211_X1 U20027 ( .C1(n16715), .C2(n16714), .A(n16713), .B(n18863), .ZN(
        n16716) );
  AOI211_X1 U20028 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16718), .A(n16717), 
        .B(n16716), .ZN(n16721) );
  NAND2_X1 U20029 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16719) );
  OAI211_X1 U20030 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16727), .B(n16719), .ZN(n16720) );
  NAND3_X1 U20031 ( .A1(n16722), .A2(n16721), .A3(n16720), .ZN(P3_U2643) );
  INV_X1 U20032 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18936) );
  AOI211_X1 U20033 ( .C1(n17678), .C2(n16724), .A(n16723), .B(n18863), .ZN(
        n16726) );
  OAI22_X1 U20034 ( .A1(n17682), .A2(n17019), .B1(n17026), .B2(n16729), .ZN(
        n16725) );
  AOI211_X1 U20035 ( .C1(n16727), .C2(n18936), .A(n16726), .B(n16725), .ZN(
        n16731) );
  OAI211_X1 U20036 ( .C1(n16733), .C2(n16729), .A(n17051), .B(n16728), .ZN(
        n16730) );
  OAI211_X1 U20037 ( .C1(n16740), .C2(n18936), .A(n16731), .B(n16730), .ZN(
        P3_U2644) );
  AOI21_X1 U20038 ( .B1(n17023), .B2(n16732), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16741) );
  AOI22_X1 U20039 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17037), .B1(
        n17052), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16739) );
  AOI211_X1 U20040 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16749), .A(n16733), .B(
        n17044), .ZN(n16737) );
  AOI211_X1 U20041 ( .C1(n17693), .C2(n16735), .A(n16734), .B(n18863), .ZN(
        n16736) );
  NOR2_X1 U20042 ( .A1(n16737), .A2(n16736), .ZN(n16738) );
  OAI211_X1 U20043 ( .C1(n16741), .C2(n16740), .A(n16739), .B(n16738), .ZN(
        P3_U2645) );
  INV_X1 U20044 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18929) );
  OAI21_X1 U20045 ( .B1(n16766), .B2(n17045), .A(n17055), .ZN(n16762) );
  AOI21_X1 U20046 ( .B1(n17023), .B2(n18929), .A(n16762), .ZN(n16753) );
  AOI211_X1 U20047 ( .C1(n16744), .C2(n16743), .A(n16742), .B(n18863), .ZN(
        n16748) );
  NAND2_X1 U20048 ( .A1(n17023), .A2(n18931), .ZN(n16745) );
  OAI22_X1 U20049 ( .A1(n17026), .A2(n16750), .B1(n16746), .B2(n16745), .ZN(
        n16747) );
  AOI211_X1 U20050 ( .C1(n17037), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16748), .B(n16747), .ZN(n16752) );
  OAI211_X1 U20051 ( .C1(n16755), .C2(n16750), .A(n17051), .B(n16749), .ZN(
        n16751) );
  OAI211_X1 U20052 ( .C1(n16753), .C2(n18931), .A(n16752), .B(n16751), .ZN(
        P3_U2646) );
  NOR2_X1 U20053 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17045), .ZN(n16754) );
  AOI22_X1 U20054 ( .A1(n17052), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16766), 
        .B2(n16754), .ZN(n16761) );
  AOI211_X1 U20055 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16771), .A(n16755), .B(
        n17044), .ZN(n16759) );
  AOI211_X1 U20056 ( .C1(n17714), .C2(n16757), .A(n16756), .B(n18863), .ZN(
        n16758) );
  AOI211_X1 U20057 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16762), .A(n16759), 
        .B(n16758), .ZN(n16760) );
  OAI211_X1 U20058 ( .C1(n17718), .C2(n17019), .A(n16761), .B(n16760), .ZN(
        P3_U2647) );
  INV_X1 U20059 ( .A(n16762), .ZN(n16774) );
  AOI211_X1 U20060 ( .C1(n16765), .C2(n16764), .A(n16763), .B(n18863), .ZN(
        n16770) );
  OR2_X1 U20061 ( .A1(n17045), .A2(n16766), .ZN(n16767) );
  OAI22_X1 U20062 ( .A1(n17026), .A2(n17061), .B1(n16768), .B2(n16767), .ZN(
        n16769) );
  AOI211_X1 U20063 ( .C1(n17037), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16770), .B(n16769), .ZN(n16773) );
  OAI211_X1 U20064 ( .C1(n16775), .C2(n17061), .A(n17051), .B(n16771), .ZN(
        n16772) );
  OAI211_X1 U20065 ( .C1(n16774), .C2(n18928), .A(n16773), .B(n16772), .ZN(
        P3_U2648) );
  AOI22_X1 U20066 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17037), .B1(
        n17052), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16782) );
  OAI221_X1 U20067 ( .B1(n17045), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17045), 
        .C2(n16800), .A(n17055), .ZN(n16788) );
  AOI211_X1 U20068 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16789), .A(n16775), .B(
        n17044), .ZN(n16779) );
  AOI211_X1 U20069 ( .C1(n17744), .C2(n16777), .A(n16776), .B(n18863), .ZN(
        n16778) );
  AOI211_X1 U20070 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16788), .A(n16779), 
        .B(n16778), .ZN(n16781) );
  INV_X1 U20071 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18925) );
  NAND4_X1 U20072 ( .A1(n17023), .A2(P3_REIP_REG_21__SCAN_IN), .A3(n16800), 
        .A4(n18925), .ZN(n16780) );
  NAND3_X1 U20073 ( .A1(n16782), .A2(n16781), .A3(n16780), .ZN(P3_U2649) );
  AOI22_X1 U20074 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17037), .B1(
        n17052), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16793) );
  AND2_X1 U20075 ( .A1(n17023), .A2(n16800), .ZN(n16787) );
  AOI211_X1 U20076 ( .C1(n16785), .C2(n16784), .A(n16783), .B(n18863), .ZN(
        n16786) );
  AOI221_X1 U20077 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16788), .C1(n16787), 
        .C2(n16788), .A(n16786), .ZN(n16792) );
  OAI211_X1 U20078 ( .C1(n16796), .C2(n16790), .A(n17051), .B(n16789), .ZN(
        n16791) );
  NAND3_X1 U20079 ( .A1(n16793), .A2(n16792), .A3(n16791), .ZN(P3_U2650) );
  AOI211_X1 U20080 ( .C1(n17768), .C2(n16795), .A(n16794), .B(n18863), .ZN(
        n16798) );
  AOI211_X1 U20081 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16814), .A(n16796), .B(
        n17044), .ZN(n16797) );
  AOI211_X1 U20082 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17052), .A(n16798), .B(
        n16797), .ZN(n16804) );
  NOR2_X1 U20083 ( .A1(n16799), .A2(n17045), .ZN(n16802) );
  OAI21_X1 U20084 ( .B1(n16800), .B2(n17045), .A(n17055), .ZN(n16801) );
  OAI21_X1 U20085 ( .B1(n16802), .B2(P3_REIP_REG_20__SCAN_IN), .A(n16801), 
        .ZN(n16803) );
  OAI211_X1 U20086 ( .C1(n17019), .C2(n10286), .A(n16804), .B(n16803), .ZN(
        P3_U2651) );
  NOR3_X1 U20087 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17045), .A3(n16805), 
        .ZN(n16819) );
  AND2_X1 U20088 ( .A1(n17023), .A2(n16805), .ZN(n16832) );
  NOR2_X1 U20089 ( .A1(n17043), .A2(n16832), .ZN(n16826) );
  INV_X1 U20090 ( .A(n16826), .ZN(n16837) );
  NOR2_X1 U20091 ( .A1(n16806), .A2(n16977), .ZN(n16822) );
  INV_X1 U20092 ( .A(n16820), .ZN(n16808) );
  OAI21_X1 U20093 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16808), .A(
        n16807), .ZN(n17780) );
  XOR2_X1 U20094 ( .A(n16822), .B(n17780), .Z(n16812) );
  NOR2_X1 U20095 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17045), .ZN(n16809) );
  AOI22_X1 U20096 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17037), .B1(
        n16810), .B2(n16809), .ZN(n16811) );
  OAI211_X1 U20097 ( .C1(n18863), .C2(n16812), .A(n16811), .B(n18339), .ZN(
        n16813) );
  AOI221_X1 U20098 ( .B1(n16819), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16837), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n16813), .ZN(n16816) );
  OAI211_X1 U20099 ( .C1(n16818), .C2(n16817), .A(n17051), .B(n16814), .ZN(
        n16815) );
  OAI211_X1 U20100 ( .C1(n16817), .C2(n17026), .A(n16816), .B(n16815), .ZN(
        P3_U2652) );
  AOI211_X1 U20101 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16838), .A(n16818), .B(
        n17044), .ZN(n16828) );
  INV_X1 U20102 ( .A(n16819), .ZN(n16825) );
  OAI21_X1 U20103 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17775), .A(
        n16820), .ZN(n17789) );
  INV_X1 U20104 ( .A(n17789), .ZN(n16823) );
  NOR2_X1 U20105 ( .A1(n17006), .A2(n18863), .ZN(n17040) );
  AOI221_X1 U20106 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16823), .C1(
        n16845), .C2(n16823), .A(n18863), .ZN(n16821) );
  OAI22_X1 U20107 ( .A1(n16823), .A2(n16822), .B1(n17040), .B2(n16821), .ZN(
        n16824) );
  OAI211_X1 U20108 ( .C1(n16826), .C2(n18917), .A(n16825), .B(n16824), .ZN(
        n16827) );
  AOI211_X1 U20109 ( .C1(n17037), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16828), .B(n16827), .ZN(n16829) );
  OAI211_X1 U20110 ( .C1(n17026), .C2(n17202), .A(n16829), .B(n18339), .ZN(
        P3_U2653) );
  AOI21_X1 U20111 ( .B1(n16830), .B2(n16843), .A(n17775), .ZN(n17807) );
  OAI21_X1 U20112 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16843), .A(
        n17006), .ZN(n16831) );
  XOR2_X1 U20113 ( .A(n17807), .B(n16831), .Z(n16835) );
  AOI22_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17037), .B1(
        n16833), .B2(n16832), .ZN(n16834) );
  OAI211_X1 U20115 ( .C1(n18863), .C2(n16835), .A(n16834), .B(n18339), .ZN(
        n16836) );
  AOI21_X1 U20116 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16837), .A(n16836), 
        .ZN(n16840) );
  OAI211_X1 U20117 ( .C1(n16844), .C2(n16841), .A(n17051), .B(n16838), .ZN(
        n16839) );
  OAI211_X1 U20118 ( .C1(n16841), .C2(n17026), .A(n16840), .B(n16839), .ZN(
        P3_U2654) );
  OR2_X1 U20119 ( .A1(n16854), .A2(n17043), .ZN(n16870) );
  OAI21_X1 U20120 ( .B1(n18911), .B2(n16870), .A(n17054), .ZN(n16855) );
  INV_X1 U20121 ( .A(n16842), .ZN(n17038) );
  AND2_X1 U20122 ( .A1(n16845), .A2(n17038), .ZN(n16865) );
  OAI21_X1 U20123 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16852), .A(
        n16843), .ZN(n17819) );
  AOI22_X1 U20124 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17037), .B1(
        n16865), .B2(n17819), .ZN(n16851) );
  AOI211_X1 U20125 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16858), .A(n16844), .B(
        n17044), .ZN(n16849) );
  AOI211_X1 U20126 ( .C1(n17006), .C2(n16845), .A(n18863), .B(n17819), .ZN(
        n16847) );
  NOR4_X1 U20127 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17045), .A3(n18911), 
        .A4(n16854), .ZN(n16846) );
  OR3_X1 U20128 ( .A1(n18357), .A2(n16847), .A3(n16846), .ZN(n16848) );
  AOI211_X1 U20129 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17052), .A(n16849), .B(
        n16848), .ZN(n16850) );
  OAI211_X1 U20130 ( .C1(n18913), .C2(n16855), .A(n16851), .B(n16850), .ZN(
        P3_U2655) );
  AOI21_X1 U20131 ( .B1(n16861), .B2(n16853), .A(n16852), .ZN(n17832) );
  INV_X1 U20132 ( .A(n17832), .ZN(n16864) );
  NOR2_X1 U20133 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18863), .ZN(
        n17039) );
  INV_X1 U20134 ( .A(n17039), .ZN(n16964) );
  INV_X1 U20135 ( .A(n17040), .ZN(n17036) );
  OAI21_X1 U20136 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n16964), .A(
        n17036), .ZN(n16863) );
  NOR2_X1 U20137 ( .A1(n17045), .A2(n16854), .ZN(n16857) );
  INV_X1 U20138 ( .A(n16855), .ZN(n16856) );
  OAI21_X1 U20139 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16857), .A(n16856), 
        .ZN(n16860) );
  OAI211_X1 U20140 ( .C1(n16868), .C2(n17236), .A(n17051), .B(n16858), .ZN(
        n16859) );
  OAI211_X1 U20141 ( .C1(n17019), .C2(n16861), .A(n16860), .B(n16859), .ZN(
        n16862) );
  AOI221_X1 U20142 ( .B1(n16865), .B2(n16864), .C1(n16863), .C2(n17832), .A(
        n16862), .ZN(n16866) );
  OAI211_X1 U20143 ( .C1(n17026), .C2(n17236), .A(n16866), .B(n18339), .ZN(
        P3_U2656) );
  INV_X1 U20144 ( .A(n16867), .ZN(n17841) );
  INV_X1 U20145 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17968) );
  NAND2_X1 U20146 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9967), .ZN(
        n16976) );
  NOR2_X1 U20147 ( .A1(n17968), .A2(n16976), .ZN(n16963) );
  NAND2_X1 U20148 ( .A1(n17841), .A2(n16963), .ZN(n16921) );
  NOR2_X1 U20149 ( .A1(n17883), .A2(n16921), .ZN(n17853) );
  INV_X1 U20150 ( .A(n17853), .ZN(n16895) );
  NOR2_X1 U20151 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16895), .ZN(
        n16896) );
  AOI21_X1 U20152 ( .B1(n17852), .B2(n16896), .A(n16977), .ZN(n16879) );
  INV_X1 U20153 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16873) );
  NAND2_X1 U20154 ( .A1(n17852), .A2(n17853), .ZN(n16878) );
  AOI21_X1 U20155 ( .B1(n16873), .B2(n16878), .A(n17816), .ZN(n17842) );
  XNOR2_X1 U20156 ( .A(n16879), .B(n17842), .ZN(n16877) );
  AOI211_X1 U20157 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16881), .A(n16868), .B(
        n17044), .ZN(n16875) );
  INV_X1 U20158 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18907) );
  NAND2_X1 U20159 ( .A1(n17023), .A2(n16869), .ZN(n16884) );
  NOR2_X1 U20160 ( .A1(n18907), .A2(n16884), .ZN(n16871) );
  OAI211_X1 U20161 ( .C1(n16871), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17054), 
        .B(n16870), .ZN(n16872) );
  OAI211_X1 U20162 ( .C1(n16873), .C2(n17019), .A(n16872), .B(n18339), .ZN(
        n16874) );
  AOI211_X1 U20163 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17052), .A(n16875), .B(
        n16874), .ZN(n16876) );
  OAI21_X1 U20164 ( .B1(n18863), .B2(n16877), .A(n16876), .ZN(P3_U2657) );
  NOR2_X1 U20165 ( .A1(n17868), .A2(n16895), .ZN(n16894) );
  OAI21_X1 U20166 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16894), .A(
        n16878), .ZN(n17856) );
  AOI21_X1 U20167 ( .B1(n16894), .B2(n17039), .A(n17040), .ZN(n16889) );
  NAND3_X1 U20168 ( .A1(n17014), .A2(n16879), .A3(n17856), .ZN(n16880) );
  OAI211_X1 U20169 ( .C1(n17858), .C2(n17019), .A(n18339), .B(n16880), .ZN(
        n16886) );
  OAI211_X1 U20170 ( .C1(n16890), .C2(n16882), .A(n17051), .B(n16881), .ZN(
        n16883) );
  OAI21_X1 U20171 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16884), .A(n16883), 
        .ZN(n16885) );
  AOI211_X1 U20172 ( .C1(n17052), .C2(P3_EBX_REG_13__SCAN_IN), .A(n16886), .B(
        n16885), .ZN(n16888) );
  NOR2_X1 U20173 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17045), .ZN(n16892) );
  OAI21_X1 U20174 ( .B1(n16893), .B2(n17045), .A(n17055), .ZN(n16902) );
  OAI21_X1 U20175 ( .B1(n16892), .B2(n16902), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16887) );
  OAI211_X1 U20176 ( .C1(n17856), .C2(n16889), .A(n16888), .B(n16887), .ZN(
        P3_U2658) );
  AOI211_X1 U20177 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16909), .A(n16890), .B(
        n17044), .ZN(n16891) );
  AOI21_X1 U20178 ( .B1(n17037), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16891), .ZN(n16901) );
  AOI22_X1 U20179 ( .A1(n17052), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16893), 
        .B2(n16892), .ZN(n16900) );
  AOI21_X1 U20180 ( .B1(n17868), .B2(n16895), .A(n16894), .ZN(n17871) );
  NOR2_X1 U20181 ( .A1(n16896), .A2(n16977), .ZN(n16897) );
  XOR2_X1 U20182 ( .A(n17871), .B(n16897), .Z(n16898) );
  AOI22_X1 U20183 ( .A1(n17014), .A2(n16898), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16902), .ZN(n16899) );
  NAND4_X1 U20184 ( .A1(n16901), .A2(n16900), .A3(n16899), .A4(n18339), .ZN(
        P3_U2659) );
  INV_X1 U20185 ( .A(n16902), .ZN(n16907) );
  NOR2_X1 U20186 ( .A1(n18901), .A2(n18899), .ZN(n16916) );
  NOR2_X1 U20187 ( .A1(n17045), .A2(n16913), .ZN(n16928) );
  AOI21_X1 U20188 ( .B1(n16916), .B2(n16928), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16906) );
  AOI21_X1 U20189 ( .B1(n17883), .B2(n16921), .A(n17853), .ZN(n17886) );
  INV_X1 U20190 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16933) );
  INV_X1 U20191 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17894) );
  NOR2_X1 U20192 ( .A1(n16933), .A2(n17894), .ZN(n16903) );
  INV_X1 U20193 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17924) );
  INV_X1 U20194 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17941) );
  OR2_X1 U20195 ( .A1(n17922), .A2(n17941), .ZN(n17921) );
  NAND2_X1 U20196 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16978), .ZN(
        n17030) );
  NOR3_X1 U20197 ( .A1(n17924), .A2(n17921), .A3(n17030), .ZN(n16930) );
  AOI21_X1 U20198 ( .B1(n16903), .B2(n16930), .A(n16977), .ZN(n16904) );
  XNOR2_X1 U20199 ( .A(n17886), .B(n16904), .ZN(n16905) );
  OAI22_X1 U20200 ( .A1(n16907), .A2(n16906), .B1(n18863), .B2(n16905), .ZN(
        n16908) );
  AOI211_X1 U20201 ( .C1(n17052), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18357), .B(
        n16908), .ZN(n16912) );
  OAI211_X1 U20202 ( .C1(n16914), .C2(n16910), .A(n17051), .B(n16909), .ZN(
        n16911) );
  OAI211_X1 U20203 ( .C1(n17019), .C2(n17883), .A(n16912), .B(n16911), .ZN(
        P3_U2660) );
  AOI21_X1 U20204 ( .B1(n16913), .B2(n17023), .A(n17043), .ZN(n16945) );
  AOI211_X1 U20205 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16915), .A(n16914), .B(
        n17044), .ZN(n16920) );
  INV_X1 U20206 ( .A(n16916), .ZN(n16917) );
  OAI211_X1 U20207 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16928), .B(n16917), .ZN(n16918) );
  OAI211_X1 U20208 ( .C1(n17894), .C2(n17019), .A(n18339), .B(n16918), .ZN(
        n16919) );
  AOI211_X1 U20209 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17052), .A(n16920), .B(
        n16919), .ZN(n16926) );
  NOR2_X1 U20210 ( .A1(n18024), .A2(n17921), .ZN(n16952) );
  NAND2_X1 U20211 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16952), .ZN(
        n16941) );
  NOR2_X1 U20212 ( .A1(n16933), .A2(n16941), .ZN(n16922) );
  OAI21_X1 U20213 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16922), .A(
        n16921), .ZN(n17908) );
  INV_X1 U20214 ( .A(n17908), .ZN(n16924) );
  AOI21_X1 U20215 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16930), .A(
        n16977), .ZN(n16931) );
  INV_X1 U20216 ( .A(n16931), .ZN(n16923) );
  OAI221_X1 U20217 ( .B1(n16924), .B2(n16931), .C1(n17908), .C2(n16923), .A(
        n17014), .ZN(n16925) );
  OAI211_X1 U20218 ( .C1(n16945), .C2(n18901), .A(n16926), .B(n16925), .ZN(
        P3_U2661) );
  AOI21_X1 U20219 ( .B1(n17051), .B2(n16927), .A(n17052), .ZN(n16939) );
  NOR2_X1 U20220 ( .A1(n16927), .A2(n17044), .ZN(n16944) );
  AOI22_X1 U20221 ( .A1(n16928), .A2(n18899), .B1(n16944), .B2(n16940), .ZN(
        n16938) );
  INV_X1 U20222 ( .A(n16945), .ZN(n16936) );
  INV_X1 U20223 ( .A(n16941), .ZN(n16929) );
  AOI22_X1 U20224 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16941), .B1(
        n16929), .B2(n16933), .ZN(n17916) );
  AOI22_X1 U20225 ( .A1(n16931), .A2(n17916), .B1(n16930), .B2(n16933), .ZN(
        n16932) );
  OAI21_X1 U20226 ( .B1(n16932), .B2(n18863), .A(n18339), .ZN(n16935) );
  OAI22_X1 U20227 ( .A1(n16933), .A2(n17019), .B1(n17916), .B2(n17036), .ZN(
        n16934) );
  AOI211_X1 U20228 ( .C1(n16936), .C2(P3_REIP_REG_9__SCAN_IN), .A(n16935), .B(
        n16934), .ZN(n16937) );
  OAI211_X1 U20229 ( .C1(n16940), .C2(n16939), .A(n16938), .B(n16937), .ZN(
        P3_U2662) );
  OAI21_X1 U20230 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16952), .A(
        n16941), .ZN(n17925) );
  OAI21_X1 U20231 ( .B1(n17921), .B2(n17030), .A(n17006), .ZN(n16942) );
  XNOR2_X1 U20232 ( .A(n17925), .B(n16942), .ZN(n16950) );
  NAND2_X1 U20233 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16959), .ZN(n16943) );
  AOI22_X1 U20234 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17037), .B1(
        n16944), .B2(n16943), .ZN(n16949) );
  AOI221_X1 U20235 ( .B1(n17045), .B2(n18898), .C1(n16946), .C2(n18898), .A(
        n16945), .ZN(n16947) );
  AOI211_X1 U20236 ( .C1(n17052), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18357), .B(
        n16947), .ZN(n16948) );
  OAI211_X1 U20237 ( .C1(n18863), .C2(n16950), .A(n16949), .B(n16948), .ZN(
        P3_U2663) );
  OAI21_X1 U20238 ( .B1(n16951), .B2(n17045), .A(n17055), .ZN(n16970) );
  INV_X1 U20239 ( .A(n16952), .ZN(n16953) );
  OAI21_X1 U20240 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16963), .A(
        n16953), .ZN(n17952) );
  OAI21_X1 U20241 ( .B1(n17922), .B2(n17030), .A(n17006), .ZN(n16955) );
  OAI21_X1 U20242 ( .B1(n17952), .B2(n16955), .A(n17014), .ZN(n16954) );
  AOI21_X1 U20243 ( .B1(n17952), .B2(n16955), .A(n16954), .ZN(n16958) );
  NOR2_X1 U20244 ( .A1(n17045), .A2(n16985), .ZN(n16971) );
  INV_X1 U20245 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18895) );
  NAND3_X1 U20246 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16971), .A3(n18895), 
        .ZN(n16956) );
  OAI211_X1 U20247 ( .C1(n17026), .C2(n16960), .A(n18339), .B(n16956), .ZN(
        n16957) );
  AOI211_X1 U20248 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16970), .A(n16958), .B(
        n16957), .ZN(n16962) );
  OAI211_X1 U20249 ( .C1(n16965), .C2(n16960), .A(n17051), .B(n16959), .ZN(
        n16961) );
  OAI211_X1 U20250 ( .C1(n17019), .C2(n17941), .A(n16962), .B(n16961), .ZN(
        P3_U2664) );
  AOI21_X1 U20251 ( .B1(n17968), .B2(n16976), .A(n16963), .ZN(n17965) );
  OAI21_X1 U20252 ( .B1(n16976), .B2(n16964), .A(n17036), .ZN(n16969) );
  AOI211_X1 U20253 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16981), .A(n16965), .B(
        n17044), .ZN(n16968) );
  INV_X1 U20254 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16966) );
  OAI22_X1 U20255 ( .A1(n17968), .A2(n17019), .B1(n17026), .B2(n16966), .ZN(
        n16967) );
  AOI211_X1 U20256 ( .C1(n17965), .C2(n16969), .A(n16968), .B(n16967), .ZN(
        n16975) );
  OAI21_X1 U20257 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16971), .A(n16970), .ZN(
        n16974) );
  INV_X1 U20258 ( .A(n17965), .ZN(n16972) );
  OAI211_X1 U20259 ( .C1(n17922), .C2(n17030), .A(n17038), .B(n16972), .ZN(
        n16973) );
  NAND4_X1 U20260 ( .A1(n16975), .A2(n18339), .A3(n16974), .A4(n16973), .ZN(
        P3_U2665) );
  NOR2_X1 U20261 ( .A1(n18024), .A2(n17976), .ZN(n16992) );
  OAI21_X1 U20262 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16992), .A(
        n16976), .ZN(n16979) );
  INV_X1 U20263 ( .A(n16979), .ZN(n17979) );
  AOI21_X1 U20264 ( .B1(n16978), .B2(n16992), .A(n16977), .ZN(n16980) );
  INV_X1 U20265 ( .A(n16980), .ZN(n16995) );
  OAI221_X1 U20266 ( .B1(n17979), .B2(n16980), .C1(n16979), .C2(n16995), .A(
        n17014), .ZN(n16983) );
  OAI211_X1 U20267 ( .C1(n16991), .C2(n16989), .A(n17051), .B(n16981), .ZN(
        n16982) );
  OAI211_X1 U20268 ( .C1(n17019), .C2(n17977), .A(n16983), .B(n16982), .ZN(
        n16984) );
  AOI211_X1 U20269 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n17043), .A(n18357), .B(
        n16984), .ZN(n16988) );
  OAI211_X1 U20270 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n16986), .A(n17023), .B(
        n16985), .ZN(n16987) );
  OAI211_X1 U20271 ( .C1(n16989), .C2(n17026), .A(n16988), .B(n16987), .ZN(
        P3_U2666) );
  AOI21_X1 U20272 ( .B1(n17023), .B2(n16990), .A(n17043), .ZN(n17009) );
  AOI211_X1 U20273 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17015), .A(n16991), .B(
        n17044), .ZN(n16994) );
  NAND2_X1 U20274 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17990), .ZN(
        n17004) );
  AOI21_X1 U20275 ( .B1(n10290), .B2(n17004), .A(n16992), .ZN(n16996) );
  INV_X1 U20276 ( .A(n16996), .ZN(n17993) );
  OAI22_X1 U20277 ( .A1(n10290), .A2(n17019), .B1(n17993), .B2(n17036), .ZN(
        n16993) );
  AOI211_X1 U20278 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17052), .A(n16994), .B(
        n16993), .ZN(n17003) );
  NAND2_X1 U20279 ( .A1(n17990), .A2(n10290), .ZN(n17985) );
  OAI22_X1 U20280 ( .A1(n16996), .A2(n16995), .B1(n17030), .B2(n17985), .ZN(
        n17001) );
  NAND2_X1 U20281 ( .A1(n16997), .A2(n19009), .ZN(n19026) );
  NAND2_X1 U20282 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17022) );
  NOR2_X1 U20283 ( .A1(n17045), .A2(n17022), .ZN(n17008) );
  NAND3_X1 U20284 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17008), .A3(n18889), 
        .ZN(n16998) );
  OAI221_X1 U20285 ( .B1(n19026), .B2(n17144), .C1(n19026), .C2(n16999), .A(
        n16998), .ZN(n17000) );
  AOI211_X1 U20286 ( .C1(n17014), .C2(n17001), .A(n18357), .B(n17000), .ZN(
        n17002) );
  OAI211_X1 U20287 ( .C1(n18889), .C2(n17009), .A(n17003), .B(n17002), .ZN(
        P3_U2667) );
  NAND2_X1 U20288 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17031) );
  INV_X1 U20289 ( .A(n17004), .ZN(n17005) );
  AOI21_X1 U20290 ( .B1(n17018), .B2(n17031), .A(n17005), .ZN(n17997) );
  OAI21_X1 U20291 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17031), .A(
        n17006), .ZN(n17007) );
  XNOR2_X1 U20292 ( .A(n17997), .B(n17007), .ZN(n17013) );
  INV_X1 U20293 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18887) );
  INV_X1 U20294 ( .A(n17008), .ZN(n17010) );
  AOI21_X1 U20295 ( .B1(n18887), .B2(n17010), .A(n17009), .ZN(n17012) );
  NOR2_X1 U20296 ( .A1(n18988), .A2(n18828), .ZN(n18812) );
  OAI21_X1 U20297 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18812), .A(
        n17144), .ZN(n18962) );
  OAI22_X1 U20298 ( .A1(n17026), .A2(n17377), .B1(n19026), .B2(n18962), .ZN(
        n17011) );
  AOI211_X1 U20299 ( .C1(n17014), .C2(n17013), .A(n17012), .B(n17011), .ZN(
        n17017) );
  OAI211_X1 U20300 ( .C1(n17020), .C2(n17377), .A(n17051), .B(n17015), .ZN(
        n17016) );
  OAI211_X1 U20301 ( .C1(n17019), .C2(n17018), .A(n17017), .B(n17016), .ZN(
        P3_U2668) );
  OAI21_X1 U20302 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17031), .ZN(n18015) );
  INV_X1 U20303 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17398) );
  INV_X1 U20304 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17392) );
  NAND2_X1 U20305 ( .A1(n17398), .A2(n17392), .ZN(n17021) );
  AOI211_X1 U20306 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17021), .A(n17020), .B(
        n17044), .ZN(n17029) );
  NAND2_X1 U20307 ( .A1(n13851), .A2(n18974), .ZN(n18810) );
  INV_X1 U20308 ( .A(n18810), .ZN(n18814) );
  NOR2_X1 U20309 ( .A1(n18812), .A2(n18814), .ZN(n18971) );
  INV_X1 U20310 ( .A(n19026), .ZN(n17053) );
  AOI22_X1 U20311 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n17043), .B1(n18971), 
        .B2(n17053), .ZN(n17025) );
  OAI211_X1 U20312 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17023), .B(n17022), .ZN(n17024) );
  OAI211_X1 U20313 ( .C1(n17027), .C2(n17026), .A(n17025), .B(n17024), .ZN(
        n17028) );
  AOI211_X1 U20314 ( .C1(n17037), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17029), .B(n17028), .ZN(n17035) );
  INV_X1 U20315 ( .A(n17030), .ZN(n17033) );
  OR2_X1 U20316 ( .A1(n17031), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17032) );
  OAI211_X1 U20317 ( .C1(n17033), .C2(n18015), .A(n17038), .B(n17032), .ZN(
        n17034) );
  OAI211_X1 U20318 ( .C1(n17036), .C2(n18015), .A(n17035), .B(n17034), .ZN(
        P3_U2669) );
  AOI211_X1 U20319 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17038), .A(
        n17037), .B(n18024), .ZN(n17050) );
  NOR3_X1 U20320 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17040), .A3(
        n17039), .ZN(n17049) );
  NOR2_X1 U20321 ( .A1(n17042), .A2(n17041), .ZN(n18979) );
  AOI22_X1 U20322 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17043), .B1(n18979), 
        .B2(n17053), .ZN(n17048) );
  OAI21_X1 U20323 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17385), .ZN(n17394) );
  OAI22_X1 U20324 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17045), .B1(n17044), 
        .B2(n17394), .ZN(n17046) );
  AOI21_X1 U20325 ( .B1(n17052), .B2(P3_EBX_REG_1__SCAN_IN), .A(n17046), .ZN(
        n17047) );
  OAI211_X1 U20326 ( .C1(n17050), .C2(n17049), .A(n17048), .B(n17047), .ZN(
        P3_U2670) );
  NOR2_X1 U20327 ( .A1(n17052), .A2(n17051), .ZN(n17058) );
  AOI22_X1 U20328 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17054), .B1(n17053), 
        .B2(n18988), .ZN(n17057) );
  NAND3_X1 U20329 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19022), .A3(
        n17055), .ZN(n17056) );
  OAI211_X1 U20330 ( .C1(n17058), .C2(n17398), .A(n17057), .B(n17056), .ZN(
        P3_U2671) );
  INV_X1 U20331 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17059) );
  NOR2_X1 U20332 ( .A1(n17059), .A2(n17186), .ZN(n17142) );
  NAND4_X1 U20333 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n17060), .ZN(n17097) );
  NOR3_X1 U20334 ( .A1(n17062), .A2(n17061), .A3(n17097), .ZN(n17063) );
  NAND4_X1 U20335 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17142), .A4(n17063), .ZN(n17066) );
  NOR2_X1 U20336 ( .A1(n17067), .A2(n17066), .ZN(n17093) );
  NAND2_X1 U20337 ( .A1(n17390), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17065) );
  NAND2_X1 U20338 ( .A1(n17093), .A2(n17445), .ZN(n17064) );
  OAI22_X1 U20339 ( .A1(n17093), .A2(n17065), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17064), .ZN(P3_U2672) );
  NAND2_X1 U20340 ( .A1(n17067), .A2(n17066), .ZN(n17068) );
  NAND2_X1 U20341 ( .A1(n17068), .A2(n17390), .ZN(n17092) );
  AOI22_X1 U20342 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20343 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20344 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17077) );
  OAI22_X1 U20345 ( .A1(n17222), .A2(n17259), .B1(n17349), .B2(n17069), .ZN(
        n17075) );
  AOI22_X1 U20346 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20347 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20348 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17071) );
  NAND2_X1 U20349 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n17070) );
  NAND4_X1 U20350 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  AOI211_X1 U20351 ( .C1(n17328), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17075), .B(n17074), .ZN(n17076) );
  NAND4_X1 U20352 ( .A1(n17079), .A2(n17078), .A3(n17077), .A4(n17076), .ZN(
        n17095) );
  NAND2_X1 U20353 ( .A1(n17096), .A2(n17095), .ZN(n17094) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17242), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17089) );
  INV_X1 U20355 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20356 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15633), .ZN(n17081) );
  AOI22_X1 U20357 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17223), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17080) );
  OAI211_X1 U20358 ( .C1(n17349), .C2(n17248), .A(n17081), .B(n17080), .ZN(
        n17087) );
  AOI22_X1 U20359 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9810), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17323), .ZN(n17085) );
  AOI22_X1 U20360 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20361 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17083) );
  NAND2_X1 U20362 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17176), .ZN(
        n17082) );
  NAND4_X1 U20363 ( .A1(n17085), .A2(n17084), .A3(n17083), .A4(n17082), .ZN(
        n17086) );
  AOI211_X1 U20364 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17087), .B(n17086), .ZN(n17088) );
  OAI211_X1 U20365 ( .C1(n17090), .C2(n17293), .A(n17089), .B(n17088), .ZN(
        n17091) );
  XOR2_X1 U20366 ( .A(n17094), .B(n17091), .Z(n17406) );
  OAI22_X1 U20367 ( .A1(n17093), .A2(n17092), .B1(n17406), .B2(n17390), .ZN(
        P3_U2673) );
  OAI21_X1 U20368 ( .B1(n17096), .B2(n17095), .A(n17094), .ZN(n17414) );
  NOR2_X1 U20369 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17097), .ZN(n17098) );
  AOI22_X1 U20370 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17099), .B1(n17125), 
        .B2(n17098), .ZN(n17100) );
  OAI21_X1 U20371 ( .B1(n17414), .B2(n17390), .A(n17100), .ZN(P3_U2674) );
  OAI21_X1 U20372 ( .B1(n17105), .B2(n17102), .A(n17101), .ZN(n17423) );
  NAND3_X1 U20373 ( .A1(n17104), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17390), 
        .ZN(n17103) );
  OAI221_X1 U20374 ( .B1(n17104), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17390), 
        .C2(n17423), .A(n17103), .ZN(P3_U2676) );
  AOI21_X1 U20375 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17390), .A(n17114), .ZN(
        n17108) );
  AOI21_X1 U20376 ( .B1(n17106), .B2(n17111), .A(n17105), .ZN(n17424) );
  INV_X1 U20377 ( .A(n17424), .ZN(n17107) );
  OAI22_X1 U20378 ( .A1(n17109), .A2(n17108), .B1(n17107), .B2(n17390), .ZN(
        P3_U2677) );
  INV_X1 U20379 ( .A(n17110), .ZN(n17119) );
  AOI21_X1 U20380 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17390), .A(n17119), .ZN(
        n17113) );
  OAI21_X1 U20381 ( .B1(n17115), .B2(n17112), .A(n17111), .ZN(n17431) );
  OAI22_X1 U20382 ( .A1(n17114), .A2(n17113), .B1(n17390), .B2(n17431), .ZN(
        P3_U2678) );
  AOI21_X1 U20383 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17390), .A(n17125), .ZN(
        n17118) );
  AOI21_X1 U20384 ( .B1(n17116), .B2(n17121), .A(n17115), .ZN(n17432) );
  INV_X1 U20385 ( .A(n17432), .ZN(n17117) );
  OAI22_X1 U20386 ( .A1(n17119), .A2(n17118), .B1(n17390), .B2(n17117), .ZN(
        P3_U2679) );
  INV_X1 U20387 ( .A(n17120), .ZN(n17141) );
  AOI21_X1 U20388 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17390), .A(n17141), .ZN(
        n17124) );
  OAI21_X1 U20389 ( .B1(n17123), .B2(n17122), .A(n17121), .ZN(n17443) );
  OAI22_X1 U20390 ( .A1(n17125), .A2(n17124), .B1(n17390), .B2(n17443), .ZN(
        P3_U2680) );
  AOI21_X1 U20391 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17390), .A(n17126), .ZN(
        n17140) );
  AOI22_X1 U20392 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20393 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17127) );
  OAI21_X1 U20394 ( .B1(n17275), .B2(n17128), .A(n17127), .ZN(n17136) );
  AOI22_X1 U20395 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17134) );
  INV_X1 U20396 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20397 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20398 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17129) );
  OAI211_X1 U20399 ( .C1(n13966), .C2(n17131), .A(n17130), .B(n17129), .ZN(
        n17132) );
  AOI21_X1 U20400 ( .B1(n17335), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17132), .ZN(n17133) );
  OAI211_X1 U20401 ( .C1(n17293), .C2(n17370), .A(n17134), .B(n17133), .ZN(
        n17135) );
  AOI211_X1 U20402 ( .C1(n17328), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17136), .B(n17135), .ZN(n17137) );
  OAI211_X1 U20403 ( .C1(n13868), .C2(n17268), .A(n17138), .B(n17137), .ZN(
        n17446) );
  INV_X1 U20404 ( .A(n17446), .ZN(n17139) );
  OAI22_X1 U20405 ( .A1(n17141), .A2(n17140), .B1(n17139), .B2(n17390), .ZN(
        P3_U2681) );
  NOR2_X1 U20406 ( .A1(n17396), .A2(n17142), .ZN(n17170) );
  AOI22_X1 U20407 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20408 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17155) );
  OAI22_X1 U20409 ( .A1(n17222), .A2(n17145), .B1(n17144), .B2(n17143), .ZN(
        n17153) );
  AOI22_X1 U20410 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20411 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20412 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17146) );
  OAI211_X1 U20413 ( .C1(n13901), .C2(n17148), .A(n17147), .B(n17146), .ZN(
        n17149) );
  AOI21_X1 U20414 ( .B1(n17335), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17149), .ZN(n17150) );
  OAI211_X1 U20415 ( .C1(n17293), .C2(n17373), .A(n17151), .B(n17150), .ZN(
        n17152) );
  AOI211_X1 U20416 ( .C1(n17176), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17153), .B(n17152), .ZN(n17154) );
  NAND3_X1 U20417 ( .A1(n17156), .A2(n17155), .A3(n17154), .ZN(n17451) );
  AOI22_X1 U20418 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17170), .B1(n17396), 
        .B2(n17451), .ZN(n17157) );
  OAI21_X1 U20419 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17158), .A(n17157), .ZN(
        P3_U2682) );
  AOI22_X1 U20420 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20421 ( .B1(n17302), .B2(n17274), .A(n17159), .ZN(n17169) );
  INV_X1 U20422 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20423 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17166) );
  OAI22_X1 U20424 ( .A1(n13934), .A2(n17277), .B1(n17293), .B2(n17381), .ZN(
        n17164) );
  AOI22_X1 U20425 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20426 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20427 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17160) );
  NAND3_X1 U20428 ( .A1(n17162), .A2(n17161), .A3(n17160), .ZN(n17163) );
  AOI211_X1 U20429 ( .C1(n17335), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17164), .B(n17163), .ZN(n17165) );
  OAI211_X1 U20430 ( .C1(n17339), .C2(n17167), .A(n17166), .B(n17165), .ZN(
        n17168) );
  AOI211_X1 U20431 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n17169), .B(n17168), .ZN(n17456) );
  OAI21_X1 U20432 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17171), .A(n17170), .ZN(
        n17172) );
  OAI21_X1 U20433 ( .B1(n17456), .B2(n17390), .A(n17172), .ZN(P3_U2683) );
  AOI22_X1 U20434 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20435 ( .B1(n17275), .B2(n17174), .A(n17173), .ZN(n17185) );
  INV_X1 U20436 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20437 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17241), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17183) );
  OAI22_X1 U20438 ( .A1(n9813), .A2(n17175), .B1(n17293), .B2(n17383), .ZN(
        n17181) );
  AOI22_X1 U20439 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17351), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20440 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20441 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17177) );
  NAND3_X1 U20442 ( .A1(n17179), .A2(n17178), .A3(n17177), .ZN(n17180) );
  AOI211_X1 U20443 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17181), .B(n17180), .ZN(n17182) );
  OAI211_X1 U20444 ( .C1(n17222), .C2(n17301), .A(n17183), .B(n17182), .ZN(
        n17184) );
  AOI211_X1 U20445 ( .C1(n17242), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17185), .B(n17184), .ZN(n17463) );
  OAI21_X1 U20446 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17187), .A(n17186), .ZN(
        n17188) );
  AOI22_X1 U20447 ( .A1(n17396), .A2(n17463), .B1(n17188), .B2(n17390), .ZN(
        P3_U2684) );
  NAND2_X1 U20448 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17189), .ZN(n17204) );
  AOI22_X1 U20449 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17190) );
  OAI21_X1 U20450 ( .B1(n13922), .B2(n17191), .A(n17190), .ZN(n17200) );
  AOI22_X1 U20451 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17198) );
  INV_X1 U20452 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18419) );
  AOI22_X1 U20453 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17192) );
  OAI21_X1 U20454 ( .B1(n13966), .B2(n18419), .A(n17192), .ZN(n17196) );
  AOI22_X1 U20455 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20456 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17193) );
  OAI211_X1 U20457 ( .C1(n17349), .C2(n17317), .A(n17194), .B(n17193), .ZN(
        n17195) );
  AOI211_X1 U20458 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17196), .B(n17195), .ZN(n17197) );
  OAI211_X1 U20459 ( .C1(n17293), .C2(n17389), .A(n17198), .B(n17197), .ZN(
        n17199) );
  AOI211_X1 U20460 ( .C1(n13852), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17200), .B(n17199), .ZN(n17468) );
  NAND2_X1 U20461 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17288), .ZN(n17272) );
  NOR2_X1 U20462 ( .A1(n17201), .A2(n17272), .ZN(n17219) );
  NAND3_X1 U20463 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17219), .A3(n17202), 
        .ZN(n17203) );
  OAI221_X1 U20464 ( .B1(n17396), .B2(n17204), .C1(n17390), .C2(n17468), .A(
        n17203), .ZN(P3_U2685) );
  AOI22_X1 U20465 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U20466 ( .B1(n13933), .B2(n17206), .A(n17205), .ZN(n17216) );
  AOI22_X1 U20467 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20468 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17207) );
  OAI21_X1 U20469 ( .B1(n13966), .B2(n18415), .A(n17207), .ZN(n17212) );
  AOI22_X1 U20470 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20471 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17208) );
  OAI211_X1 U20472 ( .C1(n13901), .C2(n17210), .A(n17209), .B(n17208), .ZN(
        n17211) );
  AOI211_X1 U20473 ( .C1(n17335), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17212), .B(n17211), .ZN(n17213) );
  OAI211_X1 U20474 ( .C1(n17339), .C2(n17332), .A(n17214), .B(n17213), .ZN(
        n17215) );
  AOI211_X1 U20475 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17216), .B(n17215), .ZN(n17472) );
  OAI211_X1 U20476 ( .C1(n17217), .C2(n18400), .A(P3_EBX_REG_17__SCAN_IN), .B(
        n17399), .ZN(n17218) );
  OAI21_X1 U20477 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17219), .A(n17218), .ZN(
        n17220) );
  OAI21_X1 U20478 ( .B1(n17472), .B2(n17390), .A(n17220), .ZN(P3_U2686) );
  OAI22_X1 U20479 ( .A1(n9813), .A2(n18689), .B1(n17222), .B2(n17221), .ZN(
        n17233) );
  AOI22_X1 U20480 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20481 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20482 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17224) );
  OAI21_X1 U20483 ( .B1(n17293), .B2(n17361), .A(n17224), .ZN(n17228) );
  AOI22_X1 U20484 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20485 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17225) );
  OAI211_X1 U20486 ( .C1(n13966), .C2(n18412), .A(n17226), .B(n17225), .ZN(
        n17227) );
  AOI211_X1 U20487 ( .C1(n17335), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17228), .B(n17227), .ZN(n17229) );
  NAND3_X1 U20488 ( .A1(n17231), .A2(n17230), .A3(n17229), .ZN(n17232) );
  AOI211_X1 U20489 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17233), .B(n17232), .ZN(n17478) );
  INV_X1 U20490 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17235) );
  NOR3_X1 U20491 ( .A1(n17235), .A2(n17384), .A3(n17234), .ZN(n17255) );
  AOI21_X1 U20492 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17255), .A(n17396), .ZN(
        n17254) );
  NOR4_X1 U20493 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17236), .A3(n17235), .A4(
        n17272), .ZN(n17237) );
  AOI21_X1 U20494 ( .B1(n17254), .B2(P3_EBX_REG_16__SCAN_IN), .A(n17237), .ZN(
        n17238) );
  OAI21_X1 U20495 ( .B1(n17478), .B2(n17390), .A(n17238), .ZN(P3_U2687) );
  AOI22_X1 U20496 ( .A1(n13852), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20497 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17350), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17324), .ZN(n17239) );
  OAI21_X1 U20498 ( .B1(n17240), .B2(n13933), .A(n17239), .ZN(n17250) );
  AOI22_X1 U20499 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17326), .B1(
        n17241), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20500 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17242), .ZN(n17244) );
  AOI22_X1 U20501 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n15633), .ZN(n17243) );
  OAI211_X1 U20502 ( .C1(n17367), .C2(n13966), .A(n17244), .B(n17243), .ZN(
        n17245) );
  AOI21_X1 U20503 ( .B1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17335), .A(
        n17245), .ZN(n17246) );
  OAI211_X1 U20504 ( .C1(n13934), .C2(n17248), .A(n17247), .B(n17246), .ZN(
        n17249) );
  AOI211_X1 U20505 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17250), .B(n17249), .ZN(n17251) );
  OAI211_X1 U20506 ( .C1(n17253), .C2(n17275), .A(n17252), .B(n17251), .ZN(
        n17479) );
  INV_X1 U20507 ( .A(n17479), .ZN(n17257) );
  OAI21_X1 U20508 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17255), .A(n17254), .ZN(
        n17256) );
  OAI21_X1 U20509 ( .B1(n17257), .B2(n17390), .A(n17256), .ZN(P3_U2688) );
  AOI22_X1 U20510 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17258) );
  OAI21_X1 U20511 ( .B1(n17275), .B2(n17259), .A(n17258), .ZN(n17270) );
  AOI22_X1 U20512 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20513 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U20514 ( .B1(n17293), .B2(n17261), .A(n17260), .ZN(n17265) );
  AOI22_X1 U20515 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20516 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17262) );
  OAI211_X1 U20517 ( .C1(n13966), .C2(n17370), .A(n17263), .B(n17262), .ZN(
        n17264) );
  AOI211_X1 U20518 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17265), .B(n17264), .ZN(n17266) );
  OAI211_X1 U20519 ( .C1(n13879), .C2(n17268), .A(n17267), .B(n17266), .ZN(
        n17269) );
  AOI211_X1 U20520 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17270), .B(n17269), .ZN(n17490) );
  NAND3_X1 U20521 ( .A1(n17272), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17390), 
        .ZN(n17271) );
  OAI221_X1 U20522 ( .B1(n17272), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17390), 
        .C2(n17490), .A(n17271), .ZN(P3_U2689) );
  OAI21_X1 U20523 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17306), .A(n17390), .ZN(
        n17287) );
  AOI22_X1 U20524 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17273) );
  OAI21_X1 U20525 ( .B1(n17275), .B2(n17274), .A(n17273), .ZN(n17286) );
  AOI22_X1 U20526 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20527 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20528 ( .B1(n13933), .B2(n17277), .A(n17276), .ZN(n17281) );
  AOI22_X1 U20529 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U20530 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17278) );
  OAI211_X1 U20531 ( .C1(n13966), .C2(n17381), .A(n17279), .B(n17278), .ZN(
        n17280) );
  AOI211_X1 U20532 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17281), .B(n17280), .ZN(n17282) );
  OAI211_X1 U20533 ( .C1(n13879), .C2(n17284), .A(n17283), .B(n17282), .ZN(
        n17285) );
  AOI211_X1 U20534 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17286), .B(n17285), .ZN(n17496) );
  OAI22_X1 U20535 ( .A1(n17288), .A2(n17287), .B1(n17496), .B2(n17390), .ZN(
        P3_U2691) );
  INV_X1 U20536 ( .A(n17318), .ZN(n17289) );
  OAI21_X1 U20537 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17289), .A(n17390), .ZN(
        n17305) );
  INV_X1 U20538 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20539 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20540 ( .B1(n13879), .B2(n17291), .A(n17290), .ZN(n17304) );
  AOI22_X1 U20541 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17300) );
  OAI22_X1 U20542 ( .A1(n17293), .A2(n17292), .B1(n13966), .B2(n17383), .ZN(
        n17298) );
  AOI22_X1 U20543 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20544 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20545 ( .A1(n17241), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17335), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17294) );
  NAND3_X1 U20546 ( .A1(n17296), .A2(n17295), .A3(n17294), .ZN(n17297) );
  AOI211_X1 U20547 ( .C1(n15618), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17298), .B(n17297), .ZN(n17299) );
  OAI211_X1 U20548 ( .C1(n17302), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        n17303) );
  AOI211_X1 U20549 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17304), .B(n17303), .ZN(n17500) );
  OAI22_X1 U20550 ( .A1(n17306), .A2(n17305), .B1(n17500), .B2(n17390), .ZN(
        P3_U2692) );
  AOI22_X1 U20551 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20552 ( .A1(n15633), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20553 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17307) );
  OAI211_X1 U20554 ( .C1(n13966), .C2(n17389), .A(n17308), .B(n17307), .ZN(
        n17314) );
  AOI22_X1 U20555 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20556 ( .A1(n13852), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20557 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15677), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17310) );
  NAND2_X1 U20558 ( .A1(n17335), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n17309) );
  NAND4_X1 U20559 ( .A1(n17312), .A2(n17311), .A3(n17310), .A4(n17309), .ZN(
        n17313) );
  AOI211_X1 U20560 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17314), .B(n17313), .ZN(n17315) );
  OAI211_X1 U20561 ( .C1(n9813), .C2(n17317), .A(n17316), .B(n17315), .ZN(
        n17504) );
  INV_X1 U20562 ( .A(n17504), .ZN(n17320) );
  OAI21_X1 U20563 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17343), .A(n17318), .ZN(
        n17319) );
  AOI22_X1 U20564 ( .A1(n17396), .A2(n17320), .B1(n17319), .B2(n17390), .ZN(
        P3_U2693) );
  INV_X1 U20565 ( .A(n17321), .ZN(n17322) );
  OAI21_X1 U20566 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17322), .A(n17390), .ZN(
        n17342) );
  AOI22_X1 U20567 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17325) );
  OAI21_X1 U20568 ( .B1(n13934), .B2(n18693), .A(n17325), .ZN(n17341) );
  INV_X1 U20569 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20570 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20571 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17327) );
  OAI21_X1 U20572 ( .B1(n13966), .B2(n17391), .A(n17327), .ZN(n17334) );
  AOI22_X1 U20573 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20574 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17330) );
  OAI211_X1 U20575 ( .C1(n13901), .C2(n17332), .A(n17331), .B(n17330), .ZN(
        n17333) );
  AOI211_X1 U20576 ( .C1(n17335), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17334), .B(n17333), .ZN(n17336) );
  OAI211_X1 U20577 ( .C1(n17339), .C2(n17338), .A(n17337), .B(n17336), .ZN(
        n17340) );
  AOI211_X1 U20578 ( .C1(n17345), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n17341), .B(n17340), .ZN(n17508) );
  OAI22_X1 U20579 ( .A1(n17343), .A2(n17342), .B1(n17508), .B2(n17390), .ZN(
        P3_U2694) );
  NAND2_X1 U20580 ( .A1(n17445), .A2(n17344), .ZN(n17363) );
  NOR2_X1 U20581 ( .A1(n17396), .A2(n17344), .ZN(n17364) );
  AOI22_X1 U20582 ( .A1(n15677), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20583 ( .A1(n17345), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U20584 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15633), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17346) );
  OAI211_X1 U20585 ( .C1(n17349), .C2(n17348), .A(n17347), .B(n17346), .ZN(
        n17358) );
  AOI22_X1 U20586 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20587 ( .A1(n17351), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20588 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17354) );
  NAND2_X1 U20589 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n17353) );
  NAND4_X1 U20590 ( .A1(n17356), .A2(n17355), .A3(n17354), .A4(n17353), .ZN(
        n17357) );
  AOI211_X1 U20591 ( .C1(n17241), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17358), .B(n17357), .ZN(n17359) );
  OAI211_X1 U20592 ( .C1(n13966), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        n17512) );
  AOI22_X1 U20593 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17364), .B1(n17396), .B2(
        n17512), .ZN(n17362) );
  OAI21_X1 U20594 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        P3_U2695) );
  INV_X1 U20595 ( .A(n17368), .ZN(n17365) );
  OAI21_X1 U20596 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17365), .A(n17364), .ZN(
        n17366) );
  OAI21_X1 U20597 ( .B1(n17390), .B2(n17367), .A(n17366), .ZN(P3_U2696) );
  OAI21_X1 U20598 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17375), .A(n17368), .ZN(
        n17369) );
  AOI22_X1 U20599 ( .A1(n17396), .A2(n17370), .B1(n17369), .B2(n17390), .ZN(
        P3_U2697) );
  NOR2_X1 U20600 ( .A1(n17384), .A2(n17371), .ZN(n17372) );
  OAI21_X1 U20601 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17372), .A(n17390), .ZN(
        n17374) );
  OAI22_X1 U20602 ( .A1(n17375), .A2(n17374), .B1(n17373), .B2(n17390), .ZN(
        P3_U2698) );
  INV_X1 U20603 ( .A(n17393), .ZN(n17395) );
  NAND2_X1 U20604 ( .A1(n17376), .A2(n17395), .ZN(n17386) );
  NOR2_X1 U20605 ( .A1(n17377), .A2(n17386), .ZN(n17379) );
  OAI21_X1 U20606 ( .B1(n17379), .B2(n17396), .A(P3_EBX_REG_4__SCAN_IN), .ZN(
        n17378) );
  OAI21_X1 U20607 ( .B1(n17379), .B2(P3_EBX_REG_4__SCAN_IN), .A(n17378), .ZN(
        n17380) );
  OAI21_X1 U20608 ( .B1(n17390), .B2(n17381), .A(n17380), .ZN(P3_U2699) );
  NAND3_X1 U20609 ( .A1(n17386), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17390), .ZN(
        n17382) );
  OAI221_X1 U20610 ( .B1(n17386), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17390), 
        .C2(n17383), .A(n17382), .ZN(P3_U2700) );
  AOI21_X1 U20611 ( .B1(n17445), .B2(n17385), .A(n17384), .ZN(n17387) );
  OAI21_X1 U20612 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17387), .A(n17386), .ZN(
        n17388) );
  AOI21_X1 U20613 ( .B1(n17396), .B2(n17389), .A(n17388), .ZN(P3_U2701) );
  OAI222_X1 U20614 ( .A1(n17394), .A2(n17393), .B1(n17392), .B2(n17399), .C1(
        n17391), .C2(n17390), .ZN(P3_U2702) );
  AOI22_X1 U20615 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17396), .B1(
        n17395), .B2(n17398), .ZN(n17397) );
  OAI21_X1 U20616 ( .B1(n17399), .B2(n17398), .A(n17397), .ZN(P3_U2703) );
  INV_X1 U20617 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17613) );
  INV_X1 U20618 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17610) );
  INV_X1 U20619 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17608) );
  INV_X1 U20620 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17606) );
  INV_X1 U20621 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17656) );
  INV_X1 U20622 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17627) );
  INV_X1 U20623 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17625) );
  NAND2_X1 U20624 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17545) );
  NAND2_X1 U20625 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17517) );
  NOR4_X1 U20626 ( .A1(n17627), .A2(n17625), .A3(n17545), .A4(n17517), .ZN(
        n17400) );
  INV_X1 U20627 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17641) );
  INV_X1 U20628 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17639) );
  INV_X1 U20629 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17637) );
  NOR3_X1 U20630 ( .A1(n17641), .A2(n17639), .A3(n17637), .ZN(n17485) );
  INV_X1 U20631 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17649) );
  INV_X1 U20632 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17646) );
  INV_X1 U20633 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17643) );
  NOR3_X1 U20634 ( .A1(n17649), .A2(n17646), .A3(n17643), .ZN(n17484) );
  INV_X1 U20635 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17600) );
  INV_X1 U20636 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17598) );
  INV_X1 U20637 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17596) );
  INV_X1 U20638 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17594) );
  NOR4_X1 U20639 ( .A1(n17600), .A2(n17598), .A3(n17596), .A4(n17594), .ZN(
        n17402) );
  NAND4_X1 U20640 ( .A1(n17444), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .A4(n17402), .ZN(n17439) );
  NAND2_X1 U20641 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17419), .ZN(n17416) );
  INV_X1 U20642 ( .A(n17416), .ZN(n17411) );
  NAND2_X1 U20643 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17411), .ZN(n17410) );
  NOR2_X1 U20644 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17410), .ZN(n17404) );
  NAND2_X1 U20645 ( .A1(n17537), .A2(n17410), .ZN(n17409) );
  OAI21_X1 U20646 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17544), .A(n17409), .ZN(
        n17403) );
  AOI22_X1 U20647 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17404), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17403), .ZN(n17405) );
  OAI21_X1 U20648 ( .B1(n19467), .B2(n17455), .A(n17405), .ZN(P3_U2704) );
  INV_X1 U20649 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17619) );
  NOR2_X2 U20650 ( .A1(n18393), .A2(n17537), .ZN(n17474) );
  OAI22_X1 U20651 ( .A1(n17406), .A2(n17549), .B1(n19460), .B2(n17455), .ZN(
        n17407) );
  AOI21_X1 U20652 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17474), .A(n17407), .ZN(
        n17408) );
  OAI221_X1 U20653 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17410), .C1(n17619), 
        .C2(n17409), .A(n17408), .ZN(P3_U2705) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17473), .ZN(n17413) );
  OAI211_X1 U20655 ( .C1(n17411), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17537), .B(
        n17410), .ZN(n17412) );
  OAI211_X1 U20656 ( .C1(n17414), .C2(n17549), .A(n17413), .B(n17412), .ZN(
        P3_U2706) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17474), .B1(n17528), .B2(
        n17415), .ZN(n17418) );
  OAI211_X1 U20658 ( .C1(n17419), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17537), .B(
        n17416), .ZN(n17417) );
  OAI211_X1 U20659 ( .C1(n17455), .C2(n19450), .A(n17418), .B(n17417), .ZN(
        P3_U2707) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17473), .ZN(n17422) );
  AOI211_X1 U20661 ( .C1(n17613), .C2(n17425), .A(n17419), .B(n17530), .ZN(
        n17420) );
  INV_X1 U20662 ( .A(n17420), .ZN(n17421) );
  OAI211_X1 U20663 ( .C1(n17423), .C2(n17549), .A(n17422), .B(n17421), .ZN(
        P3_U2708) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17474), .B1(n17528), .B2(
        n17424), .ZN(n17427) );
  OAI211_X1 U20665 ( .C1(n9924), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17537), .B(
        n17425), .ZN(n17426) );
  OAI211_X1 U20666 ( .C1(n17455), .C2(n19437), .A(n17427), .B(n17426), .ZN(
        P3_U2709) );
  AOI22_X1 U20667 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17473), .ZN(n17430) );
  AOI211_X1 U20668 ( .C1(n17610), .C2(n17434), .A(n9924), .B(n17530), .ZN(
        n17428) );
  INV_X1 U20669 ( .A(n17428), .ZN(n17429) );
  OAI211_X1 U20670 ( .C1(n17431), .C2(n17549), .A(n17430), .B(n17429), .ZN(
        P3_U2710) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17474), .B1(n17528), .B2(
        n17432), .ZN(n17437) );
  OAI21_X1 U20672 ( .B1(n17608), .B2(n17530), .A(n17433), .ZN(n17435) );
  NAND2_X1 U20673 ( .A1(n17435), .A2(n17434), .ZN(n17436) );
  OAI211_X1 U20674 ( .C1(n17455), .C2(n18375), .A(n17437), .B(n17436), .ZN(
        P3_U2711) );
  AOI211_X1 U20675 ( .C1(n17606), .C2(n17439), .A(n17530), .B(n17438), .ZN(
        n17440) );
  AOI21_X1 U20676 ( .B1(n17473), .B2(BUF2_REG_23__SCAN_IN), .A(n17440), .ZN(
        n17442) );
  NAND2_X1 U20677 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17474), .ZN(n17441) );
  OAI211_X1 U20678 ( .C1(n17443), .C2(n17549), .A(n17442), .B(n17441), .ZN(
        P3_U2712) );
  NAND3_X1 U20679 ( .A1(n17445), .A2(n17444), .A3(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17469) );
  NAND2_X1 U20680 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17464), .ZN(n17460) );
  NOR2_X1 U20681 ( .A1(n17600), .A2(n17460), .ZN(n17452) );
  NAND2_X1 U20682 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17452), .ZN(n17450) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17473), .B1(n17528), .B2(
        n17446), .ZN(n17449) );
  OR2_X1 U20684 ( .A1(n17530), .A2(n17452), .ZN(n17459) );
  OAI21_X1 U20685 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17544), .A(n17459), .ZN(
        n17447) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17474), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17447), .ZN(n17448) );
  OAI211_X1 U20687 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17450), .A(n17449), .B(
        n17448), .ZN(P3_U2713) );
  INV_X1 U20688 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17602) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17473), .B1(n17528), .B2(
        n17451), .ZN(n17454) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17474), .B1(n17452), .B2(
        n17602), .ZN(n17453) );
  OAI211_X1 U20691 ( .C1(n17602), .C2(n17459), .A(n17454), .B(n17453), .ZN(
        P3_U2714) );
  OAI22_X1 U20692 ( .A1(n17456), .A2(n17549), .B1(n18390), .B2(n17455), .ZN(
        n17457) );
  AOI21_X1 U20693 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17474), .A(n17457), .ZN(
        n17458) );
  OAI221_X1 U20694 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17460), .C1(n17600), 
        .C2(n17459), .A(n17458), .ZN(P3_U2715) );
  AOI22_X1 U20695 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17473), .ZN(n17462) );
  OAI211_X1 U20696 ( .C1(n17464), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17537), .B(
        n17460), .ZN(n17461) );
  OAI211_X1 U20697 ( .C1(n17463), .C2(n17549), .A(n17462), .B(n17461), .ZN(
        P3_U2716) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17473), .ZN(n17467) );
  AOI211_X1 U20699 ( .C1(n17596), .C2(n17469), .A(n17464), .B(n17530), .ZN(
        n17465) );
  INV_X1 U20700 ( .A(n17465), .ZN(n17466) );
  OAI211_X1 U20701 ( .C1(n17468), .C2(n17549), .A(n17467), .B(n17466), .ZN(
        P3_U2717) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17473), .ZN(n17471) );
  OAI211_X1 U20703 ( .C1(n17444), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17537), .B(
        n17469), .ZN(n17470) );
  OAI211_X1 U20704 ( .C1(n17472), .C2(n17549), .A(n17471), .B(n17470), .ZN(
        P3_U2718) );
  AOI22_X1 U20705 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17474), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17473), .ZN(n17477) );
  OAI211_X1 U20706 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17480), .A(n17537), .B(
        n17475), .ZN(n17476) );
  OAI211_X1 U20707 ( .C1(n17478), .C2(n17549), .A(n17477), .B(n17476), .ZN(
        P3_U2719) );
  AOI22_X1 U20708 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17543), .B1(n17528), .B2(
        n17479), .ZN(n17483) );
  AOI211_X1 U20709 ( .C1(n17656), .C2(n17487), .A(n17530), .B(n17480), .ZN(
        n17481) );
  INV_X1 U20710 ( .A(n17481), .ZN(n17482) );
  NAND2_X1 U20711 ( .A1(n17483), .A2(n17482), .ZN(P3_U2720) );
  INV_X1 U20712 ( .A(n17484), .ZN(n17486) );
  NOR2_X1 U20713 ( .A1(n18400), .A2(n17513), .ZN(n17520) );
  NAND2_X1 U20714 ( .A1(n17485), .A2(n17520), .ZN(n17503) );
  NOR2_X1 U20715 ( .A1(n17486), .A2(n17503), .ZN(n17493) );
  OAI211_X1 U20716 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17493), .A(n17537), .B(
        n17487), .ZN(n17489) );
  NAND2_X1 U20717 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17543), .ZN(n17488) );
  OAI211_X1 U20718 ( .C1(n17490), .C2(n17549), .A(n17489), .B(n17488), .ZN(
        P3_U2721) );
  NOR2_X1 U20719 ( .A1(n17643), .A2(n17503), .ZN(n17495) );
  AND2_X1 U20720 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17495), .ZN(n17498) );
  AOI21_X1 U20721 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17537), .A(n17498), .ZN(
        n17492) );
  OAI222_X1 U20722 ( .A1(n17541), .A2(n17494), .B1(n17493), .B2(n17492), .C1(
        n17549), .C2(n17491), .ZN(P3_U2722) );
  AOI21_X1 U20723 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17537), .A(n17495), .ZN(
        n17497) );
  OAI222_X1 U20724 ( .A1(n17541), .A2(n17499), .B1(n17498), .B2(n17497), .C1(
        n17549), .C2(n17496), .ZN(P3_U2723) );
  NAND2_X1 U20725 ( .A1(n17537), .A2(n17503), .ZN(n17506) );
  INV_X1 U20726 ( .A(n17500), .ZN(n17501) );
  AOI22_X1 U20727 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17543), .B1(n17528), .B2(
        n17501), .ZN(n17502) );
  OAI221_X1 U20728 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17503), .C1(n17643), 
        .C2(n17506), .A(n17502), .ZN(P3_U2724) );
  NAND3_X1 U20729 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17520), .ZN(n17507) );
  AOI22_X1 U20730 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17543), .B1(n17528), .B2(
        n17504), .ZN(n17505) );
  OAI221_X1 U20731 ( .B1(n17506), .B2(n17641), .C1(n17506), .C2(n17507), .A(
        n17505), .ZN(P3_U2725) );
  INV_X1 U20732 ( .A(n17507), .ZN(n17510) );
  AOI22_X1 U20733 ( .A1(n17520), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17537), .ZN(n17509) );
  OAI222_X1 U20734 ( .A1(n17541), .A2(n17511), .B1(n17510), .B2(n17509), .C1(
        n17549), .C2(n17508), .ZN(P3_U2726) );
  AOI22_X1 U20735 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17543), .B1(n17528), .B2(
        n17512), .ZN(n17516) );
  OAI221_X1 U20736 ( .B1(n17514), .B2(P3_EAX_REG_8__SCAN_IN), .C1(n17513), 
        .C2(n17637), .A(n17537), .ZN(n17515) );
  NAND2_X1 U20737 ( .A1(n17516), .A2(n17515), .ZN(P3_U2727) );
  NAND2_X1 U20738 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17540), .ZN(n17532) );
  NOR2_X1 U20739 ( .A1(n17517), .A2(n17532), .ZN(n17526) );
  AOI22_X1 U20740 ( .A1(n17526), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17537), .ZN(n17519) );
  OAI222_X1 U20741 ( .A1(n17541), .A2(n18402), .B1(n17520), .B2(n17519), .C1(
        n17549), .C2(n17518), .ZN(P3_U2728) );
  INV_X1 U20742 ( .A(n17526), .ZN(n17523) );
  NAND2_X1 U20743 ( .A1(n17523), .A2(P3_EAX_REG_6__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U20744 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17543), .B1(n17528), .B2(
        n17954), .ZN(n17521) );
  OAI221_X1 U20745 ( .B1(n17523), .B2(P3_EAX_REG_6__SCAN_IN), .C1(n17522), 
        .C2(n17530), .A(n17521), .ZN(P3_U2729) );
  INV_X1 U20746 ( .A(n17532), .ZN(n17535) );
  AOI22_X1 U20747 ( .A1(n17535), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17537), .ZN(n17525) );
  OAI222_X1 U20748 ( .A1(n17541), .A2(n18394), .B1(n17526), .B2(n17525), .C1(
        n17549), .C2(n17524), .ZN(P3_U2730) );
  NAND2_X1 U20749 ( .A1(n17532), .A2(P3_EAX_REG_4__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20750 ( .A1(n17543), .A2(BUF2_REG_4__SCAN_IN), .B1(n17528), .B2(
        n17527), .ZN(n17529) );
  OAI221_X1 U20751 ( .B1(n17532), .B2(P3_EAX_REG_4__SCAN_IN), .C1(n17531), 
        .C2(n17530), .A(n17529), .ZN(P3_U2731) );
  AOI21_X1 U20752 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17537), .A(n17540), .ZN(
        n17534) );
  OAI222_X1 U20753 ( .A1(n18386), .A2(n17541), .B1(n17535), .B2(n17534), .C1(
        n17549), .C2(n17533), .ZN(P3_U2732) );
  NOR2_X1 U20754 ( .A1(n17545), .A2(n17544), .ZN(n17536) );
  AOI21_X1 U20755 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17537), .A(n17536), .ZN(
        n17539) );
  OAI222_X1 U20756 ( .A1(n18382), .A2(n17541), .B1(n17540), .B2(n17539), .C1(
        n17549), .C2(n17538), .ZN(P3_U2733) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17543), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17542), .ZN(n17548) );
  INV_X1 U20758 ( .A(n17544), .ZN(n17546) );
  OAI211_X1 U20759 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17546), .B(n17545), .ZN(n17547) );
  OAI211_X1 U20760 ( .C1(n17550), .C2(n17549), .A(n17548), .B(n17547), .ZN(
        P3_U2734) );
  NOR2_X4 U20761 ( .A1(n17585), .A2(n17569), .ZN(n17566) );
  AND2_X1 U20762 ( .A1(n17566), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20763 ( .A1(n17585), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17566), .ZN(n17552) );
  OAI21_X1 U20764 ( .B1(n17619), .B2(n17568), .A(n17552), .ZN(P3_U2737) );
  INV_X1 U20765 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17617) );
  AOI22_X1 U20766 ( .A1(n17585), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17553) );
  OAI21_X1 U20767 ( .B1(n17617), .B2(n17568), .A(n17553), .ZN(P3_U2738) );
  INV_X1 U20768 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U20769 ( .A1(n17585), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17554) );
  OAI21_X1 U20770 ( .B1(n17615), .B2(n17568), .A(n17554), .ZN(P3_U2739) );
  AOI22_X1 U20771 ( .A1(n17585), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17555) );
  OAI21_X1 U20772 ( .B1(n17613), .B2(n17568), .A(n17555), .ZN(P3_U2740) );
  AOI22_X1 U20773 ( .A1(n17585), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17556) );
  OAI21_X1 U20774 ( .B1(n10110), .B2(n17568), .A(n17556), .ZN(P3_U2741) );
  AOI22_X1 U20775 ( .A1(n17585), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17557) );
  OAI21_X1 U20776 ( .B1(n17610), .B2(n17568), .A(n17557), .ZN(P3_U2742) );
  AOI22_X1 U20777 ( .A1(n17585), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17558) );
  OAI21_X1 U20778 ( .B1(n17608), .B2(n17568), .A(n17558), .ZN(P3_U2743) );
  INV_X2 U20779 ( .A(n19006), .ZN(n17585) );
  AOI22_X1 U20780 ( .A1(n17585), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17559) );
  OAI21_X1 U20781 ( .B1(n17606), .B2(n17568), .A(n17559), .ZN(P3_U2744) );
  INV_X1 U20782 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17604) );
  AOI22_X1 U20783 ( .A1(n17585), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17560) );
  OAI21_X1 U20784 ( .B1(n17604), .B2(n17568), .A(n17560), .ZN(P3_U2745) );
  AOI22_X1 U20785 ( .A1(n17585), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17561) );
  OAI21_X1 U20786 ( .B1(n17602), .B2(n17568), .A(n17561), .ZN(P3_U2746) );
  AOI22_X1 U20787 ( .A1(n17585), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17562) );
  OAI21_X1 U20788 ( .B1(n17600), .B2(n17568), .A(n17562), .ZN(P3_U2747) );
  AOI22_X1 U20789 ( .A1(n17585), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17563) );
  OAI21_X1 U20790 ( .B1(n17598), .B2(n17568), .A(n17563), .ZN(P3_U2748) );
  AOI22_X1 U20791 ( .A1(n17585), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17564) );
  OAI21_X1 U20792 ( .B1(n17596), .B2(n17568), .A(n17564), .ZN(P3_U2749) );
  AOI22_X1 U20793 ( .A1(n17585), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17565) );
  OAI21_X1 U20794 ( .B1(n17594), .B2(n17568), .A(n17565), .ZN(P3_U2750) );
  INV_X1 U20795 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U20796 ( .A1(n17585), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17567) );
  OAI21_X1 U20797 ( .B1(n17592), .B2(n17568), .A(n17567), .ZN(P3_U2751) );
  AOI22_X1 U20798 ( .A1(n17585), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17570) );
  OAI21_X1 U20799 ( .B1(n17656), .B2(n17587), .A(n17570), .ZN(P3_U2752) );
  INV_X1 U20800 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U20801 ( .A1(n17585), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17571) );
  OAI21_X1 U20802 ( .B1(n17651), .B2(n17587), .A(n17571), .ZN(P3_U2753) );
  AOI22_X1 U20803 ( .A1(n17585), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17572) );
  OAI21_X1 U20804 ( .B1(n17649), .B2(n17587), .A(n17572), .ZN(P3_U2754) );
  AOI22_X1 U20805 ( .A1(n17585), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17573) );
  OAI21_X1 U20806 ( .B1(n17646), .B2(n17587), .A(n17573), .ZN(P3_U2755) );
  AOI22_X1 U20807 ( .A1(n17585), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17574) );
  OAI21_X1 U20808 ( .B1(n17643), .B2(n17587), .A(n17574), .ZN(P3_U2756) );
  AOI22_X1 U20809 ( .A1(n17585), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U20810 ( .B1(n17641), .B2(n17587), .A(n17575), .ZN(P3_U2757) );
  AOI22_X1 U20811 ( .A1(n17585), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17576) );
  OAI21_X1 U20812 ( .B1(n17639), .B2(n17587), .A(n17576), .ZN(P3_U2758) );
  AOI22_X1 U20813 ( .A1(n17585), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17577) );
  OAI21_X1 U20814 ( .B1(n17637), .B2(n17587), .A(n17577), .ZN(P3_U2759) );
  INV_X1 U20815 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17635) );
  AOI22_X1 U20816 ( .A1(n17585), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17578) );
  OAI21_X1 U20817 ( .B1(n17635), .B2(n17587), .A(n17578), .ZN(P3_U2760) );
  INV_X1 U20818 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U20819 ( .A1(n17585), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17579) );
  OAI21_X1 U20820 ( .B1(n17633), .B2(n17587), .A(n17579), .ZN(P3_U2761) );
  INV_X1 U20821 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U20822 ( .A1(n17585), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17580) );
  OAI21_X1 U20823 ( .B1(n17631), .B2(n17587), .A(n17580), .ZN(P3_U2762) );
  INV_X1 U20824 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17629) );
  AOI22_X1 U20825 ( .A1(n17585), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17581) );
  OAI21_X1 U20826 ( .B1(n17629), .B2(n17587), .A(n17581), .ZN(P3_U2763) );
  AOI22_X1 U20827 ( .A1(n17585), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17582) );
  OAI21_X1 U20828 ( .B1(n17627), .B2(n17587), .A(n17582), .ZN(P3_U2764) );
  AOI22_X1 U20829 ( .A1(n17585), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17583) );
  OAI21_X1 U20830 ( .B1(n17625), .B2(n17587), .A(n17583), .ZN(P3_U2765) );
  INV_X1 U20831 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U20832 ( .A1(n17585), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17584) );
  OAI21_X1 U20833 ( .B1(n17623), .B2(n17587), .A(n17584), .ZN(P3_U2766) );
  AOI22_X1 U20834 ( .A1(n17585), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17586) );
  OAI21_X1 U20835 ( .B1(n17621), .B2(n17587), .A(n17586), .ZN(P3_U2767) );
  AND2_X1 U20836 ( .A1(n19012), .A2(n17590), .ZN(n18848) );
  AOI22_X1 U20837 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17652), .ZN(n17591) );
  OAI21_X1 U20838 ( .B1(n17592), .B2(n17655), .A(n17591), .ZN(P3_U2768) );
  AOI22_X1 U20839 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17652), .ZN(n17593) );
  OAI21_X1 U20840 ( .B1(n17594), .B2(n17655), .A(n17593), .ZN(P3_U2769) );
  AOI22_X1 U20841 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17652), .ZN(n17595) );
  OAI21_X1 U20842 ( .B1(n17596), .B2(n17655), .A(n17595), .ZN(P3_U2770) );
  AOI22_X1 U20843 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17652), .ZN(n17597) );
  OAI21_X1 U20844 ( .B1(n17598), .B2(n17655), .A(n17597), .ZN(P3_U2771) );
  AOI22_X1 U20845 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17652), .ZN(n17599) );
  OAI21_X1 U20846 ( .B1(n17600), .B2(n17655), .A(n17599), .ZN(P3_U2772) );
  AOI22_X1 U20847 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17652), .ZN(n17601) );
  OAI21_X1 U20848 ( .B1(n17602), .B2(n17655), .A(n17601), .ZN(P3_U2773) );
  AOI22_X1 U20849 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17652), .ZN(n17603) );
  OAI21_X1 U20850 ( .B1(n17604), .B2(n17655), .A(n17603), .ZN(P3_U2774) );
  AOI22_X1 U20851 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17652), .ZN(n17605) );
  OAI21_X1 U20852 ( .B1(n17606), .B2(n17655), .A(n17605), .ZN(P3_U2775) );
  AOI22_X1 U20853 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17652), .ZN(n17607) );
  OAI21_X1 U20854 ( .B1(n17608), .B2(n17655), .A(n17607), .ZN(P3_U2776) );
  AOI22_X1 U20855 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17652), .ZN(n17609) );
  OAI21_X1 U20856 ( .B1(n17610), .B2(n17655), .A(n17609), .ZN(P3_U2777) );
  AOI22_X1 U20857 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17652), .ZN(n17611) );
  OAI21_X1 U20858 ( .B1(n10110), .B2(n17655), .A(n17611), .ZN(P3_U2778) );
  AOI22_X1 U20859 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17644), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17652), .ZN(n17612) );
  OAI21_X1 U20860 ( .B1(n17613), .B2(n17655), .A(n17612), .ZN(P3_U2779) );
  AOI22_X1 U20861 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17652), .ZN(n17614) );
  OAI21_X1 U20862 ( .B1(n17615), .B2(n17655), .A(n17614), .ZN(P3_U2780) );
  AOI22_X1 U20863 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17652), .ZN(n17616) );
  OAI21_X1 U20864 ( .B1(n17617), .B2(n17655), .A(n17616), .ZN(P3_U2781) );
  AOI22_X1 U20865 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17653), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17652), .ZN(n17618) );
  OAI21_X1 U20866 ( .B1(n17619), .B2(n17655), .A(n17618), .ZN(P3_U2782) );
  AOI22_X1 U20867 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17652), .ZN(n17620) );
  OAI21_X1 U20868 ( .B1(n17621), .B2(n17655), .A(n17620), .ZN(P3_U2783) );
  AOI22_X1 U20869 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17652), .ZN(n17622) );
  OAI21_X1 U20870 ( .B1(n17623), .B2(n17655), .A(n17622), .ZN(P3_U2784) );
  AOI22_X1 U20871 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17647), .ZN(n17624) );
  OAI21_X1 U20872 ( .B1(n17625), .B2(n17655), .A(n17624), .ZN(P3_U2785) );
  AOI22_X1 U20873 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17647), .ZN(n17626) );
  OAI21_X1 U20874 ( .B1(n17627), .B2(n17655), .A(n17626), .ZN(P3_U2786) );
  AOI22_X1 U20875 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17647), .ZN(n17628) );
  OAI21_X1 U20876 ( .B1(n17629), .B2(n17655), .A(n17628), .ZN(P3_U2787) );
  AOI22_X1 U20877 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17647), .ZN(n17630) );
  OAI21_X1 U20878 ( .B1(n17631), .B2(n17655), .A(n17630), .ZN(P3_U2788) );
  AOI22_X1 U20879 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17647), .ZN(n17632) );
  OAI21_X1 U20880 ( .B1(n17633), .B2(n17655), .A(n17632), .ZN(P3_U2789) );
  AOI22_X1 U20881 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17647), .ZN(n17634) );
  OAI21_X1 U20882 ( .B1(n17635), .B2(n17655), .A(n17634), .ZN(P3_U2790) );
  AOI22_X1 U20883 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17647), .ZN(n17636) );
  OAI21_X1 U20884 ( .B1(n17637), .B2(n17655), .A(n17636), .ZN(P3_U2791) );
  AOI22_X1 U20885 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17647), .ZN(n17638) );
  OAI21_X1 U20886 ( .B1(n17639), .B2(n17655), .A(n17638), .ZN(P3_U2792) );
  AOI22_X1 U20887 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17644), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17652), .ZN(n17640) );
  OAI21_X1 U20888 ( .B1(n17641), .B2(n17655), .A(n17640), .ZN(P3_U2793) );
  AOI22_X1 U20889 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17647), .ZN(n17642) );
  OAI21_X1 U20890 ( .B1(n17643), .B2(n17655), .A(n17642), .ZN(P3_U2794) );
  AOI22_X1 U20891 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17644), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17652), .ZN(n17645) );
  OAI21_X1 U20892 ( .B1(n17646), .B2(n17655), .A(n17645), .ZN(P3_U2795) );
  AOI22_X1 U20893 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17647), .ZN(n17648) );
  OAI21_X1 U20894 ( .B1(n17649), .B2(n17655), .A(n17648), .ZN(P3_U2796) );
  AOI22_X1 U20895 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17652), .ZN(n17650) );
  OAI21_X1 U20896 ( .B1(n17651), .B2(n17655), .A(n17650), .ZN(P3_U2797) );
  AOI22_X1 U20897 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17653), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17652), .ZN(n17654) );
  OAI21_X1 U20898 ( .B1(n17656), .B2(n17655), .A(n17654), .ZN(P3_U2798) );
  OAI21_X1 U20899 ( .B1(n17657), .B2(n18029), .A(n18028), .ZN(n17658) );
  AOI21_X1 U20900 ( .B1(n17923), .B2(n17662), .A(n17658), .ZN(n17690) );
  OAI21_X1 U20901 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17802), .A(
        n17690), .ZN(n17679) );
  NOR2_X1 U20902 ( .A1(n17889), .A2(n18000), .ZN(n17769) );
  INV_X1 U20903 ( .A(n17659), .ZN(n18039) );
  OAI22_X1 U20904 ( .A1(n17660), .A2(n17938), .B1(n18039), .B2(n18033), .ZN(
        n17696) );
  NOR2_X1 U20905 ( .A1(n17686), .A2(n17696), .ZN(n17687) );
  NOR3_X1 U20906 ( .A1(n17769), .A2(n17687), .A3(n17661), .ZN(n17668) );
  NOR2_X1 U20907 ( .A1(n17777), .A2(n17662), .ZN(n17683) );
  OAI211_X1 U20908 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17683), .B(n17663), .ZN(n17665) );
  OAI211_X1 U20909 ( .C1(n17857), .C2(n17666), .A(n17665), .B(n17664), .ZN(
        n17667) );
  AOI211_X1 U20910 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17679), .A(
        n17668), .B(n17667), .ZN(n17673) );
  OAI211_X1 U20911 ( .C1(n17671), .C2(n17670), .A(n17934), .B(n17669), .ZN(
        n17672) );
  OAI211_X1 U20912 ( .C1(n17685), .C2(n17674), .A(n17673), .B(n17672), .ZN(
        P3_U2802) );
  NOR2_X1 U20913 ( .A1(n17676), .A2(n17675), .ZN(n17677) );
  XNOR2_X1 U20914 ( .A(n17677), .B(n17811), .ZN(n18047) );
  AOI22_X1 U20915 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17679), .B1(
        n17872), .B2(n17678), .ZN(n17680) );
  NAND2_X1 U20916 ( .A1(n18357), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18045) );
  OAI211_X1 U20917 ( .C1(n18047), .C2(n17893), .A(n17680), .B(n18045), .ZN(
        n17681) );
  AOI21_X1 U20918 ( .B1(n17683), .B2(n17682), .A(n17681), .ZN(n17684) );
  OAI221_X1 U20919 ( .B1(n17687), .B2(n17686), .C1(n17687), .C2(n17685), .A(
        n17684), .ZN(P3_U2803) );
  INV_X1 U20920 ( .A(n9847), .ZN(n17800) );
  NOR2_X1 U20921 ( .A1(n18058), .A2(n18059), .ZN(n18057) );
  NAND2_X1 U20922 ( .A1(n18057), .A2(n18048), .ZN(n18055) );
  INV_X1 U20923 ( .A(n17802), .ZN(n17692) );
  AOI21_X1 U20924 ( .B1(n18745), .B2(n17688), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17689) );
  INV_X1 U20925 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18933) );
  OAI22_X1 U20926 ( .A1(n17690), .A2(n17689), .B1(n18339), .B2(n18933), .ZN(
        n17691) );
  AOI221_X1 U20927 ( .B1(n17872), .B2(n17693), .C1(n17692), .C2(n17693), .A(
        n17691), .ZN(n17698) );
  OAI21_X1 U20928 ( .B1(n17695), .B2(n18048), .A(n17694), .ZN(n18051) );
  AOI22_X1 U20929 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17696), .B1(
        n17934), .B2(n18051), .ZN(n17697) );
  OAI211_X1 U20930 ( .C1(n17800), .C2(n18055), .A(n17698), .B(n17697), .ZN(
        P3_U2804) );
  NAND3_X1 U20931 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18169), .A3(
        n17713), .ZN(n17699) );
  XNOR2_X1 U20932 ( .A(n17699), .B(n18058), .ZN(n18067) );
  OAI21_X1 U20933 ( .B1(n17700), .B2(n18029), .A(n18028), .ZN(n17701) );
  AOI21_X1 U20934 ( .B1(n18745), .B2(n17702), .A(n17701), .ZN(n17731) );
  OAI21_X1 U20935 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17802), .A(
        n17731), .ZN(n17717) );
  NOR2_X1 U20936 ( .A1(n17777), .A2(n17702), .ZN(n17719) );
  OAI211_X1 U20937 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17719), .B(n17703), .ZN(n17704) );
  NAND2_X1 U20938 ( .A1(n18297), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18065) );
  OAI211_X1 U20939 ( .C1(n17857), .C2(n17705), .A(n17704), .B(n18065), .ZN(
        n17711) );
  XNOR2_X1 U20940 ( .A(n17706), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18071) );
  OAI21_X1 U20941 ( .B1(n17933), .B2(n17708), .A(n17707), .ZN(n17709) );
  XNOR2_X1 U20942 ( .A(n17709), .B(n18058), .ZN(n18066) );
  OAI22_X1 U20943 ( .A1(n17938), .A2(n18071), .B1(n17893), .B2(n18066), .ZN(
        n17710) );
  AOI211_X1 U20944 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17717), .A(
        n17711), .B(n17710), .ZN(n17712) );
  OAI21_X1 U20945 ( .B1(n18033), .B2(n18067), .A(n17712), .ZN(P3_U2805) );
  NAND2_X1 U20946 ( .A1(n17713), .A2(n18169), .ZN(n18074) );
  AOI22_X1 U20947 ( .A1(n17889), .A2(n18076), .B1(n18000), .B2(n18074), .ZN(
        n17736) );
  INV_X1 U20948 ( .A(n17714), .ZN(n17715) );
  OAI22_X1 U20949 ( .A1(n18339), .A2(n18929), .B1(n17857), .B2(n17715), .ZN(
        n17716) );
  AOI221_X1 U20950 ( .B1(n17719), .B2(n17718), .C1(n17717), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17716), .ZN(n17724) );
  OAI21_X1 U20951 ( .B1(n17721), .B2(n17725), .A(n17720), .ZN(n18073) );
  NOR2_X1 U20952 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17722), .ZN(
        n18072) );
  AOI22_X1 U20953 ( .A1(n17934), .A2(n18073), .B1(n9847), .B2(n18072), .ZN(
        n17723) );
  OAI211_X1 U20954 ( .C1(n17736), .C2(n17725), .A(n17724), .B(n17723), .ZN(
        P3_U2806) );
  NAND2_X1 U20955 ( .A1(n17726), .A2(n9847), .ZN(n17737) );
  OAI22_X1 U20956 ( .A1(n17727), .A2(n17740), .B1(n17933), .B2(n18096), .ZN(
        n17728) );
  NOR2_X1 U20957 ( .A1(n17728), .A2(n17770), .ZN(n17729) );
  XNOR2_X1 U20958 ( .A(n17729), .B(n18079), .ZN(n18092) );
  NOR2_X1 U20959 ( .A1(n18339), .A2(n18928), .ZN(n18091) );
  NOR2_X1 U20960 ( .A1(n17872), .A2(n17692), .ZN(n17733) );
  AOI21_X1 U20961 ( .B1(n18745), .B2(n9973), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17730) );
  OAI22_X1 U20962 ( .A1(n17733), .A2(n17732), .B1(n17731), .B2(n17730), .ZN(
        n17734) );
  AOI211_X1 U20963 ( .C1(n18092), .C2(n17934), .A(n18091), .B(n17734), .ZN(
        n17735) );
  OAI221_X1 U20964 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17737), 
        .C1(n18079), .C2(n17736), .A(n17735), .ZN(P3_U2807) );
  INV_X1 U20965 ( .A(n17738), .ZN(n17813) );
  INV_X1 U20966 ( .A(n17770), .ZN(n17739) );
  OAI221_X1 U20967 ( .B1(n17740), .B2(n18100), .C1(n17740), .C2(n17813), .A(
        n17739), .ZN(n17741) );
  XNOR2_X1 U20968 ( .A(n18096), .B(n17741), .ZN(n18109) );
  NOR2_X1 U20969 ( .A1(n18172), .A2(n17938), .ZN(n17837) );
  NOR2_X1 U20970 ( .A1(n18169), .A2(n18033), .ZN(n17831) );
  NOR2_X1 U20971 ( .A1(n17837), .A2(n17831), .ZN(n17821) );
  OAI21_X1 U20972 ( .B1(n18100), .B2(n17769), .A(n17821), .ZN(n17761) );
  OAI21_X1 U20973 ( .B1(n17742), .B2(n18029), .A(n18028), .ZN(n17743) );
  AOI21_X1 U20974 ( .B1(n17923), .B2(n17745), .A(n17743), .ZN(n17766) );
  OAI21_X1 U20975 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17802), .A(
        n17766), .ZN(n17754) );
  AOI22_X1 U20976 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17754), .B1(
        n17872), .B2(n17744), .ZN(n17748) );
  NOR2_X1 U20977 ( .A1(n17777), .A2(n17745), .ZN(n17756) );
  OAI211_X1 U20978 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17756), .B(n17746), .ZN(n17747) );
  OAI211_X1 U20979 ( .C1(n18925), .C2(n18339), .A(n17748), .B(n17747), .ZN(
        n17749) );
  AOI21_X1 U20980 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17761), .A(
        n17749), .ZN(n17751) );
  NAND3_X1 U20981 ( .A1(n18100), .A2(n9847), .A3(n18096), .ZN(n17750) );
  OAI211_X1 U20982 ( .C1(n17893), .C2(n18109), .A(n17751), .B(n17750), .ZN(
        P3_U2808) );
  INV_X1 U20983 ( .A(n18115), .ZN(n17759) );
  OR2_X1 U20984 ( .A1(n17759), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18119) );
  NAND2_X1 U20985 ( .A1(n18113), .A2(n9847), .ZN(n17788) );
  INV_X1 U20986 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17755) );
  INV_X1 U20987 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18924) );
  OAI22_X1 U20988 ( .A1(n18339), .A2(n18924), .B1(n17857), .B2(n17752), .ZN(
        n17753) );
  AOI221_X1 U20989 ( .B1(n17756), .B2(n17755), .C1(n17754), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17753), .ZN(n17763) );
  NAND3_X1 U20990 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17757), .ZN(n17782) );
  OAI22_X1 U20991 ( .A1(n17759), .A2(n17782), .B1(n10312), .B2(n17758), .ZN(
        n17760) );
  XOR2_X1 U20992 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17760), .Z(
        n18111) );
  AOI22_X1 U20993 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17761), .B1(
        n17934), .B2(n18111), .ZN(n17762) );
  OAI211_X1 U20994 ( .C1(n18119), .C2(n17788), .A(n17763), .B(n17762), .ZN(
        P3_U2809) );
  NAND2_X1 U20995 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17771), .ZN(
        n18128) );
  AOI21_X1 U20996 ( .B1(n18745), .B2(n17764), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17765) );
  OAI22_X1 U20997 ( .A1(n17766), .A2(n17765), .B1(n18339), .B2(n18921), .ZN(
        n17767) );
  AOI221_X1 U20998 ( .B1(n17872), .B2(n17768), .C1(n17692), .C2(n17768), .A(
        n17767), .ZN(n17774) );
  NOR2_X1 U20999 ( .A1(n18082), .A2(n17783), .ZN(n18124) );
  OAI21_X1 U21000 ( .B1(n17769), .B2(n18124), .A(n17821), .ZN(n17785) );
  AOI221_X1 U21001 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17782), 
        .C1(n17783), .C2(n17794), .A(n17770), .ZN(n17772) );
  XNOR2_X1 U21002 ( .A(n17772), .B(n17771), .ZN(n18120) );
  AOI22_X1 U21003 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17785), .B1(
        n17934), .B2(n18120), .ZN(n17773) );
  OAI211_X1 U21004 ( .C1(n17788), .C2(n18128), .A(n17774), .B(n17773), .ZN(
        P3_U2810) );
  AOI21_X1 U21005 ( .B1(n17923), .B2(n17776), .A(n17998), .ZN(n17804) );
  OAI21_X1 U21006 ( .B1(n17775), .B2(n18029), .A(n17804), .ZN(n17791) );
  NOR2_X1 U21007 ( .A1(n17777), .A2(n17776), .ZN(n17793) );
  OAI211_X1 U21008 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17793), .B(n17778), .ZN(n17779) );
  NAND2_X1 U21009 ( .A1(n18297), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18131) );
  OAI211_X1 U21010 ( .C1(n17857), .C2(n17780), .A(n17779), .B(n18131), .ZN(
        n17781) );
  AOI21_X1 U21011 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17791), .A(
        n17781), .ZN(n17787) );
  OAI21_X1 U21012 ( .B1(n10312), .B2(n17794), .A(n17782), .ZN(n17784) );
  XNOR2_X1 U21013 ( .A(n17784), .B(n17783), .ZN(n18129) );
  AOI22_X1 U21014 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17785), .B1(
        n17934), .B2(n18129), .ZN(n17786) );
  OAI211_X1 U21015 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17788), .A(
        n17787), .B(n17786), .ZN(P3_U2811) );
  NAND2_X1 U21016 ( .A1(n18142), .A2(n17795), .ZN(n18150) );
  INV_X1 U21017 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17792) );
  OAI22_X1 U21018 ( .A1(n18339), .A2(n18917), .B1(n17857), .B2(n17789), .ZN(
        n17790) );
  AOI221_X1 U21019 ( .B1(n17793), .B2(n17792), .C1(n17791), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17790), .ZN(n17799) );
  OAI21_X1 U21020 ( .B1(n18142), .B2(n17800), .A(n17821), .ZN(n17808) );
  OAI21_X1 U21021 ( .B1(n17811), .B2(n17795), .A(n17794), .ZN(n17797) );
  XNOR2_X1 U21022 ( .A(n17797), .B(n17796), .ZN(n18146) );
  AOI22_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17808), .B1(
        n17934), .B2(n18146), .ZN(n17798) );
  OAI211_X1 U21024 ( .C1(n17800), .C2(n18150), .A(n17799), .B(n17798), .ZN(
        P3_U2812) );
  AOI21_X1 U21025 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17801), .A(
        n9948), .ZN(n18158) );
  AOI21_X1 U21026 ( .B1(n17803), .B2(n18745), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17805) );
  NAND2_X1 U21027 ( .A1(n18297), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18156) );
  OAI21_X1 U21028 ( .B1(n17805), .B2(n17804), .A(n18156), .ZN(n17806) );
  AOI21_X1 U21029 ( .B1(n17807), .B2(n17996), .A(n17806), .ZN(n17810) );
  NOR2_X1 U21030 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18164), .ZN(
        n18155) );
  AOI22_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17808), .B1(
        n9847), .B2(n18155), .ZN(n17809) );
  OAI211_X1 U21032 ( .C1(n18158), .C2(n17893), .A(n17810), .B(n17809), .ZN(
        P3_U2813) );
  NAND2_X1 U21033 ( .A1(n17830), .A2(n17909), .ZN(n17827) );
  OAI22_X1 U21034 ( .A1(n17933), .A2(n17813), .B1(n17827), .B2(n18173), .ZN(
        n17814) );
  XNOR2_X1 U21035 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17814), .ZN(
        n18168) );
  AOI21_X1 U21036 ( .B1(n17923), .B2(n17815), .A(n17998), .ZN(n17850) );
  OAI21_X1 U21037 ( .B1(n17816), .B2(n18029), .A(n17850), .ZN(n17833) );
  NOR2_X1 U21038 ( .A1(n18339), .A2(n18913), .ZN(n18163) );
  NAND4_X1 U21039 ( .A1(n17854), .A2(n17852), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(n17851), .ZN(n17835) );
  OAI21_X1 U21040 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17817), .ZN(n17818) );
  OAI22_X1 U21041 ( .A1(n17857), .A2(n17819), .B1(n17835), .B2(n17818), .ZN(
        n17820) );
  AOI211_X1 U21042 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17833), .A(
        n18163), .B(n17820), .ZN(n17825) );
  INV_X1 U21043 ( .A(n17821), .ZN(n17823) );
  AOI22_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17823), .B1(
        n9847), .B2(n18164), .ZN(n17824) );
  OAI211_X1 U21045 ( .C1(n18168), .C2(n17893), .A(n17825), .B(n17824), .ZN(
        P3_U2814) );
  NAND2_X1 U21046 ( .A1(n17866), .A2(n18198), .ZN(n17828) );
  NOR2_X1 U21047 ( .A1(n17933), .A2(n17826), .ZN(n17910) );
  NAND2_X1 U21048 ( .A1(n17904), .A2(n17910), .ZN(n17879) );
  NOR2_X1 U21049 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17879), .ZN(
        n17873) );
  NAND2_X1 U21050 ( .A1(n17873), .A2(n18213), .ZN(n17861) );
  OAI21_X1 U21051 ( .B1(n17828), .B2(n17861), .A(n17827), .ZN(n17829) );
  XNOR2_X1 U21052 ( .A(n17829), .B(n18173), .ZN(n18179) );
  INV_X1 U21053 ( .A(n17830), .ZN(n18171) );
  OAI21_X1 U21054 ( .B1(n17887), .B2(n18171), .A(n18173), .ZN(n18177) );
  AOI22_X1 U21055 ( .A1(n17934), .A2(n18179), .B1(n17831), .B2(n18177), .ZN(
        n17840) );
  NAND2_X1 U21056 ( .A1(n18174), .A2(n18173), .ZN(n17838) );
  AOI22_X1 U21057 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17833), .B1(
        n17872), .B2(n17832), .ZN(n17834) );
  NAND2_X1 U21058 ( .A1(n18297), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18180) );
  OAI211_X1 U21059 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17835), .A(
        n17834), .B(n18180), .ZN(n17836) );
  AOI21_X1 U21060 ( .B1(n17838), .B2(n17837), .A(n17836), .ZN(n17839) );
  NAND2_X1 U21061 ( .A1(n17840), .A2(n17839), .ZN(P3_U2815) );
  NAND2_X1 U21062 ( .A1(n18745), .A2(n9967), .ZN(n17961) );
  NOR2_X1 U21063 ( .A1(n17968), .A2(n17961), .ZN(n17942) );
  NAND2_X1 U21064 ( .A1(n17841), .A2(n17942), .ZN(n17896) );
  NOR2_X1 U21065 ( .A1(n17883), .A2(n17896), .ZN(n17882) );
  AOI21_X1 U21066 ( .B1(n17852), .B2(n17882), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17849) );
  AOI22_X1 U21067 ( .A1(n18357), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17842), 
        .B2(n17996), .ZN(n17848) );
  NAND2_X1 U21068 ( .A1(n18183), .A2(n18224), .ZN(n18202) );
  NOR2_X1 U21069 ( .A1(n17887), .A2(n18171), .ZN(n17843) );
  AOI221_X1 U21070 ( .B1(n17866), .B2(n18198), .C1(n18202), .C2(n18198), .A(
        n17843), .ZN(n18195) );
  NAND2_X1 U21071 ( .A1(n18183), .A2(n17909), .ZN(n17862) );
  AOI22_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17862), .B1(
        n17861), .B2(n17866), .ZN(n17844) );
  XNOR2_X1 U21073 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17844), .ZN(
        n18193) );
  OAI21_X1 U21074 ( .B1(n17845), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18174), .ZN(n18192) );
  OAI22_X1 U21075 ( .A1(n18193), .A2(n17893), .B1(n17938), .B2(n18192), .ZN(
        n17846) );
  AOI21_X1 U21076 ( .B1(n18000), .B2(n18195), .A(n17846), .ZN(n17847) );
  OAI211_X1 U21077 ( .C1(n17850), .C2(n17849), .A(n17848), .B(n17847), .ZN(
        P3_U2816) );
  AOI22_X1 U21078 ( .A1(n17889), .A2(n18200), .B1(n18000), .B2(n18202), .ZN(
        n17878) );
  NAND2_X1 U21079 ( .A1(n17854), .A2(n17851), .ZN(n17869) );
  AOI211_X1 U21080 ( .C1(n17868), .C2(n17858), .A(n17852), .B(n17869), .ZN(
        n17860) );
  OAI22_X1 U21081 ( .A1(n17854), .A2(n17989), .B1(n17853), .B2(n18029), .ZN(
        n17855) );
  NOR2_X1 U21082 ( .A1(n17998), .A2(n17855), .ZN(n17867) );
  OAI22_X1 U21083 ( .A1(n17867), .A2(n17858), .B1(n17857), .B2(n17856), .ZN(
        n17859) );
  AOI211_X1 U21084 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18357), .A(n17860), 
        .B(n17859), .ZN(n17865) );
  NAND2_X1 U21085 ( .A1(n17862), .A2(n17861), .ZN(n17863) );
  XNOR2_X1 U21086 ( .A(n17863), .B(n17866), .ZN(n18209) );
  NOR2_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18213), .ZN(
        n18208) );
  NOR2_X1 U21088 ( .A1(n17920), .A2(n18207), .ZN(n17875) );
  AOI22_X1 U21089 ( .A1(n17934), .A2(n18209), .B1(n18208), .B2(n17875), .ZN(
        n17864) );
  OAI211_X1 U21090 ( .C1(n17878), .C2(n17866), .A(n17865), .B(n17864), .ZN(
        P3_U2817) );
  NAND2_X1 U21091 ( .A1(n18297), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18218) );
  OAI221_X1 U21092 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17869), .C1(
        n17868), .C2(n17867), .A(n18218), .ZN(n17870) );
  AOI21_X1 U21093 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n17877) );
  NAND2_X1 U21094 ( .A1(n18230), .A2(n17909), .ZN(n17880) );
  INV_X1 U21095 ( .A(n17880), .ZN(n17898) );
  AOI21_X1 U21096 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n17898), .A(
        n17873), .ZN(n17874) );
  XNOR2_X1 U21097 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17874), .ZN(
        n18217) );
  AOI22_X1 U21098 ( .A1(n17934), .A2(n18217), .B1(n17875), .B2(n18213), .ZN(
        n17876) );
  OAI211_X1 U21099 ( .C1(n17878), .C2(n18213), .A(n17877), .B(n17876), .ZN(
        P3_U2818) );
  NAND2_X1 U21100 ( .A1(n17880), .A2(n17879), .ZN(n17881) );
  XNOR2_X1 U21101 ( .A(n17881), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18236) );
  INV_X1 U21102 ( .A(n17953), .ZN(n18023) );
  AOI211_X1 U21103 ( .C1(n17896), .C2(n17883), .A(n18023), .B(n17882), .ZN(
        n17885) );
  NOR2_X1 U21104 ( .A1(n18339), .A2(n18903), .ZN(n17884) );
  AOI211_X1 U21105 ( .C1(n17886), .C2(n17996), .A(n17885), .B(n17884), .ZN(
        n17892) );
  AOI22_X1 U21106 ( .A1(n17889), .A2(n17888), .B1(n18000), .B2(n17887), .ZN(
        n17919) );
  OAI21_X1 U21107 ( .B1(n18230), .B2(n17920), .A(n17919), .ZN(n17890) );
  INV_X1 U21108 ( .A(n18230), .ZN(n17902) );
  NOR2_X1 U21109 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17902), .ZN(
        n18222) );
  INV_X1 U21110 ( .A(n17920), .ZN(n17901) );
  AOI22_X1 U21111 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17890), .B1(
        n18222), .B2(n17901), .ZN(n17891) );
  OAI211_X1 U21112 ( .C1(n18236), .C2(n17893), .A(n17892), .B(n17891), .ZN(
        P3_U2819) );
  NAND4_X1 U21113 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(n17942), .ZN(n17913) );
  OAI21_X1 U21114 ( .B1(n18023), .B2(n17894), .A(n17913), .ZN(n17895) );
  AOI22_X1 U21115 ( .A1(n18357), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17896), 
        .B2(n17895), .ZN(n17907) );
  NOR3_X1 U21116 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18237), .ZN(n17899) );
  AOI221_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17909), .C1(
        n18248), .C2(n17910), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17897) );
  AOI211_X1 U21118 ( .C1(n17900), .C2(n17899), .A(n17898), .B(n17897), .ZN(
        n18238) );
  NAND2_X1 U21119 ( .A1(n17902), .A2(n17901), .ZN(n17903) );
  OAI22_X1 U21120 ( .A1(n17904), .A2(n17903), .B1(n17919), .B2(n18237), .ZN(
        n17905) );
  AOI21_X1 U21121 ( .B1(n17934), .B2(n18238), .A(n17905), .ZN(n17906) );
  OAI211_X1 U21122 ( .C1(n18025), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2820) );
  NOR2_X1 U21123 ( .A1(n17910), .A2(n17909), .ZN(n17911) );
  XNOR2_X1 U21124 ( .A(n17911), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18252) );
  NAND2_X1 U21125 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17927) );
  INV_X1 U21126 ( .A(n17942), .ZN(n17912) );
  NOR2_X1 U21127 ( .A1(n17927), .A2(n17912), .ZN(n17914) );
  OAI211_X1 U21128 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17953), .B(n17913), .ZN(n17915) );
  NAND2_X1 U21129 ( .A1(n18297), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18254) );
  OAI211_X1 U21130 ( .C1(n18025), .C2(n17916), .A(n17915), .B(n18254), .ZN(
        n17917) );
  AOI21_X1 U21131 ( .B1(n17934), .B2(n18252), .A(n17917), .ZN(n17918) );
  OAI221_X1 U21132 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17920), .C1(
        n18248), .C2(n17919), .A(n17918), .ZN(P3_U2821) );
  AOI21_X1 U21133 ( .B1(n17924), .B2(n17921), .A(n18685), .ZN(n17928) );
  NOR2_X1 U21134 ( .A1(n18339), .A2(n18898), .ZN(n18267) );
  AOI21_X1 U21135 ( .B1(n17923), .B2(n17922), .A(n17998), .ZN(n17939) );
  OAI22_X1 U21136 ( .A1(n18025), .A2(n17925), .B1(n17939), .B2(n17924), .ZN(
        n17926) );
  AOI211_X1 U21137 ( .C1(n17928), .C2(n17927), .A(n18267), .B(n17926), .ZN(
        n17936) );
  AOI21_X1 U21138 ( .B1(n17931), .B2(n17930), .A(n17929), .ZN(n18268) );
  AOI21_X1 U21139 ( .B1(n17933), .B2(n17937), .A(n17932), .ZN(n18273) );
  AOI22_X1 U21140 ( .A1(n18000), .A2(n18268), .B1(n17934), .B2(n18273), .ZN(
        n17935) );
  OAI211_X1 U21141 ( .C1(n17938), .C2(n17937), .A(n17936), .B(n17935), .ZN(
        P3_U2822) );
  INV_X1 U21142 ( .A(n17939), .ZN(n17940) );
  NOR2_X1 U21143 ( .A1(n18339), .A2(n18895), .ZN(n18276) );
  AOI221_X1 U21144 ( .B1(n17942), .B2(n17941), .C1(n17940), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18276), .ZN(n17951) );
  AOI21_X1 U21145 ( .B1(n17945), .B2(n17944), .A(n17943), .ZN(n18277) );
  OAI21_X1 U21146 ( .B1(n17948), .B2(n17947), .A(n17946), .ZN(n17949) );
  XNOR2_X1 U21147 ( .A(n17949), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18278) );
  AOI22_X1 U21148 ( .A1(n18021), .A2(n18277), .B1(n18000), .B2(n18278), .ZN(
        n17950) );
  OAI211_X1 U21149 ( .C1(n18025), .C2(n17952), .A(n17951), .B(n17950), .ZN(
        P3_U2823) );
  NAND2_X1 U21150 ( .A1(n17953), .A2(n17961), .ZN(n17975) );
  AOI22_X1 U21151 ( .A1(n17955), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18285), .B2(n17954), .ZN(n17960) );
  AOI22_X1 U21152 ( .A1(n17958), .A2(n17969), .B1(n17957), .B2(n17956), .ZN(
        n17959) );
  XNOR2_X1 U21153 ( .A(n17960), .B(n17959), .ZN(n18290) );
  OAI22_X1 U21154 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17961), .B1(
        n18290), .B2(n18033), .ZN(n17962) );
  AOI21_X1 U21155 ( .B1(n18357), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17962), .ZN(
        n17967) );
  AOI21_X1 U21156 ( .B1(n9962), .B2(n17964), .A(n17963), .ZN(n18288) );
  AOI22_X1 U21157 ( .A1(n18021), .A2(n18288), .B1(n17965), .B2(n17996), .ZN(
        n17966) );
  OAI211_X1 U21158 ( .C1(n17968), .C2(n17975), .A(n17967), .B(n17966), .ZN(
        P3_U2824) );
  OAI21_X1 U21159 ( .B1(n17971), .B2(n17970), .A(n17969), .ZN(n18300) );
  AOI21_X1 U21160 ( .B1(n17974), .B2(n17973), .A(n17972), .ZN(n18296) );
  AOI22_X1 U21161 ( .A1(n18021), .A2(n18296), .B1(n18297), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17981) );
  AOI221_X1 U21162 ( .B1(n17998), .B2(n17977), .C1(n17976), .C2(n17977), .A(
        n17975), .ZN(n17978) );
  AOI21_X1 U21163 ( .B1(n17979), .B2(n17996), .A(n17978), .ZN(n17980) );
  OAI211_X1 U21164 ( .C1(n18033), .C2(n18300), .A(n17981), .B(n17980), .ZN(
        P3_U2825) );
  OAI21_X1 U21165 ( .B1(n17984), .B2(n17983), .A(n17982), .ZN(n18310) );
  OAI22_X1 U21166 ( .A1(n18033), .A2(n18310), .B1(n18685), .B2(n17985), .ZN(
        n17986) );
  AOI21_X1 U21167 ( .B1(n18357), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17986), .ZN(
        n17992) );
  AOI21_X1 U21168 ( .B1(n9968), .B2(n17988), .A(n17987), .ZN(n18301) );
  OAI21_X1 U21169 ( .B1(n17990), .B2(n17989), .A(n18028), .ZN(n17999) );
  AOI22_X1 U21170 ( .A1(n18021), .A2(n18301), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17999), .ZN(n17991) );
  OAI211_X1 U21171 ( .C1(n18025), .C2(n17993), .A(n17992), .B(n17991), .ZN(
        P3_U2826) );
  AOI21_X1 U21172 ( .B1(n18317), .B2(n17995), .A(n17994), .ZN(n18320) );
  AOI22_X1 U21173 ( .A1(n18021), .A2(n18320), .B1(n17997), .B2(n17996), .ZN(
        n18003) );
  NOR2_X1 U21174 ( .A1(n17998), .A2(n18008), .ZN(n18007) );
  OAI21_X1 U21175 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18007), .A(
        n17999), .ZN(n18002) );
  NAND2_X1 U21176 ( .A1(n18297), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18316) );
  OAI211_X1 U21177 ( .C1(n18313), .C2(n18312), .A(n18000), .B(n18311), .ZN(
        n18001) );
  NAND4_X1 U21178 ( .A1(n18003), .A2(n18002), .A3(n18316), .A4(n18001), .ZN(
        P3_U2827) );
  AOI21_X1 U21179 ( .B1(n18006), .B2(n18005), .A(n18004), .ZN(n18323) );
  AOI21_X1 U21180 ( .B1(n18685), .B2(n18008), .A(n18007), .ZN(n18013) );
  OAI21_X1 U21181 ( .B1(n18011), .B2(n18010), .A(n18009), .ZN(n18333) );
  INV_X1 U21182 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18885) );
  OAI22_X1 U21183 ( .A1(n18033), .A2(n18333), .B1(n18339), .B2(n18885), .ZN(
        n18012) );
  AOI211_X1 U21184 ( .C1(n18323), .C2(n18021), .A(n18013), .B(n18012), .ZN(
        n18014) );
  OAI21_X1 U21185 ( .B1(n18025), .B2(n18015), .A(n18014), .ZN(P3_U2828) );
  INV_X1 U21186 ( .A(n18019), .ZN(n18017) );
  AOI21_X1 U21187 ( .B1(n18017), .B2(n18027), .A(n18016), .ZN(n18344) );
  AOI21_X1 U21188 ( .B1(n18019), .B2(n18026), .A(n18018), .ZN(n18350) );
  OAI22_X1 U21189 ( .A1(n18350), .A2(n18033), .B1(n18339), .B2(n18990), .ZN(
        n18020) );
  AOI21_X1 U21190 ( .B1(n18021), .B2(n18344), .A(n18020), .ZN(n18022) );
  OAI221_X1 U21191 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18025), .C1(
        n18024), .C2(n18023), .A(n18022), .ZN(P3_U2829) );
  NAND2_X1 U21192 ( .A1(n18027), .A2(n18026), .ZN(n18360) );
  INV_X1 U21193 ( .A(n18360), .ZN(n18034) );
  NAND3_X1 U21194 ( .A1(n18970), .A2(n18029), .A3(n18028), .ZN(n18030) );
  AOI22_X1 U21195 ( .A1(n18357), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18030), .ZN(n18031) );
  OAI221_X1 U21196 ( .B1(n18034), .B2(n18033), .C1(n18360), .C2(n18032), .A(
        n18031), .ZN(P3_U2830) );
  NAND2_X1 U21197 ( .A1(n18353), .A2(n18818), .ZN(n18145) );
  AOI21_X1 U21198 ( .B1(n18036), .B2(n18145), .A(n18035), .ZN(n18038) );
  NAND2_X1 U21199 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18037) );
  NAND2_X1 U21200 ( .A1(n18813), .A2(n18985), .ZN(n18325) );
  NAND4_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18100), .A3(
        n18138), .A4(n18325), .ZN(n18075) );
  OAI21_X1 U21202 ( .B1(n18037), .B2(n18075), .A(n18145), .ZN(n18056) );
  OAI211_X1 U21203 ( .C1(n18039), .C2(n18332), .A(n18038), .B(n18056), .ZN(
        n18040) );
  AOI21_X1 U21204 ( .B1(n18201), .B2(n18041), .A(n18040), .ZN(n18049) );
  NAND2_X1 U21205 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18334), .ZN(
        n18042) );
  AOI22_X1 U21206 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18049), .B1(
        n18043), .B2(n18042), .ZN(n18044) );
  AOI21_X1 U21207 ( .B1(n18346), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18044), .ZN(n18046) );
  OAI211_X1 U21208 ( .C1(n18047), .C2(n18270), .A(n18046), .B(n18045), .ZN(
        P3_U2835) );
  INV_X1 U21209 ( .A(n18110), .ZN(n18054) );
  AOI211_X1 U21210 ( .C1(n18334), .C2(n18049), .A(n18357), .B(n18048), .ZN(
        n18050) );
  AOI21_X1 U21211 ( .B1(n18253), .B2(n18051), .A(n18050), .ZN(n18053) );
  NAND2_X1 U21212 ( .A1(n18297), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18052) );
  OAI211_X1 U21213 ( .C1(n18055), .C2(n18054), .A(n18053), .B(n18052), .ZN(
        P3_U2836) );
  INV_X1 U21214 ( .A(n18056), .ZN(n18063) );
  AOI22_X1 U21215 ( .A1(n18057), .A2(n18081), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18833), .ZN(n18062) );
  OAI21_X1 U21216 ( .B1(n18060), .B2(n18059), .A(n18058), .ZN(n18061) );
  OAI211_X1 U21217 ( .C1(n18063), .C2(n18062), .A(n18334), .B(n18061), .ZN(
        n18064) );
  NAND2_X1 U21218 ( .A1(n18065), .A2(n18064), .ZN(n18069) );
  OAI22_X1 U21219 ( .A1(n18349), .A2(n18067), .B1(n18270), .B2(n18066), .ZN(
        n18068) );
  AOI211_X1 U21220 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18346), .A(
        n18069), .B(n18068), .ZN(n18070) );
  OAI21_X1 U21221 ( .B1(n18272), .B2(n18071), .A(n18070), .ZN(P3_U2837) );
  AOI22_X1 U21222 ( .A1(n18253), .A2(n18073), .B1(n18110), .B2(n18072), .ZN(
        n18087) );
  INV_X1 U21223 ( .A(n18074), .ZN(n18078) );
  AOI22_X1 U21224 ( .A1(n18201), .A2(n18076), .B1(n18145), .B2(n18075), .ZN(
        n18077) );
  INV_X1 U21225 ( .A(n18346), .ZN(n18352) );
  OAI211_X1 U21226 ( .C1(n18078), .C2(n18332), .A(n18077), .B(n18352), .ZN(
        n18084) );
  AOI211_X1 U21227 ( .C1(n18804), .C2(n18080), .A(n18079), .B(n18084), .ZN(
        n18083) );
  INV_X1 U21228 ( .A(n18081), .ZN(n18139) );
  OAI21_X1 U21229 ( .B1(n18082), .B2(n18139), .A(n18804), .ZN(n18098) );
  AOI21_X1 U21230 ( .B1(n18083), .B2(n18098), .A(n18357), .ZN(n18089) );
  OAI211_X1 U21231 ( .C1(n18085), .C2(n18084), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18089), .ZN(n18086) );
  OAI211_X1 U21232 ( .C1(n18929), .C2(n18339), .A(n18087), .B(n18086), .ZN(
        P3_U2838) );
  NOR3_X1 U21233 ( .A1(n18346), .A2(n18097), .A3(n18088), .ZN(n18090) );
  OAI21_X1 U21234 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18090), .A(
        n18089), .ZN(n18094) );
  AOI21_X1 U21235 ( .B1(n18092), .B2(n18253), .A(n18091), .ZN(n18093) );
  NAND2_X1 U21236 ( .A1(n18094), .A2(n18093), .ZN(P3_U2839) );
  AOI221_X1 U21237 ( .B1(n18097), .B2(n18096), .C1(n18095), .C2(n18096), .A(
        n18351), .ZN(n18106) );
  OAI221_X1 U21238 ( .B1(n18353), .B2(n18138), .C1(n18353), .C2(n18124), .A(
        n18098), .ZN(n18121) );
  NOR2_X1 U21239 ( .A1(n18802), .A2(n18201), .ZN(n18229) );
  OAI22_X1 U21240 ( .A1(n18353), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18100), .B2(n18229), .ZN(n18099) );
  NOR2_X1 U21241 ( .A1(n18121), .A2(n18099), .ZN(n18114) );
  NAND2_X1 U21242 ( .A1(n18100), .A2(n18138), .ZN(n18103) );
  OAI22_X1 U21243 ( .A1(n18172), .A2(n18225), .B1(n18169), .B2(n18332), .ZN(
        n18112) );
  OAI22_X1 U21244 ( .A1(n18353), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18101), .B2(n18833), .ZN(n18102) );
  AOI211_X1 U21245 ( .C1(n18813), .C2(n18103), .A(n18112), .B(n18102), .ZN(
        n18104) );
  NAND4_X1 U21246 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18114), .A3(
        n18104), .A4(n18325), .ZN(n18105) );
  AOI22_X1 U21247 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18346), .B1(
        n18106), .B2(n18105), .ZN(n18108) );
  NAND2_X1 U21248 ( .A1(n18297), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18107) );
  OAI211_X1 U21249 ( .C1(n18109), .C2(n18270), .A(n18108), .B(n18107), .ZN(
        P3_U2840) );
  NAND2_X1 U21250 ( .A1(n18113), .A2(n18110), .ZN(n18133) );
  AOI22_X1 U21251 ( .A1(n18357), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18253), 
        .B2(n18111), .ZN(n18118) );
  NOR2_X1 U21252 ( .A1(n18351), .A2(n18112), .ZN(n18162) );
  OAI221_X1 U21253 ( .B1(n18818), .B2(n18113), .C1(n18818), .C2(n18159), .A(
        n18162), .ZN(n18122) );
  NOR2_X1 U21254 ( .A1(n18804), .A2(n18813), .ZN(n18345) );
  OAI21_X1 U21255 ( .B1(n18115), .B2(n18345), .A(n18114), .ZN(n18116) );
  OAI211_X1 U21256 ( .C1(n18122), .C2(n18116), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18339), .ZN(n18117) );
  OAI211_X1 U21257 ( .C1(n18133), .C2(n18119), .A(n18118), .B(n18117), .ZN(
        P3_U2841) );
  AOI22_X1 U21258 ( .A1(n18357), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18253), 
        .B2(n18120), .ZN(n18127) );
  NOR2_X1 U21259 ( .A1(n18122), .A2(n18121), .ZN(n18123) );
  AOI221_X1 U21260 ( .B1(n18124), .B2(n18123), .C1(n18229), .C2(n18123), .A(
        n18357), .ZN(n18130) );
  NOR3_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18345), .A3(
        n18856), .ZN(n18125) );
  OAI21_X1 U21262 ( .B1(n18130), .B2(n18125), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18126) );
  OAI211_X1 U21263 ( .C1(n18128), .C2(n18133), .A(n18127), .B(n18126), .ZN(
        P3_U2842) );
  AOI22_X1 U21264 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18130), .B1(
        n18253), .B2(n18129), .ZN(n18132) );
  OAI211_X1 U21265 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18133), .A(
        n18132), .B(n18131), .ZN(P3_U2843) );
  INV_X1 U21266 ( .A(n18327), .ZN(n18302) );
  INV_X1 U21267 ( .A(n18134), .ZN(n18326) );
  AOI22_X1 U21268 ( .A1(n18804), .A2(n18302), .B1(n18326), .B2(n18329), .ZN(
        n18315) );
  NOR2_X1 U21269 ( .A1(n18315), .A2(n18135), .ZN(n18275) );
  NAND2_X1 U21270 ( .A1(n18136), .A2(n18275), .ZN(n18188) );
  AOI21_X1 U21271 ( .B1(n18137), .B2(n18188), .A(n18351), .ZN(n18223) );
  NAND2_X1 U21272 ( .A1(n10202), .A2(n18223), .ZN(n18151) );
  NAND3_X1 U21273 ( .A1(n18138), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18325), .ZN(n18144) );
  OAI21_X1 U21274 ( .B1(n18140), .B2(n18139), .A(n18804), .ZN(n18141) );
  OAI211_X1 U21275 ( .C1(n18142), .C2(n18229), .A(n18162), .B(n18141), .ZN(
        n18143) );
  AOI21_X1 U21276 ( .B1(n18145), .B2(n18144), .A(n18143), .ZN(n18153) );
  INV_X1 U21277 ( .A(n18145), .ZN(n18324) );
  AOI221_X1 U21278 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18153), 
        .C1(n18324), .C2(n18153), .A(n18357), .ZN(n18147) );
  AOI22_X1 U21279 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18147), .B1(
        n18253), .B2(n18146), .ZN(n18149) );
  NAND2_X1 U21280 ( .A1(n18297), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18148) );
  OAI211_X1 U21281 ( .C1(n18150), .C2(n18151), .A(n18149), .B(n18148), .ZN(
        P3_U2844) );
  INV_X1 U21282 ( .A(n18151), .ZN(n18165) );
  NOR3_X1 U21283 ( .A1(n18357), .A2(n18153), .A3(n18152), .ZN(n18154) );
  AOI21_X1 U21284 ( .B1(n18155), .B2(n18165), .A(n18154), .ZN(n18157) );
  OAI211_X1 U21285 ( .C1(n18158), .C2(n18270), .A(n18157), .B(n18156), .ZN(
        P3_U2845) );
  AOI21_X1 U21286 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18818), .A(
        n18159), .ZN(n18161) );
  NAND2_X1 U21287 ( .A1(n18804), .A2(n18184), .ZN(n18228) );
  INV_X1 U21288 ( .A(n18353), .ZN(n18821) );
  NAND2_X1 U21289 ( .A1(n18821), .A2(n18160), .ZN(n18239) );
  NAND2_X1 U21290 ( .A1(n18228), .A2(n18239), .ZN(n18247) );
  AOI211_X1 U21291 ( .C1(n18204), .C2(n18171), .A(n18161), .B(n18247), .ZN(
        n18170) );
  AOI221_X1 U21292 ( .B1(n18261), .B2(n18162), .C1(n18170), .C2(n18162), .A(
        n18357), .ZN(n18166) );
  AOI221_X1 U21293 ( .B1(n18166), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .C1(n18165), .C2(n18164), .A(n18163), .ZN(n18167) );
  OAI21_X1 U21294 ( .B1(n18168), .B2(n18270), .A(n18167), .ZN(P3_U2846) );
  NOR2_X1 U21295 ( .A1(n18169), .A2(n18332), .ZN(n18178) );
  AOI221_X1 U21296 ( .B1(n18171), .B2(n18173), .C1(n18188), .C2(n18173), .A(
        n18170), .ZN(n18176) );
  AOI211_X1 U21297 ( .C1(n18174), .C2(n18173), .A(n18172), .B(n18225), .ZN(
        n18175) );
  AOI211_X1 U21298 ( .C1(n18178), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        n18182) );
  AOI22_X1 U21299 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18346), .B1(
        n18253), .B2(n18179), .ZN(n18181) );
  OAI211_X1 U21300 ( .C1(n18182), .C2(n18351), .A(n18181), .B(n18180), .ZN(
        P3_U2847) );
  INV_X1 U21301 ( .A(n18183), .ZN(n18212) );
  OAI21_X1 U21302 ( .B1(n18212), .B2(n18184), .A(n18804), .ZN(n18185) );
  OAI211_X1 U21303 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18345), .A(
        n18185), .B(n18239), .ZN(n18186) );
  AOI211_X1 U21304 ( .C1(n18821), .C2(n18189), .A(n18198), .B(n18186), .ZN(
        n18187) );
  OAI21_X1 U21305 ( .B1(n18212), .B2(n18246), .A(n18813), .ZN(n18205) );
  AOI21_X1 U21306 ( .B1(n18187), .B2(n18205), .A(n18351), .ZN(n18191) );
  OAI21_X1 U21307 ( .B1(n18189), .B2(n18188), .A(n18198), .ZN(n18190) );
  AOI22_X1 U21308 ( .A1(n18357), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18191), 
        .B2(n18190), .ZN(n18197) );
  OAI22_X1 U21309 ( .A1(n18193), .A2(n18270), .B1(n18272), .B2(n18192), .ZN(
        n18194) );
  AOI21_X1 U21310 ( .B1(n18356), .B2(n18195), .A(n18194), .ZN(n18196) );
  OAI211_X1 U21311 ( .C1(n18198), .C2(n18352), .A(n18197), .B(n18196), .ZN(
        P3_U2848) );
  INV_X1 U21312 ( .A(n18239), .ZN(n18199) );
  AOI21_X1 U21313 ( .B1(n18204), .B2(n18207), .A(n18199), .ZN(n18232) );
  AOI22_X1 U21314 ( .A1(n18802), .A2(n18202), .B1(n18201), .B2(n18200), .ZN(
        n18203) );
  NAND3_X1 U21315 ( .A1(n18232), .A2(n18203), .A3(n18228), .ZN(n18214) );
  INV_X1 U21316 ( .A(n18204), .ZN(n18241) );
  OAI211_X1 U21317 ( .C1(n18241), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18334), .B(n18205), .ZN(n18206) );
  OAI21_X1 U21318 ( .B1(n18214), .B2(n18206), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18211) );
  INV_X1 U21319 ( .A(n18223), .ZN(n18256) );
  NOR2_X1 U21320 ( .A1(n18207), .A2(n18256), .ZN(n18216) );
  AOI22_X1 U21321 ( .A1(n18253), .A2(n18209), .B1(n18208), .B2(n18216), .ZN(
        n18210) );
  OAI221_X1 U21322 ( .B1(n18357), .B2(n18211), .C1(n18339), .C2(n18907), .A(
        n18210), .ZN(P3_U2849) );
  OR2_X1 U21323 ( .A1(n18212), .A2(n18246), .ZN(n18215) );
  AOI211_X1 U21324 ( .C1(n18215), .C2(n18813), .A(n18214), .B(n18213), .ZN(
        n18221) );
  AOI21_X1 U21325 ( .B1(n18334), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18216), .ZN(n18220) );
  AOI22_X1 U21326 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18346), .B1(
        n18253), .B2(n18217), .ZN(n18219) );
  OAI211_X1 U21327 ( .C1(n18221), .C2(n18220), .A(n18219), .B(n18218), .ZN(
        P3_U2850) );
  AOI22_X1 U21328 ( .A1(n18357), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18223), 
        .B2(n18222), .ZN(n18235) );
  OAI22_X1 U21329 ( .A1(n18226), .A2(n18225), .B1(n18332), .B2(n18224), .ZN(
        n18227) );
  NOR2_X1 U21330 ( .A1(n18346), .A2(n18227), .ZN(n18250) );
  OAI211_X1 U21331 ( .C1(n18230), .C2(n18229), .A(n18250), .B(n18228), .ZN(
        n18231) );
  AOI221_X1 U21332 ( .B1(n18248), .B2(n18813), .C1(n18246), .C2(n18813), .A(
        n18231), .ZN(n18240) );
  OAI211_X1 U21333 ( .C1(n18818), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18232), .B(n18240), .ZN(n18233) );
  NAND3_X1 U21334 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18339), .A3(
        n18233), .ZN(n18234) );
  OAI211_X1 U21335 ( .C1(n18236), .C2(n18270), .A(n18235), .B(n18234), .ZN(
        P3_U2851) );
  NAND2_X1 U21336 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18237), .ZN(
        n18245) );
  AOI22_X1 U21337 ( .A1(n18357), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18253), 
        .B2(n18238), .ZN(n18244) );
  OAI211_X1 U21338 ( .C1(n18241), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18240), .B(n18239), .ZN(n18242) );
  NAND3_X1 U21339 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18339), .A3(
        n18242), .ZN(n18243) );
  OAI211_X1 U21340 ( .C1(n18245), .C2(n18256), .A(n18244), .B(n18243), .ZN(
        P3_U2852) );
  OAI21_X1 U21341 ( .B1(n18813), .B2(n18247), .A(n18246), .ZN(n18249) );
  AOI211_X1 U21342 ( .C1(n18250), .C2(n18249), .A(n18357), .B(n18248), .ZN(
        n18251) );
  AOI21_X1 U21343 ( .B1(n18253), .B2(n18252), .A(n18251), .ZN(n18255) );
  OAI211_X1 U21344 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18256), .A(
        n18255), .B(n18254), .ZN(P3_U2853) );
  INV_X1 U21345 ( .A(n18273), .ZN(n18271) );
  NAND2_X1 U21346 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18257) );
  NOR3_X1 U21347 ( .A1(n18315), .A2(n18351), .A3(n18317), .ZN(n18306) );
  NAND3_X1 U21348 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18306), .ZN(n18286) );
  NOR2_X1 U21349 ( .A1(n18257), .A2(n18286), .ZN(n18265) );
  INV_X1 U21350 ( .A(n18325), .ZN(n18304) );
  OAI22_X1 U21351 ( .A1(n18259), .A2(n18833), .B1(n18258), .B2(n18324), .ZN(
        n18260) );
  NOR2_X1 U21352 ( .A1(n18304), .A2(n18260), .ZN(n18282) );
  OAI211_X1 U21353 ( .C1(n18261), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18282), .ZN(n18274) );
  AOI21_X1 U21354 ( .B1(n18262), .B2(n18274), .A(n18346), .ZN(n18263) );
  INV_X1 U21355 ( .A(n18263), .ZN(n18264) );
  MUX2_X1 U21356 ( .A(n18265), .B(n18264), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n18266) );
  AOI211_X1 U21357 ( .C1(n18268), .C2(n18356), .A(n18267), .B(n18266), .ZN(
        n18269) );
  OAI221_X1 U21358 ( .B1(n18273), .B2(n18272), .C1(n18271), .C2(n18270), .A(
        n18269), .ZN(P3_U2854) );
  OAI221_X1 U21359 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18275), .A(n18274), .ZN(
        n18281) );
  AOI21_X1 U21360 ( .B1(n18346), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18276), .ZN(n18280) );
  AOI22_X1 U21361 ( .A1(n18356), .A2(n18278), .B1(n18343), .B2(n18277), .ZN(
        n18279) );
  OAI211_X1 U21362 ( .C1(n18351), .C2(n18281), .A(n18280), .B(n18279), .ZN(
        P3_U2855) );
  INV_X1 U21363 ( .A(n18282), .ZN(n18283) );
  OAI21_X1 U21364 ( .B1(n18351), .B2(n18283), .A(n18339), .ZN(n18292) );
  NAND2_X1 U21365 ( .A1(n18357), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18284) );
  OAI221_X1 U21366 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18286), .C1(
        n18285), .C2(n18292), .A(n18284), .ZN(n18287) );
  AOI21_X1 U21367 ( .B1(n18343), .B2(n18288), .A(n18287), .ZN(n18289) );
  OAI21_X1 U21368 ( .B1(n18290), .B2(n18349), .A(n18289), .ZN(P3_U2856) );
  INV_X1 U21369 ( .A(n18306), .ZN(n18291) );
  NOR2_X1 U21370 ( .A1(n18305), .A2(n18291), .ZN(n18294) );
  INV_X1 U21371 ( .A(n18292), .ZN(n18293) );
  MUX2_X1 U21372 ( .A(n18294), .B(n18293), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18295) );
  AOI21_X1 U21373 ( .B1(n18343), .B2(n18296), .A(n18295), .ZN(n18299) );
  NAND2_X1 U21374 ( .A1(n18297), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18298) );
  OAI211_X1 U21375 ( .C1(n18300), .C2(n18349), .A(n18299), .B(n18298), .ZN(
        P3_U2857) );
  AOI22_X1 U21376 ( .A1(n18357), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18343), 
        .B2(n18301), .ZN(n18309) );
  OAI22_X1 U21377 ( .A1(n18326), .A2(n18324), .B1(n18833), .B2(n18302), .ZN(
        n18303) );
  NOR3_X1 U21378 ( .A1(n18304), .A2(n18317), .A3(n18303), .ZN(n18314) );
  OAI21_X1 U21379 ( .B1(n18314), .B2(n18340), .A(n18352), .ZN(n18307) );
  AOI22_X1 U21380 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18307), .B1(
        n18306), .B2(n18305), .ZN(n18308) );
  OAI211_X1 U21381 ( .C1(n18349), .C2(n18310), .A(n18309), .B(n18308), .ZN(
        P3_U2858) );
  OAI21_X1 U21382 ( .B1(n18313), .B2(n18312), .A(n18311), .ZN(n18322) );
  AOI211_X1 U21383 ( .C1(n18315), .C2(n18317), .A(n18314), .B(n18351), .ZN(
        n18319) );
  OAI21_X1 U21384 ( .B1(n18352), .B2(n18317), .A(n18316), .ZN(n18318) );
  AOI211_X1 U21385 ( .C1(n18320), .C2(n18343), .A(n18319), .B(n18318), .ZN(
        n18321) );
  OAI21_X1 U21386 ( .B1(n18349), .B2(n18322), .A(n18321), .ZN(P3_U2859) );
  AOI22_X1 U21387 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18346), .B1(
        n18343), .B2(n18323), .ZN(n18338) );
  AOI211_X1 U21388 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18325), .A(
        n18324), .B(n18328), .ZN(n18336) );
  OAI221_X1 U21389 ( .B1(n18327), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n18327), .C2(n18326), .A(n18804), .ZN(n18331) );
  NAND3_X1 U21390 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18329), .A3(
        n18328), .ZN(n18330) );
  OAI211_X1 U21391 ( .C1(n18333), .C2(n18332), .A(n18331), .B(n18330), .ZN(
        n18335) );
  OAI21_X1 U21392 ( .B1(n18336), .B2(n18335), .A(n18334), .ZN(n18337) );
  OAI211_X1 U21393 ( .C1(n18885), .C2(n18339), .A(n18338), .B(n18337), .ZN(
        P3_U2860) );
  NOR2_X1 U21394 ( .A1(n18339), .A2(n18990), .ZN(n18342) );
  AOI211_X1 U21395 ( .C1(n18353), .C2(n18985), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18340), .ZN(n18341) );
  AOI211_X1 U21396 ( .C1(n18344), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        n18348) );
  NOR3_X1 U21397 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18345), .A3(
        n18351), .ZN(n18355) );
  OAI21_X1 U21398 ( .B1(n18346), .B2(n18355), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18347) );
  OAI211_X1 U21399 ( .C1(n18350), .C2(n18349), .A(n18348), .B(n18347), .ZN(
        P3_U2861) );
  AOI221_X1 U21400 ( .B1(n18353), .B2(n18352), .C1(n18351), .C2(n18352), .A(
        n18985), .ZN(n18354) );
  AOI211_X1 U21401 ( .C1(n18356), .C2(n18360), .A(n18355), .B(n18354), .ZN(
        n18359) );
  NAND2_X1 U21402 ( .A1(n18357), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18358) );
  OAI211_X1 U21403 ( .C1(n18361), .C2(n18360), .A(n18359), .B(n18358), .ZN(
        P3_U2862) );
  OAI211_X1 U21404 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18362), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18854)
         );
  INV_X1 U21405 ( .A(n18854), .ZN(n18363) );
  OAI21_X1 U21406 ( .B1(n18363), .B2(n18408), .A(n18368), .ZN(n18364) );
  OAI221_X1 U21407 ( .B1(n18822), .B2(n19004), .C1(n18822), .C2(n18368), .A(
        n18364), .ZN(P3_U2863) );
  NOR2_X1 U21408 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18373), .ZN(
        n18547) );
  NOR2_X1 U21409 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18839), .ZN(
        n18639) );
  NOR2_X1 U21410 ( .A1(n18547), .A2(n18639), .ZN(n18366) );
  OAI22_X1 U21411 ( .A1(n18367), .A2(n18839), .B1(n18366), .B2(n18365), .ZN(
        P3_U2866) );
  NOR2_X1 U21412 ( .A1(n18369), .A2(n18368), .ZN(P3_U2867) );
  NOR2_X1 U21413 ( .A1(n18371), .A2(n18370), .ZN(n18401) );
  NOR2_X1 U21414 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18826) );
  NOR2_X1 U21415 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18456) );
  NAND2_X1 U21416 ( .A1(n18826), .A2(n18456), .ZN(n18407) );
  AND2_X1 U21417 ( .A1(n18715), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18740) );
  INV_X1 U21418 ( .A(n18858), .ZN(n18739) );
  NOR2_X1 U21419 ( .A1(n18839), .A2(n18522), .ZN(n18743) );
  NOR2_X2 U21420 ( .A1(n18822), .A2(n18738), .ZN(n18737) );
  NOR2_X1 U21421 ( .A1(n18737), .A2(n18473), .ZN(n18434) );
  NOR2_X1 U21422 ( .A1(n18739), .A2(n18434), .ZN(n18403) );
  AND2_X1 U21423 ( .A1(n18745), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18746) );
  NOR2_X2 U21424 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18738), .ZN(
        n18716) );
  AOI22_X1 U21425 ( .A1(n18740), .A2(n18403), .B1(n18746), .B2(n18716), .ZN(
        n18377) );
  NOR3_X1 U21426 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18373), .A3(
        n18839), .ZN(n18744) );
  NAND2_X1 U21427 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18744), .ZN(
        n18710) );
  INV_X1 U21428 ( .A(n18710), .ZN(n18788) );
  NOR2_X1 U21429 ( .A1(n18788), .A2(n18716), .ZN(n18711) );
  OAI21_X1 U21430 ( .B1(n18822), .B2(n18960), .A(n18715), .ZN(n18615) );
  OAI22_X1 U21431 ( .A1(n18685), .A2(n18711), .B1(n18615), .B2(n18434), .ZN(
        n18374) );
  INV_X1 U21432 ( .A(n18374), .ZN(n18404) );
  NOR2_X2 U21433 ( .A1(n18375), .A2(n18685), .ZN(n18741) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18404), .B1(
        n18741), .B2(n18788), .ZN(n18376) );
  OAI211_X1 U21435 ( .C1(n18749), .C2(n18407), .A(n18377), .B(n18376), .ZN(
        P3_U2868) );
  NAND2_X1 U21436 ( .A1(n18401), .A2(n10113), .ZN(n18755) );
  AND2_X1 U21437 ( .A1(n18745), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18751) );
  AND2_X1 U21438 ( .A1(n18715), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18750) );
  AOI22_X1 U21439 ( .A1(n18751), .A2(n18716), .B1(n18750), .B2(n18403), .ZN(
        n18380) );
  NOR2_X2 U21440 ( .A1(n18378), .A2(n18685), .ZN(n18752) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18404), .B1(
        n18752), .B2(n18788), .ZN(n18379) );
  OAI211_X1 U21442 ( .C1(n18755), .C2(n18407), .A(n18380), .B(n18379), .ZN(
        P3_U2869) );
  AND2_X1 U21443 ( .A1(n18745), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18758) );
  NOR2_X2 U21444 ( .A1(n18455), .A2(n18382), .ZN(n18757) );
  AOI22_X1 U21445 ( .A1(n18758), .A2(n18716), .B1(n18757), .B2(n18403), .ZN(
        n18384) );
  NOR2_X2 U21446 ( .A1(n19437), .A2(n18685), .ZN(n18756) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18404), .B1(
        n18756), .B2(n18788), .ZN(n18383) );
  OAI211_X1 U21448 ( .C1(n18761), .C2(n18407), .A(n18384), .B(n18383), .ZN(
        P3_U2870) );
  NAND2_X1 U21449 ( .A1(n18401), .A2(n18385), .ZN(n18767) );
  NOR2_X2 U21450 ( .A1(n18455), .A2(n18386), .ZN(n18763) );
  NOR2_X2 U21451 ( .A1(n19445), .A2(n18685), .ZN(n18762) );
  AOI22_X1 U21452 ( .A1(n18763), .A2(n18403), .B1(n18762), .B2(n18788), .ZN(
        n18388) );
  AND2_X1 U21453 ( .A1(n18745), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18764) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18404), .B1(
        n18764), .B2(n18716), .ZN(n18387) );
  OAI211_X1 U21455 ( .C1(n18767), .C2(n18407), .A(n18388), .B(n18387), .ZN(
        P3_U2871) );
  NAND2_X1 U21456 ( .A1(n18401), .A2(n18389), .ZN(n18773) );
  AND2_X1 U21457 ( .A1(n18715), .A2(BUF2_REG_4__SCAN_IN), .ZN(n18768) );
  NOR2_X2 U21458 ( .A1(n19450), .A2(n18685), .ZN(n18770) );
  AOI22_X1 U21459 ( .A1(n18768), .A2(n18403), .B1(n18770), .B2(n18788), .ZN(
        n18392) );
  NOR2_X2 U21460 ( .A1(n18685), .A2(n18390), .ZN(n18769) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18404), .B1(
        n18769), .B2(n18716), .ZN(n18391) );
  OAI211_X1 U21462 ( .C1(n18773), .C2(n18407), .A(n18392), .B(n18391), .ZN(
        P3_U2872) );
  NAND2_X1 U21463 ( .A1(n18401), .A2(n18393), .ZN(n18779) );
  NOR2_X2 U21464 ( .A1(n19456), .A2(n18685), .ZN(n18776) );
  NOR2_X2 U21465 ( .A1(n18394), .A2(n18455), .ZN(n18775) );
  AOI22_X1 U21466 ( .A1(n18776), .A2(n18788), .B1(n18775), .B2(n18403), .ZN(
        n18396) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18404), .B1(
        n18774), .B2(n18716), .ZN(n18395) );
  OAI211_X1 U21468 ( .C1(n18779), .C2(n18407), .A(n18396), .B(n18395), .ZN(
        P3_U2873) );
  AND2_X1 U21469 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18715), .ZN(n18780) );
  AND2_X1 U21470 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18745), .ZN(n18782) );
  AOI22_X1 U21471 ( .A1(n18780), .A2(n18403), .B1(n18782), .B2(n18716), .ZN(
        n18399) );
  NOR2_X2 U21472 ( .A1(n19460), .A2(n18685), .ZN(n18781) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18404), .B1(
        n18781), .B2(n18788), .ZN(n18398) );
  OAI211_X1 U21474 ( .C1(n18785), .C2(n18407), .A(n18399), .B(n18398), .ZN(
        P3_U2874) );
  NAND2_X1 U21475 ( .A1(n18401), .A2(n18400), .ZN(n18796) );
  NOR2_X2 U21476 ( .A1(n18402), .A2(n18455), .ZN(n18787) );
  AOI22_X1 U21477 ( .A1(n18789), .A2(n18716), .B1(n18787), .B2(n18403), .ZN(
        n18406) );
  NOR2_X2 U21478 ( .A1(n18685), .A2(n19467), .ZN(n18791) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18404), .B1(
        n18791), .B2(n18788), .ZN(n18405) );
  OAI211_X1 U21480 ( .C1(n18796), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2875) );
  INV_X1 U21481 ( .A(n18456), .ZN(n18409) );
  NOR2_X1 U21482 ( .A1(n18408), .A2(n18455), .ZN(n18742) );
  NAND2_X1 U21483 ( .A1(n18742), .A2(n18823), .ZN(n18682) );
  OAI22_X1 U21484 ( .A1(n18685), .A2(n18738), .B1(n18409), .B2(n18682), .ZN(
        n18420) );
  NAND2_X1 U21485 ( .A1(n18823), .A2(n18858), .ZN(n18591) );
  NOR2_X1 U21486 ( .A1(n18409), .A2(n18591), .ZN(n18429) );
  AOI22_X1 U21487 ( .A1(n18740), .A2(n18429), .B1(n18746), .B2(n18737), .ZN(
        n18411) );
  NAND2_X1 U21488 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18823), .ZN(
        n18500) );
  NOR2_X2 U21489 ( .A1(n18500), .A2(n18409), .ZN(n18495) );
  INV_X1 U21490 ( .A(n18749), .ZN(n18686) );
  AOI22_X1 U21491 ( .A1(n18741), .A2(n18716), .B1(n18495), .B2(n18686), .ZN(
        n18410) );
  OAI211_X1 U21492 ( .C1(n18412), .C2(n18420), .A(n18411), .B(n18410), .ZN(
        P3_U2876) );
  AOI22_X1 U21493 ( .A1(n18752), .A2(n18716), .B1(n18750), .B2(n18429), .ZN(
        n18414) );
  INV_X1 U21494 ( .A(n18755), .ZN(n18690) );
  AOI22_X1 U21495 ( .A1(n18495), .A2(n18690), .B1(n18751), .B2(n18737), .ZN(
        n18413) );
  OAI211_X1 U21496 ( .C1(n18415), .C2(n18420), .A(n18414), .B(n18413), .ZN(
        P3_U2877) );
  AOI22_X1 U21497 ( .A1(n18757), .A2(n18429), .B1(n18756), .B2(n18716), .ZN(
        n18418) );
  INV_X1 U21498 ( .A(n18761), .ZN(n18416) );
  AOI22_X1 U21499 ( .A1(n18495), .A2(n18416), .B1(n18758), .B2(n18737), .ZN(
        n18417) );
  OAI211_X1 U21500 ( .C1(n18419), .C2(n18420), .A(n18418), .B(n18417), .ZN(
        P3_U2878) );
  INV_X1 U21501 ( .A(n18495), .ZN(n18433) );
  AOI22_X1 U21502 ( .A1(n18763), .A2(n18429), .B1(n18762), .B2(n18716), .ZN(
        n18422) );
  INV_X1 U21503 ( .A(n18420), .ZN(n18430) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18430), .B1(
        n18764), .B2(n18737), .ZN(n18421) );
  OAI211_X1 U21505 ( .C1(n18433), .C2(n18767), .A(n18422), .B(n18421), .ZN(
        P3_U2879) );
  AOI22_X1 U21506 ( .A1(n18768), .A2(n18429), .B1(n18770), .B2(n18716), .ZN(
        n18424) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18430), .B1(
        n18769), .B2(n18737), .ZN(n18423) );
  OAI211_X1 U21508 ( .C1(n18433), .C2(n18773), .A(n18424), .B(n18423), .ZN(
        P3_U2880) );
  AOI22_X1 U21509 ( .A1(n18776), .A2(n18716), .B1(n18775), .B2(n18429), .ZN(
        n18426) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18430), .B1(
        n18774), .B2(n18737), .ZN(n18425) );
  OAI211_X1 U21511 ( .C1(n18433), .C2(n18779), .A(n18426), .B(n18425), .ZN(
        P3_U2881) );
  AOI22_X1 U21512 ( .A1(n18781), .A2(n18716), .B1(n18780), .B2(n18429), .ZN(
        n18428) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18430), .B1(
        n18782), .B2(n18737), .ZN(n18427) );
  OAI211_X1 U21514 ( .C1(n18433), .C2(n18785), .A(n18428), .B(n18427), .ZN(
        P3_U2882) );
  AOI22_X1 U21515 ( .A1(n18791), .A2(n18716), .B1(n18787), .B2(n18429), .ZN(
        n18432) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18430), .B1(
        n18789), .B2(n18737), .ZN(n18431) );
  OAI211_X1 U21517 ( .C1(n18433), .C2(n18796), .A(n18432), .B(n18431), .ZN(
        P3_U2883) );
  NAND2_X1 U21518 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18456), .ZN(
        n18457) );
  NOR2_X2 U21519 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18457), .ZN(
        n18518) );
  INV_X1 U21520 ( .A(n18518), .ZN(n18454) );
  NOR2_X1 U21521 ( .A1(n18495), .A2(n18518), .ZN(n18478) );
  NOR2_X1 U21522 ( .A1(n18739), .A2(n18478), .ZN(n18450) );
  AOI22_X1 U21523 ( .A1(n18741), .A2(n18737), .B1(n18740), .B2(n18450), .ZN(
        n18437) );
  OAI21_X1 U21524 ( .B1(n18434), .B2(n18712), .A(n18478), .ZN(n18435) );
  OAI211_X1 U21525 ( .C1(n18518), .C2(n18960), .A(n18715), .B(n18435), .ZN(
        n18451) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18451), .B1(
        n18746), .B2(n18473), .ZN(n18436) );
  OAI211_X1 U21527 ( .C1(n18454), .C2(n18749), .A(n18437), .B(n18436), .ZN(
        P3_U2884) );
  AOI22_X1 U21528 ( .A1(n18752), .A2(n18737), .B1(n18750), .B2(n18450), .ZN(
        n18439) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18451), .B1(
        n18751), .B2(n18473), .ZN(n18438) );
  OAI211_X1 U21530 ( .C1(n18454), .C2(n18755), .A(n18439), .B(n18438), .ZN(
        P3_U2885) );
  AOI22_X1 U21531 ( .A1(n18757), .A2(n18450), .B1(n18756), .B2(n18737), .ZN(
        n18441) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18451), .B1(
        n18758), .B2(n18473), .ZN(n18440) );
  OAI211_X1 U21533 ( .C1(n18454), .C2(n18761), .A(n18441), .B(n18440), .ZN(
        P3_U2886) );
  AOI22_X1 U21534 ( .A1(n18763), .A2(n18450), .B1(n18762), .B2(n18737), .ZN(
        n18443) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18451), .B1(
        n18764), .B2(n18473), .ZN(n18442) );
  OAI211_X1 U21536 ( .C1(n18454), .C2(n18767), .A(n18443), .B(n18442), .ZN(
        P3_U2887) );
  AOI22_X1 U21537 ( .A1(n18769), .A2(n18473), .B1(n18768), .B2(n18450), .ZN(
        n18445) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18451), .B1(
        n18770), .B2(n18737), .ZN(n18444) );
  OAI211_X1 U21539 ( .C1(n18454), .C2(n18773), .A(n18445), .B(n18444), .ZN(
        P3_U2888) );
  AOI22_X1 U21540 ( .A1(n18775), .A2(n18450), .B1(n18774), .B2(n18473), .ZN(
        n18447) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18451), .B1(
        n18776), .B2(n18737), .ZN(n18446) );
  OAI211_X1 U21542 ( .C1(n18454), .C2(n18779), .A(n18447), .B(n18446), .ZN(
        P3_U2889) );
  AOI22_X1 U21543 ( .A1(n18781), .A2(n18737), .B1(n18780), .B2(n18450), .ZN(
        n18449) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18451), .B1(
        n18782), .B2(n18473), .ZN(n18448) );
  OAI211_X1 U21545 ( .C1(n18454), .C2(n18785), .A(n18449), .B(n18448), .ZN(
        P3_U2890) );
  AOI22_X1 U21546 ( .A1(n18789), .A2(n18473), .B1(n18787), .B2(n18450), .ZN(
        n18453) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18451), .B1(
        n18791), .B2(n18737), .ZN(n18452) );
  OAI211_X1 U21548 ( .C1(n18454), .C2(n18796), .A(n18453), .B(n18452), .ZN(
        P3_U2891) );
  INV_X1 U21549 ( .A(n18457), .ZN(n18502) );
  NAND2_X1 U21550 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18502), .ZN(
        n18477) );
  AOI21_X1 U21551 ( .B1(n18823), .B2(n18712), .A(n18455), .ZN(n18546) );
  OAI211_X1 U21552 ( .C1(n18541), .C2(n18960), .A(n18456), .B(n18546), .ZN(
        n18474) );
  NOR2_X1 U21553 ( .A1(n18739), .A2(n18457), .ZN(n18472) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18474), .B1(
        n18740), .B2(n18472), .ZN(n18459) );
  AOI22_X1 U21555 ( .A1(n18741), .A2(n18473), .B1(n18495), .B2(n18746), .ZN(
        n18458) );
  OAI211_X1 U21556 ( .C1(n18477), .C2(n18749), .A(n18459), .B(n18458), .ZN(
        P3_U2892) );
  AOI22_X1 U21557 ( .A1(n18752), .A2(n18473), .B1(n18750), .B2(n18472), .ZN(
        n18461) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18474), .B1(
        n18495), .B2(n18751), .ZN(n18460) );
  OAI211_X1 U21559 ( .C1(n18477), .C2(n18755), .A(n18461), .B(n18460), .ZN(
        P3_U2893) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18474), .B1(
        n18757), .B2(n18472), .ZN(n18463) );
  AOI22_X1 U21561 ( .A1(n18495), .A2(n18758), .B1(n18756), .B2(n18473), .ZN(
        n18462) );
  OAI211_X1 U21562 ( .C1(n18477), .C2(n18761), .A(n18463), .B(n18462), .ZN(
        P3_U2894) );
  AOI22_X1 U21563 ( .A1(n18495), .A2(n18764), .B1(n18763), .B2(n18472), .ZN(
        n18465) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18474), .B1(
        n18762), .B2(n18473), .ZN(n18464) );
  OAI211_X1 U21565 ( .C1(n18477), .C2(n18767), .A(n18465), .B(n18464), .ZN(
        P3_U2895) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18474), .B1(
        n18768), .B2(n18472), .ZN(n18467) );
  AOI22_X1 U21567 ( .A1(n18495), .A2(n18769), .B1(n18770), .B2(n18473), .ZN(
        n18466) );
  OAI211_X1 U21568 ( .C1(n18477), .C2(n18773), .A(n18467), .B(n18466), .ZN(
        P3_U2896) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18474), .B1(
        n18775), .B2(n18472), .ZN(n18469) );
  AOI22_X1 U21570 ( .A1(n18495), .A2(n18774), .B1(n18776), .B2(n18473), .ZN(
        n18468) );
  OAI211_X1 U21571 ( .C1(n18477), .C2(n18779), .A(n18469), .B(n18468), .ZN(
        P3_U2897) );
  AOI22_X1 U21572 ( .A1(n18781), .A2(n18473), .B1(n18780), .B2(n18472), .ZN(
        n18471) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18474), .B1(
        n18495), .B2(n18782), .ZN(n18470) );
  OAI211_X1 U21574 ( .C1(n18477), .C2(n18785), .A(n18471), .B(n18470), .ZN(
        P3_U2898) );
  AOI22_X1 U21575 ( .A1(n18791), .A2(n18473), .B1(n18787), .B2(n18472), .ZN(
        n18476) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18474), .B1(
        n18495), .B2(n18789), .ZN(n18475) );
  OAI211_X1 U21577 ( .C1(n18477), .C2(n18796), .A(n18476), .B(n18475), .ZN(
        P3_U2899) );
  NAND2_X1 U21578 ( .A1(n18826), .A2(n18547), .ZN(n18499) );
  AOI21_X1 U21579 ( .B1(n18499), .B2(n18477), .A(n18739), .ZN(n18494) );
  AOI22_X1 U21580 ( .A1(n18518), .A2(n18746), .B1(n18740), .B2(n18494), .ZN(
        n18481) );
  INV_X1 U21581 ( .A(n18499), .ZN(n18564) );
  AOI221_X1 U21582 ( .B1(n18478), .B2(n18477), .C1(n18712), .C2(n18477), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18479) );
  OAI21_X1 U21583 ( .B1(n18564), .B2(n18479), .A(n18715), .ZN(n18496) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18496), .B1(
        n18741), .B2(n18495), .ZN(n18480) );
  OAI211_X1 U21585 ( .C1(n18499), .C2(n18749), .A(n18481), .B(n18480), .ZN(
        P3_U2900) );
  AOI22_X1 U21586 ( .A1(n18518), .A2(n18751), .B1(n18494), .B2(n18750), .ZN(
        n18483) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18496), .B1(
        n18495), .B2(n18752), .ZN(n18482) );
  OAI211_X1 U21588 ( .C1(n18499), .C2(n18755), .A(n18483), .B(n18482), .ZN(
        P3_U2901) );
  AOI22_X1 U21589 ( .A1(n18495), .A2(n18756), .B1(n18494), .B2(n18757), .ZN(
        n18485) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18496), .B1(
        n18518), .B2(n18758), .ZN(n18484) );
  OAI211_X1 U21591 ( .C1(n18499), .C2(n18761), .A(n18485), .B(n18484), .ZN(
        P3_U2902) );
  AOI22_X1 U21592 ( .A1(n18495), .A2(n18762), .B1(n18494), .B2(n18763), .ZN(
        n18487) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18496), .B1(
        n18518), .B2(n18764), .ZN(n18486) );
  OAI211_X1 U21594 ( .C1(n18499), .C2(n18767), .A(n18487), .B(n18486), .ZN(
        P3_U2903) );
  AOI22_X1 U21595 ( .A1(n18495), .A2(n18770), .B1(n18494), .B2(n18768), .ZN(
        n18489) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18496), .B1(
        n18518), .B2(n18769), .ZN(n18488) );
  OAI211_X1 U21597 ( .C1(n18499), .C2(n18773), .A(n18489), .B(n18488), .ZN(
        P3_U2904) );
  AOI22_X1 U21598 ( .A1(n18518), .A2(n18774), .B1(n18494), .B2(n18775), .ZN(
        n18491) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18496), .B1(
        n18495), .B2(n18776), .ZN(n18490) );
  OAI211_X1 U21600 ( .C1(n18499), .C2(n18779), .A(n18491), .B(n18490), .ZN(
        P3_U2905) );
  AOI22_X1 U21601 ( .A1(n18518), .A2(n18782), .B1(n18494), .B2(n18780), .ZN(
        n18493) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18496), .B1(
        n18495), .B2(n18781), .ZN(n18492) );
  OAI211_X1 U21603 ( .C1(n18499), .C2(n18785), .A(n18493), .B(n18492), .ZN(
        P3_U2906) );
  AOI22_X1 U21604 ( .A1(n18495), .A2(n18791), .B1(n18494), .B2(n18787), .ZN(
        n18498) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18496), .B1(
        n18518), .B2(n18789), .ZN(n18497) );
  OAI211_X1 U21606 ( .C1(n18499), .C2(n18796), .A(n18498), .B(n18497), .ZN(
        P3_U2907) );
  INV_X1 U21607 ( .A(n18500), .ZN(n18590) );
  NAND2_X1 U21608 ( .A1(n18590), .A2(n18547), .ZN(n18523) );
  INV_X1 U21609 ( .A(n18547), .ZN(n18501) );
  NOR2_X1 U21610 ( .A1(n18501), .A2(n18591), .ZN(n18517) );
  AOI22_X1 U21611 ( .A1(n18541), .A2(n18746), .B1(n18740), .B2(n18517), .ZN(
        n18504) );
  INV_X1 U21612 ( .A(n18682), .ZN(n18592) );
  AOI22_X1 U21613 ( .A1(n18745), .A2(n18502), .B1(n18547), .B2(n18592), .ZN(
        n18519) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18519), .B1(
        n18741), .B2(n18518), .ZN(n18503) );
  OAI211_X1 U21615 ( .C1(n18749), .C2(n18523), .A(n18504), .B(n18503), .ZN(
        P3_U2908) );
  AOI22_X1 U21616 ( .A1(n18541), .A2(n18751), .B1(n18750), .B2(n18517), .ZN(
        n18506) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18519), .B1(
        n18518), .B2(n18752), .ZN(n18505) );
  OAI211_X1 U21618 ( .C1(n18755), .C2(n18523), .A(n18506), .B(n18505), .ZN(
        P3_U2909) );
  AOI22_X1 U21619 ( .A1(n18518), .A2(n18756), .B1(n18757), .B2(n18517), .ZN(
        n18508) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18519), .B1(
        n18541), .B2(n18758), .ZN(n18507) );
  OAI211_X1 U21621 ( .C1(n18761), .C2(n18523), .A(n18508), .B(n18507), .ZN(
        P3_U2910) );
  AOI22_X1 U21622 ( .A1(n18518), .A2(n18762), .B1(n18763), .B2(n18517), .ZN(
        n18510) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18519), .B1(
        n18541), .B2(n18764), .ZN(n18509) );
  OAI211_X1 U21624 ( .C1(n18767), .C2(n18523), .A(n18510), .B(n18509), .ZN(
        P3_U2911) );
  AOI22_X1 U21625 ( .A1(n18518), .A2(n18770), .B1(n18768), .B2(n18517), .ZN(
        n18512) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18519), .B1(
        n18541), .B2(n18769), .ZN(n18511) );
  OAI211_X1 U21627 ( .C1(n18773), .C2(n18523), .A(n18512), .B(n18511), .ZN(
        P3_U2912) );
  AOI22_X1 U21628 ( .A1(n18541), .A2(n18774), .B1(n18775), .B2(n18517), .ZN(
        n18514) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18519), .B1(
        n18518), .B2(n18776), .ZN(n18513) );
  OAI211_X1 U21630 ( .C1(n18779), .C2(n18523), .A(n18514), .B(n18513), .ZN(
        P3_U2913) );
  AOI22_X1 U21631 ( .A1(n18541), .A2(n18782), .B1(n18780), .B2(n18517), .ZN(
        n18516) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18519), .B1(
        n18518), .B2(n18781), .ZN(n18515) );
  OAI211_X1 U21633 ( .C1(n18785), .C2(n18523), .A(n18516), .B(n18515), .ZN(
        P3_U2914) );
  AOI22_X1 U21634 ( .A1(n18541), .A2(n18789), .B1(n18787), .B2(n18517), .ZN(
        n18521) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18519), .B1(
        n18518), .B2(n18791), .ZN(n18520) );
  OAI211_X1 U21636 ( .C1(n18796), .C2(n18523), .A(n18521), .B(n18520), .ZN(
        P3_U2915) );
  NOR2_X1 U21637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18522), .ZN(
        n18593) );
  NAND2_X1 U21638 ( .A1(n18593), .A2(n18822), .ZN(n18545) );
  NOR2_X1 U21639 ( .A1(n18585), .A2(n18609), .ZN(n18568) );
  NOR2_X1 U21640 ( .A1(n18739), .A2(n18568), .ZN(n18540) );
  AOI22_X1 U21641 ( .A1(n18564), .A2(n18746), .B1(n18740), .B2(n18540), .ZN(
        n18527) );
  NOR2_X1 U21642 ( .A1(n18564), .A2(n18541), .ZN(n18524) );
  OAI21_X1 U21643 ( .B1(n18524), .B2(n18712), .A(n18568), .ZN(n18525) );
  OAI211_X1 U21644 ( .C1(n18609), .C2(n18960), .A(n18715), .B(n18525), .ZN(
        n18542) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18542), .B1(
        n18741), .B2(n18541), .ZN(n18526) );
  OAI211_X1 U21646 ( .C1(n18749), .C2(n18545), .A(n18527), .B(n18526), .ZN(
        P3_U2916) );
  AOI22_X1 U21647 ( .A1(n18564), .A2(n18751), .B1(n18750), .B2(n18540), .ZN(
        n18529) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18752), .ZN(n18528) );
  OAI211_X1 U21649 ( .C1(n18755), .C2(n18545), .A(n18529), .B(n18528), .ZN(
        P3_U2917) );
  AOI22_X1 U21650 ( .A1(n18541), .A2(n18756), .B1(n18757), .B2(n18540), .ZN(
        n18531) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18542), .B1(
        n18564), .B2(n18758), .ZN(n18530) );
  OAI211_X1 U21652 ( .C1(n18761), .C2(n18545), .A(n18531), .B(n18530), .ZN(
        P3_U2918) );
  AOI22_X1 U21653 ( .A1(n18564), .A2(n18764), .B1(n18763), .B2(n18540), .ZN(
        n18533) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18762), .ZN(n18532) );
  OAI211_X1 U21655 ( .C1(n18767), .C2(n18545), .A(n18533), .B(n18532), .ZN(
        P3_U2919) );
  AOI22_X1 U21656 ( .A1(n18564), .A2(n18769), .B1(n18768), .B2(n18540), .ZN(
        n18535) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18770), .ZN(n18534) );
  OAI211_X1 U21658 ( .C1(n18773), .C2(n18545), .A(n18535), .B(n18534), .ZN(
        P3_U2920) );
  AOI22_X1 U21659 ( .A1(n18541), .A2(n18776), .B1(n18775), .B2(n18540), .ZN(
        n18537) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18542), .B1(
        n18564), .B2(n18774), .ZN(n18536) );
  OAI211_X1 U21661 ( .C1(n18779), .C2(n18545), .A(n18537), .B(n18536), .ZN(
        P3_U2921) );
  AOI22_X1 U21662 ( .A1(n18564), .A2(n18782), .B1(n18780), .B2(n18540), .ZN(
        n18539) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18781), .ZN(n18538) );
  OAI211_X1 U21664 ( .C1(n18785), .C2(n18545), .A(n18539), .B(n18538), .ZN(
        P3_U2922) );
  AOI22_X1 U21665 ( .A1(n18541), .A2(n18791), .B1(n18787), .B2(n18540), .ZN(
        n18544) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18542), .B1(
        n18564), .B2(n18789), .ZN(n18543) );
  OAI211_X1 U21667 ( .C1(n18796), .C2(n18545), .A(n18544), .B(n18543), .ZN(
        P3_U2923) );
  NAND2_X1 U21668 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18593), .ZN(
        n18567) );
  OAI211_X1 U21669 ( .C1(n18633), .C2(n18960), .A(n18547), .B(n18546), .ZN(
        n18563) );
  AND2_X1 U21670 ( .A1(n18858), .A2(n18593), .ZN(n18562) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18563), .B1(
        n18740), .B2(n18562), .ZN(n18549) );
  AOI22_X1 U21672 ( .A1(n18741), .A2(n18564), .B1(n18746), .B2(n18585), .ZN(
        n18548) );
  OAI211_X1 U21673 ( .C1(n18749), .C2(n18567), .A(n18549), .B(n18548), .ZN(
        P3_U2924) );
  AOI22_X1 U21674 ( .A1(n18564), .A2(n18752), .B1(n18750), .B2(n18562), .ZN(
        n18551) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18563), .B1(
        n18751), .B2(n18585), .ZN(n18550) );
  OAI211_X1 U21676 ( .C1(n18755), .C2(n18567), .A(n18551), .B(n18550), .ZN(
        P3_U2925) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18563), .B1(
        n18757), .B2(n18562), .ZN(n18553) );
  AOI22_X1 U21678 ( .A1(n18564), .A2(n18756), .B1(n18758), .B2(n18585), .ZN(
        n18552) );
  OAI211_X1 U21679 ( .C1(n18761), .C2(n18567), .A(n18553), .B(n18552), .ZN(
        P3_U2926) );
  AOI22_X1 U21680 ( .A1(n18764), .A2(n18585), .B1(n18763), .B2(n18562), .ZN(
        n18555) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18563), .B1(
        n18564), .B2(n18762), .ZN(n18554) );
  OAI211_X1 U21682 ( .C1(n18767), .C2(n18567), .A(n18555), .B(n18554), .ZN(
        P3_U2927) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18563), .B1(
        n18768), .B2(n18562), .ZN(n18557) );
  AOI22_X1 U21684 ( .A1(n18564), .A2(n18770), .B1(n18769), .B2(n18585), .ZN(
        n18556) );
  OAI211_X1 U21685 ( .C1(n18773), .C2(n18567), .A(n18557), .B(n18556), .ZN(
        P3_U2928) );
  AOI22_X1 U21686 ( .A1(n18564), .A2(n18776), .B1(n18775), .B2(n18562), .ZN(
        n18559) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18563), .B1(
        n18774), .B2(n18585), .ZN(n18558) );
  OAI211_X1 U21688 ( .C1(n18779), .C2(n18567), .A(n18559), .B(n18558), .ZN(
        P3_U2929) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18563), .B1(
        n18780), .B2(n18562), .ZN(n18561) );
  AOI22_X1 U21690 ( .A1(n18564), .A2(n18781), .B1(n18782), .B2(n18585), .ZN(
        n18560) );
  OAI211_X1 U21691 ( .C1(n18785), .C2(n18567), .A(n18561), .B(n18560), .ZN(
        P3_U2930) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18563), .B1(
        n18787), .B2(n18562), .ZN(n18566) );
  AOI22_X1 U21693 ( .A1(n18564), .A2(n18791), .B1(n18789), .B2(n18585), .ZN(
        n18565) );
  OAI211_X1 U21694 ( .C1(n18796), .C2(n18567), .A(n18566), .B(n18565), .ZN(
        P3_U2931) );
  NAND2_X1 U21695 ( .A1(n18826), .A2(n18639), .ZN(n18589) );
  NOR2_X1 U21696 ( .A1(n18633), .A2(n18655), .ZN(n18616) );
  NOR2_X1 U21697 ( .A1(n18739), .A2(n18616), .ZN(n18584) );
  AOI22_X1 U21698 ( .A1(n18741), .A2(n18585), .B1(n18740), .B2(n18584), .ZN(
        n18571) );
  OAI21_X1 U21699 ( .B1(n18568), .B2(n18712), .A(n18616), .ZN(n18569) );
  OAI211_X1 U21700 ( .C1(n18655), .C2(n18960), .A(n18715), .B(n18569), .ZN(
        n18586) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18586), .B1(
        n18746), .B2(n18609), .ZN(n18570) );
  OAI211_X1 U21702 ( .C1(n18749), .C2(n18589), .A(n18571), .B(n18570), .ZN(
        P3_U2932) );
  AOI22_X1 U21703 ( .A1(n18751), .A2(n18609), .B1(n18750), .B2(n18584), .ZN(
        n18573) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18586), .B1(
        n18752), .B2(n18585), .ZN(n18572) );
  OAI211_X1 U21705 ( .C1(n18755), .C2(n18589), .A(n18573), .B(n18572), .ZN(
        P3_U2933) );
  AOI22_X1 U21706 ( .A1(n18757), .A2(n18584), .B1(n18756), .B2(n18585), .ZN(
        n18575) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18586), .B1(
        n18758), .B2(n18609), .ZN(n18574) );
  OAI211_X1 U21708 ( .C1(n18761), .C2(n18589), .A(n18575), .B(n18574), .ZN(
        P3_U2934) );
  AOI22_X1 U21709 ( .A1(n18763), .A2(n18584), .B1(n18762), .B2(n18585), .ZN(
        n18577) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18586), .B1(
        n18764), .B2(n18609), .ZN(n18576) );
  OAI211_X1 U21711 ( .C1(n18767), .C2(n18589), .A(n18577), .B(n18576), .ZN(
        P3_U2935) );
  AOI22_X1 U21712 ( .A1(n18769), .A2(n18609), .B1(n18768), .B2(n18584), .ZN(
        n18579) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18586), .B1(
        n18770), .B2(n18585), .ZN(n18578) );
  OAI211_X1 U21714 ( .C1(n18773), .C2(n18589), .A(n18579), .B(n18578), .ZN(
        P3_U2936) );
  AOI22_X1 U21715 ( .A1(n18776), .A2(n18585), .B1(n18775), .B2(n18584), .ZN(
        n18581) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18586), .B1(
        n18774), .B2(n18609), .ZN(n18580) );
  OAI211_X1 U21717 ( .C1(n18779), .C2(n18589), .A(n18581), .B(n18580), .ZN(
        P3_U2937) );
  AOI22_X1 U21718 ( .A1(n18780), .A2(n18584), .B1(n18782), .B2(n18609), .ZN(
        n18583) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18586), .B1(
        n18781), .B2(n18585), .ZN(n18582) );
  OAI211_X1 U21720 ( .C1(n18785), .C2(n18589), .A(n18583), .B(n18582), .ZN(
        P3_U2938) );
  AOI22_X1 U21721 ( .A1(n18789), .A2(n18609), .B1(n18787), .B2(n18584), .ZN(
        n18588) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18586), .B1(
        n18791), .B2(n18585), .ZN(n18587) );
  OAI211_X1 U21723 ( .C1(n18796), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P3_U2939) );
  NAND2_X1 U21724 ( .A1(n18590), .A2(n18639), .ZN(n18614) );
  INV_X1 U21725 ( .A(n18639), .ZN(n18613) );
  NOR2_X1 U21726 ( .A1(n18613), .A2(n18591), .ZN(n18608) );
  AOI22_X1 U21727 ( .A1(n18740), .A2(n18608), .B1(n18746), .B2(n18633), .ZN(
        n18595) );
  AOI22_X1 U21728 ( .A1(n18745), .A2(n18593), .B1(n18639), .B2(n18592), .ZN(
        n18610) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18610), .B1(
        n18741), .B2(n18609), .ZN(n18594) );
  OAI211_X1 U21730 ( .C1(n18749), .C2(n18614), .A(n18595), .B(n18594), .ZN(
        P3_U2940) );
  AOI22_X1 U21731 ( .A1(n18752), .A2(n18609), .B1(n18750), .B2(n18608), .ZN(
        n18597) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18610), .B1(
        n18751), .B2(n18633), .ZN(n18596) );
  OAI211_X1 U21733 ( .C1(n18755), .C2(n18614), .A(n18597), .B(n18596), .ZN(
        P3_U2941) );
  AOI22_X1 U21734 ( .A1(n18757), .A2(n18608), .B1(n18756), .B2(n18609), .ZN(
        n18599) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18610), .B1(
        n18758), .B2(n18633), .ZN(n18598) );
  OAI211_X1 U21736 ( .C1(n18761), .C2(n18614), .A(n18599), .B(n18598), .ZN(
        P3_U2942) );
  AOI22_X1 U21737 ( .A1(n18764), .A2(n18633), .B1(n18763), .B2(n18608), .ZN(
        n18601) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18610), .B1(
        n18762), .B2(n18609), .ZN(n18600) );
  OAI211_X1 U21739 ( .C1(n18767), .C2(n18614), .A(n18601), .B(n18600), .ZN(
        P3_U2943) );
  AOI22_X1 U21740 ( .A1(n18768), .A2(n18608), .B1(n18770), .B2(n18609), .ZN(
        n18603) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18610), .B1(
        n18769), .B2(n18633), .ZN(n18602) );
  OAI211_X1 U21742 ( .C1(n18773), .C2(n18614), .A(n18603), .B(n18602), .ZN(
        P3_U2944) );
  AOI22_X1 U21743 ( .A1(n18775), .A2(n18608), .B1(n18774), .B2(n18633), .ZN(
        n18605) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18610), .B1(
        n18776), .B2(n18609), .ZN(n18604) );
  OAI211_X1 U21745 ( .C1(n18779), .C2(n18614), .A(n18605), .B(n18604), .ZN(
        P3_U2945) );
  AOI22_X1 U21746 ( .A1(n18781), .A2(n18609), .B1(n18780), .B2(n18608), .ZN(
        n18607) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18610), .B1(
        n18782), .B2(n18633), .ZN(n18606) );
  OAI211_X1 U21748 ( .C1(n18785), .C2(n18614), .A(n18607), .B(n18606), .ZN(
        P3_U2946) );
  AOI22_X1 U21749 ( .A1(n18789), .A2(n18633), .B1(n18787), .B2(n18608), .ZN(
        n18612) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18610), .B1(
        n18791), .B2(n18609), .ZN(n18611) );
  OAI211_X1 U21751 ( .C1(n18796), .C2(n18614), .A(n18612), .B(n18611), .ZN(
        P3_U2947) );
  NOR2_X1 U21752 ( .A1(n18823), .A2(n18613), .ZN(n18638) );
  NAND2_X1 U21753 ( .A1(n18638), .A2(n18822), .ZN(n18637) );
  NOR2_X1 U21754 ( .A1(n18677), .A2(n18706), .ZN(n18660) );
  NOR2_X1 U21755 ( .A1(n18739), .A2(n18660), .ZN(n18632) );
  AOI22_X1 U21756 ( .A1(n18740), .A2(n18632), .B1(n18746), .B2(n18655), .ZN(
        n18619) );
  AOI221_X1 U21757 ( .B1(n18660), .B2(n18712), .C1(n18660), .C2(n18616), .A(
        n18615), .ZN(n18617) );
  INV_X1 U21758 ( .A(n18617), .ZN(n18634) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18634), .B1(
        n18741), .B2(n18633), .ZN(n18618) );
  OAI211_X1 U21760 ( .C1(n18749), .C2(n18637), .A(n18619), .B(n18618), .ZN(
        P3_U2948) );
  AOI22_X1 U21761 ( .A1(n18751), .A2(n18655), .B1(n18750), .B2(n18632), .ZN(
        n18621) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18634), .B1(
        n18752), .B2(n18633), .ZN(n18620) );
  OAI211_X1 U21763 ( .C1(n18755), .C2(n18637), .A(n18621), .B(n18620), .ZN(
        P3_U2949) );
  AOI22_X1 U21764 ( .A1(n18757), .A2(n18632), .B1(n18756), .B2(n18633), .ZN(
        n18623) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18634), .B1(
        n18758), .B2(n18655), .ZN(n18622) );
  OAI211_X1 U21766 ( .C1(n18761), .C2(n18637), .A(n18623), .B(n18622), .ZN(
        P3_U2950) );
  AOI22_X1 U21767 ( .A1(n18764), .A2(n18655), .B1(n18763), .B2(n18632), .ZN(
        n18625) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18634), .B1(
        n18762), .B2(n18633), .ZN(n18624) );
  OAI211_X1 U21769 ( .C1(n18767), .C2(n18637), .A(n18625), .B(n18624), .ZN(
        P3_U2951) );
  AOI22_X1 U21770 ( .A1(n18769), .A2(n18655), .B1(n18768), .B2(n18632), .ZN(
        n18627) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18634), .B1(
        n18770), .B2(n18633), .ZN(n18626) );
  OAI211_X1 U21772 ( .C1(n18773), .C2(n18637), .A(n18627), .B(n18626), .ZN(
        P3_U2952) );
  AOI22_X1 U21773 ( .A1(n18776), .A2(n18633), .B1(n18775), .B2(n18632), .ZN(
        n18629) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18634), .B1(
        n18774), .B2(n18655), .ZN(n18628) );
  OAI211_X1 U21775 ( .C1(n18779), .C2(n18637), .A(n18629), .B(n18628), .ZN(
        P3_U2953) );
  AOI22_X1 U21776 ( .A1(n18781), .A2(n18633), .B1(n18780), .B2(n18632), .ZN(
        n18631) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18634), .B1(
        n18782), .B2(n18655), .ZN(n18630) );
  OAI211_X1 U21778 ( .C1(n18785), .C2(n18637), .A(n18631), .B(n18630), .ZN(
        P3_U2954) );
  AOI22_X1 U21779 ( .A1(n18791), .A2(n18633), .B1(n18787), .B2(n18632), .ZN(
        n18636) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18634), .B1(
        n18789), .B2(n18655), .ZN(n18635) );
  OAI211_X1 U21781 ( .C1(n18796), .C2(n18637), .A(n18636), .B(n18635), .ZN(
        P3_U2955) );
  NAND2_X1 U21782 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18638), .ZN(
        n18659) );
  INV_X1 U21783 ( .A(n18638), .ZN(n18684) );
  NOR2_X1 U21784 ( .A1(n18739), .A2(n18684), .ZN(n18654) );
  AOI22_X1 U21785 ( .A1(n18741), .A2(n18655), .B1(n18740), .B2(n18654), .ZN(
        n18641) );
  AOI22_X1 U21786 ( .A1(n18745), .A2(n18639), .B1(n18742), .B2(n18638), .ZN(
        n18656) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18656), .B1(
        n18746), .B2(n18677), .ZN(n18640) );
  OAI211_X1 U21788 ( .C1(n18749), .C2(n18659), .A(n18641), .B(n18640), .ZN(
        P3_U2956) );
  AOI22_X1 U21789 ( .A1(n18752), .A2(n18655), .B1(n18750), .B2(n18654), .ZN(
        n18643) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18656), .B1(
        n18751), .B2(n18677), .ZN(n18642) );
  OAI211_X1 U21791 ( .C1(n18755), .C2(n18659), .A(n18643), .B(n18642), .ZN(
        P3_U2957) );
  AOI22_X1 U21792 ( .A1(n18758), .A2(n18677), .B1(n18757), .B2(n18654), .ZN(
        n18645) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18656), .B1(
        n18756), .B2(n18655), .ZN(n18644) );
  OAI211_X1 U21794 ( .C1(n18761), .C2(n18659), .A(n18645), .B(n18644), .ZN(
        P3_U2958) );
  AOI22_X1 U21795 ( .A1(n18764), .A2(n18677), .B1(n18763), .B2(n18654), .ZN(
        n18647) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18656), .B1(
        n18762), .B2(n18655), .ZN(n18646) );
  OAI211_X1 U21797 ( .C1(n18767), .C2(n18659), .A(n18647), .B(n18646), .ZN(
        P3_U2959) );
  AOI22_X1 U21798 ( .A1(n18768), .A2(n18654), .B1(n18770), .B2(n18655), .ZN(
        n18649) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18656), .B1(
        n18769), .B2(n18677), .ZN(n18648) );
  OAI211_X1 U21800 ( .C1(n18773), .C2(n18659), .A(n18649), .B(n18648), .ZN(
        P3_U2960) );
  AOI22_X1 U21801 ( .A1(n18776), .A2(n18655), .B1(n18775), .B2(n18654), .ZN(
        n18651) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18656), .B1(
        n18774), .B2(n18677), .ZN(n18650) );
  OAI211_X1 U21803 ( .C1(n18779), .C2(n18659), .A(n18651), .B(n18650), .ZN(
        P3_U2961) );
  AOI22_X1 U21804 ( .A1(n18781), .A2(n18655), .B1(n18780), .B2(n18654), .ZN(
        n18653) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18656), .B1(
        n18782), .B2(n18677), .ZN(n18652) );
  OAI211_X1 U21806 ( .C1(n18785), .C2(n18659), .A(n18653), .B(n18652), .ZN(
        P3_U2962) );
  AOI22_X1 U21807 ( .A1(n18789), .A2(n18677), .B1(n18787), .B2(n18654), .ZN(
        n18658) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18656), .B1(
        n18791), .B2(n18655), .ZN(n18657) );
  OAI211_X1 U21809 ( .C1(n18796), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        P3_U2963) );
  NAND2_X1 U21810 ( .A1(n18744), .A2(n18822), .ZN(n18681) );
  INV_X1 U21811 ( .A(n18659), .ZN(n18732) );
  INV_X1 U21812 ( .A(n18681), .ZN(n18790) );
  NOR2_X1 U21813 ( .A1(n18732), .A2(n18790), .ZN(n18713) );
  NOR2_X1 U21814 ( .A1(n18739), .A2(n18713), .ZN(n18676) );
  AOI22_X1 U21815 ( .A1(n18741), .A2(n18677), .B1(n18740), .B2(n18676), .ZN(
        n18663) );
  OAI21_X1 U21816 ( .B1(n18660), .B2(n18712), .A(n18713), .ZN(n18661) );
  OAI211_X1 U21817 ( .C1(n18790), .C2(n18960), .A(n18715), .B(n18661), .ZN(
        n18678) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18678), .B1(
        n18746), .B2(n18706), .ZN(n18662) );
  OAI211_X1 U21819 ( .C1(n18749), .C2(n18681), .A(n18663), .B(n18662), .ZN(
        P3_U2964) );
  AOI22_X1 U21820 ( .A1(n18752), .A2(n18677), .B1(n18750), .B2(n18676), .ZN(
        n18665) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18678), .B1(
        n18751), .B2(n18706), .ZN(n18664) );
  OAI211_X1 U21822 ( .C1(n18755), .C2(n18681), .A(n18665), .B(n18664), .ZN(
        P3_U2965) );
  AOI22_X1 U21823 ( .A1(n18757), .A2(n18676), .B1(n18756), .B2(n18677), .ZN(
        n18667) );
  AOI22_X1 U21824 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18678), .B1(
        n18758), .B2(n18706), .ZN(n18666) );
  OAI211_X1 U21825 ( .C1(n18761), .C2(n18681), .A(n18667), .B(n18666), .ZN(
        P3_U2966) );
  AOI22_X1 U21826 ( .A1(n18764), .A2(n18706), .B1(n18763), .B2(n18676), .ZN(
        n18669) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18678), .B1(
        n18762), .B2(n18677), .ZN(n18668) );
  OAI211_X1 U21828 ( .C1(n18767), .C2(n18681), .A(n18669), .B(n18668), .ZN(
        P3_U2967) );
  AOI22_X1 U21829 ( .A1(n18769), .A2(n18706), .B1(n18768), .B2(n18676), .ZN(
        n18671) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18678), .B1(
        n18770), .B2(n18677), .ZN(n18670) );
  OAI211_X1 U21831 ( .C1(n18773), .C2(n18681), .A(n18671), .B(n18670), .ZN(
        P3_U2968) );
  AOI22_X1 U21832 ( .A1(n18775), .A2(n18676), .B1(n18774), .B2(n18706), .ZN(
        n18673) );
  AOI22_X1 U21833 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18678), .B1(
        n18776), .B2(n18677), .ZN(n18672) );
  OAI211_X1 U21834 ( .C1(n18779), .C2(n18681), .A(n18673), .B(n18672), .ZN(
        P3_U2969) );
  AOI22_X1 U21835 ( .A1(n18780), .A2(n18676), .B1(n18782), .B2(n18706), .ZN(
        n18675) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18678), .B1(
        n18781), .B2(n18677), .ZN(n18674) );
  OAI211_X1 U21837 ( .C1(n18785), .C2(n18681), .A(n18675), .B(n18674), .ZN(
        P3_U2970) );
  AOI22_X1 U21838 ( .A1(n18791), .A2(n18677), .B1(n18787), .B2(n18676), .ZN(
        n18680) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18678), .B1(
        n18789), .B2(n18706), .ZN(n18679) );
  OAI211_X1 U21840 ( .C1(n18796), .C2(n18681), .A(n18680), .B(n18679), .ZN(
        P3_U2971) );
  NAND2_X1 U21841 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18683) );
  OAI22_X1 U21842 ( .A1(n18685), .A2(n18684), .B1(n18683), .B2(n18682), .ZN(
        n18694) );
  AND2_X1 U21843 ( .A1(n18858), .A2(n18744), .ZN(n18705) );
  AOI22_X1 U21844 ( .A1(n18740), .A2(n18705), .B1(n18746), .B2(n18732), .ZN(
        n18688) );
  AOI22_X1 U21845 ( .A1(n18741), .A2(n18706), .B1(n18686), .B2(n18788), .ZN(
        n18687) );
  OAI211_X1 U21846 ( .C1(n18689), .C2(n18694), .A(n18688), .B(n18687), .ZN(
        P3_U2972) );
  AOI22_X1 U21847 ( .A1(n18751), .A2(n18732), .B1(n18750), .B2(n18705), .ZN(
        n18692) );
  AOI22_X1 U21848 ( .A1(n18752), .A2(n18706), .B1(n18690), .B2(n18788), .ZN(
        n18691) );
  OAI211_X1 U21849 ( .C1(n18693), .C2(n18694), .A(n18692), .B(n18691), .ZN(
        P3_U2973) );
  AOI22_X1 U21850 ( .A1(n18758), .A2(n18732), .B1(n18757), .B2(n18705), .ZN(
        n18696) );
  INV_X1 U21851 ( .A(n18694), .ZN(n18707) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18707), .B1(
        n18756), .B2(n18706), .ZN(n18695) );
  OAI211_X1 U21853 ( .C1(n18761), .C2(n18710), .A(n18696), .B(n18695), .ZN(
        P3_U2974) );
  AOI22_X1 U21854 ( .A1(n18763), .A2(n18705), .B1(n18762), .B2(n18706), .ZN(
        n18698) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18707), .B1(
        n18764), .B2(n18732), .ZN(n18697) );
  OAI211_X1 U21856 ( .C1(n18767), .C2(n18710), .A(n18698), .B(n18697), .ZN(
        P3_U2975) );
  AOI22_X1 U21857 ( .A1(n18769), .A2(n18732), .B1(n18768), .B2(n18705), .ZN(
        n18700) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18707), .B1(
        n18770), .B2(n18706), .ZN(n18699) );
  OAI211_X1 U21859 ( .C1(n18773), .C2(n18710), .A(n18700), .B(n18699), .ZN(
        P3_U2976) );
  AOI22_X1 U21860 ( .A1(n18775), .A2(n18705), .B1(n18774), .B2(n18732), .ZN(
        n18702) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18707), .B1(
        n18776), .B2(n18706), .ZN(n18701) );
  OAI211_X1 U21862 ( .C1(n18779), .C2(n18710), .A(n18702), .B(n18701), .ZN(
        P3_U2977) );
  AOI22_X1 U21863 ( .A1(n18780), .A2(n18705), .B1(n18782), .B2(n18732), .ZN(
        n18704) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18707), .B1(
        n18781), .B2(n18706), .ZN(n18703) );
  OAI211_X1 U21865 ( .C1(n18785), .C2(n18710), .A(n18704), .B(n18703), .ZN(
        P3_U2978) );
  AOI22_X1 U21866 ( .A1(n18791), .A2(n18706), .B1(n18787), .B2(n18705), .ZN(
        n18709) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18707), .B1(
        n18789), .B2(n18732), .ZN(n18708) );
  OAI211_X1 U21868 ( .C1(n18796), .C2(n18710), .A(n18709), .B(n18708), .ZN(
        P3_U2979) );
  INV_X1 U21869 ( .A(n18716), .ZN(n18736) );
  NOR2_X1 U21870 ( .A1(n18739), .A2(n18711), .ZN(n18731) );
  AOI22_X1 U21871 ( .A1(n18741), .A2(n18732), .B1(n18740), .B2(n18731), .ZN(
        n18718) );
  OAI21_X1 U21872 ( .B1(n18713), .B2(n18712), .A(n18711), .ZN(n18714) );
  OAI211_X1 U21873 ( .C1(n18716), .C2(n18960), .A(n18715), .B(n18714), .ZN(
        n18733) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18733), .B1(
        n18746), .B2(n18790), .ZN(n18717) );
  OAI211_X1 U21875 ( .C1(n18749), .C2(n18736), .A(n18718), .B(n18717), .ZN(
        P3_U2980) );
  AOI22_X1 U21876 ( .A1(n18752), .A2(n18732), .B1(n18750), .B2(n18731), .ZN(
        n18720) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18733), .B1(
        n18751), .B2(n18790), .ZN(n18719) );
  OAI211_X1 U21878 ( .C1(n18755), .C2(n18736), .A(n18720), .B(n18719), .ZN(
        P3_U2981) );
  AOI22_X1 U21879 ( .A1(n18758), .A2(n18790), .B1(n18757), .B2(n18731), .ZN(
        n18722) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18733), .B1(
        n18756), .B2(n18732), .ZN(n18721) );
  OAI211_X1 U21881 ( .C1(n18761), .C2(n18736), .A(n18722), .B(n18721), .ZN(
        P3_U2982) );
  AOI22_X1 U21882 ( .A1(n18763), .A2(n18731), .B1(n18762), .B2(n18732), .ZN(
        n18724) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18733), .B1(
        n18764), .B2(n18790), .ZN(n18723) );
  OAI211_X1 U21884 ( .C1(n18767), .C2(n18736), .A(n18724), .B(n18723), .ZN(
        P3_U2983) );
  AOI22_X1 U21885 ( .A1(n18768), .A2(n18731), .B1(n18770), .B2(n18732), .ZN(
        n18726) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18733), .B1(
        n18769), .B2(n18790), .ZN(n18725) );
  OAI211_X1 U21887 ( .C1(n18773), .C2(n18736), .A(n18726), .B(n18725), .ZN(
        P3_U2984) );
  AOI22_X1 U21888 ( .A1(n18775), .A2(n18731), .B1(n18774), .B2(n18790), .ZN(
        n18728) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18733), .B1(
        n18776), .B2(n18732), .ZN(n18727) );
  OAI211_X1 U21890 ( .C1(n18779), .C2(n18736), .A(n18728), .B(n18727), .ZN(
        P3_U2985) );
  AOI22_X1 U21891 ( .A1(n18780), .A2(n18731), .B1(n18782), .B2(n18790), .ZN(
        n18730) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18733), .B1(
        n18781), .B2(n18732), .ZN(n18729) );
  OAI211_X1 U21893 ( .C1(n18785), .C2(n18736), .A(n18730), .B(n18729), .ZN(
        P3_U2986) );
  AOI22_X1 U21894 ( .A1(n18789), .A2(n18790), .B1(n18787), .B2(n18731), .ZN(
        n18735) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18733), .B1(
        n18791), .B2(n18732), .ZN(n18734) );
  OAI211_X1 U21896 ( .C1(n18796), .C2(n18736), .A(n18735), .B(n18734), .ZN(
        P3_U2987) );
  INV_X1 U21897 ( .A(n18737), .ZN(n18795) );
  NOR2_X1 U21898 ( .A1(n18739), .A2(n18738), .ZN(n18786) );
  AOI22_X1 U21899 ( .A1(n18741), .A2(n18790), .B1(n18740), .B2(n18786), .ZN(
        n18748) );
  AOI22_X1 U21900 ( .A1(n18745), .A2(n18744), .B1(n18743), .B2(n18742), .ZN(
        n18792) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18792), .B1(
        n18746), .B2(n18788), .ZN(n18747) );
  OAI211_X1 U21902 ( .C1(n18749), .C2(n18795), .A(n18748), .B(n18747), .ZN(
        P3_U2988) );
  AOI22_X1 U21903 ( .A1(n18751), .A2(n18788), .B1(n18750), .B2(n18786), .ZN(
        n18754) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18792), .B1(
        n18752), .B2(n18790), .ZN(n18753) );
  OAI211_X1 U21905 ( .C1(n18755), .C2(n18795), .A(n18754), .B(n18753), .ZN(
        P3_U2989) );
  AOI22_X1 U21906 ( .A1(n18757), .A2(n18786), .B1(n18756), .B2(n18790), .ZN(
        n18760) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18792), .B1(
        n18758), .B2(n18788), .ZN(n18759) );
  OAI211_X1 U21908 ( .C1(n18761), .C2(n18795), .A(n18760), .B(n18759), .ZN(
        P3_U2990) );
  AOI22_X1 U21909 ( .A1(n18763), .A2(n18786), .B1(n18762), .B2(n18790), .ZN(
        n18766) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18792), .B1(
        n18764), .B2(n18788), .ZN(n18765) );
  OAI211_X1 U21911 ( .C1(n18767), .C2(n18795), .A(n18766), .B(n18765), .ZN(
        P3_U2991) );
  AOI22_X1 U21912 ( .A1(n18769), .A2(n18788), .B1(n18768), .B2(n18786), .ZN(
        n18772) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18792), .B1(
        n18770), .B2(n18790), .ZN(n18771) );
  OAI211_X1 U21914 ( .C1(n18773), .C2(n18795), .A(n18772), .B(n18771), .ZN(
        P3_U2992) );
  AOI22_X1 U21915 ( .A1(n18775), .A2(n18786), .B1(n18774), .B2(n18788), .ZN(
        n18778) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18792), .B1(
        n18776), .B2(n18790), .ZN(n18777) );
  OAI211_X1 U21917 ( .C1(n18779), .C2(n18795), .A(n18778), .B(n18777), .ZN(
        P3_U2993) );
  AOI22_X1 U21918 ( .A1(n18781), .A2(n18790), .B1(n18780), .B2(n18786), .ZN(
        n18784) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18792), .B1(
        n18782), .B2(n18788), .ZN(n18783) );
  OAI211_X1 U21920 ( .C1(n18785), .C2(n18795), .A(n18784), .B(n18783), .ZN(
        P3_U2994) );
  AOI22_X1 U21921 ( .A1(n18789), .A2(n18788), .B1(n18787), .B2(n18786), .ZN(
        n18794) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18792), .B1(
        n18791), .B2(n18790), .ZN(n18793) );
  OAI211_X1 U21923 ( .C1(n18796), .C2(n18795), .A(n18794), .B(n18793), .ZN(
        P3_U2995) );
  OAI22_X1 U21924 ( .A1(n18800), .A2(n18799), .B1(n18798), .B2(n18797), .ZN(
        n18801) );
  AOI221_X1 U21925 ( .B1(n18804), .B2(n18803), .C1(n18802), .C2(n18803), .A(
        n18801), .ZN(n19002) );
  AOI211_X1 U21926 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18835), .A(
        n18806), .B(n18805), .ZN(n18846) );
  OAI21_X1 U21927 ( .B1(n18809), .B2(n18808), .A(n18807), .ZN(n18830) );
  AOI21_X1 U21928 ( .B1(n18828), .B2(n18821), .A(n18830), .ZN(n18811) );
  OAI21_X1 U21929 ( .B1(n18812), .B2(n18811), .A(n18810), .ZN(n18966) );
  NOR2_X1 U21930 ( .A1(n18835), .A2(n18966), .ZN(n18816) );
  AOI21_X1 U21931 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18813), .A(
        n18821), .ZN(n18819) );
  OAI22_X1 U21932 ( .A1(n18814), .A2(n18833), .B1(n18828), .B2(n18819), .ZN(
        n18963) );
  NAND2_X1 U21933 ( .A1(n18967), .A2(n18963), .ZN(n18815) );
  OAI22_X1 U21934 ( .A1(n18816), .A2(n18967), .B1(n18835), .B2(n18815), .ZN(
        n18842) );
  NAND2_X1 U21935 ( .A1(n18818), .A2(n18817), .ZN(n18820) );
  INV_X1 U21936 ( .A(n18819), .ZN(n18829) );
  AOI22_X1 U21937 ( .A1(n18979), .A2(n18820), .B1(n18829), .B2(n13850), .ZN(
        n18975) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18821), .B1(
        n18820), .B2(n18988), .ZN(n18824) );
  INV_X1 U21939 ( .A(n18824), .ZN(n18983) );
  NOR3_X1 U21940 ( .A1(n18823), .A2(n18822), .A3(n18983), .ZN(n18825) );
  OAI22_X1 U21941 ( .A1(n18975), .A2(n18825), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18824), .ZN(n18827) );
  INV_X1 U21942 ( .A(n18835), .ZN(n18834) );
  AOI21_X1 U21943 ( .B1(n18827), .B2(n18834), .A(n18826), .ZN(n18837) );
  OAI211_X1 U21944 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18829), .B(n18828), .ZN(
        n18832) );
  NAND3_X1 U21945 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13851), .A3(
        n18830), .ZN(n18831) );
  OAI211_X1 U21946 ( .C1(n18971), .C2(n18833), .A(n18832), .B(n18831), .ZN(
        n18972) );
  AOI22_X1 U21947 ( .A1(n18835), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18972), .B2(n18834), .ZN(n18838) );
  OR2_X1 U21948 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18838), .ZN(
        n18836) );
  AOI221_X1 U21949 ( .B1(n18837), .B2(n18836), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18838), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18841) );
  OAI21_X1 U21950 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18838), .ZN(n18840) );
  AOI222_X1 U21951 ( .A1(n18842), .A2(n18841), .B1(n18842), .B2(n18840), .C1(
        n18841), .C2(n18839), .ZN(n18845) );
  OAI21_X1 U21952 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18843), .ZN(n18844) );
  NAND4_X1 U21953 ( .A1(n19002), .A2(n18846), .A3(n18845), .A4(n18844), .ZN(
        n18852) );
  AOI211_X1 U21954 ( .C1(n18849), .C2(n18848), .A(n18847), .B(n18852), .ZN(
        n18958) );
  AOI21_X1 U21955 ( .B1(n19007), .B2(n18856), .A(n18958), .ZN(n18859) );
  NOR2_X1 U21956 ( .A1(n18857), .A2(n18858), .ZN(n18851) );
  NOR2_X1 U21957 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19015) );
  NOR2_X1 U21958 ( .A1(n19013), .A2(n19006), .ZN(n18855) );
  AOI211_X1 U21959 ( .C1(n18982), .C2(n19015), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18855), .ZN(n18850) );
  AOI211_X1 U21960 ( .C1(n19005), .C2(n18852), .A(n18851), .B(n18850), .ZN(
        n18853) );
  OAI221_X1 U21961 ( .B1(n18957), .B2(n18859), .C1(n18957), .C2(n18854), .A(
        n18853), .ZN(P3_U2996) );
  INV_X1 U21962 ( .A(n18855), .ZN(n18862) );
  NAND4_X1 U21963 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19007), .A4(n18856), .ZN(n18864) );
  INV_X1 U21964 ( .A(n18857), .ZN(n18860) );
  NAND3_X1 U21965 ( .A1(n18860), .A2(n18859), .A3(n18858), .ZN(n18861) );
  NAND4_X1 U21966 ( .A1(n18863), .A2(n18862), .A3(n18864), .A4(n18861), .ZN(
        P3_U2997) );
  INV_X1 U21967 ( .A(n19015), .ZN(n18866) );
  AND4_X1 U21968 ( .A1(n18866), .A2(n18865), .A3(n18864), .A4(n18959), .ZN(
        P3_U2998) );
  AND2_X1 U21969 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n9798), .ZN(P3_U2999) );
  AND2_X1 U21970 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n9797), .ZN(P3_U3000) );
  AND2_X1 U21971 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n9798), .ZN(P3_U3001) );
  AND2_X1 U21972 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n9797), .ZN(P3_U3002) );
  AND2_X1 U21973 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n9798), .ZN(P3_U3003) );
  AND2_X1 U21974 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n9797), .ZN(P3_U3004) );
  AND2_X1 U21975 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n9798), .ZN(P3_U3005) );
  AND2_X1 U21976 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n9797), .ZN(P3_U3006) );
  AND2_X1 U21977 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n9797), .ZN(P3_U3007) );
  AND2_X1 U21978 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n9798), .ZN(P3_U3008) );
  AND2_X1 U21979 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n9797), .ZN(P3_U3009) );
  AND2_X1 U21980 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n9798), .ZN(P3_U3010) );
  AND2_X1 U21981 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n9797), .ZN(P3_U3011) );
  AND2_X1 U21982 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n9798), .ZN(P3_U3012) );
  AND2_X1 U21983 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n9797), .ZN(P3_U3013) );
  AND2_X1 U21984 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n9798), .ZN(P3_U3014) );
  AND2_X1 U21985 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n9797), .ZN(P3_U3015) );
  AND2_X1 U21986 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n9798), .ZN(P3_U3016) );
  AND2_X1 U21987 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n9798), .ZN(P3_U3017) );
  AND2_X1 U21988 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n9797), .ZN(P3_U3018) );
  AND2_X1 U21989 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n9798), .ZN(P3_U3019) );
  AND2_X1 U21990 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n9797), .ZN(P3_U3020) );
  AND2_X1 U21991 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n9797), .ZN(P3_U3021)
         );
  AND2_X1 U21992 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n9798), .ZN(P3_U3022)
         );
  AND2_X1 U21993 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n9797), .ZN(P3_U3023)
         );
  AND2_X1 U21994 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n9798), .ZN(P3_U3024)
         );
  AND2_X1 U21995 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n9797), .ZN(P3_U3025)
         );
  AND2_X1 U21996 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n9798), .ZN(P3_U3026)
         );
  AND2_X1 U21997 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n9797), .ZN(P3_U3027)
         );
  AND2_X1 U21998 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n9798), .ZN(P3_U3028)
         );
  INV_X1 U21999 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18868) );
  AOI21_X1 U22000 ( .B1(HOLD), .B2(n18869), .A(n18868), .ZN(n18872) );
  AOI21_X1 U22001 ( .B1(n19007), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18880), 
        .ZN(n18882) );
  INV_X1 U22002 ( .A(NA), .ZN(n21117) );
  OAI21_X1 U22003 ( .B1(n21117), .B2(n18870), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18881) );
  INV_X1 U22004 ( .A(n18881), .ZN(n18871) );
  OAI22_X1 U22005 ( .A1(n18999), .A2(n18872), .B1(n18882), .B2(n18871), .ZN(
        P3_U3029) );
  AOI21_X1 U22006 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18873) );
  AOI21_X1 U22007 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18873), .ZN(
        n18874) );
  AOI22_X1 U22008 ( .A1(n19007), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18874), .ZN(n18875) );
  NAND2_X1 U22009 ( .A1(n18875), .A2(n19010), .ZN(P3_U3030) );
  NOR2_X1 U22010 ( .A1(n18883), .A2(n21254), .ZN(n18878) );
  NAND2_X1 U22011 ( .A1(n19007), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18876) );
  OAI22_X1 U22012 ( .A1(NA), .A2(n18876), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18877) );
  OAI22_X1 U22013 ( .A1(n18878), .A2(n18877), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18879) );
  OAI22_X1 U22014 ( .A1(n18882), .A2(n18881), .B1(n18880), .B2(n18879), .ZN(
        P3_U3031) );
  OAI222_X1 U22015 ( .A1(n18990), .A2(n18945), .B1(n18884), .B2(n18999), .C1(
        n18885), .C2(n18935), .ZN(P3_U3032) );
  OAI222_X1 U22016 ( .A1(n18935), .A2(n18887), .B1(n18886), .B2(n18999), .C1(
        n18885), .C2(n18945), .ZN(P3_U3033) );
  OAI222_X1 U22017 ( .A1(n18935), .A2(n18889), .B1(n18888), .B2(n18999), .C1(
        n18887), .C2(n18945), .ZN(P3_U3034) );
  INV_X1 U22018 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18891) );
  OAI222_X1 U22019 ( .A1(n18935), .A2(n18891), .B1(n18890), .B2(n18999), .C1(
        n18889), .C2(n18945), .ZN(P3_U3035) );
  OAI222_X1 U22020 ( .A1(n18935), .A2(n18893), .B1(n18892), .B2(n18999), .C1(
        n18891), .C2(n18945), .ZN(P3_U3036) );
  OAI222_X1 U22021 ( .A1(n18935), .A2(n18895), .B1(n18894), .B2(n18999), .C1(
        n18893), .C2(n18945), .ZN(P3_U3037) );
  OAI222_X1 U22022 ( .A1(n18935), .A2(n18898), .B1(n18896), .B2(n18999), .C1(
        n18895), .C2(n18945), .ZN(P3_U3038) );
  OAI222_X1 U22023 ( .A1(n18898), .A2(n18945), .B1(n18897), .B2(n18999), .C1(
        n18899), .C2(n18935), .ZN(P3_U3039) );
  OAI222_X1 U22024 ( .A1(n18935), .A2(n18901), .B1(n18900), .B2(n18999), .C1(
        n18899), .C2(n18945), .ZN(P3_U3040) );
  OAI222_X1 U22025 ( .A1(n18935), .A2(n18903), .B1(n18902), .B2(n18999), .C1(
        n18901), .C2(n18945), .ZN(P3_U3041) );
  INV_X1 U22026 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18905) );
  OAI222_X1 U22027 ( .A1(n18935), .A2(n18905), .B1(n18904), .B2(n18999), .C1(
        n18903), .C2(n18945), .ZN(P3_U3042) );
  OAI222_X1 U22028 ( .A1(n18935), .A2(n18907), .B1(n18906), .B2(n18999), .C1(
        n18905), .C2(n18945), .ZN(P3_U3043) );
  INV_X1 U22029 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18909) );
  OAI222_X1 U22030 ( .A1(n18935), .A2(n18909), .B1(n18908), .B2(n18999), .C1(
        n18907), .C2(n18945), .ZN(P3_U3044) );
  OAI222_X1 U22031 ( .A1(n18935), .A2(n18911), .B1(n18910), .B2(n18999), .C1(
        n18909), .C2(n18945), .ZN(P3_U3045) );
  OAI222_X1 U22032 ( .A1(n18935), .A2(n18913), .B1(n18912), .B2(n18999), .C1(
        n18911), .C2(n18945), .ZN(P3_U3046) );
  INV_X1 U22033 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18915) );
  OAI222_X1 U22034 ( .A1(n18935), .A2(n18915), .B1(n18914), .B2(n18999), .C1(
        n18913), .C2(n18945), .ZN(P3_U3047) );
  OAI222_X1 U22035 ( .A1(n18935), .A2(n18917), .B1(n18916), .B2(n18999), .C1(
        n18915), .C2(n18945), .ZN(P3_U3048) );
  INV_X1 U22036 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18920) );
  OAI222_X1 U22037 ( .A1(n18935), .A2(n18920), .B1(n18918), .B2(n18999), .C1(
        n18917), .C2(n18945), .ZN(P3_U3049) );
  OAI222_X1 U22038 ( .A1(n18920), .A2(n18945), .B1(n18919), .B2(n18999), .C1(
        n18921), .C2(n18935), .ZN(P3_U3050) );
  OAI222_X1 U22039 ( .A1(n18935), .A2(n18924), .B1(n18922), .B2(n18999), .C1(
        n18921), .C2(n18945), .ZN(P3_U3051) );
  OAI222_X1 U22040 ( .A1(n18924), .A2(n18945), .B1(n18923), .B2(n18999), .C1(
        n18925), .C2(n18935), .ZN(P3_U3052) );
  OAI222_X1 U22041 ( .A1(n18935), .A2(n18928), .B1(n18926), .B2(n18999), .C1(
        n18925), .C2(n18945), .ZN(P3_U3053) );
  OAI222_X1 U22042 ( .A1(n18928), .A2(n18945), .B1(n18927), .B2(n18999), .C1(
        n18929), .C2(n18935), .ZN(P3_U3054) );
  OAI222_X1 U22043 ( .A1(n18935), .A2(n18931), .B1(n18930), .B2(n18999), .C1(
        n18929), .C2(n18945), .ZN(P3_U3055) );
  OAI222_X1 U22044 ( .A1(n18935), .A2(n18933), .B1(n18932), .B2(n18999), .C1(
        n18931), .C2(n18945), .ZN(P3_U3056) );
  OAI222_X1 U22045 ( .A1(n18935), .A2(n18936), .B1(n18934), .B2(n18999), .C1(
        n18933), .C2(n18945), .ZN(P3_U3057) );
  INV_X1 U22046 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18939) );
  OAI222_X1 U22047 ( .A1(n18935), .A2(n18939), .B1(n18937), .B2(n18999), .C1(
        n18936), .C2(n18945), .ZN(P3_U3058) );
  OAI222_X1 U22048 ( .A1(n18939), .A2(n18945), .B1(n18938), .B2(n18999), .C1(
        n18940), .C2(n18935), .ZN(P3_U3059) );
  OAI222_X1 U22049 ( .A1(n18935), .A2(n18944), .B1(n18941), .B2(n18999), .C1(
        n18940), .C2(n18945), .ZN(P3_U3060) );
  INV_X1 U22050 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18943) );
  OAI222_X1 U22051 ( .A1(n18945), .A2(n18944), .B1(n18943), .B2(n18999), .C1(
        n18942), .C2(n18935), .ZN(P3_U3061) );
  INV_X1 U22052 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18946) );
  AOI22_X1 U22053 ( .A1(n18999), .A2(n18947), .B1(n18946), .B2(n19020), .ZN(
        P3_U3274) );
  INV_X1 U22054 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18993) );
  INV_X1 U22055 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18948) );
  AOI22_X1 U22056 ( .A1(n18999), .A2(n18993), .B1(n18948), .B2(n19020), .ZN(
        P3_U3275) );
  INV_X1 U22057 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18949) );
  AOI22_X1 U22058 ( .A1(n18999), .A2(n18950), .B1(n18949), .B2(n19020), .ZN(
        P3_U3276) );
  INV_X1 U22059 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18996) );
  INV_X1 U22060 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18951) );
  AOI22_X1 U22061 ( .A1(n18999), .A2(n18996), .B1(n18951), .B2(n19020), .ZN(
        P3_U3277) );
  INV_X1 U22062 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18953) );
  AOI21_X1 U22063 ( .B1(n9798), .B2(n18953), .A(n18952), .ZN(P3_U3280) );
  OAI21_X1 U22064 ( .B1(n18956), .B2(n18955), .A(n18954), .ZN(P3_U3281) );
  NOR2_X1 U22065 ( .A1(n18958), .A2(n18957), .ZN(n18961) );
  OAI21_X1 U22066 ( .B1(n18961), .B2(n18960), .A(n18959), .ZN(P3_U3282) );
  INV_X1 U22067 ( .A(n18962), .ZN(n18965) );
  NOR2_X1 U22068 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19022), .ZN(
        n18964) );
  AOI22_X1 U22069 ( .A1(n18982), .A2(n18965), .B1(n18964), .B2(n18963), .ZN(
        n18969) );
  AOI21_X1 U22070 ( .B1(n18984), .B2(n18966), .A(n18989), .ZN(n18968) );
  OAI22_X1 U22071 ( .A1(n18989), .A2(n18969), .B1(n18968), .B2(n18967), .ZN(
        P3_U3285) );
  NOR2_X1 U22072 ( .A1(n18970), .A2(n18985), .ZN(n18977) );
  AOI22_X1 U22073 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n15673), .B2(n16482), .ZN(
        n18976) );
  AOI222_X1 U22074 ( .A1(n18972), .A2(n18984), .B1(n18977), .B2(n18976), .C1(
        n18982), .C2(n18971), .ZN(n18973) );
  AOI22_X1 U22075 ( .A1(n18989), .A2(n18974), .B1(n18973), .B2(n18986), .ZN(
        P3_U3288) );
  INV_X1 U22076 ( .A(n18975), .ZN(n18980) );
  INV_X1 U22077 ( .A(n18976), .ZN(n18978) );
  AOI222_X1 U22078 ( .A1(n18980), .A2(n18984), .B1(n18982), .B2(n18979), .C1(
        n18978), .C2(n18977), .ZN(n18981) );
  AOI22_X1 U22079 ( .A1(n18989), .A2(n13850), .B1(n18981), .B2(n18986), .ZN(
        P3_U3289) );
  AOI222_X1 U22080 ( .A1(n18985), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18984), 
        .B2(n18983), .C1(n18988), .C2(n18982), .ZN(n18987) );
  AOI22_X1 U22081 ( .A1(n18989), .A2(n18988), .B1(n18987), .B2(n18986), .ZN(
        P3_U3290) );
  AOI21_X1 U22082 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18991) );
  AOI22_X1 U22083 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18991), .B2(n18990), .ZN(n18994) );
  AOI22_X1 U22084 ( .A1(n18997), .A2(n18994), .B1(n18993), .B2(n18992), .ZN(
        P3_U3292) );
  OAI21_X1 U22085 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18997), .ZN(n18995) );
  OAI21_X1 U22086 ( .B1(n18997), .B2(n18996), .A(n18995), .ZN(P3_U3293) );
  INV_X1 U22087 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18998) );
  AOI22_X1 U22088 ( .A1(n18999), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18998), 
        .B2(n19020), .ZN(P3_U3294) );
  INV_X1 U22089 ( .A(n19000), .ZN(n19003) );
  NAND2_X1 U22090 ( .A1(n19003), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19001) );
  OAI21_X1 U22091 ( .B1(n19003), .B2(n19002), .A(n19001), .ZN(P3_U3295) );
  OAI22_X1 U22092 ( .A1(n19007), .A2(n19006), .B1(n19005), .B2(n19004), .ZN(
        n19008) );
  NOR2_X1 U22093 ( .A1(n19009), .A2(n19008), .ZN(n19019) );
  AOI21_X1 U22094 ( .B1(n19012), .B2(n19011), .A(n19010), .ZN(n19014) );
  OAI211_X1 U22095 ( .C1(n19014), .C2(n19024), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19013), .ZN(n19016) );
  AOI21_X1 U22096 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19016), .A(n19015), 
        .ZN(n19018) );
  NAND2_X1 U22097 ( .A1(n19019), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19017) );
  OAI21_X1 U22098 ( .B1(n19019), .B2(n19018), .A(n19017), .ZN(P3_U3296) );
  OAI22_X1 U22099 ( .A1(n19020), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18999), .ZN(n19021) );
  INV_X1 U22100 ( .A(n19021), .ZN(P3_U3297) );
  OAI21_X1 U22101 ( .B1(n19022), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19023), 
        .ZN(n19027) );
  OAI22_X1 U22102 ( .A1(n19024), .A2(n19023), .B1(n19027), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n19025) );
  INV_X1 U22103 ( .A(n19025), .ZN(P3_U3298) );
  OAI21_X1 U22104 ( .B1(n19027), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19026), 
        .ZN(n19028) );
  INV_X1 U22105 ( .A(n19028), .ZN(P3_U3299) );
  INV_X1 U22106 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19030) );
  INV_X1 U22107 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19978) );
  NAND2_X1 U22108 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19978), .ZN(n19969) );
  NOR2_X1 U22109 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19965) );
  INV_X1 U22110 ( .A(n19965), .ZN(n19029) );
  OAI21_X1 U22111 ( .B1(n19959), .B2(n19969), .A(n19029), .ZN(n20052) );
  OAI21_X1 U22112 ( .B1(n19959), .B2(n19030), .A(n19957), .ZN(P2_U2815) );
  INV_X1 U22113 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19031) );
  OAI22_X1 U22114 ( .A1(n19034), .A2(n19033), .B1(n19032), .B2(n19031), .ZN(
        P2_U2816) );
  NAND2_X1 U22115 ( .A1(n20100), .A2(n19971), .ZN(n19960) );
  AOI21_X1 U22116 ( .B1(n19959), .B2(n19960), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19035) );
  AOI21_X1 U22117 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20036), .A(n19035), 
        .ZN(P2_U2817) );
  OAI21_X1 U22118 ( .B1(n19036), .B2(BS16), .A(n20052), .ZN(n20050) );
  OAI21_X1 U22119 ( .B1(n20052), .B2(n19627), .A(n20050), .ZN(P2_U2818) );
  NOR4_X1 U22120 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19040) );
  NOR4_X1 U22121 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19039) );
  NOR4_X1 U22122 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19038) );
  NOR4_X1 U22123 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19037) );
  NAND4_X1 U22124 ( .A1(n19040), .A2(n19039), .A3(n19038), .A4(n19037), .ZN(
        n19046) );
  NOR4_X1 U22125 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19044) );
  AOI211_X1 U22126 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19043) );
  NOR4_X1 U22127 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19042) );
  NOR4_X1 U22128 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19041) );
  NAND4_X1 U22129 ( .A1(n19044), .A2(n19043), .A3(n19042), .A4(n19041), .ZN(
        n19045) );
  NOR2_X1 U22130 ( .A1(n19046), .A2(n19045), .ZN(n19053) );
  INV_X1 U22131 ( .A(n19053), .ZN(n19052) );
  NOR2_X1 U22132 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19052), .ZN(n19047) );
  INV_X1 U22133 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20048) );
  AOI22_X1 U22134 ( .A1(n19047), .A2(n11840), .B1(n19052), .B2(n20048), .ZN(
        P2_U2820) );
  OR3_X1 U22135 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19051) );
  INV_X1 U22136 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20046) );
  AOI22_X1 U22137 ( .A1(n19047), .A2(n19051), .B1(n19052), .B2(n20046), .ZN(
        P2_U2821) );
  INV_X1 U22138 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20051) );
  NAND2_X1 U22139 ( .A1(n19047), .A2(n20051), .ZN(n19050) );
  INV_X1 U22140 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19979) );
  OAI21_X1 U22141 ( .B1(n11840), .B2(n19979), .A(n19053), .ZN(n19048) );
  OAI21_X1 U22142 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19053), .A(n19048), 
        .ZN(n19049) );
  OAI221_X1 U22143 ( .B1(n19050), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19050), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19049), .ZN(P2_U2822) );
  INV_X1 U22144 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20044) );
  OAI221_X1 U22145 ( .B1(n19053), .B2(n20044), .C1(n19052), .C2(n19051), .A(
        n19050), .ZN(P2_U2823) );
  AOI211_X1 U22146 ( .C1(n19055), .C2(n10344), .A(n19054), .B(n19953), .ZN(
        n19061) );
  AOI22_X1 U22147 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19248), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19244), .ZN(n19058) );
  AOI22_X1 U22148 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19245), .B1(
        n19056), .B2(n19247), .ZN(n19057) );
  OAI211_X1 U22149 ( .C1(n19059), .C2(n19232), .A(n19058), .B(n19057), .ZN(
        n19060) );
  AOI211_X1 U22150 ( .C1(n19249), .C2(n19062), .A(n19061), .B(n19060), .ZN(
        n19063) );
  INV_X1 U22151 ( .A(n19063), .ZN(P2_U2835) );
  AOI211_X1 U22152 ( .C1(n19066), .C2(n19065), .A(n19064), .B(n19953), .ZN(
        n19071) );
  AOI21_X1 U22153 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n19248), .A(n19412), 
        .ZN(n19068) );
  AOI22_X1 U22154 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19245), .ZN(n19067) );
  OAI211_X1 U22155 ( .C1(n19069), .C2(n19233), .A(n19068), .B(n19067), .ZN(
        n19070) );
  AOI211_X1 U22156 ( .C1(n19249), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        n19073) );
  OAI21_X1 U22157 ( .B1(n19074), .B2(n19232), .A(n19073), .ZN(P2_U2836) );
  AOI211_X1 U22158 ( .C1(n19076), .C2(n19090), .A(n19075), .B(n19953), .ZN(
        n19081) );
  AOI21_X1 U22159 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n19248), .A(n19412), 
        .ZN(n19078) );
  AOI22_X1 U22160 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19244), .ZN(n19077) );
  OAI211_X1 U22161 ( .C1(n19079), .C2(n19233), .A(n19078), .B(n19077), .ZN(
        n19080) );
  AOI211_X1 U22162 ( .C1(n19249), .C2(n19082), .A(n19081), .B(n19080), .ZN(
        n19083) );
  OAI21_X1 U22163 ( .B1(n19084), .B2(n19232), .A(n19083), .ZN(P2_U2837) );
  INV_X1 U22164 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20011) );
  AOI22_X1 U22165 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19245), .ZN(n19085) );
  OAI211_X1 U22166 ( .C1(n20011), .C2(n19183), .A(n19085), .B(n16334), .ZN(
        n19088) );
  OAI22_X1 U22167 ( .A1(n19086), .A2(n19233), .B1(n19091), .B2(n19141), .ZN(
        n19087) );
  AOI211_X1 U22168 ( .C1(n19089), .C2(n19251), .A(n19088), .B(n19087), .ZN(
        n19094) );
  OAI211_X1 U22169 ( .C1(n19092), .C2(n19091), .A(n19226), .B(n19090), .ZN(
        n19093) );
  OAI211_X1 U22170 ( .C1(n19230), .C2(n19095), .A(n19094), .B(n19093), .ZN(
        P2_U2838) );
  INV_X1 U22171 ( .A(n19096), .ZN(n19101) );
  INV_X1 U22172 ( .A(n19097), .ZN(n19103) );
  OAI211_X1 U22173 ( .C1(n9835), .C2(n19103), .A(n19226), .B(n19098), .ZN(
        n19100) );
  AOI22_X1 U22174 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19244), .ZN(n19099) );
  OAI211_X1 U22175 ( .C1(n19101), .C2(n19233), .A(n19100), .B(n19099), .ZN(
        n19102) );
  AOI211_X1 U22176 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19248), .A(n19412), 
        .B(n19102), .ZN(n19107) );
  NOR3_X1 U22177 ( .A1(n9835), .A2(n19103), .A3(n19953), .ZN(n19115) );
  AOI22_X1 U22178 ( .A1(n19105), .A2(n19249), .B1(n19115), .B2(n19104), .ZN(
        n19106) );
  OAI211_X1 U22179 ( .C1(n19108), .C2(n19232), .A(n19107), .B(n19106), .ZN(
        P2_U2839) );
  OAI22_X1 U22180 ( .A1(n19110), .A2(n12744), .B1(n19109), .B2(n19185), .ZN(
        n19111) );
  AOI211_X1 U22181 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19248), .A(n19412), 
        .B(n19111), .ZN(n19121) );
  AOI22_X1 U22182 ( .A1(n19113), .A2(n19247), .B1(n19112), .B2(n19256), .ZN(
        n19120) );
  AOI22_X1 U22183 ( .A1(n19114), .A2(n19249), .B1(n19271), .B2(n19251), .ZN(
        n19119) );
  OAI21_X1 U22184 ( .B1(n19117), .B2(n19116), .A(n19115), .ZN(n19118) );
  NAND4_X1 U22185 ( .A1(n19121), .A2(n19120), .A3(n19119), .A4(n19118), .ZN(
        P2_U2840) );
  AOI22_X1 U22186 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19245), .B1(
        n19122), .B2(n19247), .ZN(n19123) );
  OAI211_X1 U22187 ( .C1(n20005), .C2(n19183), .A(n19123), .B(n16334), .ZN(
        n19124) );
  AOI21_X1 U22188 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19189), .A(n19124), .ZN(
        n19130) );
  NAND2_X1 U22189 ( .A1(n9831), .A2(n19131), .ZN(n19125) );
  XNOR2_X1 U22190 ( .A(n19126), .B(n19125), .ZN(n19127) );
  AOI22_X1 U22191 ( .A1(n19128), .A2(n19249), .B1(n19226), .B2(n19127), .ZN(
        n19129) );
  OAI211_X1 U22192 ( .C1(n19274), .C2(n19232), .A(n19130), .B(n19129), .ZN(
        P2_U2841) );
  AOI22_X1 U22193 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19245), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19244), .ZN(n19135) );
  NOR2_X1 U22194 ( .A1(n9835), .A2(n19953), .ZN(n19132) );
  OAI211_X1 U22195 ( .C1(n19133), .C2(n19142), .A(n19132), .B(n19131), .ZN(
        n19134) );
  OAI211_X1 U22196 ( .C1(n19233), .C2(n19136), .A(n19135), .B(n19134), .ZN(
        n19137) );
  AOI211_X1 U22197 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19248), .A(n19412), 
        .B(n19137), .ZN(n19140) );
  AOI22_X1 U22198 ( .A1(n19138), .A2(n19249), .B1(n19275), .B2(n19251), .ZN(
        n19139) );
  OAI211_X1 U22199 ( .C1(n19142), .C2(n19141), .A(n19140), .B(n19139), .ZN(
        P2_U2842) );
  AOI22_X1 U22200 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19245), .B1(
        n19143), .B2(n19247), .ZN(n19144) );
  OAI211_X1 U22201 ( .C1(n20001), .C2(n19183), .A(n19144), .B(n16334), .ZN(
        n19145) );
  AOI21_X1 U22202 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19189), .A(n19145), .ZN(
        n19152) );
  NAND2_X1 U22203 ( .A1(n9831), .A2(n19146), .ZN(n19147) );
  XNOR2_X1 U22204 ( .A(n19148), .B(n19147), .ZN(n19149) );
  AOI22_X1 U22205 ( .A1(n19150), .A2(n19249), .B1(n19226), .B2(n19149), .ZN(
        n19151) );
  OAI211_X1 U22206 ( .C1(n19277), .C2(n19232), .A(n19152), .B(n19151), .ZN(
        P2_U2843) );
  AOI22_X1 U22207 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19244), .ZN(n19153) );
  OAI21_X1 U22208 ( .B1(n19154), .B2(n19233), .A(n19153), .ZN(n19155) );
  AOI211_X1 U22209 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19248), .A(n19412), 
        .B(n19155), .ZN(n19161) );
  NOR2_X1 U22210 ( .A1(n9835), .A2(n19156), .ZN(n19158) );
  XNOR2_X1 U22211 ( .A(n19158), .B(n19157), .ZN(n19159) );
  AOI22_X1 U22212 ( .A1(n19279), .A2(n19251), .B1(n19226), .B2(n19159), .ZN(
        n19160) );
  OAI211_X1 U22213 ( .C1(n19162), .C2(n19230), .A(n19161), .B(n19160), .ZN(
        P2_U2844) );
  AOI22_X1 U22214 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19245), .B1(
        n19163), .B2(n19247), .ZN(n19164) );
  OAI211_X1 U22215 ( .C1(n19997), .C2(n19183), .A(n19164), .B(n16334), .ZN(
        n19165) );
  AOI21_X1 U22216 ( .B1(P2_EBX_REG_10__SCAN_IN), .B2(n19189), .A(n19165), .ZN(
        n19172) );
  NAND2_X1 U22217 ( .A1(n9831), .A2(n19166), .ZN(n19167) );
  XNOR2_X1 U22218 ( .A(n19168), .B(n19167), .ZN(n19169) );
  AOI22_X1 U22219 ( .A1(n19170), .A2(n19249), .B1(n19226), .B2(n19169), .ZN(
        n19171) );
  OAI211_X1 U22220 ( .C1(n19281), .C2(n19232), .A(n19172), .B(n19171), .ZN(
        P2_U2845) );
  AOI22_X1 U22221 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_9__SCAN_IN), .B2(n19244), .ZN(n19173) );
  OAI21_X1 U22222 ( .B1(n19174), .B2(n19233), .A(n19173), .ZN(n19175) );
  AOI211_X1 U22223 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19248), .A(n19412), .B(
        n19175), .ZN(n19181) );
  NOR2_X1 U22224 ( .A1(n9835), .A2(n19176), .ZN(n19178) );
  XNOR2_X1 U22225 ( .A(n19178), .B(n19177), .ZN(n19179) );
  AOI22_X1 U22226 ( .A1(n19251), .A2(n19283), .B1(n19226), .B2(n19179), .ZN(
        n19180) );
  OAI211_X1 U22227 ( .C1(n19230), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        P2_U2846) );
  OAI21_X1 U22228 ( .B1(n19993), .B2(n19183), .A(n16334), .ZN(n19188) );
  OAI22_X1 U22229 ( .A1(n19186), .A2(n19185), .B1(n19184), .B2(n19233), .ZN(
        n19187) );
  AOI211_X1 U22230 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19189), .A(n19188), .B(
        n19187), .ZN(n19196) );
  NAND2_X1 U22231 ( .A1(n9831), .A2(n19190), .ZN(n19191) );
  XNOR2_X1 U22232 ( .A(n19192), .B(n19191), .ZN(n19194) );
  AOI22_X1 U22233 ( .A1(n19226), .A2(n19194), .B1(n19249), .B2(n19193), .ZN(
        n19195) );
  OAI211_X1 U22234 ( .C1(n19232), .C2(n19288), .A(n19196), .B(n19195), .ZN(
        P2_U2847) );
  AOI22_X1 U22235 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_7__SCAN_IN), .B2(n19244), .ZN(n19197) );
  OAI21_X1 U22236 ( .B1(n19198), .B2(n19233), .A(n19197), .ZN(n19199) );
  AOI211_X1 U22237 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n19248), .A(n19412), .B(
        n19199), .ZN(n19205) );
  NOR2_X1 U22238 ( .A1(n9835), .A2(n19200), .ZN(n19202) );
  XNOR2_X1 U22239 ( .A(n19202), .B(n19201), .ZN(n19203) );
  AOI22_X1 U22240 ( .A1(n19251), .A2(n19290), .B1(n19226), .B2(n19203), .ZN(
        n19204) );
  OAI211_X1 U22241 ( .C1(n19230), .C2(n19206), .A(n19205), .B(n19204), .ZN(
        P2_U2848) );
  AOI22_X1 U22242 ( .A1(P2_EBX_REG_6__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19245), .ZN(n19207) );
  OAI21_X1 U22243 ( .B1(n19208), .B2(n19233), .A(n19207), .ZN(n19209) );
  AOI211_X1 U22244 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19248), .A(n19412), .B(
        n19209), .ZN(n19215) );
  NAND2_X1 U22245 ( .A1(n9831), .A2(n19210), .ZN(n19211) );
  XNOR2_X1 U22246 ( .A(n19212), .B(n19211), .ZN(n19213) );
  AOI22_X1 U22247 ( .A1(n19251), .A2(n19292), .B1(n19226), .B2(n19213), .ZN(
        n19214) );
  OAI211_X1 U22248 ( .C1(n19230), .C2(n19216), .A(n19215), .B(n19214), .ZN(
        P2_U2849) );
  AOI22_X1 U22249 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19217), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19244), .ZN(n19218) );
  OAI21_X1 U22250 ( .B1(n19219), .B2(n19233), .A(n19218), .ZN(n19220) );
  AOI211_X1 U22251 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19248), .A(n19412), .B(
        n19220), .ZN(n19228) );
  NOR2_X1 U22252 ( .A1(n9835), .A2(n19221), .ZN(n19224) );
  XNOR2_X1 U22253 ( .A(n19224), .B(n19223), .ZN(n19225) );
  AOI22_X1 U22254 ( .A1(n19251), .A2(n19295), .B1(n19226), .B2(n19225), .ZN(
        n19227) );
  OAI211_X1 U22255 ( .C1(n19230), .C2(n19229), .A(n19228), .B(n19227), .ZN(
        P2_U2850) );
  AOI22_X1 U22256 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19244), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19245), .ZN(n19243) );
  OAI22_X1 U22257 ( .A1(n19234), .A2(n19233), .B1(n19232), .B2(n19231), .ZN(
        n19235) );
  AOI211_X1 U22258 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19248), .A(n19412), .B(
        n19235), .ZN(n19242) );
  INV_X1 U22259 ( .A(n19236), .ZN(n19296) );
  AOI22_X1 U22260 ( .A1(n19296), .A2(n19258), .B1(n19419), .B2(n19249), .ZN(
        n19241) );
  AND2_X1 U22261 ( .A1(n9831), .A2(n19237), .ZN(n19239) );
  AOI21_X1 U22262 ( .B1(n19410), .B2(n19239), .A(n19953), .ZN(n19238) );
  OAI21_X1 U22263 ( .B1(n19410), .B2(n19239), .A(n19238), .ZN(n19240) );
  NAND4_X1 U22264 ( .A1(n19243), .A2(n19242), .A3(n19241), .A4(n19240), .ZN(
        P2_U2851) );
  AOI22_X1 U22265 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19245), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19244), .ZN(n19255) );
  AOI22_X1 U22266 ( .A1(n19248), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n19247), 
        .B2(n19246), .ZN(n19254) );
  NAND2_X1 U22267 ( .A1(n19250), .A2(n19249), .ZN(n19253) );
  NAND2_X1 U22268 ( .A1(n19251), .A2(n20076), .ZN(n19252) );
  AND4_X1 U22269 ( .A1(n19255), .A2(n19254), .A3(n19253), .A4(n19252), .ZN(
        n19260) );
  AOI22_X1 U22270 ( .A1(n20072), .A2(n19258), .B1(n19257), .B2(n19256), .ZN(
        n19259) );
  OAI211_X1 U22271 ( .C1(n19953), .C2(n19261), .A(n19260), .B(n19259), .ZN(
        P2_U2854) );
  AOI22_X1 U22272 ( .A1(n19263), .A2(n19318), .B1(n19262), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19266) );
  AOI22_X1 U22273 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19264), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19317), .ZN(n19265) );
  NAND2_X1 U22274 ( .A1(n19266), .A2(n19265), .ZN(P2_U2888) );
  AOI22_X1 U22275 ( .A1(n19268), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19267), .ZN(n19409) );
  AOI22_X1 U22276 ( .A1(n19271), .A2(n19294), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n19317), .ZN(n19272) );
  OAI21_X1 U22277 ( .B1(n19325), .B2(n19409), .A(n19272), .ZN(P2_U2904) );
  AOI22_X1 U22278 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19317), .B1(n19382), 
        .B2(n19285), .ZN(n19273) );
  OAI21_X1 U22279 ( .B1(n19289), .B2(n19274), .A(n19273), .ZN(P2_U2905) );
  INV_X1 U22280 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19341) );
  AOI22_X1 U22281 ( .A1(n19275), .A2(n19294), .B1(n19380), .B2(n19285), .ZN(
        n19276) );
  OAI21_X1 U22282 ( .B1(n19282), .B2(n19341), .A(n19276), .ZN(P2_U2906) );
  INV_X1 U22283 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19343) );
  OAI222_X1 U22284 ( .A1(n19343), .A2(n19282), .B1(n19277), .B2(n19289), .C1(
        n19325), .C2(n19400), .ZN(P2_U2907) );
  AOI22_X1 U22285 ( .A1(n19279), .A2(n19294), .B1(n19278), .B2(n19285), .ZN(
        n19280) );
  OAI21_X1 U22286 ( .B1(n19282), .B2(n12564), .A(n19280), .ZN(P2_U2908) );
  INV_X1 U22287 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19346) );
  OAI222_X1 U22288 ( .A1(n19346), .A2(n19282), .B1(n19281), .B2(n19289), .C1(
        n19325), .C2(n19398), .ZN(P2_U2909) );
  AOI22_X1 U22289 ( .A1(n19283), .A2(n19294), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19317), .ZN(n19284) );
  OAI21_X1 U22290 ( .B1(n19396), .B2(n19325), .A(n19284), .ZN(P2_U2910) );
  AOI22_X1 U22291 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19317), .B1(n19286), .B2(
        n19285), .ZN(n19287) );
  OAI21_X1 U22292 ( .B1(n19289), .B2(n19288), .A(n19287), .ZN(P2_U2911) );
  AOI22_X1 U22293 ( .A1(n19290), .A2(n19294), .B1(P2_EAX_REG_7__SCAN_IN), .B2(
        n19317), .ZN(n19291) );
  OAI21_X1 U22294 ( .B1(n19472), .B2(n19325), .A(n19291), .ZN(P2_U2912) );
  AOI22_X1 U22295 ( .A1(n19292), .A2(n19294), .B1(P2_EAX_REG_6__SCAN_IN), .B2(
        n19317), .ZN(n19293) );
  OAI21_X1 U22296 ( .B1(n19461), .B2(n19325), .A(n19293), .ZN(P2_U2913) );
  AOI22_X1 U22297 ( .A1(n19295), .A2(n19294), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19317), .ZN(n19299) );
  NAND3_X1 U22298 ( .A1(n19297), .A2(n19296), .A3(n19319), .ZN(n19298) );
  OAI211_X1 U22299 ( .C1(n19457), .C2(n19325), .A(n19299), .B(n19298), .ZN(
        P2_U2914) );
  AOI22_X1 U22300 ( .A1(n19318), .A2(n20058), .B1(n19317), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19305) );
  OAI21_X1 U22301 ( .B1(n19302), .B2(n19301), .A(n19300), .ZN(n19303) );
  NAND2_X1 U22302 ( .A1(n19303), .A2(n19319), .ZN(n19304) );
  OAI211_X1 U22303 ( .C1(n19446), .C2(n19325), .A(n19305), .B(n19304), .ZN(
        P2_U2916) );
  AOI22_X1 U22304 ( .A1(n19318), .A2(n20067), .B1(n19317), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19311) );
  OAI21_X1 U22305 ( .B1(n19308), .B2(n19307), .A(n19306), .ZN(n19309) );
  NAND2_X1 U22306 ( .A1(n19309), .A2(n19319), .ZN(n19310) );
  OAI211_X1 U22307 ( .C1(n19440), .C2(n19325), .A(n19311), .B(n19310), .ZN(
        P2_U2917) );
  AOI22_X1 U22308 ( .A1(n19318), .A2(n20076), .B1(n19317), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19316) );
  OAI21_X1 U22309 ( .B1(n19313), .B2(n19320), .A(n19312), .ZN(n19314) );
  NAND2_X1 U22310 ( .A1(n19314), .A2(n19319), .ZN(n19315) );
  OAI211_X1 U22311 ( .C1(n19388), .C2(n19325), .A(n19316), .B(n19315), .ZN(
        P2_U2918) );
  AOI22_X1 U22312 ( .A1(n19318), .A2(n19321), .B1(n19317), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19324) );
  OAI211_X1 U22313 ( .C1(n19322), .C2(n19321), .A(n19320), .B(n19319), .ZN(
        n19323) );
  OAI211_X1 U22314 ( .C1(n19386), .C2(n19325), .A(n19324), .B(n19323), .ZN(
        P2_U2919) );
  NOR2_X1 U22315 ( .A1(n19333), .A2(n19326), .ZN(P2_U2920) );
  INV_X1 U22316 ( .A(n19327), .ZN(n19330) );
  AOI22_X1 U22317 ( .A1(n19330), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19366), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19328) );
  OAI21_X1 U22318 ( .B1(n19329), .B2(n19333), .A(n19328), .ZN(P2_U2921) );
  AOI22_X1 U22319 ( .A1(n19330), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19366), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19331) );
  OAI21_X1 U22320 ( .B1(n19333), .B2(n19332), .A(n19331), .ZN(P2_U2922) );
  INV_X1 U22321 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19337) );
  AOI22_X1 U22322 ( .A1(n19335), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19336) );
  OAI21_X1 U22323 ( .B1(n19337), .B2(n19368), .A(n19336), .ZN(P2_U2936) );
  INV_X1 U22324 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19339) );
  AOI22_X1 U22325 ( .A1(n19366), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19338) );
  OAI21_X1 U22326 ( .B1(n19339), .B2(n19368), .A(n19338), .ZN(P2_U2937) );
  AOI22_X1 U22327 ( .A1(n19366), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19340) );
  OAI21_X1 U22328 ( .B1(n19341), .B2(n19368), .A(n19340), .ZN(P2_U2938) );
  AOI22_X1 U22329 ( .A1(n19366), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19342) );
  OAI21_X1 U22330 ( .B1(n19343), .B2(n19368), .A(n19342), .ZN(P2_U2939) );
  AOI22_X1 U22331 ( .A1(n19366), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19344) );
  OAI21_X1 U22332 ( .B1(n12564), .B2(n19368), .A(n19344), .ZN(P2_U2940) );
  AOI22_X1 U22333 ( .A1(n19366), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19345) );
  OAI21_X1 U22334 ( .B1(n19346), .B2(n19368), .A(n19345), .ZN(P2_U2941) );
  INV_X1 U22335 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19348) );
  AOI22_X1 U22336 ( .A1(n19366), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19347) );
  OAI21_X1 U22337 ( .B1(n19348), .B2(n19368), .A(n19347), .ZN(P2_U2942) );
  AOI22_X1 U22338 ( .A1(n19366), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19349) );
  OAI21_X1 U22339 ( .B1(n19350), .B2(n19368), .A(n19349), .ZN(P2_U2943) );
  INV_X1 U22340 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19352) );
  AOI22_X1 U22341 ( .A1(n19366), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19351) );
  OAI21_X1 U22342 ( .B1(n19352), .B2(n19368), .A(n19351), .ZN(P2_U2944) );
  INV_X1 U22343 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19354) );
  AOI22_X1 U22344 ( .A1(n19366), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19353) );
  OAI21_X1 U22345 ( .B1(n19354), .B2(n19368), .A(n19353), .ZN(P2_U2945) );
  INV_X1 U22346 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19356) );
  AOI22_X1 U22347 ( .A1(n19366), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19355) );
  OAI21_X1 U22348 ( .B1(n19356), .B2(n19368), .A(n19355), .ZN(P2_U2946) );
  INV_X1 U22349 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19358) );
  AOI22_X1 U22350 ( .A1(n19366), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19357) );
  OAI21_X1 U22351 ( .B1(n19358), .B2(n19368), .A(n19357), .ZN(P2_U2947) );
  INV_X1 U22352 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19360) );
  AOI22_X1 U22353 ( .A1(n19366), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19359) );
  OAI21_X1 U22354 ( .B1(n19360), .B2(n19368), .A(n19359), .ZN(P2_U2948) );
  INV_X1 U22355 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19362) );
  AOI22_X1 U22356 ( .A1(n19366), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19361) );
  OAI21_X1 U22357 ( .B1(n19362), .B2(n19368), .A(n19361), .ZN(P2_U2949) );
  INV_X1 U22358 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19365) );
  AOI22_X1 U22359 ( .A1(n19366), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19364) );
  OAI21_X1 U22360 ( .B1(n19365), .B2(n19368), .A(n19364), .ZN(P2_U2950) );
  AOI22_X1 U22361 ( .A1(n19366), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19363), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19367) );
  OAI21_X1 U22362 ( .B1(n12449), .B2(n19368), .A(n19367), .ZN(P2_U2951) );
  AOI22_X1 U22363 ( .A1(n19406), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n19369) );
  OAI21_X1 U22364 ( .B1(n19386), .B2(n19408), .A(n19369), .ZN(P2_U2952) );
  AOI22_X1 U22365 ( .A1(n19406), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19405), .ZN(n19370) );
  OAI21_X1 U22366 ( .B1(n19388), .B2(n19408), .A(n19370), .ZN(P2_U2953) );
  AOI22_X1 U22367 ( .A1(n19406), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n19371) );
  OAI21_X1 U22368 ( .B1(n19440), .B2(n19408), .A(n19371), .ZN(P2_U2954) );
  AOI22_X1 U22369 ( .A1(n19406), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19405), .ZN(n19372) );
  OAI21_X1 U22370 ( .B1(n19446), .B2(n19408), .A(n19372), .ZN(P2_U2955) );
  AOI22_X1 U22371 ( .A1(n19406), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n19373) );
  OAI21_X1 U22372 ( .B1(n19453), .B2(n19408), .A(n19373), .ZN(P2_U2956) );
  AOI22_X1 U22373 ( .A1(n19406), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19405), .ZN(n19374) );
  OAI21_X1 U22374 ( .B1(n19457), .B2(n19408), .A(n19374), .ZN(P2_U2957) );
  AOI22_X1 U22375 ( .A1(n19406), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n19375) );
  OAI21_X1 U22376 ( .B1(n19461), .B2(n19408), .A(n19375), .ZN(P2_U2958) );
  AOI22_X1 U22377 ( .A1(n19406), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19405), .ZN(n19376) );
  OAI21_X1 U22378 ( .B1(n19472), .B2(n19408), .A(n19376), .ZN(P2_U2959) );
  AOI22_X1 U22379 ( .A1(n19406), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19405), .ZN(n19377) );
  OAI21_X1 U22380 ( .B1(n19396), .B2(n19408), .A(n19377), .ZN(P2_U2961) );
  AOI22_X1 U22381 ( .A1(n19406), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n19405), .ZN(n19378) );
  OAI21_X1 U22382 ( .B1(n19398), .B2(n19408), .A(n19378), .ZN(P2_U2962) );
  AOI22_X1 U22383 ( .A1(n19406), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19405), .ZN(n19379) );
  OAI21_X1 U22384 ( .B1(n19400), .B2(n19408), .A(n19379), .ZN(P2_U2964) );
  AOI22_X1 U22385 ( .A1(n19406), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19405), .ZN(n19381) );
  NAND2_X1 U22386 ( .A1(n19383), .A2(n19380), .ZN(n19401) );
  NAND2_X1 U22387 ( .A1(n19381), .A2(n19401), .ZN(P2_U2965) );
  AOI22_X1 U22388 ( .A1(n19406), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19405), .ZN(n19384) );
  NAND2_X1 U22389 ( .A1(n19383), .A2(n19382), .ZN(n19403) );
  NAND2_X1 U22390 ( .A1(n19384), .A2(n19403), .ZN(P2_U2966) );
  AOI22_X1 U22391 ( .A1(n19406), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19405), .ZN(n19385) );
  OAI21_X1 U22392 ( .B1(n19386), .B2(n19408), .A(n19385), .ZN(P2_U2967) );
  AOI22_X1 U22393 ( .A1(n19406), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n19405), .ZN(n19387) );
  OAI21_X1 U22394 ( .B1(n19388), .B2(n19408), .A(n19387), .ZN(P2_U2968) );
  AOI22_X1 U22395 ( .A1(n19406), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19405), .ZN(n19389) );
  OAI21_X1 U22396 ( .B1(n19440), .B2(n19408), .A(n19389), .ZN(P2_U2969) );
  AOI22_X1 U22397 ( .A1(n19406), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19405), .ZN(n19390) );
  OAI21_X1 U22398 ( .B1(n19446), .B2(n19408), .A(n19390), .ZN(P2_U2970) );
  AOI22_X1 U22399 ( .A1(n19406), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19405), .ZN(n19391) );
  OAI21_X1 U22400 ( .B1(n19453), .B2(n19408), .A(n19391), .ZN(P2_U2971) );
  AOI22_X1 U22401 ( .A1(n19406), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19405), .ZN(n19392) );
  OAI21_X1 U22402 ( .B1(n19457), .B2(n19408), .A(n19392), .ZN(P2_U2972) );
  AOI22_X1 U22403 ( .A1(n19406), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n19405), .ZN(n19393) );
  OAI21_X1 U22404 ( .B1(n19461), .B2(n19408), .A(n19393), .ZN(P2_U2973) );
  AOI22_X1 U22405 ( .A1(n19406), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n19405), .ZN(n19394) );
  OAI21_X1 U22406 ( .B1(n19472), .B2(n19408), .A(n19394), .ZN(P2_U2974) );
  AOI22_X1 U22407 ( .A1(n19406), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19405), .ZN(n19395) );
  OAI21_X1 U22408 ( .B1(n19396), .B2(n19408), .A(n19395), .ZN(P2_U2976) );
  AOI22_X1 U22409 ( .A1(n19406), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n19405), .ZN(n19397) );
  OAI21_X1 U22410 ( .B1(n19398), .B2(n19408), .A(n19397), .ZN(P2_U2977) );
  AOI22_X1 U22411 ( .A1(n19406), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19405), .ZN(n19399) );
  OAI21_X1 U22412 ( .B1(n19400), .B2(n19408), .A(n19399), .ZN(P2_U2979) );
  AOI22_X1 U22413 ( .A1(n19406), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n19402) );
  NAND2_X1 U22414 ( .A1(n19402), .A2(n19401), .ZN(P2_U2980) );
  AOI22_X1 U22415 ( .A1(n19406), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19405), .ZN(n19404) );
  NAND2_X1 U22416 ( .A1(n19404), .A2(n19403), .ZN(P2_U2981) );
  AOI22_X1 U22417 ( .A1(n19406), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19405), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n19407) );
  OAI21_X1 U22418 ( .B1(n19409), .B2(n19408), .A(n19407), .ZN(P2_U2982) );
  AOI22_X1 U22419 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19412), .B1(n19411), 
        .B2(n19410), .ZN(n19422) );
  INV_X1 U22420 ( .A(n19413), .ZN(n19417) );
  OAI22_X1 U22421 ( .A1(n19417), .A2(n19416), .B1(n19415), .B2(n19414), .ZN(
        n19418) );
  AOI21_X1 U22422 ( .B1(n19420), .B2(n19419), .A(n19418), .ZN(n19421) );
  OAI211_X1 U22423 ( .C1(n19424), .C2(n19423), .A(n19422), .B(n19421), .ZN(
        P2_U3010) );
  NAND2_X1 U22424 ( .A1(n19538), .A2(n20078), .ZN(n19482) );
  NOR2_X1 U22425 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19482), .ZN(
        n19471) );
  AOI22_X1 U22426 ( .A1(n19832), .A2(n19942), .B1(n19856), .B2(n19471), .ZN(
        n19434) );
  AOI21_X1 U22427 ( .B1(n19926), .B2(n19486), .A(n19627), .ZN(n19425) );
  NOR2_X1 U22428 ( .A1(n19425), .A2(n19861), .ZN(n19429) );
  INV_X1 U22429 ( .A(n13648), .ZN(n19430) );
  OAI21_X1 U22430 ( .B1(n19430), .B2(n19822), .A(n20079), .ZN(n19426) );
  AOI21_X1 U22431 ( .B1(n19429), .B2(n19427), .A(n19426), .ZN(n19428) );
  OAI21_X1 U22432 ( .B1(n19428), .B2(n19471), .A(n19863), .ZN(n19474) );
  OAI21_X1 U22433 ( .B1(n19938), .B2(n19471), .A(n19429), .ZN(n19432) );
  OAI21_X1 U22434 ( .B1(n19430), .B2(n19471), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19431) );
  NAND2_X1 U22435 ( .A1(n19432), .A2(n19431), .ZN(n19473) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19474), .B1(
        n13210), .B2(n19473), .ZN(n19433) );
  OAI211_X1 U22437 ( .C1(n19835), .C2(n19486), .A(n19434), .B(n19433), .ZN(
        P2_U3048) );
  AOI22_X1 U22438 ( .A1(n19900), .A2(n19942), .B1(n19899), .B2(n19471), .ZN(
        n19436) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19474), .B1(
        n13231), .B2(n19473), .ZN(n19435) );
  OAI211_X1 U22440 ( .C1(n19903), .C2(n19486), .A(n19436), .B(n19435), .ZN(
        P2_U3049) );
  AOI22_X1 U22441 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19464), .ZN(n19841) );
  OAI22_X2 U22442 ( .A1(n19438), .A2(n19468), .B1(n19437), .B2(n19466), .ZN(
        n19838) );
  NOR2_X2 U22443 ( .A1(n19439), .A2(n19470), .ZN(n19904) );
  AOI22_X1 U22444 ( .A1(n19838), .A2(n19942), .B1(n19904), .B2(n19471), .ZN(
        n19443) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19474), .B1(
        n19441), .B2(n19473), .ZN(n19442) );
  OAI211_X1 U22446 ( .C1(n19841), .C2(n19486), .A(n19443), .B(n19442), .ZN(
        P2_U3050) );
  AOI22_X1 U22447 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19464), .ZN(n19878) );
  OAI22_X2 U22448 ( .A1(n19445), .A2(n19466), .B1(n19444), .B2(n19468), .ZN(
        n19910) );
  NOR2_X2 U22449 ( .A1(n11792), .A2(n19470), .ZN(n19909) );
  AOI22_X1 U22450 ( .A1(n19910), .A2(n19942), .B1(n19909), .B2(n19471), .ZN(
        n19449) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19474), .B1(
        n19447), .B2(n19473), .ZN(n19448) );
  OAI211_X1 U22452 ( .C1(n19878), .C2(n19486), .A(n19449), .B(n19448), .ZN(
        P2_U3051) );
  AOI22_X1 U22453 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19464), .ZN(n19882) );
  NOR2_X2 U22454 ( .A1(n19452), .A2(n19470), .ZN(n19915) );
  AOI22_X1 U22455 ( .A1(n19879), .A2(n19942), .B1(n19915), .B2(n19471), .ZN(
        n19455) );
  NOR2_X2 U22456 ( .A1(n19453), .A2(n19826), .ZN(n19916) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19474), .B1(
        n19916), .B2(n19473), .ZN(n19454) );
  OAI211_X1 U22458 ( .C1(n19882), .C2(n19486), .A(n19455), .B(n19454), .ZN(
        P2_U3052) );
  AOI22_X1 U22459 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19464), .ZN(n19927) );
  OAI22_X2 U22460 ( .A1(n20364), .A2(n19468), .B1(n19456), .B2(n19466), .ZN(
        n19923) );
  NOR2_X2 U22461 ( .A1(n12683), .A2(n19470), .ZN(n19921) );
  AOI22_X1 U22462 ( .A1(n19923), .A2(n19942), .B1(n19921), .B2(n19471), .ZN(
        n19459) );
  NOR2_X2 U22463 ( .A1(n19457), .A2(n19826), .ZN(n19922) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19474), .B1(
        n19922), .B2(n19473), .ZN(n19458) );
  OAI211_X1 U22465 ( .C1(n19927), .C2(n19486), .A(n19459), .B(n19458), .ZN(
        P2_U3053) );
  AOI22_X1 U22466 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19464), .ZN(n19890) );
  OAI22_X2 U22467 ( .A1(n19460), .A2(n19466), .B1(n20372), .B2(n19468), .ZN(
        n19930) );
  NOR2_X2 U22468 ( .A1(n11868), .A2(n19470), .ZN(n19928) );
  AOI22_X1 U22469 ( .A1(n19930), .A2(n19942), .B1(n19928), .B2(n19471), .ZN(
        n19463) );
  NOR2_X2 U22470 ( .A1(n19461), .A2(n19826), .ZN(n19929) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19474), .B1(
        n19929), .B2(n19473), .ZN(n19462) );
  OAI211_X1 U22472 ( .C1(n19890), .C2(n19486), .A(n19463), .B(n19462), .ZN(
        P2_U3054) );
  AOI22_X1 U22473 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19465), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19464), .ZN(n19898) );
  OAI22_X2 U22474 ( .A1(n19469), .A2(n19468), .B1(n19467), .B2(n19466), .ZN(
        n19893) );
  NOR2_X2 U22475 ( .A1(n11744), .A2(n19470), .ZN(n19937) );
  AOI22_X1 U22476 ( .A1(n19893), .A2(n19942), .B1(n19937), .B2(n19471), .ZN(
        n19476) );
  NOR2_X2 U22477 ( .A1(n19472), .A2(n19826), .ZN(n19940) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19474), .B1(
        n19940), .B2(n19473), .ZN(n19475) );
  OAI211_X1 U22479 ( .C1(n19898), .C2(n19486), .A(n19476), .B(n19475), .ZN(
        P2_U3055) );
  INV_X1 U22480 ( .A(n19478), .ZN(n19480) );
  NOR2_X1 U22481 ( .A1(n19479), .A2(n19540), .ZN(n19501) );
  OAI21_X1 U22482 ( .B1(n19480), .B2(n19501), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19481) );
  OAI21_X1 U22483 ( .B1(n19482), .B2(n19861), .A(n19481), .ZN(n19502) );
  AOI22_X1 U22484 ( .A1(n19502), .A2(n13210), .B1(n19856), .B2(n19501), .ZN(
        n19488) );
  AOI21_X1 U22485 ( .B1(n19478), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19485) );
  OAI21_X1 U22486 ( .B1(n19660), .B2(n19483), .A(n19482), .ZN(n19484) );
  OAI211_X1 U22487 ( .C1(n19501), .C2(n19485), .A(n19484), .B(n19863), .ZN(
        n19504) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19832), .ZN(n19487) );
  OAI211_X1 U22489 ( .C1(n19835), .C2(n19536), .A(n19488), .B(n19487), .ZN(
        P2_U3056) );
  AOI22_X1 U22490 ( .A1(n19502), .A2(n13231), .B1(n19899), .B2(n19501), .ZN(
        n19490) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19900), .ZN(n19489) );
  OAI211_X1 U22492 ( .C1(n19903), .C2(n19536), .A(n19490), .B(n19489), .ZN(
        P2_U3057) );
  AOI22_X1 U22493 ( .A1(n19502), .A2(n19441), .B1(n19904), .B2(n19501), .ZN(
        n19492) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19838), .ZN(n19491) );
  OAI211_X1 U22495 ( .C1(n19841), .C2(n19536), .A(n19492), .B(n19491), .ZN(
        P2_U3058) );
  AOI22_X1 U22496 ( .A1(n19502), .A2(n19447), .B1(n19909), .B2(n19501), .ZN(
        n19494) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19910), .ZN(n19493) );
  OAI211_X1 U22498 ( .C1(n19878), .C2(n19536), .A(n19494), .B(n19493), .ZN(
        P2_U3059) );
  AOI22_X1 U22499 ( .A1(n19502), .A2(n19916), .B1(n19915), .B2(n19501), .ZN(
        n19496) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19879), .ZN(n19495) );
  OAI211_X1 U22501 ( .C1(n19882), .C2(n19536), .A(n19496), .B(n19495), .ZN(
        P2_U3060) );
  AOI22_X1 U22502 ( .A1(n19502), .A2(n19922), .B1(n19921), .B2(n19501), .ZN(
        n19498) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19923), .ZN(n19497) );
  OAI211_X1 U22504 ( .C1(n19927), .C2(n19536), .A(n19498), .B(n19497), .ZN(
        P2_U3061) );
  AOI22_X1 U22505 ( .A1(n19502), .A2(n19929), .B1(n19928), .B2(n19501), .ZN(
        n19500) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19930), .ZN(n19499) );
  OAI211_X1 U22507 ( .C1(n19890), .C2(n19536), .A(n19500), .B(n19499), .ZN(
        P2_U3062) );
  AOI22_X1 U22508 ( .A1(n19940), .A2(n19502), .B1(n19937), .B2(n19501), .ZN(
        n19506) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19893), .ZN(n19505) );
  OAI211_X1 U22510 ( .C1(n19898), .C2(n19536), .A(n19506), .B(n19505), .ZN(
        P2_U3063) );
  NOR2_X1 U22511 ( .A1(n19508), .A2(n19540), .ZN(n19531) );
  OAI21_X1 U22512 ( .B1(n13398), .B2(n19531), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19511) );
  NOR2_X1 U22513 ( .A1(n19509), .A2(n19540), .ZN(n19512) );
  INV_X1 U22514 ( .A(n19512), .ZN(n19510) );
  NAND2_X1 U22515 ( .A1(n19511), .A2(n19510), .ZN(n19532) );
  AOI22_X1 U22516 ( .A1(n19532), .A2(n13210), .B1(n19856), .B2(n19531), .ZN(
        n19518) );
  AOI21_X1 U22517 ( .B1(n13398), .B2(n20079), .A(n19531), .ZN(n19515) );
  AOI21_X1 U22518 ( .B1(n19573), .B2(n19536), .A(n19627), .ZN(n19513) );
  NOR2_X1 U22519 ( .A1(n19513), .A2(n19512), .ZN(n19514) );
  MUX2_X1 U22520 ( .A(n19515), .B(n19514), .S(n20057), .Z(n19516) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19857), .ZN(n19517) );
  OAI211_X1 U22522 ( .C1(n19871), .C2(n19536), .A(n19518), .B(n19517), .ZN(
        P2_U3064) );
  AOI22_X1 U22523 ( .A1(n19532), .A2(n13231), .B1(n19899), .B2(n19531), .ZN(
        n19520) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19798), .ZN(n19519) );
  OAI211_X1 U22525 ( .C1(n19801), .C2(n19536), .A(n19520), .B(n19519), .ZN(
        P2_U3065) );
  AOI22_X1 U22526 ( .A1(n19532), .A2(n19441), .B1(n19904), .B2(n19531), .ZN(
        n19522) );
  INV_X1 U22527 ( .A(n19841), .ZN(n19905) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19905), .ZN(n19521) );
  OAI211_X1 U22529 ( .C1(n19908), .C2(n19536), .A(n19522), .B(n19521), .ZN(
        P2_U3066) );
  AOI22_X1 U22530 ( .A1(n19532), .A2(n19447), .B1(n19909), .B2(n19531), .ZN(
        n19524) );
  INV_X1 U22531 ( .A(n19878), .ZN(n19911) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19911), .ZN(n19523) );
  OAI211_X1 U22533 ( .C1(n19806), .C2(n19536), .A(n19524), .B(n19523), .ZN(
        P2_U3067) );
  INV_X1 U22534 ( .A(n19879), .ZN(n19920) );
  AOI22_X1 U22535 ( .A1(n19532), .A2(n19916), .B1(n19915), .B2(n19531), .ZN(
        n19526) );
  INV_X1 U22536 ( .A(n19882), .ZN(n19917) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19917), .ZN(n19525) );
  OAI211_X1 U22538 ( .C1(n19920), .C2(n19536), .A(n19526), .B(n19525), .ZN(
        P2_U3068) );
  INV_X1 U22539 ( .A(n19923), .ZN(n19887) );
  AOI22_X1 U22540 ( .A1(n19532), .A2(n19922), .B1(n19921), .B2(n19531), .ZN(
        n19528) );
  INV_X1 U22541 ( .A(n19927), .ZN(n19883) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19883), .ZN(n19527) );
  OAI211_X1 U22543 ( .C1(n19887), .C2(n19536), .A(n19528), .B(n19527), .ZN(
        P2_U3069) );
  INV_X1 U22544 ( .A(n19930), .ZN(n19813) );
  AOI22_X1 U22545 ( .A1(n19532), .A2(n19929), .B1(n19928), .B2(n19531), .ZN(
        n19530) );
  INV_X1 U22546 ( .A(n19890), .ZN(n19932) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19932), .ZN(n19529) );
  OAI211_X1 U22548 ( .C1(n19813), .C2(n19536), .A(n19530), .B(n19529), .ZN(
        P2_U3070) );
  INV_X1 U22549 ( .A(n19893), .ZN(n19947) );
  AOI22_X1 U22550 ( .A1(n19940), .A2(n19532), .B1(n19937), .B2(n19531), .ZN(
        n19535) );
  INV_X1 U22551 ( .A(n19898), .ZN(n19941) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19533), .B1(
        n19562), .B2(n19941), .ZN(n19534) );
  OAI211_X1 U22553 ( .C1(n19947), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P2_U3071) );
  OAI21_X1 U22554 ( .B1(n19660), .B2(n19537), .A(n20057), .ZN(n19549) );
  NAND2_X1 U22555 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19538), .ZN(
        n19548) );
  INV_X1 U22556 ( .A(n19548), .ZN(n19539) );
  OR2_X1 U22557 ( .A1(n19549), .A2(n19539), .ZN(n19545) );
  NOR2_X1 U22558 ( .A1(n19756), .A2(n19540), .ZN(n19568) );
  INV_X1 U22559 ( .A(n19568), .ZN(n19541) );
  OAI211_X1 U22560 ( .C1(n19542), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19861), 
        .B(n19541), .ZN(n19543) );
  AND2_X1 U22561 ( .A1(n19543), .A2(n19863), .ZN(n19544) );
  AND2_X1 U22562 ( .A1(n19545), .A2(n19544), .ZN(n19553) );
  AOI22_X1 U22563 ( .A1(n19857), .A2(n19599), .B1(n19856), .B2(n19568), .ZN(
        n19551) );
  OAI21_X1 U22564 ( .B1(n19546), .B2(n19568), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19547) );
  OAI21_X1 U22565 ( .B1(n19549), .B2(n19548), .A(n19547), .ZN(n19569) );
  AOI22_X1 U22566 ( .A1(n13210), .A2(n19569), .B1(n19562), .B2(n19832), .ZN(
        n19550) );
  OAI211_X1 U22567 ( .C1(n19553), .C2(n19552), .A(n19551), .B(n19550), .ZN(
        P2_U3072) );
  AOI22_X1 U22568 ( .A1(n19798), .A2(n19599), .B1(n19899), .B2(n19568), .ZN(
        n19555) );
  INV_X1 U22569 ( .A(n19553), .ZN(n19570) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19570), .B1(
        n13231), .B2(n19569), .ZN(n19554) );
  OAI211_X1 U22571 ( .C1(n19801), .C2(n19573), .A(n19555), .B(n19554), .ZN(
        P2_U3073) );
  INV_X1 U22572 ( .A(n19599), .ZN(n19565) );
  AOI22_X1 U22573 ( .A1(n19838), .A2(n19562), .B1(n19568), .B2(n19904), .ZN(
        n19557) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19570), .B1(
        n19441), .B2(n19569), .ZN(n19556) );
  OAI211_X1 U22575 ( .C1(n19841), .C2(n19565), .A(n19557), .B(n19556), .ZN(
        P2_U3074) );
  AOI22_X1 U22576 ( .A1(n19911), .A2(n19599), .B1(n19568), .B2(n19909), .ZN(
        n19559) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19570), .B1(
        n19447), .B2(n19569), .ZN(n19558) );
  OAI211_X1 U22578 ( .C1(n19806), .C2(n19573), .A(n19559), .B(n19558), .ZN(
        P2_U3075) );
  AOI22_X1 U22579 ( .A1(n19917), .A2(n19599), .B1(n19568), .B2(n19915), .ZN(
        n19561) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19570), .B1(
        n19916), .B2(n19569), .ZN(n19560) );
  OAI211_X1 U22581 ( .C1(n19920), .C2(n19573), .A(n19561), .B(n19560), .ZN(
        P2_U3076) );
  AOI22_X1 U22582 ( .A1(n19923), .A2(n19562), .B1(n19568), .B2(n19921), .ZN(
        n19564) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19570), .B1(
        n19922), .B2(n19569), .ZN(n19563) );
  OAI211_X1 U22584 ( .C1(n19927), .C2(n19565), .A(n19564), .B(n19563), .ZN(
        P2_U3077) );
  AOI22_X1 U22585 ( .A1(n19932), .A2(n19599), .B1(n19568), .B2(n19928), .ZN(
        n19567) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19570), .B1(
        n19929), .B2(n19569), .ZN(n19566) );
  OAI211_X1 U22587 ( .C1(n19813), .C2(n19573), .A(n19567), .B(n19566), .ZN(
        P2_U3078) );
  AOI22_X1 U22588 ( .A1(n19941), .A2(n19599), .B1(n19568), .B2(n19937), .ZN(
        n19572) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19570), .B1(
        n19940), .B2(n19569), .ZN(n19571) );
  OAI211_X1 U22590 ( .C1(n19947), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P2_U3079) );
  NOR2_X1 U22591 ( .A1(n19575), .A2(n19574), .ZN(n19785) );
  NAND2_X1 U22592 ( .A1(n19785), .A2(n20062), .ZN(n19581) );
  NOR2_X1 U22593 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19577), .ZN(
        n19597) );
  OAI21_X1 U22594 ( .B1(n9809), .B2(n19597), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19578) );
  OAI21_X1 U22595 ( .B1(n19581), .B2(n19861), .A(n19578), .ZN(n19598) );
  AOI22_X1 U22596 ( .A1(n19598), .A2(n13210), .B1(n19856), .B2(n19597), .ZN(
        n19584) );
  OAI21_X1 U22597 ( .B1(n19599), .B2(n19618), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19580) );
  AOI211_X1 U22598 ( .C1(n9809), .C2(n20079), .A(n20057), .B(n19597), .ZN(
        n19579) );
  AOI211_X1 U22599 ( .C1(n19581), .C2(n19580), .A(n19826), .B(n19579), .ZN(
        n19582) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19832), .ZN(n19583) );
  OAI211_X1 U22601 ( .C1(n19835), .C2(n19611), .A(n19584), .B(n19583), .ZN(
        P2_U3080) );
  AOI22_X1 U22602 ( .A1(n19598), .A2(n13231), .B1(n19899), .B2(n19597), .ZN(
        n19586) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19900), .ZN(n19585) );
  OAI211_X1 U22604 ( .C1(n19903), .C2(n19611), .A(n19586), .B(n19585), .ZN(
        P2_U3081) );
  AOI22_X1 U22605 ( .A1(n19598), .A2(n19441), .B1(n19904), .B2(n19597), .ZN(
        n19588) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19838), .ZN(n19587) );
  OAI211_X1 U22607 ( .C1(n19841), .C2(n19611), .A(n19588), .B(n19587), .ZN(
        P2_U3082) );
  AOI22_X1 U22608 ( .A1(n19598), .A2(n19447), .B1(n19909), .B2(n19597), .ZN(
        n19590) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19910), .ZN(n19589) );
  OAI211_X1 U22610 ( .C1(n19878), .C2(n19611), .A(n19590), .B(n19589), .ZN(
        P2_U3083) );
  AOI22_X1 U22611 ( .A1(n19598), .A2(n19916), .B1(n19915), .B2(n19597), .ZN(
        n19592) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19879), .ZN(n19591) );
  OAI211_X1 U22613 ( .C1(n19882), .C2(n19611), .A(n19592), .B(n19591), .ZN(
        P2_U3084) );
  AOI22_X1 U22614 ( .A1(n19598), .A2(n19922), .B1(n19921), .B2(n19597), .ZN(
        n19594) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19923), .ZN(n19593) );
  OAI211_X1 U22616 ( .C1(n19927), .C2(n19611), .A(n19594), .B(n19593), .ZN(
        P2_U3085) );
  AOI22_X1 U22617 ( .A1(n19598), .A2(n19929), .B1(n19928), .B2(n19597), .ZN(
        n19596) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19930), .ZN(n19595) );
  OAI211_X1 U22619 ( .C1(n19890), .C2(n19611), .A(n19596), .B(n19595), .ZN(
        P2_U3086) );
  AOI22_X1 U22620 ( .A1(n19940), .A2(n19598), .B1(n19937), .B2(n19597), .ZN(
        n19602) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19893), .ZN(n19601) );
  OAI211_X1 U22622 ( .C1(n19898), .C2(n19611), .A(n19602), .B(n19601), .ZN(
        P2_U3087) );
  AOI22_X1 U22623 ( .A1(n19900), .A2(n19618), .B1(n19899), .B2(n19629), .ZN(
        n19604) );
  AOI22_X1 U22624 ( .A1(n13231), .A2(n19619), .B1(n19649), .B2(n19798), .ZN(
        n19603) );
  OAI211_X1 U22625 ( .C1(n19608), .C2(n13388), .A(n19604), .B(n19603), .ZN(
        P2_U3089) );
  INV_X1 U22626 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19607) );
  AOI22_X1 U22627 ( .A1(n19838), .A2(n19618), .B1(n19629), .B2(n19904), .ZN(
        n19606) );
  AOI22_X1 U22628 ( .A1(n19441), .A2(n19619), .B1(n19649), .B2(n19905), .ZN(
        n19605) );
  OAI211_X1 U22629 ( .C1(n19608), .C2(n19607), .A(n19606), .B(n19605), .ZN(
        P2_U3090) );
  AOI22_X1 U22630 ( .A1(n19911), .A2(n19649), .B1(n19629), .B2(n19909), .ZN(
        n19610) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19620), .B1(
        n19447), .B2(n19619), .ZN(n19609) );
  OAI211_X1 U22632 ( .C1(n19806), .C2(n19611), .A(n19610), .B(n19609), .ZN(
        P2_U3091) );
  AOI22_X1 U22633 ( .A1(n19879), .A2(n19618), .B1(n19629), .B2(n19915), .ZN(
        n19613) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19620), .B1(
        n19916), .B2(n19619), .ZN(n19612) );
  OAI211_X1 U22635 ( .C1(n19882), .C2(n19646), .A(n19613), .B(n19612), .ZN(
        P2_U3092) );
  AOI22_X1 U22636 ( .A1(n19923), .A2(n19618), .B1(n19629), .B2(n19921), .ZN(
        n19615) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19620), .B1(
        n19922), .B2(n19619), .ZN(n19614) );
  OAI211_X1 U22638 ( .C1(n19927), .C2(n19646), .A(n19615), .B(n19614), .ZN(
        P2_U3093) );
  AOI22_X1 U22639 ( .A1(n19930), .A2(n19618), .B1(n19629), .B2(n19928), .ZN(
        n19617) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19620), .B1(
        n19929), .B2(n19619), .ZN(n19616) );
  OAI211_X1 U22641 ( .C1(n19890), .C2(n19646), .A(n19617), .B(n19616), .ZN(
        P2_U3094) );
  AOI22_X1 U22642 ( .A1(n19893), .A2(n19618), .B1(n19629), .B2(n19937), .ZN(
        n19622) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19620), .B1(
        n19940), .B2(n19619), .ZN(n19621) );
  OAI211_X1 U22644 ( .C1(n19898), .C2(n19646), .A(n19622), .B(n19621), .ZN(
        P2_U3095) );
  NAND2_X1 U22645 ( .A1(n19623), .A2(n19655), .ZN(n19653) );
  NOR2_X1 U22646 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19855), .ZN(
        n19664) );
  INV_X1 U22647 ( .A(n19664), .ZN(n19658) );
  NOR2_X1 U22648 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19658), .ZN(
        n19647) );
  NOR2_X1 U22649 ( .A1(n19629), .A2(n19647), .ZN(n19626) );
  INV_X1 U22650 ( .A(n19948), .ZN(n19657) );
  INV_X1 U22651 ( .A(n19624), .ZN(n19625) );
  INV_X1 U22652 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19822) );
  NOR3_X1 U22653 ( .A1(n19625), .A2(n19647), .A3(n19822), .ZN(n19630) );
  AOI211_X2 U22654 ( .C1(n19626), .C2(n19822), .A(n19657), .B(n19630), .ZN(
        n19648) );
  AOI22_X1 U22655 ( .A1(n19648), .A2(n13210), .B1(n19856), .B2(n19647), .ZN(
        n19633) );
  AOI21_X1 U22656 ( .B1(n19646), .B2(n19653), .A(n19627), .ZN(n19628) );
  AOI221_X1 U22657 ( .B1(n20079), .B2(n19629), .C1(n20079), .C2(n19628), .A(
        n19647), .ZN(n19631) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19650), .B1(
        n19649), .B2(n19832), .ZN(n19632) );
  OAI211_X1 U22659 ( .C1(n19835), .C2(n19653), .A(n19633), .B(n19632), .ZN(
        P2_U3096) );
  AOI22_X1 U22660 ( .A1(n19648), .A2(n13231), .B1(n19899), .B2(n19647), .ZN(
        n19635) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19650), .B1(
        n19680), .B2(n19798), .ZN(n19634) );
  OAI211_X1 U22662 ( .C1(n19801), .C2(n19646), .A(n19635), .B(n19634), .ZN(
        P2_U3097) );
  AOI22_X1 U22663 ( .A1(n19648), .A2(n19441), .B1(n19904), .B2(n19647), .ZN(
        n19637) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19650), .B1(
        n19649), .B2(n19838), .ZN(n19636) );
  OAI211_X1 U22665 ( .C1(n19841), .C2(n19653), .A(n19637), .B(n19636), .ZN(
        P2_U3098) );
  AOI22_X1 U22666 ( .A1(n19648), .A2(n19447), .B1(n19909), .B2(n19647), .ZN(
        n19639) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19650), .B1(
        n19680), .B2(n19911), .ZN(n19638) );
  OAI211_X1 U22668 ( .C1(n19806), .C2(n19646), .A(n19639), .B(n19638), .ZN(
        P2_U3099) );
  AOI22_X1 U22669 ( .A1(n19648), .A2(n19916), .B1(n19915), .B2(n19647), .ZN(
        n19641) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19650), .B1(
        n19680), .B2(n19917), .ZN(n19640) );
  OAI211_X1 U22671 ( .C1(n19920), .C2(n19646), .A(n19641), .B(n19640), .ZN(
        P2_U3100) );
  AOI22_X1 U22672 ( .A1(n19648), .A2(n19922), .B1(n19921), .B2(n19647), .ZN(
        n19643) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19650), .B1(
        n19649), .B2(n19923), .ZN(n19642) );
  OAI211_X1 U22674 ( .C1(n19927), .C2(n19653), .A(n19643), .B(n19642), .ZN(
        P2_U3101) );
  AOI22_X1 U22675 ( .A1(n19648), .A2(n19929), .B1(n19928), .B2(n19647), .ZN(
        n19645) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19650), .B1(
        n19680), .B2(n19932), .ZN(n19644) );
  OAI211_X1 U22677 ( .C1(n19813), .C2(n19646), .A(n19645), .B(n19644), .ZN(
        P2_U3102) );
  AOI22_X1 U22678 ( .A1(n19648), .A2(n19940), .B1(n19937), .B2(n19647), .ZN(
        n19652) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19650), .B1(
        n19649), .B2(n19893), .ZN(n19651) );
  OAI211_X1 U22680 ( .C1(n19898), .C2(n19653), .A(n19652), .B(n19651), .ZN(
        P2_U3103) );
  INV_X1 U22681 ( .A(n13639), .ZN(n19656) );
  NAND2_X1 U22682 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19664), .ZN(
        n19662) );
  INV_X1 U22683 ( .A(n19662), .ZN(n19687) );
  NOR3_X1 U22684 ( .A1(n19656), .A2(n19687), .A3(n19822), .ZN(n19661) );
  AOI211_X2 U22685 ( .C1(n19658), .C2(n19822), .A(n19657), .B(n19661), .ZN(
        n19679) );
  AOI22_X1 U22686 ( .A1(n19679), .A2(n13210), .B1(n19856), .B2(n19687), .ZN(
        n19666) );
  NOR2_X1 U22687 ( .A1(n19660), .A2(n19659), .ZN(n20056) );
  AOI211_X1 U22688 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19662), .A(n19826), 
        .B(n19661), .ZN(n19663) );
  OAI21_X1 U22689 ( .B1(n19664), .B2(n20056), .A(n19663), .ZN(n19681) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19832), .ZN(n19665) );
  OAI211_X1 U22691 ( .C1(n19835), .C2(n19715), .A(n19666), .B(n19665), .ZN(
        P2_U3104) );
  AOI22_X1 U22692 ( .A1(n19679), .A2(n13231), .B1(n19899), .B2(n19687), .ZN(
        n19668) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19900), .ZN(n19667) );
  OAI211_X1 U22694 ( .C1(n19903), .C2(n19715), .A(n19668), .B(n19667), .ZN(
        P2_U3105) );
  AOI22_X1 U22695 ( .A1(n19679), .A2(n19441), .B1(n19904), .B2(n19687), .ZN(
        n19670) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19838), .ZN(n19669) );
  OAI211_X1 U22697 ( .C1(n19841), .C2(n19715), .A(n19670), .B(n19669), .ZN(
        P2_U3106) );
  AOI22_X1 U22698 ( .A1(n19679), .A2(n19447), .B1(n19909), .B2(n19687), .ZN(
        n19672) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19910), .ZN(n19671) );
  OAI211_X1 U22700 ( .C1(n19878), .C2(n19715), .A(n19672), .B(n19671), .ZN(
        P2_U3107) );
  AOI22_X1 U22701 ( .A1(n19679), .A2(n19916), .B1(n19915), .B2(n19687), .ZN(
        n19674) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19879), .ZN(n19673) );
  OAI211_X1 U22703 ( .C1(n19882), .C2(n19715), .A(n19674), .B(n19673), .ZN(
        P2_U3108) );
  AOI22_X1 U22704 ( .A1(n19679), .A2(n19922), .B1(n19921), .B2(n19687), .ZN(
        n19676) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19923), .ZN(n19675) );
  OAI211_X1 U22706 ( .C1(n19927), .C2(n19715), .A(n19676), .B(n19675), .ZN(
        P2_U3109) );
  AOI22_X1 U22707 ( .A1(n19679), .A2(n19929), .B1(n19928), .B2(n19687), .ZN(
        n19678) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19930), .ZN(n19677) );
  OAI211_X1 U22709 ( .C1(n19890), .C2(n19715), .A(n19678), .B(n19677), .ZN(
        P2_U3110) );
  AOI22_X1 U22710 ( .A1(n19679), .A2(n19940), .B1(n19937), .B2(n19687), .ZN(
        n19683) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19681), .B1(
        n19680), .B2(n19893), .ZN(n19682) );
  OAI211_X1 U22712 ( .C1(n19898), .C2(n19715), .A(n19683), .B(n19682), .ZN(
        P2_U3111) );
  NOR2_X1 U22713 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19684), .ZN(
        n19710) );
  AOI22_X1 U22714 ( .A1(n19857), .A2(n19728), .B1(n19856), .B2(n19710), .ZN(
        n19697) );
  INV_X1 U22715 ( .A(n19715), .ZN(n19685) );
  OAI21_X1 U22716 ( .B1(n19728), .B2(n19685), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19686) );
  NAND2_X1 U22717 ( .A1(n19686), .A2(n20057), .ZN(n19695) );
  NOR2_X1 U22718 ( .A1(n19710), .A2(n19687), .ZN(n19693) );
  INV_X1 U22719 ( .A(n19693), .ZN(n19690) );
  INV_X1 U22720 ( .A(n19710), .ZN(n19688) );
  OAI211_X1 U22721 ( .C1(n19691), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19861), 
        .B(n19688), .ZN(n19689) );
  OAI211_X1 U22722 ( .C1(n19695), .C2(n19690), .A(n19863), .B(n19689), .ZN(
        n19712) );
  INV_X1 U22723 ( .A(n19691), .ZN(n19692) );
  OAI21_X1 U22724 ( .B1(n19692), .B2(n19710), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19694) );
  AOI22_X1 U22725 ( .A1(n19695), .A2(n19694), .B1(n19693), .B2(n19822), .ZN(
        n19711) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19712), .B1(
        n13210), .B2(n19711), .ZN(n19696) );
  OAI211_X1 U22727 ( .C1(n19871), .C2(n19715), .A(n19697), .B(n19696), .ZN(
        P2_U3112) );
  AOI22_X1 U22728 ( .A1(n19798), .A2(n19728), .B1(n19899), .B2(n19710), .ZN(
        n19699) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19712), .B1(
        n13231), .B2(n19711), .ZN(n19698) );
  OAI211_X1 U22730 ( .C1(n19801), .C2(n19715), .A(n19699), .B(n19698), .ZN(
        P2_U3113) );
  AOI22_X1 U22731 ( .A1(n19905), .A2(n19728), .B1(n19904), .B2(n19710), .ZN(
        n19701) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19712), .B1(
        n19441), .B2(n19711), .ZN(n19700) );
  OAI211_X1 U22733 ( .C1(n19908), .C2(n19715), .A(n19701), .B(n19700), .ZN(
        P2_U3114) );
  AOI22_X1 U22734 ( .A1(n19911), .A2(n19728), .B1(n19909), .B2(n19710), .ZN(
        n19703) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19712), .B1(
        n19447), .B2(n19711), .ZN(n19702) );
  OAI211_X1 U22736 ( .C1(n19806), .C2(n19715), .A(n19703), .B(n19702), .ZN(
        P2_U3115) );
  AOI22_X1 U22737 ( .A1(n19917), .A2(n19728), .B1(n19915), .B2(n19710), .ZN(
        n19705) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19712), .B1(
        n19916), .B2(n19711), .ZN(n19704) );
  OAI211_X1 U22739 ( .C1(n19920), .C2(n19715), .A(n19705), .B(n19704), .ZN(
        P2_U3116) );
  AOI22_X1 U22740 ( .A1(n19883), .A2(n19728), .B1(n19921), .B2(n19710), .ZN(
        n19707) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19712), .B1(
        n19922), .B2(n19711), .ZN(n19706) );
  OAI211_X1 U22742 ( .C1(n19887), .C2(n19715), .A(n19707), .B(n19706), .ZN(
        P2_U3117) );
  AOI22_X1 U22743 ( .A1(n19932), .A2(n19728), .B1(n19928), .B2(n19710), .ZN(
        n19709) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19712), .B1(
        n19929), .B2(n19711), .ZN(n19708) );
  OAI211_X1 U22745 ( .C1(n19813), .C2(n19715), .A(n19709), .B(n19708), .ZN(
        P2_U3118) );
  AOI22_X1 U22746 ( .A1(n19941), .A2(n19728), .B1(n19937), .B2(n19710), .ZN(
        n19714) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19712), .B1(
        n19940), .B2(n19711), .ZN(n19713) );
  OAI211_X1 U22748 ( .C1(n19947), .C2(n19715), .A(n19714), .B(n19713), .ZN(
        P2_U3119) );
  AOI22_X1 U22749 ( .A1(n19905), .A2(n19751), .B1(n19727), .B2(n19904), .ZN(
        n19717) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19730), .B1(
        n19441), .B2(n19729), .ZN(n19716) );
  OAI211_X1 U22751 ( .C1(n19908), .C2(n19724), .A(n19717), .B(n19716), .ZN(
        P2_U3122) );
  INV_X1 U22752 ( .A(n19751), .ZN(n19733) );
  AOI22_X1 U22753 ( .A1(n19910), .A2(n19728), .B1(n19727), .B2(n19909), .ZN(
        n19719) );
  AOI22_X1 U22754 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19730), .B1(
        n19447), .B2(n19729), .ZN(n19718) );
  OAI211_X1 U22755 ( .C1(n19878), .C2(n19733), .A(n19719), .B(n19718), .ZN(
        P2_U3123) );
  AOI22_X1 U22756 ( .A1(n19917), .A2(n19751), .B1(n19727), .B2(n19915), .ZN(
        n19721) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19730), .B1(
        n19916), .B2(n19729), .ZN(n19720) );
  OAI211_X1 U22758 ( .C1(n19920), .C2(n19724), .A(n19721), .B(n19720), .ZN(
        P2_U3124) );
  AOI22_X1 U22759 ( .A1(n19883), .A2(n19751), .B1(n19727), .B2(n19921), .ZN(
        n19723) );
  AOI22_X1 U22760 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19730), .B1(
        n19922), .B2(n19729), .ZN(n19722) );
  OAI211_X1 U22761 ( .C1(n19887), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3125) );
  AOI22_X1 U22762 ( .A1(n19930), .A2(n19728), .B1(n19727), .B2(n19928), .ZN(
        n19726) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19730), .B1(
        n19929), .B2(n19729), .ZN(n19725) );
  OAI211_X1 U22764 ( .C1(n19890), .C2(n19733), .A(n19726), .B(n19725), .ZN(
        P2_U3126) );
  AOI22_X1 U22765 ( .A1(n19893), .A2(n19728), .B1(n19727), .B2(n19937), .ZN(
        n19732) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19730), .B1(
        n19940), .B2(n19729), .ZN(n19731) );
  OAI211_X1 U22767 ( .C1(n19898), .C2(n19733), .A(n19732), .B(n19731), .ZN(
        P2_U3127) );
  INV_X1 U22768 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U22769 ( .A1(n19750), .A2(n13210), .B1(n19749), .B2(n19856), .ZN(
        n19735) );
  AOI22_X1 U22770 ( .A1(n19751), .A2(n19832), .B1(n19781), .B2(n19857), .ZN(
        n19734) );
  OAI211_X1 U22771 ( .C1(n19755), .C2(n19736), .A(n19735), .B(n19734), .ZN(
        P2_U3128) );
  INV_X1 U22772 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U22773 ( .A1(n19750), .A2(n19441), .B1(n19749), .B2(n19904), .ZN(
        n19738) );
  AOI22_X1 U22774 ( .A1(n19751), .A2(n19838), .B1(n19781), .B2(n19905), .ZN(
        n19737) );
  OAI211_X1 U22775 ( .C1(n19755), .C2(n19739), .A(n19738), .B(n19737), .ZN(
        P2_U3130) );
  AOI22_X1 U22776 ( .A1(n19750), .A2(n19447), .B1(n19749), .B2(n19909), .ZN(
        n19741) );
  AOI22_X1 U22777 ( .A1(n19751), .A2(n19910), .B1(n19781), .B2(n19911), .ZN(
        n19740) );
  OAI211_X1 U22778 ( .C1(n19755), .C2(n13427), .A(n19741), .B(n19740), .ZN(
        P2_U3131) );
  INV_X1 U22779 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U22780 ( .A1(n19750), .A2(n19916), .B1(n19749), .B2(n19915), .ZN(
        n19743) );
  AOI22_X1 U22781 ( .A1(n19751), .A2(n19879), .B1(n19781), .B2(n19917), .ZN(
        n19742) );
  OAI211_X1 U22782 ( .C1(n19755), .C2(n19744), .A(n19743), .B(n19742), .ZN(
        P2_U3132) );
  AOI22_X1 U22783 ( .A1(n19750), .A2(n19922), .B1(n19749), .B2(n19921), .ZN(
        n19746) );
  AOI22_X1 U22784 ( .A1(n19751), .A2(n19923), .B1(n19781), .B2(n19883), .ZN(
        n19745) );
  OAI211_X1 U22785 ( .C1(n19755), .C2(n13659), .A(n19746), .B(n19745), .ZN(
        P2_U3133) );
  AOI22_X1 U22786 ( .A1(n19750), .A2(n19929), .B1(n19749), .B2(n19928), .ZN(
        n19748) );
  AOI22_X1 U22787 ( .A1(n19751), .A2(n19930), .B1(n19781), .B2(n19932), .ZN(
        n19747) );
  OAI211_X1 U22788 ( .C1(n19755), .C2(n14894), .A(n19748), .B(n19747), .ZN(
        P2_U3134) );
  INV_X1 U22789 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U22790 ( .A1(n19940), .A2(n19750), .B1(n19749), .B2(n19937), .ZN(
        n19753) );
  AOI22_X1 U22791 ( .A1(n19751), .A2(n19893), .B1(n19781), .B2(n19941), .ZN(
        n19752) );
  OAI211_X1 U22792 ( .C1(n19755), .C2(n19754), .A(n19753), .B(n19752), .ZN(
        P2_U3135) );
  NOR2_X1 U22793 ( .A1(n19756), .A2(n19758), .ZN(n19779) );
  NOR2_X1 U22794 ( .A1(n20078), .A2(n19758), .ZN(n19764) );
  INV_X1 U22795 ( .A(n19764), .ZN(n19759) );
  OAI21_X1 U22796 ( .B1(n19759), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19822), 
        .ZN(n19760) );
  AND2_X1 U22797 ( .A1(n19761), .A2(n19760), .ZN(n19780) );
  AOI22_X1 U22798 ( .A1(n19780), .A2(n13210), .B1(n19856), .B2(n19779), .ZN(
        n19766) );
  OAI211_X1 U22799 ( .C1(n19779), .C2(n20079), .A(n19761), .B(n19863), .ZN(
        n19762) );
  INV_X1 U22800 ( .A(n19762), .ZN(n19763) );
  OAI221_X1 U22801 ( .B1(n19764), .B2(n20053), .C1(n19764), .C2(n19829), .A(
        n19763), .ZN(n19782) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19832), .ZN(n19765) );
  OAI211_X1 U22803 ( .C1(n19835), .C2(n19819), .A(n19766), .B(n19765), .ZN(
        P2_U3136) );
  AOI22_X1 U22804 ( .A1(n19780), .A2(n13231), .B1(n19899), .B2(n19779), .ZN(
        n19768) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19900), .ZN(n19767) );
  OAI211_X1 U22806 ( .C1(n19903), .C2(n19819), .A(n19768), .B(n19767), .ZN(
        P2_U3137) );
  AOI22_X1 U22807 ( .A1(n19780), .A2(n19441), .B1(n19904), .B2(n19779), .ZN(
        n19770) );
  AOI22_X1 U22808 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19838), .ZN(n19769) );
  OAI211_X1 U22809 ( .C1(n19841), .C2(n19819), .A(n19770), .B(n19769), .ZN(
        P2_U3138) );
  AOI22_X1 U22810 ( .A1(n19780), .A2(n19447), .B1(n19909), .B2(n19779), .ZN(
        n19772) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19910), .ZN(n19771) );
  OAI211_X1 U22812 ( .C1(n19878), .C2(n19819), .A(n19772), .B(n19771), .ZN(
        P2_U3139) );
  AOI22_X1 U22813 ( .A1(n19780), .A2(n19916), .B1(n19915), .B2(n19779), .ZN(
        n19774) );
  AOI22_X1 U22814 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19879), .ZN(n19773) );
  OAI211_X1 U22815 ( .C1(n19882), .C2(n19819), .A(n19774), .B(n19773), .ZN(
        P2_U3140) );
  AOI22_X1 U22816 ( .A1(n19780), .A2(n19922), .B1(n19921), .B2(n19779), .ZN(
        n19776) );
  AOI22_X1 U22817 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19923), .ZN(n19775) );
  OAI211_X1 U22818 ( .C1(n19927), .C2(n19819), .A(n19776), .B(n19775), .ZN(
        P2_U3141) );
  AOI22_X1 U22819 ( .A1(n19780), .A2(n19929), .B1(n19928), .B2(n19779), .ZN(
        n19778) );
  AOI22_X1 U22820 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19930), .ZN(n19777) );
  OAI211_X1 U22821 ( .C1(n19890), .C2(n19819), .A(n19778), .B(n19777), .ZN(
        P2_U3142) );
  AOI22_X1 U22822 ( .A1(n19940), .A2(n19780), .B1(n19937), .B2(n19779), .ZN(
        n19784) );
  AOI22_X1 U22823 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19893), .ZN(n19783) );
  OAI211_X1 U22824 ( .C1(n19898), .C2(n19819), .A(n19784), .B(n19783), .ZN(
        P2_U3143) );
  NAND2_X1 U22825 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19785), .ZN(
        n19793) );
  OR2_X1 U22826 ( .A1(n19793), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19788) );
  INV_X1 U22827 ( .A(n19786), .ZN(n19787) );
  NOR3_X1 U22828 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20069), .A3(
        n20062), .ZN(n19831) );
  INV_X1 U22829 ( .A(n19831), .ZN(n19821) );
  NOR2_X1 U22830 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19821), .ZN(
        n19814) );
  NOR3_X1 U22831 ( .A1(n19787), .A2(n19814), .A3(n19822), .ZN(n19792) );
  AOI21_X1 U22832 ( .B1(n19822), .B2(n19788), .A(n19792), .ZN(n19815) );
  AOI22_X1 U22833 ( .A1(n19815), .A2(n13210), .B1(n19856), .B2(n19814), .ZN(
        n19797) );
  NOR2_X2 U22834 ( .A1(n19790), .A2(n19789), .ZN(n19851) );
  INV_X1 U22835 ( .A(n19819), .ZN(n19791) );
  OAI21_X1 U22836 ( .B1(n19851), .B2(n19791), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19794) );
  AOI211_X1 U22837 ( .C1(n19794), .C2(n19793), .A(n19826), .B(n19792), .ZN(
        n19795) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19857), .ZN(n19796) );
  OAI211_X1 U22839 ( .C1(n19871), .C2(n19819), .A(n19797), .B(n19796), .ZN(
        P2_U3144) );
  AOI22_X1 U22840 ( .A1(n19815), .A2(n13231), .B1(n19899), .B2(n19814), .ZN(
        n19800) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19798), .ZN(n19799) );
  OAI211_X1 U22842 ( .C1(n19801), .C2(n19819), .A(n19800), .B(n19799), .ZN(
        P2_U3145) );
  AOI22_X1 U22843 ( .A1(n19815), .A2(n19441), .B1(n19904), .B2(n19814), .ZN(
        n19803) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19905), .ZN(n19802) );
  OAI211_X1 U22845 ( .C1(n19908), .C2(n19819), .A(n19803), .B(n19802), .ZN(
        P2_U3146) );
  AOI22_X1 U22846 ( .A1(n19815), .A2(n19447), .B1(n19909), .B2(n19814), .ZN(
        n19805) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19911), .ZN(n19804) );
  OAI211_X1 U22848 ( .C1(n19806), .C2(n19819), .A(n19805), .B(n19804), .ZN(
        P2_U3147) );
  AOI22_X1 U22849 ( .A1(n19815), .A2(n19916), .B1(n19915), .B2(n19814), .ZN(
        n19808) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19917), .ZN(n19807) );
  OAI211_X1 U22851 ( .C1(n19920), .C2(n19819), .A(n19808), .B(n19807), .ZN(
        P2_U3148) );
  AOI22_X1 U22852 ( .A1(n19815), .A2(n19922), .B1(n19921), .B2(n19814), .ZN(
        n19810) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19883), .ZN(n19809) );
  OAI211_X1 U22854 ( .C1(n19887), .C2(n19819), .A(n19810), .B(n19809), .ZN(
        P2_U3149) );
  AOI22_X1 U22855 ( .A1(n19815), .A2(n19929), .B1(n19928), .B2(n19814), .ZN(
        n19812) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19932), .ZN(n19811) );
  OAI211_X1 U22857 ( .C1(n19813), .C2(n19819), .A(n19812), .B(n19811), .ZN(
        P2_U3150) );
  AOI22_X1 U22858 ( .A1(n19815), .A2(n19940), .B1(n19937), .B2(n19814), .ZN(
        n19818) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19816), .B1(
        n19851), .B2(n19941), .ZN(n19817) );
  OAI211_X1 U22860 ( .C1(n19947), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        P2_U3151) );
  OR2_X1 U22861 ( .A1(n19821), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19824) );
  NAND2_X1 U22862 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n19827) );
  INV_X1 U22863 ( .A(n19827), .ZN(n19859) );
  NOR3_X1 U22864 ( .A1(n19823), .A2(n19859), .A3(n19822), .ZN(n19825) );
  AOI21_X1 U22865 ( .B1(n19822), .B2(n19824), .A(n19825), .ZN(n19850) );
  AOI22_X1 U22866 ( .A1(n19850), .A2(n13210), .B1(n19856), .B2(n19859), .ZN(
        n19834) );
  AOI211_X1 U22867 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19827), .A(n19826), 
        .B(n19825), .ZN(n19828) );
  OAI221_X1 U22868 ( .B1(n19831), .B2(n19830), .C1(n19831), .C2(n19829), .A(
        n19828), .ZN(n19852) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19832), .ZN(n19833) );
  OAI211_X1 U22870 ( .C1(n19835), .C2(n19886), .A(n19834), .B(n19833), .ZN(
        P2_U3152) );
  AOI22_X1 U22871 ( .A1(n19850), .A2(n13231), .B1(n19899), .B2(n19859), .ZN(
        n19837) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19900), .ZN(n19836) );
  OAI211_X1 U22873 ( .C1(n19903), .C2(n19886), .A(n19837), .B(n19836), .ZN(
        P2_U3153) );
  AOI22_X1 U22874 ( .A1(n19850), .A2(n19441), .B1(n19904), .B2(n19859), .ZN(
        n19840) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19838), .ZN(n19839) );
  OAI211_X1 U22876 ( .C1(n19841), .C2(n19886), .A(n19840), .B(n19839), .ZN(
        P2_U3154) );
  AOI22_X1 U22877 ( .A1(n19850), .A2(n19447), .B1(n19909), .B2(n19859), .ZN(
        n19843) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19910), .ZN(n19842) );
  OAI211_X1 U22879 ( .C1(n19878), .C2(n19886), .A(n19843), .B(n19842), .ZN(
        P2_U3155) );
  AOI22_X1 U22880 ( .A1(n19850), .A2(n19916), .B1(n19915), .B2(n19859), .ZN(
        n19845) );
  AOI22_X1 U22881 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19879), .ZN(n19844) );
  OAI211_X1 U22882 ( .C1(n19882), .C2(n19886), .A(n19845), .B(n19844), .ZN(
        P2_U3156) );
  AOI22_X1 U22883 ( .A1(n19850), .A2(n19922), .B1(n19921), .B2(n19859), .ZN(
        n19847) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19923), .ZN(n19846) );
  OAI211_X1 U22885 ( .C1(n19927), .C2(n19886), .A(n19847), .B(n19846), .ZN(
        P2_U3157) );
  AOI22_X1 U22886 ( .A1(n19850), .A2(n19929), .B1(n19928), .B2(n19859), .ZN(
        n19849) );
  AOI22_X1 U22887 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19930), .ZN(n19848) );
  OAI211_X1 U22888 ( .C1(n19890), .C2(n19886), .A(n19849), .B(n19848), .ZN(
        P2_U3158) );
  AOI22_X1 U22889 ( .A1(n19850), .A2(n19940), .B1(n19937), .B2(n19859), .ZN(
        n19854) );
  AOI22_X1 U22890 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19852), .B1(
        n19851), .B2(n19893), .ZN(n19853) );
  OAI211_X1 U22891 ( .C1(n19898), .C2(n19886), .A(n19854), .B(n19853), .ZN(
        P2_U3159) );
  NOR3_X2 U22892 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20062), .A3(
        n19855), .ZN(n19891) );
  AOI22_X1 U22893 ( .A1(n19857), .A2(n19931), .B1(n19856), .B2(n19891), .ZN(
        n19870) );
  OAI21_X1 U22894 ( .B1(n19892), .B2(n19931), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19858) );
  NAND2_X1 U22895 ( .A1(n19858), .A2(n20057), .ZN(n19868) );
  NOR2_X1 U22896 ( .A1(n19891), .A2(n19859), .ZN(n19867) );
  INV_X1 U22897 ( .A(n19867), .ZN(n19864) );
  INV_X1 U22898 ( .A(n19891), .ZN(n19860) );
  OAI211_X1 U22899 ( .C1(n13654), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19861), 
        .B(n19860), .ZN(n19862) );
  OAI211_X1 U22900 ( .C1(n19868), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        n19895) );
  INV_X1 U22901 ( .A(n13654), .ZN(n19865) );
  OAI21_X1 U22902 ( .B1(n19865), .B2(n19891), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19866) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19895), .B1(
        n13210), .B2(n19894), .ZN(n19869) );
  OAI211_X1 U22904 ( .C1(n19871), .C2(n19886), .A(n19870), .B(n19869), .ZN(
        P2_U3160) );
  AOI22_X1 U22905 ( .A1(n19900), .A2(n19892), .B1(n19899), .B2(n19891), .ZN(
        n19873) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19895), .B1(
        n13231), .B2(n19894), .ZN(n19872) );
  OAI211_X1 U22907 ( .C1(n19903), .C2(n19946), .A(n19873), .B(n19872), .ZN(
        P2_U3161) );
  AOI22_X1 U22908 ( .A1(n19905), .A2(n19931), .B1(n19904), .B2(n19891), .ZN(
        n19875) );
  AOI22_X1 U22909 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19895), .B1(
        n19441), .B2(n19894), .ZN(n19874) );
  OAI211_X1 U22910 ( .C1(n19908), .C2(n19886), .A(n19875), .B(n19874), .ZN(
        P2_U3162) );
  AOI22_X1 U22911 ( .A1(n19910), .A2(n19892), .B1(n19909), .B2(n19891), .ZN(
        n19877) );
  AOI22_X1 U22912 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19895), .B1(
        n19447), .B2(n19894), .ZN(n19876) );
  OAI211_X1 U22913 ( .C1(n19878), .C2(n19946), .A(n19877), .B(n19876), .ZN(
        P2_U3163) );
  AOI22_X1 U22914 ( .A1(n19879), .A2(n19892), .B1(n19915), .B2(n19891), .ZN(
        n19881) );
  AOI22_X1 U22915 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19895), .B1(
        n19916), .B2(n19894), .ZN(n19880) );
  OAI211_X1 U22916 ( .C1(n19882), .C2(n19946), .A(n19881), .B(n19880), .ZN(
        P2_U3164) );
  AOI22_X1 U22917 ( .A1(n19883), .A2(n19931), .B1(n19921), .B2(n19891), .ZN(
        n19885) );
  AOI22_X1 U22918 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19895), .B1(
        n19922), .B2(n19894), .ZN(n19884) );
  OAI211_X1 U22919 ( .C1(n19887), .C2(n19886), .A(n19885), .B(n19884), .ZN(
        P2_U3165) );
  AOI22_X1 U22920 ( .A1(n19930), .A2(n19892), .B1(n19928), .B2(n19891), .ZN(
        n19889) );
  AOI22_X1 U22921 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19895), .B1(
        n19929), .B2(n19894), .ZN(n19888) );
  OAI211_X1 U22922 ( .C1(n19890), .C2(n19946), .A(n19889), .B(n19888), .ZN(
        P2_U3166) );
  AOI22_X1 U22923 ( .A1(n19893), .A2(n19892), .B1(n19937), .B2(n19891), .ZN(
        n19897) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19895), .B1(
        n19940), .B2(n19894), .ZN(n19896) );
  OAI211_X1 U22925 ( .C1(n19898), .C2(n19946), .A(n19897), .B(n19896), .ZN(
        P2_U3167) );
  AOI22_X1 U22926 ( .A1(n19939), .A2(n13231), .B1(n19938), .B2(n19899), .ZN(
        n19902) );
  INV_X1 U22927 ( .A(n19936), .ZN(n19943) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19943), .B1(
        n19931), .B2(n19900), .ZN(n19901) );
  OAI211_X1 U22929 ( .C1(n19903), .C2(n19926), .A(n19902), .B(n19901), .ZN(
        P2_U3169) );
  AOI22_X1 U22930 ( .A1(n19939), .A2(n19441), .B1(n19938), .B2(n19904), .ZN(
        n19907) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19905), .ZN(n19906) );
  OAI211_X1 U22932 ( .C1(n19908), .C2(n19946), .A(n19907), .B(n19906), .ZN(
        P2_U3170) );
  AOI22_X1 U22933 ( .A1(n19939), .A2(n19447), .B1(n19938), .B2(n19909), .ZN(
        n19913) );
  AOI22_X1 U22934 ( .A1(n19942), .A2(n19911), .B1(n19931), .B2(n19910), .ZN(
        n19912) );
  OAI211_X1 U22935 ( .C1(n19936), .C2(n19914), .A(n19913), .B(n19912), .ZN(
        P2_U3171) );
  AOI22_X1 U22936 ( .A1(n19939), .A2(n19916), .B1(n19938), .B2(n19915), .ZN(
        n19919) );
  AOI22_X1 U22937 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19917), .ZN(n19918) );
  OAI211_X1 U22938 ( .C1(n19920), .C2(n19946), .A(n19919), .B(n19918), .ZN(
        P2_U3172) );
  AOI22_X1 U22939 ( .A1(n19939), .A2(n19922), .B1(n19938), .B2(n19921), .ZN(
        n19925) );
  AOI22_X1 U22940 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19943), .B1(
        n19931), .B2(n19923), .ZN(n19924) );
  OAI211_X1 U22941 ( .C1(n19927), .C2(n19926), .A(n19925), .B(n19924), .ZN(
        P2_U3173) );
  AOI22_X1 U22942 ( .A1(n19939), .A2(n19929), .B1(n19938), .B2(n19928), .ZN(
        n19934) );
  AOI22_X1 U22943 ( .A1(n19942), .A2(n19932), .B1(n19931), .B2(n19930), .ZN(
        n19933) );
  OAI211_X1 U22944 ( .C1(n19936), .C2(n19935), .A(n19934), .B(n19933), .ZN(
        P2_U3174) );
  AOI22_X1 U22945 ( .A1(n19940), .A2(n19939), .B1(n19938), .B2(n19937), .ZN(
        n19945) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n19941), .ZN(n19944) );
  OAI211_X1 U22947 ( .C1(n19947), .C2(n19946), .A(n19945), .B(n19944), .ZN(
        P2_U3175) );
  OAI211_X1 U22948 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19950), .A(n19949), 
        .B(n19948), .ZN(n19955) );
  OAI21_X1 U22949 ( .B1(n19952), .B2(n19951), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19954) );
  OAI211_X1 U22950 ( .C1(n19956), .C2(n19955), .A(n19954), .B(n19953), .ZN(
        P2_U3177) );
  AND2_X1 U22951 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19957), .ZN(
        P2_U3179) );
  AND2_X1 U22952 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19957), .ZN(
        P2_U3180) );
  AND2_X1 U22953 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19957), .ZN(
        P2_U3181) );
  AND2_X1 U22954 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19957), .ZN(
        P2_U3182) );
  AND2_X1 U22955 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19957), .ZN(
        P2_U3183) );
  AND2_X1 U22956 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19957), .ZN(
        P2_U3184) );
  AND2_X1 U22957 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19957), .ZN(
        P2_U3185) );
  AND2_X1 U22958 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19957), .ZN(
        P2_U3186) );
  AND2_X1 U22959 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19957), .ZN(
        P2_U3187) );
  AND2_X1 U22960 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19957), .ZN(
        P2_U3188) );
  AND2_X1 U22961 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19957), .ZN(
        P2_U3189) );
  AND2_X1 U22962 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19957), .ZN(
        P2_U3190) );
  AND2_X1 U22963 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19957), .ZN(
        P2_U3191) );
  AND2_X1 U22964 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19957), .ZN(
        P2_U3192) );
  AND2_X1 U22965 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19957), .ZN(
        P2_U3193) );
  AND2_X1 U22966 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19957), .ZN(
        P2_U3194) );
  AND2_X1 U22967 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19957), .ZN(
        P2_U3195) );
  AND2_X1 U22968 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19957), .ZN(
        P2_U3196) );
  AND2_X1 U22969 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19957), .ZN(
        P2_U3197) );
  AND2_X1 U22970 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19957), .ZN(
        P2_U3198) );
  AND2_X1 U22971 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19957), .ZN(
        P2_U3199) );
  AND2_X1 U22972 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19957), .ZN(
        P2_U3200) );
  AND2_X1 U22973 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19957), .ZN(P2_U3201) );
  AND2_X1 U22974 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19957), .ZN(P2_U3202) );
  AND2_X1 U22975 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19957), .ZN(P2_U3203) );
  AND2_X1 U22976 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19957), .ZN(P2_U3204) );
  AND2_X1 U22977 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19957), .ZN(P2_U3205) );
  AND2_X1 U22978 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19957), .ZN(P2_U3206) );
  AND2_X1 U22979 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19957), .ZN(P2_U3207) );
  AND2_X1 U22980 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19957), .ZN(P2_U3208) );
  NAND2_X1 U22981 ( .A1(n19958), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19970) );
  INV_X1 U22982 ( .A(n19970), .ZN(n19975) );
  INV_X1 U22983 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19964) );
  NOR3_X1 U22984 ( .A1(n19975), .A2(n19964), .A3(n19959), .ZN(n19963) );
  AOI21_X1 U22985 ( .B1(n21254), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n19960), .ZN(n19961) );
  INV_X1 U22986 ( .A(n19961), .ZN(n19962) );
  NAND2_X1 U22987 ( .A1(NA), .A2(n19965), .ZN(n19973) );
  OAI211_X1 U22988 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19963), .A(n19962), 
        .B(n19973), .ZN(P2_U3209) );
  NAND2_X1 U22989 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21254), .ZN(n19974) );
  AOI211_X1 U22990 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19974), .A(n19965), 
        .B(n19964), .ZN(n19966) );
  NOR3_X1 U22991 ( .A1(n19967), .A2(n19975), .A3(n19966), .ZN(n19968) );
  OAI21_X1 U22992 ( .B1(n21254), .B2(n19969), .A(n19968), .ZN(P2_U3210) );
  OAI22_X1 U22993 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19971), .B1(NA), 
        .B2(n19970), .ZN(n19972) );
  OAI211_X1 U22994 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19972), .ZN(n19977) );
  OAI211_X1 U22995 ( .C1(n19975), .C2(n19974), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n19973), .ZN(n19976) );
  NAND2_X1 U22996 ( .A1(n19977), .A2(n19976), .ZN(P2_U3211) );
  OAI222_X1 U22997 ( .A1(n20042), .A2(n19982), .B1(n19980), .B2(n20036), .C1(
        n19979), .C2(n20038), .ZN(P2_U3212) );
  OAI222_X1 U22998 ( .A1(n20038), .A2(n19982), .B1(n19981), .B2(n20036), .C1(
        n19984), .C2(n20042), .ZN(P2_U3213) );
  OAI222_X1 U22999 ( .A1(n20038), .A2(n19984), .B1(n19983), .B2(n20036), .C1(
        n19985), .C2(n20042), .ZN(P2_U3214) );
  INV_X1 U23000 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19987) );
  OAI222_X1 U23001 ( .A1(n20042), .A2(n19987), .B1(n19986), .B2(n20036), .C1(
        n19985), .C2(n20038), .ZN(P2_U3215) );
  INV_X1 U23002 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19989) );
  OAI222_X1 U23003 ( .A1(n20042), .A2(n19989), .B1(n19988), .B2(n20036), .C1(
        n19987), .C2(n20038), .ZN(P2_U3216) );
  INV_X1 U23004 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19991) );
  OAI222_X1 U23005 ( .A1(n20042), .A2(n19991), .B1(n19990), .B2(n20036), .C1(
        n19989), .C2(n20038), .ZN(P2_U3217) );
  OAI222_X1 U23006 ( .A1(n20042), .A2(n19993), .B1(n19992), .B2(n20036), .C1(
        n19991), .C2(n20038), .ZN(P2_U3218) );
  INV_X1 U23007 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19995) );
  OAI222_X1 U23008 ( .A1(n20042), .A2(n19995), .B1(n19994), .B2(n20036), .C1(
        n19993), .C2(n20038), .ZN(P2_U3219) );
  OAI222_X1 U23009 ( .A1(n20042), .A2(n19997), .B1(n19996), .B2(n20036), .C1(
        n19995), .C2(n20038), .ZN(P2_U3220) );
  INV_X1 U23010 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19999) );
  OAI222_X1 U23011 ( .A1(n20042), .A2(n19999), .B1(n19998), .B2(n20036), .C1(
        n19997), .C2(n20038), .ZN(P2_U3221) );
  OAI222_X1 U23012 ( .A1(n20042), .A2(n20001), .B1(n20000), .B2(n20036), .C1(
        n19999), .C2(n20038), .ZN(P2_U3222) );
  OAI222_X1 U23013 ( .A1(n20042), .A2(n20003), .B1(n20002), .B2(n20036), .C1(
        n20001), .C2(n20038), .ZN(P2_U3223) );
  OAI222_X1 U23014 ( .A1(n20042), .A2(n20005), .B1(n20004), .B2(n20036), .C1(
        n20003), .C2(n20038), .ZN(P2_U3224) );
  INV_X1 U23015 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U23016 ( .A1(n20042), .A2(n20007), .B1(n20006), .B2(n20036), .C1(
        n20005), .C2(n20038), .ZN(P2_U3225) );
  OAI222_X1 U23017 ( .A1(n20042), .A2(n20009), .B1(n20008), .B2(n20036), .C1(
        n20007), .C2(n20038), .ZN(P2_U3226) );
  OAI222_X1 U23018 ( .A1(n20042), .A2(n20011), .B1(n20010), .B2(n20036), .C1(
        n20009), .C2(n20038), .ZN(P2_U3227) );
  OAI222_X1 U23019 ( .A1(n20042), .A2(n20013), .B1(n20012), .B2(n20036), .C1(
        n20011), .C2(n20038), .ZN(P2_U3228) );
  OAI222_X1 U23020 ( .A1(n20042), .A2(n20015), .B1(n20014), .B2(n20036), .C1(
        n20013), .C2(n20038), .ZN(P2_U3229) );
  OAI222_X1 U23021 ( .A1(n20042), .A2(n20017), .B1(n20016), .B2(n20036), .C1(
        n20015), .C2(n20038), .ZN(P2_U3230) );
  OAI222_X1 U23022 ( .A1(n20042), .A2(n20019), .B1(n20018), .B2(n20036), .C1(
        n20017), .C2(n20038), .ZN(P2_U3231) );
  OAI222_X1 U23023 ( .A1(n20042), .A2(n20021), .B1(n20020), .B2(n20036), .C1(
        n20019), .C2(n20038), .ZN(P2_U3232) );
  OAI222_X1 U23024 ( .A1(n20042), .A2(n20023), .B1(n20022), .B2(n20036), .C1(
        n20021), .C2(n20038), .ZN(P2_U3233) );
  OAI222_X1 U23025 ( .A1(n20042), .A2(n20025), .B1(n20024), .B2(n20036), .C1(
        n20023), .C2(n20038), .ZN(P2_U3234) );
  INV_X1 U23026 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20027) );
  OAI222_X1 U23027 ( .A1(n20042), .A2(n20027), .B1(n20026), .B2(n20036), .C1(
        n20025), .C2(n20038), .ZN(P2_U3235) );
  INV_X1 U23028 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20029) );
  OAI222_X1 U23029 ( .A1(n20042), .A2(n20029), .B1(n20028), .B2(n20036), .C1(
        n20027), .C2(n20038), .ZN(P2_U3236) );
  INV_X1 U23030 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20032) );
  OAI222_X1 U23031 ( .A1(n20042), .A2(n20032), .B1(n20030), .B2(n20036), .C1(
        n20029), .C2(n20038), .ZN(P2_U3237) );
  OAI222_X1 U23032 ( .A1(n20038), .A2(n20032), .B1(n20031), .B2(n20036), .C1(
        n20033), .C2(n20042), .ZN(P2_U3238) );
  INV_X1 U23033 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20035) );
  OAI222_X1 U23034 ( .A1(n20042), .A2(n20035), .B1(n20034), .B2(n20036), .C1(
        n20033), .C2(n20038), .ZN(P2_U3239) );
  INV_X1 U23035 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20039) );
  OAI222_X1 U23036 ( .A1(n20042), .A2(n20039), .B1(n20037), .B2(n20036), .C1(
        n20035), .C2(n20038), .ZN(P2_U3240) );
  INV_X1 U23037 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20041) );
  INV_X1 U23038 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20040) );
  OAI222_X1 U23039 ( .A1(n20042), .A2(n20041), .B1(n20040), .B2(n20036), .C1(
        n20039), .C2(n20038), .ZN(P2_U3241) );
  INV_X1 U23040 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20043) );
  AOI22_X1 U23041 ( .A1(n20036), .A2(n20044), .B1(n20043), .B2(n20100), .ZN(
        P2_U3585) );
  MUX2_X1 U23042 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20036), .Z(P2_U3586) );
  INV_X1 U23043 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U23044 ( .A1(n20036), .A2(n20046), .B1(n20045), .B2(n20100), .ZN(
        P2_U3587) );
  INV_X1 U23045 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U23046 ( .A1(n20036), .A2(n20048), .B1(n20047), .B2(n20100), .ZN(
        P2_U3588) );
  OAI21_X1 U23047 ( .B1(n20052), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20050), 
        .ZN(n20049) );
  INV_X1 U23048 ( .A(n20049), .ZN(P2_U3591) );
  OAI21_X1 U23049 ( .B1(n20052), .B2(n20051), .A(n20050), .ZN(P2_U3592) );
  AND2_X1 U23050 ( .A1(n20057), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20074) );
  NAND2_X1 U23051 ( .A1(n20053), .A2(n20074), .ZN(n20063) );
  NAND3_X1 U23052 ( .A1(n20072), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20054), 
        .ZN(n20055) );
  NAND2_X1 U23053 ( .A1(n20055), .A2(n20070), .ZN(n20064) );
  NAND2_X1 U23054 ( .A1(n20063), .A2(n20064), .ZN(n20060) );
  AOI222_X1 U23055 ( .A1(n20060), .A2(n20059), .B1(n20058), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n20057), .C2(n20056), .ZN(n20061) );
  AOI22_X1 U23056 ( .A1(n20087), .A2(n20062), .B1(n20061), .B2(n20084), .ZN(
        P2_U3602) );
  OAI21_X1 U23057 ( .B1(n20065), .B2(n20064), .A(n20063), .ZN(n20066) );
  AOI21_X1 U23058 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20067), .A(n20066), 
        .ZN(n20068) );
  AOI22_X1 U23059 ( .A1(n20087), .A2(n20069), .B1(n20068), .B2(n20084), .ZN(
        P2_U3603) );
  INV_X1 U23060 ( .A(n20070), .ZN(n20080) );
  NOR2_X1 U23061 ( .A1(n20080), .A2(n20071), .ZN(n20073) );
  MUX2_X1 U23062 ( .A(n20074), .B(n20073), .S(n20072), .Z(n20075) );
  AOI21_X1 U23063 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20076), .A(n20075), 
        .ZN(n20077) );
  AOI22_X1 U23064 ( .A1(n20087), .A2(n20078), .B1(n20077), .B2(n20084), .ZN(
        P2_U3604) );
  OAI22_X1 U23065 ( .A1(n20081), .A2(n20080), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20079), .ZN(n20082) );
  AOI21_X1 U23066 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20083), .A(n20082), 
        .ZN(n20085) );
  AOI22_X1 U23067 ( .A1(n20087), .A2(n20086), .B1(n20085), .B2(n20084), .ZN(
        P2_U3605) );
  INV_X1 U23068 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20088) );
  AOI22_X1 U23069 ( .A1(n20036), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20088), 
        .B2(n20100), .ZN(P2_U3608) );
  INV_X1 U23070 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20099) );
  INV_X1 U23071 ( .A(n20089), .ZN(n20098) );
  INV_X1 U23072 ( .A(n20090), .ZN(n20094) );
  AOI22_X1 U23073 ( .A1(n20094), .A2(n20093), .B1(n20092), .B2(n20091), .ZN(
        n20097) );
  NOR2_X1 U23074 ( .A1(n20098), .A2(n20095), .ZN(n20096) );
  AOI22_X1 U23075 ( .A1(n20099), .A2(n20098), .B1(n20097), .B2(n20096), .ZN(
        P2_U3609) );
  INV_X1 U23076 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20101) );
  AOI22_X1 U23077 ( .A1(n20036), .A2(n20102), .B1(n20101), .B2(n20100), .ZN(
        P2_U3611) );
  NAND2_X1 U23078 ( .A1(n20920), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21023) );
  AOI21_X1 U23079 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20924), .A(n20972), 
        .ZN(n20984) );
  AOI21_X1 U23080 ( .B1(n21023), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20984), .ZN(
        n20103) );
  INV_X1 U23081 ( .A(n20103), .ZN(P1_U2802) );
  NOR2_X1 U23082 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20105) );
  OAI21_X1 U23083 ( .B1(n20105), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21023), .ZN(
        n20104) );
  OAI21_X1 U23084 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21023), .A(n20104), 
        .ZN(P1_U2804) );
  OAI21_X1 U23085 ( .B1(BS16), .B2(n20105), .A(n20984), .ZN(n20982) );
  OAI21_X1 U23086 ( .B1(n20984), .B2(n21346), .A(n20982), .ZN(P1_U2805) );
  NAND2_X1 U23087 ( .A1(n20107), .A2(n20106), .ZN(n21002) );
  INV_X1 U23088 ( .A(n21002), .ZN(n21004) );
  OAI21_X1 U23089 ( .B1(n21004), .B2(n21213), .A(n20108), .ZN(P1_U2806) );
  NOR4_X1 U23090 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20112) );
  NOR4_X1 U23091 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20111) );
  NOR4_X1 U23092 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20110) );
  NOR4_X1 U23093 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20109) );
  NAND4_X1 U23094 ( .A1(n20112), .A2(n20111), .A3(n20110), .A4(n20109), .ZN(
        n20118) );
  NOR4_X1 U23095 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20116) );
  AOI211_X1 U23096 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20115) );
  NOR4_X1 U23097 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20114) );
  NOR4_X1 U23098 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20113) );
  NAND4_X1 U23099 ( .A1(n20116), .A2(n20115), .A3(n20114), .A4(n20113), .ZN(
        n20117) );
  NOR2_X1 U23100 ( .A1(n20118), .A2(n20117), .ZN(n20999) );
  INV_X1 U23101 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21190) );
  NOR3_X1 U23102 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20120) );
  OAI21_X1 U23103 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20120), .A(n20999), .ZN(
        n20119) );
  OAI21_X1 U23104 ( .B1(n20999), .B2(n21190), .A(n20119), .ZN(P1_U2807) );
  INV_X1 U23105 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20983) );
  AOI21_X1 U23106 ( .B1(n21352), .B2(n20983), .A(n20120), .ZN(n20121) );
  INV_X1 U23107 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21167) );
  INV_X1 U23108 ( .A(n20999), .ZN(n21001) );
  AOI22_X1 U23109 ( .A1(n20999), .A2(n20121), .B1(n21167), .B2(n21001), .ZN(
        P1_U2808) );
  NAND2_X1 U23110 ( .A1(n20123), .A2(n20122), .ZN(n20138) );
  AOI22_X1 U23111 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20177), .B1(n20186), .B2(
        n20203), .ZN(n20124) );
  OAI21_X1 U23112 ( .B1(n21219), .B2(n20138), .A(n20124), .ZN(n20125) );
  AOI211_X1 U23113 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20153), .B(n20125), .ZN(n20128) );
  AOI22_X1 U23114 ( .A1(n20204), .A2(n20155), .B1(n20191), .B2(n20126), .ZN(
        n20127) );
  OAI211_X1 U23115 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20129), .A(n20128), .B(
        n20127), .ZN(P1_U2831) );
  NOR2_X1 U23116 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n9954), .ZN(n20139) );
  OAI22_X1 U23117 ( .A1(n21250), .A2(n20201), .B1(n20174), .B2(n20130), .ZN(
        n20131) );
  AOI211_X1 U23118 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20153), .B(n20131), .ZN(n20137) );
  OAI22_X1 U23119 ( .A1(n20134), .A2(n20133), .B1(n20132), .B2(n20184), .ZN(
        n20135) );
  INV_X1 U23120 ( .A(n20135), .ZN(n20136) );
  OAI211_X1 U23121 ( .C1(n20139), .C2(n20138), .A(n20137), .B(n20136), .ZN(
        P1_U2832) );
  AOI22_X1 U23122 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20177), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n10498), .ZN(n20141) );
  OAI211_X1 U23123 ( .C1(n20172), .C2(n20142), .A(n20170), .B(n20141), .ZN(
        n20143) );
  AOI21_X1 U23124 ( .B1(n20144), .B2(n20186), .A(n20143), .ZN(n20145) );
  OAI21_X1 U23125 ( .B1(n20146), .B2(P1_REIP_REG_7__SCAN_IN), .A(n20145), .ZN(
        n20147) );
  AOI21_X1 U23126 ( .B1(n20148), .B2(n20155), .A(n20147), .ZN(n20149) );
  OAI21_X1 U23127 ( .B1(n20150), .B2(n20184), .A(n20149), .ZN(P1_U2833) );
  OAI22_X1 U23128 ( .A1(n21334), .A2(n20201), .B1(n20174), .B2(n20151), .ZN(
        n20152) );
  AOI211_X1 U23129 ( .C1(n20190), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20153), .B(n20152), .ZN(n20158) );
  INV_X1 U23130 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21368) );
  NAND2_X1 U23131 ( .A1(n20179), .A2(n20162), .ZN(n20164) );
  OAI21_X1 U23132 ( .B1(n21368), .B2(n20164), .A(n13564), .ZN(n20154) );
  AOI22_X1 U23133 ( .A1(n20156), .A2(n20155), .B1(n10498), .B2(n20154), .ZN(
        n20157) );
  OAI211_X1 U23134 ( .C1(n20159), .C2(n20184), .A(n20158), .B(n20157), .ZN(
        P1_U2834) );
  INV_X1 U23135 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20210) );
  AOI21_X1 U23136 ( .B1(n20162), .B2(n20161), .A(n20160), .ZN(n20180) );
  AOI22_X1 U23137 ( .A1(n20186), .A2(n9951), .B1(P1_REIP_REG_5__SCAN_IN), .B2(
        n20180), .ZN(n20163) );
  OAI211_X1 U23138 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20164), .A(n20170), .B(
        n20163), .ZN(n20165) );
  AOI21_X1 U23139 ( .B1(n20190), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20165), .ZN(n20166) );
  OAI21_X1 U23140 ( .B1(n20201), .B2(n20210), .A(n20166), .ZN(n20167) );
  AOI21_X1 U23141 ( .B1(n20208), .B2(n20197), .A(n20167), .ZN(n20168) );
  OAI21_X1 U23142 ( .B1(n20169), .B2(n20184), .A(n20168), .ZN(P1_U2835) );
  INV_X1 U23143 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20171) );
  OAI21_X1 U23144 ( .B1(n20172), .B2(n20171), .A(n20170), .ZN(n20176) );
  OAI22_X1 U23145 ( .A1(n20174), .A2(n20306), .B1(n20173), .B2(n20187), .ZN(
        n20175) );
  AOI211_X1 U23146 ( .C1(P1_EBX_REG_4__SCAN_IN), .C2(n20177), .A(n20176), .B(
        n20175), .ZN(n20183) );
  INV_X1 U23147 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21187) );
  NAND2_X1 U23148 ( .A1(n20179), .A2(n20178), .ZN(n20194) );
  INV_X1 U23149 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21375) );
  OAI21_X1 U23150 ( .B1(n21187), .B2(n20194), .A(n21375), .ZN(n20181) );
  AOI22_X1 U23151 ( .A1(n20297), .A2(n20197), .B1(n20181), .B2(n20180), .ZN(
        n20182) );
  OAI211_X1 U23152 ( .C1(n20301), .C2(n20184), .A(n20183), .B(n20182), .ZN(
        P1_U2836) );
  AOI22_X1 U23153 ( .A1(n20186), .A2(n20315), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20185), .ZN(n20200) );
  INV_X1 U23154 ( .A(n20594), .ZN(n20188) );
  NOR2_X1 U23155 ( .A1(n20188), .A2(n20187), .ZN(n20196) );
  INV_X1 U23156 ( .A(n20189), .ZN(n20192) );
  AOI22_X1 U23157 ( .A1(n20192), .A2(n20191), .B1(n20190), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20193) );
  OAI21_X1 U23158 ( .B1(n20194), .B2(P1_REIP_REG_3__SCAN_IN), .A(n20193), .ZN(
        n20195) );
  AOI211_X1 U23159 ( .C1(n20198), .C2(n20197), .A(n20196), .B(n20195), .ZN(
        n20199) );
  OAI211_X1 U23160 ( .C1(n20202), .C2(n20201), .A(n20200), .B(n20199), .ZN(
        P1_U2837) );
  INV_X1 U23161 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21381) );
  AOI22_X1 U23162 ( .A1(n20204), .A2(n20207), .B1(n20206), .B2(n20203), .ZN(
        n20205) );
  OAI21_X1 U23163 ( .B1(n20211), .B2(n21381), .A(n20205), .ZN(P1_U2863) );
  AOI22_X1 U23164 ( .A1(n20208), .A2(n20207), .B1(n20206), .B2(n9951), .ZN(
        n20209) );
  OAI21_X1 U23165 ( .B1(n20211), .B2(n20210), .A(n20209), .ZN(P1_U2867) );
  AOI22_X1 U23166 ( .A1(n20241), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20213) );
  OAI21_X1 U23167 ( .B1(n20214), .B2(n20243), .A(n20213), .ZN(P1_U2921) );
  INV_X1 U23168 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U23169 ( .A1(n20241), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20215) );
  OAI21_X1 U23170 ( .B1(n20216), .B2(n20243), .A(n20215), .ZN(P1_U2922) );
  INV_X1 U23171 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U23172 ( .A1(n20241), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20217) );
  OAI21_X1 U23173 ( .B1(n20218), .B2(n20243), .A(n20217), .ZN(P1_U2923) );
  AOI22_X1 U23174 ( .A1(n20241), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20219) );
  OAI21_X1 U23175 ( .B1(n14381), .B2(n20243), .A(n20219), .ZN(P1_U2924) );
  INV_X1 U23176 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20221) );
  AOI22_X1 U23177 ( .A1(n20241), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20220) );
  OAI21_X1 U23178 ( .B1(n20221), .B2(n20243), .A(n20220), .ZN(P1_U2925) );
  INV_X1 U23179 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20223) );
  AOI22_X1 U23180 ( .A1(n20241), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20222) );
  OAI21_X1 U23181 ( .B1(n20223), .B2(n20243), .A(n20222), .ZN(P1_U2926) );
  INV_X1 U23182 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20226) );
  AOI22_X1 U23183 ( .A1(n20241), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20225) );
  OAI21_X1 U23184 ( .B1(n20226), .B2(n20243), .A(n20225), .ZN(P1_U2927) );
  AOI22_X1 U23185 ( .A1(n20241), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20227) );
  OAI21_X1 U23186 ( .B1(n20228), .B2(n20243), .A(n20227), .ZN(P1_U2928) );
  AOI22_X1 U23187 ( .A1(n20241), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20229) );
  OAI21_X1 U23188 ( .B1(n20230), .B2(n20243), .A(n20229), .ZN(P1_U2929) );
  AOI22_X1 U23189 ( .A1(n20241), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20231) );
  OAI21_X1 U23190 ( .B1(n10981), .B2(n20243), .A(n20231), .ZN(P1_U2930) );
  AOI22_X1 U23191 ( .A1(n20241), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20232) );
  OAI21_X1 U23192 ( .B1(n10962), .B2(n20243), .A(n20232), .ZN(P1_U2931) );
  AOI22_X1 U23193 ( .A1(n20241), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20233) );
  OAI21_X1 U23194 ( .B1(n20234), .B2(n20243), .A(n20233), .ZN(P1_U2932) );
  AOI22_X1 U23195 ( .A1(n20241), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20235) );
  OAI21_X1 U23196 ( .B1(n20236), .B2(n20243), .A(n20235), .ZN(P1_U2933) );
  AOI22_X1 U23197 ( .A1(n20241), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20237) );
  OAI21_X1 U23198 ( .B1(n20238), .B2(n20243), .A(n20237), .ZN(P1_U2934) );
  AOI22_X1 U23199 ( .A1(n20241), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20239) );
  OAI21_X1 U23200 ( .B1(n20240), .B2(n20243), .A(n20239), .ZN(P1_U2935) );
  AOI22_X1 U23201 ( .A1(n20241), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20224), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20242) );
  OAI21_X1 U23202 ( .B1(n20244), .B2(n20243), .A(n20242), .ZN(P1_U2936) );
  AOI22_X1 U23203 ( .A1(n20287), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20286), .ZN(n20246) );
  OAI21_X1 U23204 ( .B1(n20255), .B2(n20289), .A(n20246), .ZN(P1_U2937) );
  AOI22_X1 U23205 ( .A1(n20287), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20286), .ZN(n20247) );
  OAI21_X1 U23206 ( .B1(n20357), .B2(n20289), .A(n20247), .ZN(P1_U2938) );
  AOI22_X1 U23207 ( .A1(n20287), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20286), .ZN(n20248) );
  OAI21_X1 U23208 ( .B1(n20258), .B2(n20289), .A(n20248), .ZN(P1_U2939) );
  AOI22_X1 U23209 ( .A1(n20287), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20286), .ZN(n20249) );
  OAI21_X1 U23210 ( .B1(n20260), .B2(n20289), .A(n20249), .ZN(P1_U2940) );
  AOI22_X1 U23211 ( .A1(n20287), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20286), .ZN(n20250) );
  OAI21_X1 U23212 ( .B1(n20262), .B2(n20289), .A(n20250), .ZN(P1_U2941) );
  AOI22_X1 U23213 ( .A1(n20287), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20286), .ZN(n20251) );
  OAI21_X1 U23214 ( .B1(n20367), .B2(n20289), .A(n20251), .ZN(P1_U2942) );
  AOI22_X1 U23215 ( .A1(n20287), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20286), .ZN(n20252) );
  OAI21_X1 U23216 ( .B1(n20376), .B2(n20289), .A(n20252), .ZN(P1_U2943) );
  AOI22_X1 U23217 ( .A1(n20287), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20286), .ZN(n20253) );
  OAI21_X1 U23218 ( .B1(n20266), .B2(n20289), .A(n20253), .ZN(P1_U2944) );
  AOI22_X1 U23219 ( .A1(n20287), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20286), .ZN(n20254) );
  OAI21_X1 U23220 ( .B1(n20255), .B2(n20289), .A(n20254), .ZN(P1_U2952) );
  AOI22_X1 U23221 ( .A1(n20287), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20286), .ZN(n20256) );
  OAI21_X1 U23222 ( .B1(n20357), .B2(n20289), .A(n20256), .ZN(P1_U2953) );
  AOI22_X1 U23223 ( .A1(n20287), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20286), .ZN(n20257) );
  OAI21_X1 U23224 ( .B1(n20258), .B2(n20289), .A(n20257), .ZN(P1_U2954) );
  AOI22_X1 U23225 ( .A1(n20287), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20286), .ZN(n20259) );
  OAI21_X1 U23226 ( .B1(n20260), .B2(n20289), .A(n20259), .ZN(P1_U2955) );
  AOI22_X1 U23227 ( .A1(n20287), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20286), .ZN(n20261) );
  OAI21_X1 U23228 ( .B1(n20262), .B2(n20289), .A(n20261), .ZN(P1_U2956) );
  AOI22_X1 U23229 ( .A1(n20287), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20286), .ZN(n20263) );
  OAI21_X1 U23230 ( .B1(n20367), .B2(n20289), .A(n20263), .ZN(P1_U2957) );
  AOI22_X1 U23231 ( .A1(n20287), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20286), .ZN(n20264) );
  OAI21_X1 U23232 ( .B1(n20376), .B2(n20289), .A(n20264), .ZN(P1_U2958) );
  AOI22_X1 U23233 ( .A1(n20287), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20286), .ZN(n20265) );
  OAI21_X1 U23234 ( .B1(n20266), .B2(n20289), .A(n20265), .ZN(P1_U2959) );
  AOI22_X1 U23235 ( .A1(n20287), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20286), .ZN(n20269) );
  NAND2_X1 U23236 ( .A1(n20283), .A2(n20267), .ZN(n20268) );
  NAND2_X1 U23237 ( .A1(n20269), .A2(n20268), .ZN(P1_U2961) );
  AOI22_X1 U23238 ( .A1(n20287), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20286), .ZN(n20272) );
  NAND2_X1 U23239 ( .A1(n20283), .A2(n20270), .ZN(n20271) );
  NAND2_X1 U23240 ( .A1(n20272), .A2(n20271), .ZN(P1_U2962) );
  AOI22_X1 U23241 ( .A1(n20287), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20286), .ZN(n20275) );
  NAND2_X1 U23242 ( .A1(n20283), .A2(n20273), .ZN(n20274) );
  NAND2_X1 U23243 ( .A1(n20275), .A2(n20274), .ZN(P1_U2963) );
  AOI22_X1 U23244 ( .A1(n20287), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20286), .ZN(n20278) );
  NAND2_X1 U23245 ( .A1(n20283), .A2(n20276), .ZN(n20277) );
  NAND2_X1 U23246 ( .A1(n20278), .A2(n20277), .ZN(P1_U2964) );
  AOI22_X1 U23247 ( .A1(n20287), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20286), .ZN(n20281) );
  NAND2_X1 U23248 ( .A1(n20283), .A2(n20279), .ZN(n20280) );
  NAND2_X1 U23249 ( .A1(n20281), .A2(n20280), .ZN(P1_U2965) );
  AOI22_X1 U23250 ( .A1(n20287), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20286), .ZN(n20285) );
  NAND2_X1 U23251 ( .A1(n20283), .A2(n20282), .ZN(n20284) );
  NAND2_X1 U23252 ( .A1(n20285), .A2(n20284), .ZN(P1_U2966) );
  AOI22_X1 U23253 ( .A1(n20287), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n20286), .ZN(n20288) );
  OAI21_X1 U23254 ( .B1(n20290), .B2(n20289), .A(n20288), .ZN(P1_U2967) );
  AOI22_X1 U23255 ( .A1(n20291), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20317), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20300) );
  OAI21_X1 U23256 ( .B1(n20294), .B2(n20293), .A(n20292), .ZN(n20295) );
  INV_X1 U23257 ( .A(n20295), .ZN(n20310) );
  AOI22_X1 U23258 ( .A1(n20310), .A2(n20298), .B1(n20297), .B2(n20296), .ZN(
        n20299) );
  OAI211_X1 U23259 ( .C1(n20302), .C2(n20301), .A(n20300), .B(n20299), .ZN(
        P1_U2995) );
  INV_X1 U23260 ( .A(n20303), .ZN(n20305) );
  NOR2_X1 U23261 ( .A1(n20323), .A2(n20304), .ZN(n20331) );
  AOI211_X1 U23262 ( .C1(n20327), .C2(n20305), .A(n20331), .B(n20325), .ZN(
        n20319) );
  OAI22_X1 U23263 ( .A1(n20344), .A2(n20306), .B1(n21375), .B2(n20342), .ZN(
        n20309) );
  AOI211_X1 U23264 ( .C1(n20312), .C2(n20320), .A(n20307), .B(n20321), .ZN(
        n20308) );
  AOI211_X1 U23265 ( .C1(n20310), .C2(n20332), .A(n20309), .B(n20308), .ZN(
        n20311) );
  OAI21_X1 U23266 ( .B1(n20319), .B2(n20312), .A(n20311), .ZN(P1_U3027) );
  INV_X1 U23267 ( .A(n20313), .ZN(n20314) );
  AOI222_X1 U23268 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20317), .B1(n20316), 
        .B2(n20315), .C1(n20332), .C2(n20314), .ZN(n20318) );
  OAI221_X1 U23269 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20321), .C1(
        n20320), .C2(n20319), .A(n20318), .ZN(P1_U3028) );
  NAND2_X1 U23270 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20322), .ZN(
        n20337) );
  NOR3_X1 U23271 ( .A1(n20324), .A2(n20350), .A3(n20323), .ZN(n20326) );
  AOI211_X1 U23272 ( .C1(n20350), .C2(n20327), .A(n20326), .B(n20325), .ZN(
        n20335) );
  INV_X1 U23273 ( .A(n20328), .ZN(n20333) );
  OAI22_X1 U23274 ( .A1(n20344), .A2(n20329), .B1(n20935), .B2(n20342), .ZN(
        n20330) );
  AOI211_X1 U23275 ( .C1(n20333), .C2(n20332), .A(n20331), .B(n20330), .ZN(
        n20334) );
  OAI221_X1 U23276 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20337), .C1(
        n20336), .C2(n20335), .A(n20334), .ZN(P1_U3029) );
  NAND2_X1 U23277 ( .A1(n20339), .A2(n20338), .ZN(n20351) );
  NOR2_X1 U23278 ( .A1(n20341), .A2(n20340), .ZN(n20347) );
  OAI22_X1 U23279 ( .A1(n20344), .A2(n20343), .B1(n21352), .B2(n20342), .ZN(
        n20345) );
  AOI21_X1 U23280 ( .B1(n20347), .B2(n20346), .A(n20345), .ZN(n20348) );
  OAI221_X1 U23281 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20351), .C1(
        n20350), .C2(n20349), .A(n20348), .ZN(P1_U3030) );
  NOR2_X1 U23282 ( .A1(n20353), .A2(n20352), .ZN(P1_U3032) );
  INV_X1 U23283 ( .A(DATAI_25_), .ZN(n21165) );
  OAI22_X2 U23284 ( .A1(n20354), .A2(n20377), .B1(n21165), .B2(n20379), .ZN(
        n20866) );
  NOR2_X2 U23285 ( .A1(n20365), .A2(n20355), .ZN(n20865) );
  AOI22_X1 U23286 ( .A1(n20911), .A2(n20866), .B1(n20356), .B2(n20865), .ZN(
        n20361) );
  INV_X1 U23287 ( .A(DATAI_17_), .ZN(n20358) );
  OAI22_X1 U23288 ( .A1(n20359), .A2(n20377), .B1(n20358), .B2(n20379), .ZN(
        n20777) );
  AOI22_X1 U23289 ( .A1(n20864), .A2(n20380), .B1(n20407), .B2(n20777), .ZN(
        n20360) );
  OAI211_X1 U23290 ( .C1(n20384), .C2(n20362), .A(n20361), .B(n20360), .ZN(
        P1_U3034) );
  INV_X1 U23291 ( .A(DATAI_29_), .ZN(n20363) );
  OAI22_X1 U23292 ( .A1(n20364), .A2(n20377), .B1(n20363), .B2(n20379), .ZN(
        n20833) );
  INV_X1 U23293 ( .A(n20833), .ZN(n20897) );
  NOR2_X2 U23294 ( .A1(n20365), .A2(n9845), .ZN(n20893) );
  INV_X1 U23295 ( .A(n20893), .ZN(n20747) );
  OAI22_X1 U23296 ( .A1(n20904), .A2(n20897), .B1(n20374), .B2(n20747), .ZN(
        n20366) );
  INV_X1 U23297 ( .A(n20366), .ZN(n20370) );
  INV_X1 U23298 ( .A(DATAI_21_), .ZN(n21350) );
  OAI22_X2 U23299 ( .A1(n21350), .A2(n20379), .B1(n20368), .B2(n20377), .ZN(
        n20894) );
  AOI22_X1 U23300 ( .A1(n20892), .A2(n20380), .B1(n20407), .B2(n20894), .ZN(
        n20369) );
  OAI211_X1 U23301 ( .C1(n20384), .C2(n20371), .A(n20370), .B(n20369), .ZN(
        P1_U3038) );
  INV_X1 U23302 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20383) );
  INV_X1 U23303 ( .A(DATAI_30_), .ZN(n21054) );
  INV_X1 U23304 ( .A(n20900), .ZN(n20792) );
  NAND2_X1 U23305 ( .A1(n20373), .A2(n10694), .ZN(n20752) );
  OAI22_X1 U23306 ( .A1(n20904), .A2(n20792), .B1(n20374), .B2(n20752), .ZN(
        n20375) );
  INV_X1 U23307 ( .A(n20375), .ZN(n20382) );
  INV_X1 U23308 ( .A(DATAI_22_), .ZN(n21225) );
  OAI22_X1 U23309 ( .A1(n21225), .A2(n20379), .B1(n20378), .B2(n20377), .ZN(
        n20789) );
  AOI22_X1 U23310 ( .A1(n20898), .A2(n20380), .B1(n20407), .B2(n20789), .ZN(
        n20381) );
  OAI211_X1 U23311 ( .C1(n20384), .C2(n20383), .A(n20382), .B(n20381), .ZN(
        P1_U3039) );
  INV_X1 U23312 ( .A(n20773), .ZN(n20863) );
  INV_X1 U23313 ( .A(n20446), .ZN(n20386) );
  INV_X1 U23314 ( .A(n20385), .ZN(n20767) );
  NOR2_X1 U23315 ( .A1(n20766), .A2(n20387), .ZN(n20405) );
  AOI21_X1 U23316 ( .B1(n20386), .B2(n20767), .A(n20405), .ZN(n20388) );
  OAI22_X1 U23317 ( .A1(n20388), .A2(n20804), .B1(n20387), .B2(n20625), .ZN(
        n20406) );
  AOI22_X1 U23318 ( .A1(n20406), .A2(n20805), .B1(n20806), .B2(n20405), .ZN(
        n20392) );
  INV_X1 U23319 ( .A(n20387), .ZN(n20390) );
  OAI21_X1 U23320 ( .B1(n20455), .B2(n21346), .A(n20388), .ZN(n20389) );
  OAI221_X1 U23321 ( .B1(n20848), .B2(n20390), .C1(n20804), .C2(n20389), .A(
        n20858), .ZN(n20408) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20860), .ZN(n20391) );
  OAI211_X1 U23323 ( .C1(n20863), .C2(n20437), .A(n20392), .B(n20391), .ZN(
        P1_U3041) );
  INV_X1 U23324 ( .A(n20777), .ZN(n20869) );
  AOI22_X1 U23325 ( .A1(n20406), .A2(n20864), .B1(n20865), .B2(n20405), .ZN(
        n20394) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20866), .ZN(n20393) );
  OAI211_X1 U23327 ( .C1(n20869), .C2(n20437), .A(n20394), .B(n20393), .ZN(
        P1_U3042) );
  INV_X1 U23328 ( .A(n20873), .ZN(n20821) );
  AOI22_X1 U23329 ( .A1(n20406), .A2(n20816), .B1(n20817), .B2(n20405), .ZN(
        n20396) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20818), .ZN(n20395) );
  OAI211_X1 U23331 ( .C1(n20821), .C2(n20437), .A(n20396), .B(n20395), .ZN(
        P1_U3043) );
  AOI22_X1 U23332 ( .A1(n20406), .A2(n20822), .B1(n20823), .B2(n20405), .ZN(
        n20398) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20824), .ZN(n20397) );
  OAI211_X1 U23334 ( .C1(n20827), .C2(n20437), .A(n20398), .B(n20397), .ZN(
        P1_U3044) );
  AOI22_X1 U23335 ( .A1(n20406), .A2(n20828), .B1(n20829), .B2(n20405), .ZN(
        n20400) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20830), .ZN(n20399) );
  OAI211_X1 U23337 ( .C1(n9977), .C2(n20437), .A(n20400), .B(n20399), .ZN(
        P1_U3045) );
  INV_X1 U23338 ( .A(n20894), .ZN(n20836) );
  AOI22_X1 U23339 ( .A1(n20406), .A2(n20892), .B1(n20893), .B2(n20405), .ZN(
        n20402) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20833), .ZN(n20401) );
  OAI211_X1 U23341 ( .C1(n20836), .C2(n20437), .A(n20402), .B(n20401), .ZN(
        P1_U3046) );
  INV_X1 U23342 ( .A(n20789), .ZN(n20905) );
  AOI22_X1 U23343 ( .A1(n20406), .A2(n20898), .B1(n20899), .B2(n20405), .ZN(
        n20404) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20900), .ZN(n20403) );
  OAI211_X1 U23345 ( .C1(n20905), .C2(n20437), .A(n20404), .B(n20403), .ZN(
        P1_U3047) );
  AOI22_X1 U23346 ( .A1(n20406), .A2(n20907), .B1(n20909), .B2(n20405), .ZN(
        n20410) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20408), .B1(
        n20407), .B2(n20841), .ZN(n20409) );
  OAI211_X1 U23348 ( .C1(n20846), .C2(n20437), .A(n20410), .B(n20409), .ZN(
        P1_U3048) );
  NAND2_X1 U23349 ( .A1(n20437), .A2(n20848), .ZN(n20411) );
  NAND2_X1 U23350 ( .A1(n20848), .A2(n21346), .ZN(n20717) );
  OAI21_X1 U23351 ( .B1(n20471), .B2(n20411), .A(n20717), .ZN(n20414) );
  NOR2_X1 U23352 ( .A1(n20446), .A2(n20595), .ZN(n20412) );
  NOR3_X1 U23353 ( .A1(n20723), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20450) );
  AND2_X1 U23354 ( .A1(n20766), .A2(n20450), .ZN(n20426) );
  AOI22_X1 U23355 ( .A1(n20471), .A2(n20773), .B1(n20806), .B2(n20426), .ZN(
        n20417) );
  INV_X1 U23356 ( .A(n20412), .ZN(n20413) );
  NOR2_X1 U23357 ( .A1(n10492), .A2(n20625), .ZN(n20535) );
  INV_X1 U23358 ( .A(n20604), .ZN(n20659) );
  AOI211_X1 U23359 ( .C1(n20414), .C2(n20413), .A(n20535), .B(n20659), .ZN(
        n20415) );
  INV_X1 U23360 ( .A(n20437), .ZN(n20427) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20439), .B1(
        n20427), .B2(n20860), .ZN(n20416) );
  OAI211_X1 U23362 ( .C1(n20442), .C2(n20852), .A(n20417), .B(n20416), .ZN(
        P1_U3049) );
  INV_X1 U23363 ( .A(n20864), .ZN(n20737) );
  AOI22_X1 U23364 ( .A1(n20471), .A2(n20777), .B1(n20865), .B2(n20426), .ZN(
        n20419) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20439), .B1(
        n20427), .B2(n20866), .ZN(n20418) );
  OAI211_X1 U23366 ( .C1(n20442), .C2(n20737), .A(n20419), .B(n20418), .ZN(
        P1_U3050) );
  INV_X1 U23367 ( .A(n20816), .ZN(n20870) );
  INV_X1 U23368 ( .A(n20426), .ZN(n20436) );
  OAI22_X1 U23369 ( .A1(n20437), .A2(n20876), .B1(n20871), .B2(n20436), .ZN(
        n20420) );
  INV_X1 U23370 ( .A(n20420), .ZN(n20422) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20439), .B1(
        n20471), .B2(n20873), .ZN(n20421) );
  OAI211_X1 U23372 ( .C1(n20442), .C2(n20870), .A(n20422), .B(n20421), .ZN(
        P1_U3051) );
  OAI22_X1 U23373 ( .A1(n20437), .A2(n20883), .B1(n20878), .B2(n20436), .ZN(
        n20423) );
  INV_X1 U23374 ( .A(n20423), .ZN(n20425) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20439), .B1(
        n20471), .B2(n20880), .ZN(n20424) );
  OAI211_X1 U23376 ( .C1(n20442), .C2(n20877), .A(n20425), .B(n20424), .ZN(
        P1_U3052) );
  INV_X1 U23377 ( .A(n20828), .ZN(n20884) );
  AOI22_X1 U23378 ( .A1(n20471), .A2(n20889), .B1(n20829), .B2(n20426), .ZN(
        n20429) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20439), .B1(
        n20427), .B2(n20830), .ZN(n20428) );
  OAI211_X1 U23380 ( .C1(n20442), .C2(n20884), .A(n20429), .B(n20428), .ZN(
        P1_U3053) );
  OAI22_X1 U23381 ( .A1(n20437), .A2(n20897), .B1(n20436), .B2(n20747), .ZN(
        n20430) );
  INV_X1 U23382 ( .A(n20430), .ZN(n20432) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20439), .B1(
        n20471), .B2(n20894), .ZN(n20431) );
  OAI211_X1 U23384 ( .C1(n20442), .C2(n20751), .A(n20432), .B(n20431), .ZN(
        P1_U3054) );
  INV_X1 U23385 ( .A(n20898), .ZN(n20756) );
  OAI22_X1 U23386 ( .A1(n20437), .A2(n20792), .B1(n20436), .B2(n20752), .ZN(
        n20433) );
  INV_X1 U23387 ( .A(n20433), .ZN(n20435) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20439), .B1(
        n20471), .B2(n20789), .ZN(n20434) );
  OAI211_X1 U23389 ( .C1(n20442), .C2(n20756), .A(n20435), .B(n20434), .ZN(
        P1_U3055) );
  INV_X1 U23390 ( .A(n20907), .ZN(n20764) );
  OAI22_X1 U23391 ( .A1(n20437), .A2(n20916), .B1(n20758), .B2(n20436), .ZN(
        n20438) );
  INV_X1 U23392 ( .A(n20438), .ZN(n20441) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20439), .B1(
        n20471), .B2(n20910), .ZN(n20440) );
  OAI211_X1 U23394 ( .C1(n20442), .C2(n20764), .A(n20441), .B(n20440), .ZN(
        P1_U3056) );
  INV_X1 U23395 ( .A(n20455), .ZN(n20444) );
  OAI21_X1 U23396 ( .B1(n20444), .B2(n20804), .A(n20443), .ZN(n20453) );
  NAND2_X1 U23397 ( .A1(n10883), .A2(n20445), .ZN(n20561) );
  OR2_X1 U23398 ( .A1(n20446), .A2(n20561), .ZN(n20448) );
  NOR2_X1 U23399 ( .A1(n20687), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20470) );
  INV_X1 U23400 ( .A(n20470), .ZN(n20447) );
  INV_X1 U23401 ( .A(n20452), .ZN(n20449) );
  AOI22_X1 U23402 ( .A1(n20471), .A2(n20860), .B1(n20806), .B2(n20470), .ZN(
        n20457) );
  OAI21_X1 U23403 ( .B1(n20848), .B2(n20450), .A(n20858), .ZN(n20451) );
  AOI21_X1 U23404 ( .B1(n20453), .B2(n20452), .A(n20451), .ZN(n20454) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20472), .B1(
        n20501), .B2(n20773), .ZN(n20456) );
  OAI211_X1 U23406 ( .C1(n20475), .C2(n20852), .A(n20457), .B(n20456), .ZN(
        P1_U3057) );
  AOI22_X1 U23407 ( .A1(n20501), .A2(n20777), .B1(n20865), .B2(n20470), .ZN(
        n20459) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20472), .B1(
        n20471), .B2(n20866), .ZN(n20458) );
  OAI211_X1 U23409 ( .C1(n20475), .C2(n20737), .A(n20459), .B(n20458), .ZN(
        P1_U3058) );
  AOI22_X1 U23410 ( .A1(n20501), .A2(n20873), .B1(n20817), .B2(n20470), .ZN(
        n20461) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20472), .B1(
        n20471), .B2(n20818), .ZN(n20460) );
  OAI211_X1 U23412 ( .C1(n20475), .C2(n20870), .A(n20461), .B(n20460), .ZN(
        P1_U3059) );
  AOI22_X1 U23413 ( .A1(n20501), .A2(n20880), .B1(n20823), .B2(n20470), .ZN(
        n20463) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20472), .B1(
        n20471), .B2(n20824), .ZN(n20462) );
  OAI211_X1 U23415 ( .C1(n20475), .C2(n20877), .A(n20463), .B(n20462), .ZN(
        P1_U3060) );
  AOI22_X1 U23416 ( .A1(n20471), .A2(n20830), .B1(n20829), .B2(n20470), .ZN(
        n20465) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20472), .B1(
        n20501), .B2(n20889), .ZN(n20464) );
  OAI211_X1 U23418 ( .C1(n20475), .C2(n20884), .A(n20465), .B(n20464), .ZN(
        P1_U3061) );
  AOI22_X1 U23419 ( .A1(n20471), .A2(n20833), .B1(n20470), .B2(n20893), .ZN(
        n20467) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20472), .B1(
        n20501), .B2(n20894), .ZN(n20466) );
  OAI211_X1 U23421 ( .C1(n20475), .C2(n20751), .A(n20467), .B(n20466), .ZN(
        P1_U3062) );
  AOI22_X1 U23422 ( .A1(n20471), .A2(n20900), .B1(n20470), .B2(n20899), .ZN(
        n20469) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20472), .B1(
        n20501), .B2(n20789), .ZN(n20468) );
  OAI211_X1 U23424 ( .C1(n20475), .C2(n20756), .A(n20469), .B(n20468), .ZN(
        P1_U3063) );
  AOI22_X1 U23425 ( .A1(n20501), .A2(n20910), .B1(n20909), .B2(n20470), .ZN(
        n20474) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20472), .B1(
        n20471), .B2(n20841), .ZN(n20473) );
  OAI211_X1 U23427 ( .C1(n20475), .C2(n20764), .A(n20474), .B(n20473), .ZN(
        P1_U3064) );
  NAND3_X1 U23428 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20653), .A3(
        n20723), .ZN(n20506) );
  NOR2_X1 U23429 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20506), .ZN(
        n20500) );
  INV_X1 U23430 ( .A(n20722), .ZN(n20802) );
  OR2_X1 U23431 ( .A1(n20720), .A2(n20477), .ZN(n20564) );
  INV_X1 U23432 ( .A(n20564), .ZN(n20505) );
  NAND3_X1 U23433 ( .A1(n20505), .A2(n20848), .A3(n20595), .ZN(n20478) );
  OAI21_X1 U23434 ( .B1(n20802), .B2(n20479), .A(n20478), .ZN(n20499) );
  AOI22_X1 U23435 ( .A1(n20806), .A2(n20500), .B1(n20805), .B2(n20499), .ZN(
        n20486) );
  INV_X1 U23436 ( .A(n20501), .ZN(n20480) );
  AOI21_X1 U23437 ( .B1(n20480), .B2(n20529), .A(n21346), .ZN(n20481) );
  AOI21_X1 U23438 ( .B1(n20505), .B2(n20595), .A(n20481), .ZN(n20482) );
  NOR2_X1 U23439 ( .A1(n20482), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20484) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20860), .ZN(n20485) );
  OAI211_X1 U23441 ( .C1(n20863), .C2(n20529), .A(n20486), .B(n20485), .ZN(
        P1_U3065) );
  AOI22_X1 U23442 ( .A1(n20865), .A2(n20500), .B1(n20864), .B2(n20499), .ZN(
        n20488) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20866), .ZN(n20487) );
  OAI211_X1 U23444 ( .C1(n20869), .C2(n20529), .A(n20488), .B(n20487), .ZN(
        P1_U3066) );
  AOI22_X1 U23445 ( .A1(n20817), .A2(n20500), .B1(n20816), .B2(n20499), .ZN(
        n20490) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20818), .ZN(n20489) );
  OAI211_X1 U23447 ( .C1(n20821), .C2(n20529), .A(n20490), .B(n20489), .ZN(
        P1_U3067) );
  AOI22_X1 U23448 ( .A1(n20823), .A2(n20500), .B1(n20822), .B2(n20499), .ZN(
        n20492) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20824), .ZN(n20491) );
  OAI211_X1 U23450 ( .C1(n20827), .C2(n20529), .A(n20492), .B(n20491), .ZN(
        P1_U3068) );
  AOI22_X1 U23451 ( .A1(n20829), .A2(n20500), .B1(n20828), .B2(n20499), .ZN(
        n20494) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20830), .ZN(n20493) );
  OAI211_X1 U23453 ( .C1(n9977), .C2(n20529), .A(n20494), .B(n20493), .ZN(
        P1_U3069) );
  AOI22_X1 U23454 ( .A1(n20893), .A2(n20500), .B1(n20892), .B2(n20499), .ZN(
        n20496) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20833), .ZN(n20495) );
  OAI211_X1 U23456 ( .C1(n20836), .C2(n20529), .A(n20496), .B(n20495), .ZN(
        P1_U3070) );
  AOI22_X1 U23457 ( .A1(n20899), .A2(n20500), .B1(n20898), .B2(n20499), .ZN(
        n20498) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20900), .ZN(n20497) );
  OAI211_X1 U23459 ( .C1(n20905), .C2(n20529), .A(n20498), .B(n20497), .ZN(
        P1_U3071) );
  AOI22_X1 U23460 ( .A1(n20909), .A2(n20500), .B1(n20907), .B2(n20499), .ZN(
        n20504) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20841), .ZN(n20503) );
  OAI211_X1 U23462 ( .C1(n20846), .C2(n20529), .A(n20504), .B(n20503), .ZN(
        P1_U3072) );
  NOR2_X1 U23463 ( .A1(n20766), .A2(n20506), .ZN(n20525) );
  AOI21_X1 U23464 ( .B1(n20505), .B2(n20767), .A(n20525), .ZN(n20507) );
  OAI22_X1 U23465 ( .A1(n20507), .A2(n20804), .B1(n20506), .B2(n20625), .ZN(
        n20524) );
  AOI22_X1 U23466 ( .A1(n20806), .A2(n20525), .B1(n20524), .B2(n20805), .ZN(
        n20511) );
  INV_X1 U23467 ( .A(n20506), .ZN(n20509) );
  OAI21_X1 U23468 ( .B1(n20532), .B2(n21346), .A(n20507), .ZN(n20508) );
  OAI221_X1 U23469 ( .B1(n20848), .B2(n20509), .C1(n20804), .C2(n20508), .A(
        n20858), .ZN(n20526) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20773), .ZN(n20510) );
  OAI211_X1 U23471 ( .C1(n20776), .C2(n20529), .A(n20511), .B(n20510), .ZN(
        P1_U3073) );
  INV_X1 U23472 ( .A(n20866), .ZN(n20780) );
  AOI22_X1 U23473 ( .A1(n20524), .A2(n20864), .B1(n20865), .B2(n20525), .ZN(
        n20513) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20777), .ZN(n20512) );
  OAI211_X1 U23475 ( .C1(n20780), .C2(n20529), .A(n20513), .B(n20512), .ZN(
        P1_U3074) );
  AOI22_X1 U23476 ( .A1(n20817), .A2(n20525), .B1(n20524), .B2(n20816), .ZN(
        n20515) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20873), .ZN(n20514) );
  OAI211_X1 U23478 ( .C1(n20876), .C2(n20529), .A(n20515), .B(n20514), .ZN(
        P1_U3075) );
  AOI22_X1 U23479 ( .A1(n20823), .A2(n20525), .B1(n20524), .B2(n20822), .ZN(
        n20517) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20880), .ZN(n20516) );
  OAI211_X1 U23481 ( .C1(n20883), .C2(n20529), .A(n20517), .B(n20516), .ZN(
        P1_U3076) );
  AOI22_X1 U23482 ( .A1(n20829), .A2(n20525), .B1(n20524), .B2(n20828), .ZN(
        n20519) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20889), .ZN(n20518) );
  OAI211_X1 U23484 ( .C1(n9980), .C2(n20529), .A(n20519), .B(n20518), .ZN(
        P1_U3077) );
  AOI22_X1 U23485 ( .A1(n20524), .A2(n20892), .B1(n20893), .B2(n20525), .ZN(
        n20521) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20894), .ZN(n20520) );
  OAI211_X1 U23487 ( .C1(n20897), .C2(n20529), .A(n20521), .B(n20520), .ZN(
        P1_U3078) );
  AOI22_X1 U23488 ( .A1(n20899), .A2(n20525), .B1(n20524), .B2(n20898), .ZN(
        n20523) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20789), .ZN(n20522) );
  OAI211_X1 U23490 ( .C1(n20792), .C2(n20529), .A(n20523), .B(n20522), .ZN(
        P1_U3079) );
  AOI22_X1 U23491 ( .A1(n20909), .A2(n20525), .B1(n20524), .B2(n20907), .ZN(
        n20528) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20526), .B1(
        n20554), .B2(n20910), .ZN(n20527) );
  OAI211_X1 U23493 ( .C1(n20916), .C2(n20529), .A(n20528), .B(n20527), .ZN(
        P1_U3080) );
  INV_X1 U23494 ( .A(n20554), .ZN(n20530) );
  NAND2_X1 U23495 ( .A1(n20530), .A2(n20848), .ZN(n20533) );
  OAI21_X1 U23496 ( .B1(n20533), .B2(n20589), .A(n20717), .ZN(n20537) );
  NOR2_X1 U23497 ( .A1(n20564), .A2(n20595), .ZN(n20534) );
  INV_X1 U23498 ( .A(n20567), .ZN(n20562) );
  NOR2_X1 U23499 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20562), .ZN(
        n20553) );
  AOI22_X1 U23500 ( .A1(n20589), .A2(n20773), .B1(n20806), .B2(n20553), .ZN(
        n20540) );
  INV_X1 U23501 ( .A(n20534), .ZN(n20536) );
  AOI21_X1 U23502 ( .B1(n20537), .B2(n20536), .A(n20535), .ZN(n20538) );
  OAI211_X1 U23503 ( .C1(n20553), .C2(n20985), .A(n20810), .B(n20538), .ZN(
        n20555) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20860), .ZN(n20539) );
  OAI211_X1 U23505 ( .C1(n20558), .C2(n20852), .A(n20540), .B(n20539), .ZN(
        P1_U3081) );
  AOI22_X1 U23506 ( .A1(n20589), .A2(n20777), .B1(n20865), .B2(n20553), .ZN(
        n20542) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20866), .ZN(n20541) );
  OAI211_X1 U23508 ( .C1(n20558), .C2(n20737), .A(n20542), .B(n20541), .ZN(
        P1_U3082) );
  AOI22_X1 U23509 ( .A1(n20589), .A2(n20873), .B1(n20817), .B2(n20553), .ZN(
        n20544) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20818), .ZN(n20543) );
  OAI211_X1 U23511 ( .C1(n20558), .C2(n20870), .A(n20544), .B(n20543), .ZN(
        P1_U3083) );
  AOI22_X1 U23512 ( .A1(n20589), .A2(n20880), .B1(n20823), .B2(n20553), .ZN(
        n20546) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20824), .ZN(n20545) );
  OAI211_X1 U23514 ( .C1(n20558), .C2(n20877), .A(n20546), .B(n20545), .ZN(
        P1_U3084) );
  AOI22_X1 U23515 ( .A1(n20554), .A2(n20830), .B1(n20829), .B2(n20553), .ZN(
        n20548) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20555), .B1(
        n20889), .B2(n20589), .ZN(n20547) );
  OAI211_X1 U23517 ( .C1(n20558), .C2(n20884), .A(n20548), .B(n20547), .ZN(
        P1_U3085) );
  AOI22_X1 U23518 ( .A1(n20589), .A2(n20894), .B1(n20893), .B2(n20553), .ZN(
        n20550) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20833), .ZN(n20549) );
  OAI211_X1 U23520 ( .C1(n20558), .C2(n20751), .A(n20550), .B(n20549), .ZN(
        P1_U3086) );
  AOI22_X1 U23521 ( .A1(n20554), .A2(n20900), .B1(n20899), .B2(n20553), .ZN(
        n20552) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20555), .B1(
        n20589), .B2(n20789), .ZN(n20551) );
  OAI211_X1 U23523 ( .C1(n20558), .C2(n20756), .A(n20552), .B(n20551), .ZN(
        P1_U3087) );
  AOI22_X1 U23524 ( .A1(n20589), .A2(n20910), .B1(n20909), .B2(n20553), .ZN(
        n20557) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20555), .B1(
        n20554), .B2(n20841), .ZN(n20556) );
  OAI211_X1 U23526 ( .C1(n20558), .C2(n20764), .A(n20557), .B(n20556), .ZN(
        P1_U3088) );
  OR2_X1 U23527 ( .A1(n20561), .A2(n20804), .ZN(n20850) );
  INV_X1 U23528 ( .A(n20579), .ZN(n20588) );
  AOI22_X1 U23529 ( .A1(n20848), .A2(n20588), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20567), .ZN(n20563) );
  OAI21_X1 U23530 ( .B1(n20564), .B2(n20850), .A(n20563), .ZN(n20587) );
  INV_X1 U23531 ( .A(n20587), .ZN(n20578) );
  OAI22_X1 U23532 ( .A1(n20853), .A2(n20579), .B1(n20578), .B2(n20852), .ZN(
        n20565) );
  INV_X1 U23533 ( .A(n20565), .ZN(n20569) );
  OAI21_X1 U23534 ( .B1(n20567), .B2(n20566), .A(n20858), .ZN(n20590) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20860), .ZN(n20568) );
  OAI211_X1 U23536 ( .C1(n20863), .C2(n20599), .A(n20569), .B(n20568), .ZN(
        P1_U3089) );
  AOI22_X1 U23537 ( .A1(n20865), .A2(n20588), .B1(n20864), .B2(n20587), .ZN(
        n20571) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20866), .ZN(n20570) );
  OAI211_X1 U23539 ( .C1(n20869), .C2(n20599), .A(n20571), .B(n20570), .ZN(
        P1_U3090) );
  OAI22_X1 U23540 ( .A1(n20871), .A2(n20579), .B1(n20578), .B2(n20870), .ZN(
        n20572) );
  INV_X1 U23541 ( .A(n20572), .ZN(n20574) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20818), .ZN(n20573) );
  OAI211_X1 U23543 ( .C1(n20821), .C2(n20599), .A(n20574), .B(n20573), .ZN(
        P1_U3091) );
  OAI22_X1 U23544 ( .A1(n20878), .A2(n20579), .B1(n20578), .B2(n20877), .ZN(
        n20575) );
  INV_X1 U23545 ( .A(n20575), .ZN(n20577) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20824), .ZN(n20576) );
  OAI211_X1 U23547 ( .C1(n20827), .C2(n20599), .A(n20577), .B(n20576), .ZN(
        P1_U3092) );
  OAI22_X1 U23548 ( .A1(n20887), .A2(n20579), .B1(n20578), .B2(n20884), .ZN(
        n20580) );
  INV_X1 U23549 ( .A(n20580), .ZN(n20582) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20830), .ZN(n20581) );
  OAI211_X1 U23551 ( .C1(n9977), .C2(n20599), .A(n20582), .B(n20581), .ZN(
        P1_U3093) );
  AOI22_X1 U23552 ( .A1(n20893), .A2(n20588), .B1(n20892), .B2(n20587), .ZN(
        n20584) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20833), .ZN(n20583) );
  OAI211_X1 U23554 ( .C1(n20836), .C2(n20599), .A(n20584), .B(n20583), .ZN(
        P1_U3094) );
  AOI22_X1 U23555 ( .A1(n20899), .A2(n20588), .B1(n20898), .B2(n20587), .ZN(
        n20586) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20900), .ZN(n20585) );
  OAI211_X1 U23557 ( .C1(n20905), .C2(n20599), .A(n20586), .B(n20585), .ZN(
        P1_U3095) );
  AOI22_X1 U23558 ( .A1(n20909), .A2(n20588), .B1(n20907), .B2(n20587), .ZN(
        n20592) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20841), .ZN(n20591) );
  OAI211_X1 U23560 ( .C1(n20846), .C2(n20599), .A(n20592), .B(n20591), .ZN(
        P1_U3096) );
  AND2_X1 U23561 ( .A1(n20594), .A2(n20720), .ZN(n20689) );
  NAND3_X1 U23562 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11313), .A3(
        n20723), .ZN(n20626) );
  NOR2_X1 U23563 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20626), .ZN(
        n20619) );
  AOI21_X1 U23564 ( .B1(n20689), .B2(n20595), .A(n20619), .ZN(n20601) );
  INV_X1 U23565 ( .A(n20654), .ZN(n20596) );
  NOR2_X1 U23566 ( .A1(n20597), .A2(n20596), .ZN(n20721) );
  INV_X1 U23567 ( .A(n20721), .ZN(n20726) );
  OAI22_X1 U23568 ( .A1(n20601), .A2(n20804), .B1(n20598), .B2(n20726), .ZN(
        n20620) );
  AOI22_X1 U23569 ( .A1(n20620), .A2(n20805), .B1(n20806), .B2(n20619), .ZN(
        n20606) );
  INV_X1 U23570 ( .A(n20649), .ZN(n20600) );
  OAI21_X1 U23571 ( .B1(n20600), .B2(n20621), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20602) );
  NAND2_X1 U23572 ( .A1(n20602), .A2(n20601), .ZN(n20603) );
  OAI211_X1 U23573 ( .C1(n20619), .C2(n20985), .A(n20604), .B(n20603), .ZN(
        n20622) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20860), .ZN(n20605) );
  OAI211_X1 U23575 ( .C1(n20863), .C2(n20649), .A(n20606), .B(n20605), .ZN(
        P1_U3097) );
  AOI22_X1 U23576 ( .A1(n20620), .A2(n20864), .B1(n20865), .B2(n20619), .ZN(
        n20608) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20866), .ZN(n20607) );
  OAI211_X1 U23578 ( .C1(n20869), .C2(n20649), .A(n20608), .B(n20607), .ZN(
        P1_U3098) );
  AOI22_X1 U23579 ( .A1(n20620), .A2(n20816), .B1(n20817), .B2(n20619), .ZN(
        n20610) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20818), .ZN(n20609) );
  OAI211_X1 U23581 ( .C1(n20821), .C2(n20649), .A(n20610), .B(n20609), .ZN(
        P1_U3099) );
  AOI22_X1 U23582 ( .A1(n20620), .A2(n20822), .B1(n20823), .B2(n20619), .ZN(
        n20612) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20824), .ZN(n20611) );
  OAI211_X1 U23584 ( .C1(n20827), .C2(n20649), .A(n20612), .B(n20611), .ZN(
        P1_U3100) );
  AOI22_X1 U23585 ( .A1(n20620), .A2(n20828), .B1(n20829), .B2(n20619), .ZN(
        n20614) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20830), .ZN(n20613) );
  OAI211_X1 U23587 ( .C1(n9977), .C2(n20649), .A(n20614), .B(n20613), .ZN(
        P1_U3101) );
  AOI22_X1 U23588 ( .A1(n20620), .A2(n20892), .B1(n20893), .B2(n20619), .ZN(
        n20616) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20833), .ZN(n20615) );
  OAI211_X1 U23590 ( .C1(n20836), .C2(n20649), .A(n20616), .B(n20615), .ZN(
        P1_U3102) );
  AOI22_X1 U23591 ( .A1(n20620), .A2(n20898), .B1(n20899), .B2(n20619), .ZN(
        n20618) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20900), .ZN(n20617) );
  OAI211_X1 U23593 ( .C1(n20905), .C2(n20649), .A(n20618), .B(n20617), .ZN(
        P1_U3103) );
  AOI22_X1 U23594 ( .A1(n20620), .A2(n20907), .B1(n20909), .B2(n20619), .ZN(
        n20624) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20841), .ZN(n20623) );
  OAI211_X1 U23596 ( .C1(n20846), .C2(n20649), .A(n20624), .B(n20623), .ZN(
        P1_U3104) );
  NOR2_X1 U23597 ( .A1(n20766), .A2(n20626), .ZN(n20644) );
  AOI21_X1 U23598 ( .B1(n20689), .B2(n20767), .A(n20644), .ZN(n20627) );
  OAI22_X1 U23599 ( .A1(n20627), .A2(n20804), .B1(n20626), .B2(n20625), .ZN(
        n20645) );
  AOI22_X1 U23600 ( .A1(n20645), .A2(n20805), .B1(n20806), .B2(n20644), .ZN(
        n20631) );
  INV_X1 U23601 ( .A(n20626), .ZN(n20629) );
  OAI21_X1 U23602 ( .B1(n20695), .B2(n21346), .A(n20627), .ZN(n20628) );
  OAI221_X1 U23603 ( .B1(n20848), .B2(n20629), .C1(n20804), .C2(n20628), .A(
        n20858), .ZN(n20646) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20773), .ZN(n20630) );
  OAI211_X1 U23605 ( .C1(n20776), .C2(n20649), .A(n20631), .B(n20630), .ZN(
        P1_U3105) );
  AOI22_X1 U23606 ( .A1(n20645), .A2(n20864), .B1(n20865), .B2(n20644), .ZN(
        n20633) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20777), .ZN(n20632) );
  OAI211_X1 U23608 ( .C1(n20780), .C2(n20649), .A(n20633), .B(n20632), .ZN(
        P1_U3106) );
  AOI22_X1 U23609 ( .A1(n20645), .A2(n20816), .B1(n20817), .B2(n20644), .ZN(
        n20635) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20873), .ZN(n20634) );
  OAI211_X1 U23611 ( .C1(n20876), .C2(n20649), .A(n20635), .B(n20634), .ZN(
        P1_U3107) );
  AOI22_X1 U23612 ( .A1(n20645), .A2(n20822), .B1(n20823), .B2(n20644), .ZN(
        n20637) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20880), .ZN(n20636) );
  OAI211_X1 U23614 ( .C1(n20883), .C2(n20649), .A(n20637), .B(n20636), .ZN(
        P1_U3108) );
  AOI22_X1 U23615 ( .A1(n20645), .A2(n20828), .B1(n20829), .B2(n20644), .ZN(
        n20639) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20889), .ZN(n20638) );
  OAI211_X1 U23617 ( .C1(n9980), .C2(n20649), .A(n20639), .B(n20638), .ZN(
        P1_U3109) );
  AOI22_X1 U23618 ( .A1(n20645), .A2(n20892), .B1(n20893), .B2(n20644), .ZN(
        n20641) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20894), .ZN(n20640) );
  OAI211_X1 U23620 ( .C1(n20897), .C2(n20649), .A(n20641), .B(n20640), .ZN(
        P1_U3110) );
  AOI22_X1 U23621 ( .A1(n20645), .A2(n20898), .B1(n20899), .B2(n20644), .ZN(
        n20643) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20789), .ZN(n20642) );
  OAI211_X1 U23623 ( .C1(n20792), .C2(n20649), .A(n20643), .B(n20642), .ZN(
        P1_U3111) );
  AOI22_X1 U23624 ( .A1(n20645), .A2(n20907), .B1(n20909), .B2(n20644), .ZN(
        n20648) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20646), .B1(
        n20681), .B2(n20910), .ZN(n20647) );
  OAI211_X1 U23626 ( .C1(n20916), .C2(n20649), .A(n20648), .B(n20647), .ZN(
        P1_U3112) );
  INV_X1 U23627 ( .A(n20681), .ZN(n20651) );
  NAND3_X1 U23628 ( .A1(n20651), .A2(n20848), .A3(n20715), .ZN(n20652) );
  NAND2_X1 U23629 ( .A1(n20652), .A2(n20717), .ZN(n20661) );
  AND2_X1 U23630 ( .A1(n20689), .A2(n10856), .ZN(n20657) );
  OR2_X1 U23631 ( .A1(n20654), .A2(n20653), .ZN(n20803) );
  INV_X1 U23632 ( .A(n20803), .ZN(n20655) );
  NAND3_X1 U23633 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n11313), .ZN(n20692) );
  NOR2_X1 U23634 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20692), .ZN(
        n20680) );
  AOI22_X1 U23635 ( .A1(n20681), .A2(n20860), .B1(n20806), .B2(n20680), .ZN(
        n20664) );
  INV_X1 U23636 ( .A(n20657), .ZN(n20660) );
  NAND2_X1 U23637 ( .A1(n20803), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20809) );
  INV_X1 U23638 ( .A(n20809), .ZN(n20658) );
  AOI211_X1 U23639 ( .C1(n20661), .C2(n20660), .A(n20659), .B(n20658), .ZN(
        n20662) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20773), .ZN(n20663) );
  OAI211_X1 U23641 ( .C1(n20686), .C2(n20852), .A(n20664), .B(n20663), .ZN(
        P1_U3113) );
  AOI22_X1 U23642 ( .A1(n20681), .A2(n20866), .B1(n20865), .B2(n20680), .ZN(
        n20666) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20777), .ZN(n20665) );
  OAI211_X1 U23644 ( .C1(n20686), .C2(n20737), .A(n20666), .B(n20665), .ZN(
        P1_U3114) );
  INV_X1 U23645 ( .A(n20680), .ZN(n20676) );
  OAI22_X1 U23646 ( .A1(n20715), .A2(n20821), .B1(n20871), .B2(n20676), .ZN(
        n20667) );
  INV_X1 U23647 ( .A(n20667), .ZN(n20669) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20683), .B1(
        n20681), .B2(n20818), .ZN(n20668) );
  OAI211_X1 U23649 ( .C1(n20686), .C2(n20870), .A(n20669), .B(n20668), .ZN(
        P1_U3115) );
  AOI22_X1 U23650 ( .A1(n20681), .A2(n20824), .B1(n20823), .B2(n20680), .ZN(
        n20671) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20880), .ZN(n20670) );
  OAI211_X1 U23652 ( .C1(n20686), .C2(n20877), .A(n20671), .B(n20670), .ZN(
        P1_U3116) );
  AOI22_X1 U23653 ( .A1(n20681), .A2(n20830), .B1(n20829), .B2(n20680), .ZN(
        n20673) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20889), .ZN(n20672) );
  OAI211_X1 U23655 ( .C1(n20686), .C2(n20884), .A(n20673), .B(n20672), .ZN(
        P1_U3117) );
  AOI22_X1 U23656 ( .A1(n20681), .A2(n20833), .B1(n20893), .B2(n20680), .ZN(
        n20675) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20894), .ZN(n20674) );
  OAI211_X1 U23658 ( .C1(n20686), .C2(n20751), .A(n20675), .B(n20674), .ZN(
        P1_U3118) );
  OAI22_X1 U23659 ( .A1(n20715), .A2(n20905), .B1(n20752), .B2(n20676), .ZN(
        n20677) );
  INV_X1 U23660 ( .A(n20677), .ZN(n20679) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20683), .B1(
        n20681), .B2(n20900), .ZN(n20678) );
  OAI211_X1 U23662 ( .C1(n20686), .C2(n20756), .A(n20679), .B(n20678), .ZN(
        P1_U3119) );
  AOI22_X1 U23663 ( .A1(n20681), .A2(n20841), .B1(n20909), .B2(n20680), .ZN(
        n20685) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20910), .ZN(n20684) );
  OAI211_X1 U23665 ( .C1(n20686), .C2(n20764), .A(n20685), .B(n20684), .ZN(
        P1_U3120) );
  INV_X1 U23666 ( .A(n20687), .ZN(n20688) );
  NAND2_X1 U23667 ( .A1(n20688), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20690) );
  INV_X1 U23668 ( .A(n20690), .ZN(n20711) );
  INV_X1 U23669 ( .A(n20689), .ZN(n20691) );
  OAI222_X1 U23670 ( .A1(n20850), .A2(n20691), .B1(n20625), .B2(n20692), .C1(
        n20804), .C2(n20690), .ZN(n20710) );
  AOI22_X1 U23671 ( .A1(n20806), .A2(n20711), .B1(n20710), .B2(n20805), .ZN(
        n20697) );
  OAI21_X1 U23672 ( .B1(n20695), .B2(n20856), .A(n20692), .ZN(n20693) );
  NAND2_X1 U23673 ( .A1(n20693), .A2(n20858), .ZN(n20712) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20773), .ZN(n20696) );
  OAI211_X1 U23675 ( .C1(n20776), .C2(n20715), .A(n20697), .B(n20696), .ZN(
        P1_U3121) );
  AOI22_X1 U23676 ( .A1(n20710), .A2(n20864), .B1(n20865), .B2(n20711), .ZN(
        n20699) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20777), .ZN(n20698) );
  OAI211_X1 U23678 ( .C1(n20780), .C2(n20715), .A(n20699), .B(n20698), .ZN(
        P1_U3122) );
  AOI22_X1 U23679 ( .A1(n20817), .A2(n20711), .B1(n20710), .B2(n20816), .ZN(
        n20701) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20873), .ZN(n20700) );
  OAI211_X1 U23681 ( .C1(n20876), .C2(n20715), .A(n20701), .B(n20700), .ZN(
        P1_U3123) );
  AOI22_X1 U23682 ( .A1(n20823), .A2(n20711), .B1(n20710), .B2(n20822), .ZN(
        n20703) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20880), .ZN(n20702) );
  OAI211_X1 U23684 ( .C1(n20883), .C2(n20715), .A(n20703), .B(n20702), .ZN(
        P1_U3124) );
  AOI22_X1 U23685 ( .A1(n20829), .A2(n20711), .B1(n20710), .B2(n20828), .ZN(
        n20705) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20889), .ZN(n20704) );
  OAI211_X1 U23687 ( .C1(n9980), .C2(n20715), .A(n20705), .B(n20704), .ZN(
        P1_U3125) );
  AOI22_X1 U23688 ( .A1(n20710), .A2(n20892), .B1(n20893), .B2(n20711), .ZN(
        n20707) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20894), .ZN(n20706) );
  OAI211_X1 U23690 ( .C1(n20897), .C2(n20715), .A(n20707), .B(n20706), .ZN(
        P1_U3126) );
  AOI22_X1 U23691 ( .A1(n20899), .A2(n20711), .B1(n20710), .B2(n20898), .ZN(
        n20709) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20789), .ZN(n20708) );
  OAI211_X1 U23693 ( .C1(n20792), .C2(n20715), .A(n20709), .B(n20708), .ZN(
        P1_U3127) );
  AOI22_X1 U23694 ( .A1(n20909), .A2(n20711), .B1(n20710), .B2(n20907), .ZN(
        n20714) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20712), .B1(
        n20760), .B2(n20910), .ZN(n20713) );
  OAI211_X1 U23696 ( .C1(n20916), .C2(n20715), .A(n20714), .B(n20713), .ZN(
        P1_U3128) );
  NAND2_X1 U23697 ( .A1(n20798), .A2(n20848), .ZN(n20718) );
  OAI21_X1 U23698 ( .B1(n20760), .B2(n20718), .A(n20717), .ZN(n20728) );
  OR2_X1 U23699 ( .A1(n20720), .A2(n20719), .ZN(n20851) );
  NOR2_X1 U23700 ( .A1(n20851), .A2(n10856), .ZN(n20725) );
  NAND3_X1 U23701 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20723), .ZN(n20768) );
  NOR2_X1 U23702 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20768), .ZN(
        n20730) );
  INV_X1 U23703 ( .A(n20730), .ZN(n20757) );
  OAI22_X1 U23704 ( .A1(n20798), .A2(n20863), .B1(n20853), .B2(n20757), .ZN(
        n20724) );
  INV_X1 U23705 ( .A(n20724), .ZN(n20732) );
  INV_X1 U23706 ( .A(n20725), .ZN(n20727) );
  AOI22_X1 U23707 ( .A1(n20728), .A2(n20727), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20726), .ZN(n20729) );
  OAI211_X1 U23708 ( .C1(n20730), .C2(n20985), .A(n20810), .B(n20729), .ZN(
        n20761) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20860), .ZN(n20731) );
  OAI211_X1 U23710 ( .C1(n20765), .C2(n20852), .A(n20732), .B(n20731), .ZN(
        P1_U3129) );
  INV_X1 U23711 ( .A(n20865), .ZN(n20733) );
  OAI22_X1 U23712 ( .A1(n20798), .A2(n20869), .B1(n20733), .B2(n20757), .ZN(
        n20734) );
  INV_X1 U23713 ( .A(n20734), .ZN(n20736) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20866), .ZN(n20735) );
  OAI211_X1 U23715 ( .C1(n20765), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P1_U3130) );
  OAI22_X1 U23716 ( .A1(n20798), .A2(n20821), .B1(n20871), .B2(n20757), .ZN(
        n20738) );
  INV_X1 U23717 ( .A(n20738), .ZN(n20740) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20818), .ZN(n20739) );
  OAI211_X1 U23719 ( .C1(n20765), .C2(n20870), .A(n20740), .B(n20739), .ZN(
        P1_U3131) );
  OAI22_X1 U23720 ( .A1(n20798), .A2(n20827), .B1(n20878), .B2(n20757), .ZN(
        n20741) );
  INV_X1 U23721 ( .A(n20741), .ZN(n20743) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20824), .ZN(n20742) );
  OAI211_X1 U23723 ( .C1(n20765), .C2(n20877), .A(n20743), .B(n20742), .ZN(
        P1_U3132) );
  OAI22_X1 U23724 ( .A1(n20798), .A2(n9977), .B1(n20887), .B2(n20757), .ZN(
        n20744) );
  INV_X1 U23725 ( .A(n20744), .ZN(n20746) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20830), .ZN(n20745) );
  OAI211_X1 U23727 ( .C1(n20765), .C2(n20884), .A(n20746), .B(n20745), .ZN(
        P1_U3133) );
  OAI22_X1 U23728 ( .A1(n20798), .A2(n20836), .B1(n20747), .B2(n20757), .ZN(
        n20748) );
  INV_X1 U23729 ( .A(n20748), .ZN(n20750) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20833), .ZN(n20749) );
  OAI211_X1 U23731 ( .C1(n20765), .C2(n20751), .A(n20750), .B(n20749), .ZN(
        P1_U3134) );
  OAI22_X1 U23732 ( .A1(n20798), .A2(n20905), .B1(n20752), .B2(n20757), .ZN(
        n20753) );
  INV_X1 U23733 ( .A(n20753), .ZN(n20755) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20900), .ZN(n20754) );
  OAI211_X1 U23735 ( .C1(n20765), .C2(n20756), .A(n20755), .B(n20754), .ZN(
        P1_U3135) );
  OAI22_X1 U23736 ( .A1(n20798), .A2(n20846), .B1(n20758), .B2(n20757), .ZN(
        n20759) );
  INV_X1 U23737 ( .A(n20759), .ZN(n20763) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20761), .B1(
        n20760), .B2(n20841), .ZN(n20762) );
  OAI211_X1 U23739 ( .C1(n20765), .C2(n20764), .A(n20763), .B(n20762), .ZN(
        P1_U3136) );
  NOR2_X1 U23740 ( .A1(n20766), .A2(n20768), .ZN(n20794) );
  INV_X1 U23741 ( .A(n20851), .ZN(n20801) );
  AOI21_X1 U23742 ( .B1(n20801), .B2(n20767), .A(n20794), .ZN(n20769) );
  OAI22_X1 U23743 ( .A1(n20769), .A2(n20804), .B1(n20768), .B2(n20625), .ZN(
        n20793) );
  AOI22_X1 U23744 ( .A1(n20806), .A2(n20794), .B1(n20793), .B2(n20805), .ZN(
        n20775) );
  INV_X1 U23745 ( .A(n20768), .ZN(n20771) );
  OAI21_X1 U23746 ( .B1(n20857), .B2(n21346), .A(n20769), .ZN(n20770) );
  OAI221_X1 U23747 ( .B1(n20848), .B2(n20771), .C1(n20804), .C2(n20770), .A(
        n20858), .ZN(n20795) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20773), .ZN(n20774) );
  OAI211_X1 U23749 ( .C1(n20776), .C2(n20798), .A(n20775), .B(n20774), .ZN(
        P1_U3137) );
  AOI22_X1 U23750 ( .A1(n20793), .A2(n20864), .B1(n20865), .B2(n20794), .ZN(
        n20779) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20777), .ZN(n20778) );
  OAI211_X1 U23752 ( .C1(n20780), .C2(n20798), .A(n20779), .B(n20778), .ZN(
        P1_U3138) );
  AOI22_X1 U23753 ( .A1(n20817), .A2(n20794), .B1(n20793), .B2(n20816), .ZN(
        n20782) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20873), .ZN(n20781) );
  OAI211_X1 U23755 ( .C1(n20876), .C2(n20798), .A(n20782), .B(n20781), .ZN(
        P1_U3139) );
  AOI22_X1 U23756 ( .A1(n20823), .A2(n20794), .B1(n20793), .B2(n20822), .ZN(
        n20784) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20880), .ZN(n20783) );
  OAI211_X1 U23758 ( .C1(n20883), .C2(n20798), .A(n20784), .B(n20783), .ZN(
        P1_U3140) );
  AOI22_X1 U23759 ( .A1(n20829), .A2(n20794), .B1(n20793), .B2(n20828), .ZN(
        n20786) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20889), .ZN(n20785) );
  OAI211_X1 U23761 ( .C1(n9980), .C2(n20798), .A(n20786), .B(n20785), .ZN(
        P1_U3141) );
  AOI22_X1 U23762 ( .A1(n20793), .A2(n20892), .B1(n20893), .B2(n20794), .ZN(
        n20788) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20894), .ZN(n20787) );
  OAI211_X1 U23764 ( .C1(n20897), .C2(n20798), .A(n20788), .B(n20787), .ZN(
        P1_U3142) );
  AOI22_X1 U23765 ( .A1(n20899), .A2(n20794), .B1(n20793), .B2(n20898), .ZN(
        n20791) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20789), .ZN(n20790) );
  OAI211_X1 U23767 ( .C1(n20792), .C2(n20798), .A(n20791), .B(n20790), .ZN(
        P1_U3143) );
  AOI22_X1 U23768 ( .A1(n20909), .A2(n20794), .B1(n20793), .B2(n20907), .ZN(
        n20797) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20795), .B1(
        n20842), .B2(n20910), .ZN(n20796) );
  OAI211_X1 U23770 ( .C1(n20916), .C2(n20798), .A(n20797), .B(n20796), .ZN(
        P1_U3144) );
  NOR2_X1 U23771 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20855), .ZN(
        n20840) );
  NAND2_X1 U23772 ( .A1(n20801), .A2(n10856), .ZN(n20807) );
  OAI22_X1 U23773 ( .A1(n20807), .A2(n20804), .B1(n20803), .B2(n20802), .ZN(
        n20839) );
  AOI22_X1 U23774 ( .A1(n20806), .A2(n20840), .B1(n20805), .B2(n20839), .ZN(
        n20813) );
  INV_X1 U23775 ( .A(n20915), .ZN(n20901) );
  OAI21_X1 U23776 ( .B1(n20901), .B2(n20842), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20808) );
  AOI21_X1 U23777 ( .B1(n20808), .B2(n20807), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20811) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20860), .ZN(n20812) );
  OAI211_X1 U23779 ( .C1(n20863), .C2(n20915), .A(n20813), .B(n20812), .ZN(
        P1_U3145) );
  AOI22_X1 U23780 ( .A1(n20865), .A2(n20840), .B1(n20839), .B2(n20864), .ZN(
        n20815) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20866), .ZN(n20814) );
  OAI211_X1 U23782 ( .C1(n20869), .C2(n20915), .A(n20815), .B(n20814), .ZN(
        P1_U3146) );
  AOI22_X1 U23783 ( .A1(n20817), .A2(n20840), .B1(n20816), .B2(n20839), .ZN(
        n20820) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20818), .ZN(n20819) );
  OAI211_X1 U23785 ( .C1(n20821), .C2(n20915), .A(n20820), .B(n20819), .ZN(
        P1_U3147) );
  AOI22_X1 U23786 ( .A1(n20823), .A2(n20840), .B1(n20822), .B2(n20839), .ZN(
        n20826) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20824), .ZN(n20825) );
  OAI211_X1 U23788 ( .C1(n20827), .C2(n20915), .A(n20826), .B(n20825), .ZN(
        P1_U3148) );
  AOI22_X1 U23789 ( .A1(n20829), .A2(n20840), .B1(n20828), .B2(n20839), .ZN(
        n20832) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20830), .ZN(n20831) );
  OAI211_X1 U23791 ( .C1(n9977), .C2(n20915), .A(n20832), .B(n20831), .ZN(
        P1_U3149) );
  AOI22_X1 U23792 ( .A1(n20893), .A2(n20840), .B1(n20839), .B2(n20892), .ZN(
        n20835) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20833), .ZN(n20834) );
  OAI211_X1 U23794 ( .C1(n20836), .C2(n20915), .A(n20835), .B(n20834), .ZN(
        P1_U3150) );
  AOI22_X1 U23795 ( .A1(n20899), .A2(n20840), .B1(n20898), .B2(n20839), .ZN(
        n20838) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20900), .ZN(n20837) );
  OAI211_X1 U23797 ( .C1(n20905), .C2(n20915), .A(n20838), .B(n20837), .ZN(
        P1_U3151) );
  AOI22_X1 U23798 ( .A1(n20909), .A2(n20840), .B1(n20907), .B2(n20839), .ZN(
        n20845) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20841), .ZN(n20844) );
  OAI211_X1 U23800 ( .C1(n20846), .C2(n20915), .A(n20845), .B(n20844), .ZN(
        P1_U3152) );
  INV_X1 U23801 ( .A(n20886), .ZN(n20908) );
  AOI22_X1 U23802 ( .A1(n20848), .A2(n20908), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20847), .ZN(n20849) );
  OAI21_X1 U23803 ( .B1(n20851), .B2(n20850), .A(n20849), .ZN(n20906) );
  INV_X1 U23804 ( .A(n20906), .ZN(n20885) );
  OAI22_X1 U23805 ( .A1(n20853), .A2(n20886), .B1(n20885), .B2(n20852), .ZN(
        n20854) );
  INV_X1 U23806 ( .A(n20854), .ZN(n20862) );
  OAI21_X1 U23807 ( .B1(n20857), .B2(n20856), .A(n20855), .ZN(n20859) );
  NAND2_X1 U23808 ( .A1(n20859), .A2(n20858), .ZN(n20912) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20912), .B1(
        n20901), .B2(n20860), .ZN(n20861) );
  OAI211_X1 U23810 ( .C1(n20863), .C2(n20904), .A(n20862), .B(n20861), .ZN(
        P1_U3153) );
  AOI22_X1 U23811 ( .A1(n20865), .A2(n20908), .B1(n20864), .B2(n20906), .ZN(
        n20868) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20912), .B1(
        n20901), .B2(n20866), .ZN(n20867) );
  OAI211_X1 U23813 ( .C1(n20869), .C2(n20904), .A(n20868), .B(n20867), .ZN(
        P1_U3154) );
  OAI22_X1 U23814 ( .A1(n20871), .A2(n20886), .B1(n20885), .B2(n20870), .ZN(
        n20872) );
  INV_X1 U23815 ( .A(n20872), .ZN(n20875) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20912), .B1(
        n20911), .B2(n20873), .ZN(n20874) );
  OAI211_X1 U23817 ( .C1(n20876), .C2(n20915), .A(n20875), .B(n20874), .ZN(
        P1_U3155) );
  OAI22_X1 U23818 ( .A1(n20878), .A2(n20886), .B1(n20885), .B2(n20877), .ZN(
        n20879) );
  INV_X1 U23819 ( .A(n20879), .ZN(n20882) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20912), .B1(
        n20911), .B2(n20880), .ZN(n20881) );
  OAI211_X1 U23821 ( .C1(n20883), .C2(n20915), .A(n20882), .B(n20881), .ZN(
        P1_U3156) );
  OAI22_X1 U23822 ( .A1(n20887), .A2(n20886), .B1(n20885), .B2(n20884), .ZN(
        n20888) );
  INV_X1 U23823 ( .A(n20888), .ZN(n20891) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20912), .B1(
        n20911), .B2(n20889), .ZN(n20890) );
  OAI211_X1 U23825 ( .C1(n9980), .C2(n20915), .A(n20891), .B(n20890), .ZN(
        P1_U3157) );
  AOI22_X1 U23826 ( .A1(n20893), .A2(n20908), .B1(n20892), .B2(n20906), .ZN(
        n20896) );
  AOI22_X1 U23827 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20912), .B1(
        n20911), .B2(n20894), .ZN(n20895) );
  OAI211_X1 U23828 ( .C1(n20897), .C2(n20915), .A(n20896), .B(n20895), .ZN(
        P1_U3158) );
  AOI22_X1 U23829 ( .A1(n20899), .A2(n20908), .B1(n20898), .B2(n20906), .ZN(
        n20903) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20912), .B1(
        n20901), .B2(n20900), .ZN(n20902) );
  OAI211_X1 U23831 ( .C1(n20905), .C2(n20904), .A(n20903), .B(n20902), .ZN(
        P1_U3159) );
  AOI22_X1 U23832 ( .A1(n20909), .A2(n20908), .B1(n20907), .B2(n20906), .ZN(
        n20914) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20912), .B1(
        n20911), .B2(n20910), .ZN(n20913) );
  OAI211_X1 U23834 ( .C1(n20916), .C2(n20915), .A(n20914), .B(n20913), .ZN(
        P1_U3160) );
  OAI221_X1 U23835 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20919), .C1(n20625), 
        .C2(n20918), .A(n20917), .ZN(P1_U3163) );
  AND2_X1 U23836 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20980), .ZN(
        P1_U3164) );
  AND2_X1 U23837 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20980), .ZN(
        P1_U3165) );
  AND2_X1 U23838 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20980), .ZN(
        P1_U3166) );
  AND2_X1 U23839 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20980), .ZN(
        P1_U3167) );
  AND2_X1 U23840 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20980), .ZN(
        P1_U3168) );
  AND2_X1 U23841 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20980), .ZN(
        P1_U3169) );
  AND2_X1 U23842 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20980), .ZN(
        P1_U3170) );
  AND2_X1 U23843 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20980), .ZN(
        P1_U3171) );
  AND2_X1 U23844 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20980), .ZN(
        P1_U3172) );
  AND2_X1 U23845 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20980), .ZN(
        P1_U3173) );
  AND2_X1 U23846 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20980), .ZN(
        P1_U3174) );
  AND2_X1 U23847 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20980), .ZN(
        P1_U3175) );
  AND2_X1 U23848 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20980), .ZN(
        P1_U3176) );
  AND2_X1 U23849 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20980), .ZN(
        P1_U3177) );
  AND2_X1 U23850 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20980), .ZN(
        P1_U3178) );
  AND2_X1 U23851 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20980), .ZN(
        P1_U3179) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20980), .ZN(
        P1_U3180) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20980), .ZN(
        P1_U3181) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20980), .ZN(
        P1_U3182) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20980), .ZN(
        P1_U3183) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20980), .ZN(
        P1_U3184) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20980), .ZN(
        P1_U3185) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20980), .ZN(P1_U3186) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20980), .ZN(P1_U3187) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20980), .ZN(P1_U3188) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20980), .ZN(P1_U3189) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20980), .ZN(P1_U3190) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20980), .ZN(P1_U3191) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20980), .ZN(P1_U3192) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20980), .ZN(P1_U3193) );
  AOI21_X1 U23866 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21005), .A(n20920), 
        .ZN(n20929) );
  NOR2_X1 U23867 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20921) );
  OAI22_X1 U23868 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21117), .B1(n20921), 
        .B2(n21254), .ZN(n20922) );
  NOR2_X1 U23869 ( .A1(n21022), .A2(n20922), .ZN(n20923) );
  OAI22_X1 U23870 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20929), .B1(n20972), 
        .B2(n20923), .ZN(P1_U3194) );
  AOI21_X1 U23871 ( .B1(n21005), .B2(n21117), .A(n20924), .ZN(n20931) );
  OAI211_X1 U23872 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21022), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20930) );
  INV_X1 U23873 ( .A(n20925), .ZN(n20926) );
  AOI221_X1 U23874 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21117), .C1(n20927), 
        .C2(n21117), .A(n20926), .ZN(n20928) );
  OAI22_X1 U23875 ( .A1(n20931), .A2(n20930), .B1(n20929), .B2(n20928), .ZN(
        P1_U3196) );
  INV_X2 U23876 ( .A(n20951), .ZN(n20974) );
  INV_X1 U23877 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20933) );
  AND2_X1 U23878 ( .A1(n20972), .A2(n20932), .ZN(n20949) );
  INV_X2 U23879 ( .A(n20949), .ZN(n20970) );
  OAI222_X1 U23880 ( .A1(n20974), .A2(n21352), .B1(n20933), .B2(n20972), .C1(
        n20935), .C2(n20970), .ZN(P1_U3197) );
  INV_X1 U23881 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20934) );
  OAI222_X1 U23882 ( .A1(n20974), .A2(n20935), .B1(n20934), .B2(n20972), .C1(
        n21187), .C2(n20970), .ZN(P1_U3198) );
  OAI222_X1 U23883 ( .A1(n20970), .A2(n21375), .B1(n20936), .B2(n20972), .C1(
        n21187), .C2(n20974), .ZN(P1_U3199) );
  INV_X1 U23884 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20937) );
  OAI222_X1 U23885 ( .A1(n20974), .A2(n21375), .B1(n20937), .B2(n20972), .C1(
        n21368), .C2(n20970), .ZN(P1_U3200) );
  INV_X1 U23886 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20938) );
  OAI222_X1 U23887 ( .A1(n20974), .A2(n21368), .B1(n20938), .B2(n20972), .C1(
        n13564), .C2(n20970), .ZN(P1_U3201) );
  INV_X1 U23888 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20939) );
  OAI222_X1 U23889 ( .A1(n20974), .A2(n13564), .B1(n20939), .B2(n20972), .C1(
        n20941), .C2(n20970), .ZN(P1_U3202) );
  INV_X1 U23890 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20940) );
  INV_X1 U23891 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21226) );
  OAI222_X1 U23892 ( .A1(n20974), .A2(n20941), .B1(n20940), .B2(n20972), .C1(
        n21226), .C2(n20970), .ZN(P1_U3203) );
  INV_X1 U23893 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20942) );
  OAI222_X1 U23894 ( .A1(n20970), .A2(n21219), .B1(n20942), .B2(n20972), .C1(
        n21226), .C2(n20974), .ZN(P1_U3204) );
  INV_X1 U23895 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20943) );
  OAI222_X1 U23896 ( .A1(n20970), .A2(n21364), .B1(n20943), .B2(n20972), .C1(
        n21219), .C2(n20974), .ZN(P1_U3205) );
  INV_X1 U23897 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20944) );
  OAI222_X1 U23898 ( .A1(n20974), .A2(n21364), .B1(n20944), .B2(n20972), .C1(
        n20946), .C2(n20970), .ZN(P1_U3206) );
  INV_X1 U23899 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20945) );
  OAI222_X1 U23900 ( .A1(n20974), .A2(n20946), .B1(n20945), .B2(n20972), .C1(
        n21376), .C2(n20970), .ZN(P1_U3207) );
  INV_X1 U23901 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20947) );
  OAI222_X1 U23902 ( .A1(n20970), .A2(n21363), .B1(n20947), .B2(n20972), .C1(
        n21376), .C2(n20974), .ZN(P1_U3208) );
  INV_X1 U23903 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20948) );
  INV_X1 U23904 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21126) );
  OAI222_X1 U23905 ( .A1(n20974), .A2(n21363), .B1(n20948), .B2(n20972), .C1(
        n21126), .C2(n20970), .ZN(P1_U3209) );
  AOI22_X1 U23906 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21023), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20949), .ZN(n20950) );
  OAI21_X1 U23907 ( .B1(n21126), .B2(n20974), .A(n20950), .ZN(P1_U3210) );
  AOI22_X1 U23908 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21023), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20951), .ZN(n20952) );
  OAI21_X1 U23909 ( .B1(n14637), .B2(n20970), .A(n20952), .ZN(P1_U3211) );
  INV_X1 U23910 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20953) );
  INV_X1 U23911 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21119) );
  OAI222_X1 U23912 ( .A1(n20974), .A2(n14637), .B1(n20953), .B2(n20972), .C1(
        n21119), .C2(n20970), .ZN(P1_U3212) );
  INV_X1 U23913 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20954) );
  OAI222_X1 U23914 ( .A1(n20974), .A2(n21119), .B1(n20954), .B2(n20972), .C1(
        n21128), .C2(n20970), .ZN(P1_U3213) );
  INV_X1 U23915 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21366) );
  INV_X1 U23916 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20955) );
  OAI222_X1 U23917 ( .A1(n20970), .A2(n21366), .B1(n20955), .B2(n20972), .C1(
        n21128), .C2(n20974), .ZN(P1_U3214) );
  INV_X1 U23918 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20956) );
  OAI222_X1 U23919 ( .A1(n20974), .A2(n21366), .B1(n20956), .B2(n20972), .C1(
        n21246), .C2(n20970), .ZN(P1_U3215) );
  INV_X1 U23920 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20957) );
  OAI222_X1 U23921 ( .A1(n20970), .A2(n21273), .B1(n20957), .B2(n20972), .C1(
        n21246), .C2(n20974), .ZN(P1_U3216) );
  INV_X1 U23922 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20958) );
  INV_X1 U23923 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20960) );
  OAI222_X1 U23924 ( .A1(n20974), .A2(n21273), .B1(n20958), .B2(n20972), .C1(
        n20960), .C2(n20970), .ZN(P1_U3217) );
  INV_X1 U23925 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20959) );
  INV_X1 U23926 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21355) );
  OAI222_X1 U23927 ( .A1(n20974), .A2(n20960), .B1(n20959), .B2(n20972), .C1(
        n21355), .C2(n20970), .ZN(P1_U3218) );
  INV_X1 U23928 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20961) );
  OAI222_X1 U23929 ( .A1(n20974), .A2(n21355), .B1(n20961), .B2(n20972), .C1(
        n20962), .C2(n20970), .ZN(P1_U3219) );
  INV_X1 U23930 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20963) );
  OAI222_X1 U23931 ( .A1(n20970), .A2(n21120), .B1(n20963), .B2(n20972), .C1(
        n20962), .C2(n20974), .ZN(P1_U3220) );
  INV_X1 U23932 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20965) );
  INV_X1 U23933 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20964) );
  OAI222_X1 U23934 ( .A1(n20970), .A2(n20965), .B1(n20964), .B2(n20972), .C1(
        n21120), .C2(n20974), .ZN(P1_U3221) );
  INV_X1 U23935 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20966) );
  OAI222_X1 U23936 ( .A1(n20970), .A2(n21384), .B1(n20966), .B2(n20972), .C1(
        n20965), .C2(n20974), .ZN(P1_U3222) );
  INV_X1 U23937 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20967) );
  OAI222_X1 U23938 ( .A1(n20974), .A2(n21384), .B1(n20967), .B2(n20972), .C1(
        n21220), .C2(n20970), .ZN(P1_U3223) );
  INV_X1 U23939 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20968) );
  OAI222_X1 U23940 ( .A1(n20974), .A2(n21220), .B1(n20968), .B2(n20972), .C1(
        n21249), .C2(n20970), .ZN(P1_U3224) );
  INV_X1 U23941 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20969) );
  OAI222_X1 U23942 ( .A1(n20974), .A2(n21249), .B1(n20969), .B2(n20972), .C1(
        n21178), .C2(n20970), .ZN(P1_U3225) );
  INV_X1 U23943 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20973) );
  OAI222_X1 U23944 ( .A1(n20974), .A2(n21178), .B1(n20973), .B2(n20972), .C1(
        n20971), .C2(n20970), .ZN(P1_U3226) );
  INV_X1 U23945 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U23946 ( .A1(n20972), .A2(n21167), .B1(n20975), .B2(n21023), .ZN(
        P1_U3458) );
  INV_X1 U23947 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20997) );
  INV_X1 U23948 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U23949 ( .A1(n20972), .A2(n20997), .B1(n20976), .B2(n21023), .ZN(
        P1_U3459) );
  INV_X1 U23950 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20977) );
  AOI22_X1 U23951 ( .A1(n20972), .A2(n21190), .B1(n20977), .B2(n21023), .ZN(
        P1_U3460) );
  INV_X1 U23952 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21131) );
  INV_X1 U23953 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20978) );
  AOI22_X1 U23954 ( .A1(n20972), .A2(n21131), .B1(n20978), .B2(n21023), .ZN(
        P1_U3461) );
  INV_X1 U23955 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20981) );
  INV_X1 U23956 ( .A(n20982), .ZN(n20979) );
  AOI21_X1 U23957 ( .B1(n20981), .B2(n20980), .A(n20979), .ZN(P1_U3464) );
  OAI21_X1 U23958 ( .B1(n20984), .B2(n20983), .A(n20982), .ZN(P1_U3465) );
  AOI21_X1 U23959 ( .B1(n20986), .B2(n20985), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n20988) );
  OAI22_X1 U23960 ( .A1(n20989), .A2(n20988), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20987), .ZN(n20991) );
  AOI22_X1 U23961 ( .A1(n20992), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20991), .B2(n20990), .ZN(n20993) );
  OAI21_X1 U23962 ( .B1(n20995), .B2(n20994), .A(n20993), .ZN(P1_U3474) );
  AOI21_X1 U23963 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20996) );
  AOI22_X1 U23964 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20996), .B2(n21352), .ZN(n20998) );
  AOI22_X1 U23965 ( .A1(n20999), .A2(n20998), .B1(n20997), .B2(n21001), .ZN(
        P1_U3481) );
  INV_X1 U23966 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21169) );
  NOR2_X1 U23967 ( .A1(n21001), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U23968 ( .A1(n21131), .A2(n21001), .B1(n21169), .B2(n21000), .ZN(
        P1_U3482) );
  AOI22_X1 U23969 ( .A1(n20972), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21104), 
        .B2(n21023), .ZN(P1_U3483) );
  AOI22_X1 U23970 ( .A1(n21004), .A2(n21003), .B1(n21222), .B2(n21002), .ZN(
        P1_U3484) );
  NOR2_X1 U23971 ( .A1(n21005), .A2(n20625), .ZN(n21013) );
  AOI211_X1 U23972 ( .C1(n21008), .C2(n21013), .A(n21007), .B(n21006), .ZN(
        n21021) );
  INV_X1 U23973 ( .A(n21009), .ZN(n21017) );
  OAI21_X1 U23974 ( .B1(n21011), .B2(n21346), .A(n21010), .ZN(n21014) );
  AOI21_X1 U23975 ( .B1(n21014), .B2(n21013), .A(n21012), .ZN(n21015) );
  AOI21_X1 U23976 ( .B1(n21017), .B2(n21016), .A(n21015), .ZN(n21020) );
  NOR2_X1 U23977 ( .A1(n21021), .A2(n21018), .ZN(n21019) );
  AOI22_X1 U23978 ( .A1(n21022), .A2(n21021), .B1(n21020), .B2(n21019), .ZN(
        P1_U3485) );
  INV_X1 U23979 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21024) );
  AOI22_X1 U23980 ( .A1(n20972), .A2(n21024), .B1(n21140), .B2(n21023), .ZN(
        P1_U3486) );
  OAI22_X1 U23981 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        DATAI_4_), .B2(keyinput_g28), .ZN(n21025) );
  AOI221_X1 U23982 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .C1(
        keyinput_g28), .C2(DATAI_4_), .A(n21025), .ZN(n21032) );
  OAI22_X1 U23983 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_g124), .B1(
        keyinput_g82), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n21026) );
  AOI221_X1 U23984 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_g124), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_g82), .A(n21026), .ZN(n21031) );
  OAI22_X1 U23985 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g84), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n21027) );
  AOI221_X1 U23986 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_g84), .A(n21027), .ZN(n21030) );
  OAI22_X1 U23987 ( .A1(DATAI_27_), .A2(keyinput_g5), .B1(keyinput_g31), .B2(
        DATAI_1_), .ZN(n21028) );
  AOI221_X1 U23988 ( .B1(DATAI_27_), .B2(keyinput_g5), .C1(DATAI_1_), .C2(
        keyinput_g31), .A(n21028), .ZN(n21029) );
  NAND4_X1 U23989 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21064) );
  OAI22_X1 U23990 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(keyinput_g78), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n21033) );
  AOI221_X1 U23991 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(keyinput_g78), .C1(
        keyinput_g61), .C2(P1_REIP_REG_22__SCAN_IN), .A(n21033), .ZN(n21040)
         );
  OAI22_X1 U23992 ( .A1(READY1), .A2(keyinput_g36), .B1(keyinput_g43), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21034) );
  AOI221_X1 U23993 ( .B1(READY1), .B2(keyinput_g36), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g43), .A(n21034), .ZN(
        n21039) );
  OAI22_X1 U23994 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_g87), .B1(
        keyinput_g22), .B2(DATAI_10_), .ZN(n21035) );
  AOI221_X1 U23995 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_g87), .C1(
        DATAI_10_), .C2(keyinput_g22), .A(n21035), .ZN(n21038) );
  OAI22_X1 U23996 ( .A1(DATAI_13_), .A2(keyinput_g19), .B1(keyinput_g39), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n21036) );
  AOI221_X1 U23997 ( .B1(DATAI_13_), .B2(keyinput_g19), .C1(
        P1_ADS_N_REG_SCAN_IN), .C2(keyinput_g39), .A(n21036), .ZN(n21037) );
  NAND4_X1 U23998 ( .A1(n21040), .A2(n21039), .A3(n21038), .A4(n21037), .ZN(
        n21063) );
  OAI22_X1 U23999 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        DATAI_29_), .B2(keyinput_g3), .ZN(n21041) );
  AOI221_X1 U24000 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        keyinput_g3), .C2(DATAI_29_), .A(n21041), .ZN(n21048) );
  OAI22_X1 U24001 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_g123), .B1(
        DATAI_8_), .B2(keyinput_g24), .ZN(n21042) );
  AOI221_X1 U24002 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_g123), .C1(
        keyinput_g24), .C2(DATAI_8_), .A(n21042), .ZN(n21047) );
  OAI22_X1 U24003 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_g110), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(keyinput_g81), .ZN(n21043) );
  AOI221_X1 U24004 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g81), .C2(P1_REIP_REG_2__SCAN_IN), .A(n21043), .ZN(n21046) );
  OAI22_X1 U24005 ( .A1(DATAI_28_), .A2(keyinput_g4), .B1(keyinput_g29), .B2(
        DATAI_3_), .ZN(n21044) );
  AOI221_X1 U24006 ( .B1(DATAI_28_), .B2(keyinput_g4), .C1(DATAI_3_), .C2(
        keyinput_g29), .A(n21044), .ZN(n21045) );
  NAND4_X1 U24007 ( .A1(n21048), .A2(n21047), .A3(n21046), .A4(n21045), .ZN(
        n21062) );
  AOI22_X1 U24008 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(n11679), .B2(
        keyinput_g1), .ZN(n21049) );
  OAI221_X1 U24009 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(n11679), .C2(
        keyinput_g1), .A(n21049), .ZN(n21060) );
  AOI22_X1 U24010 ( .A1(n14280), .A2(keyinput_g96), .B1(keyinput_g13), .B2(
        n21051), .ZN(n21050) );
  OAI221_X1 U24011 ( .B1(n14280), .B2(keyinput_g96), .C1(n21051), .C2(
        keyinput_g13), .A(n21050), .ZN(n21059) );
  AOI22_X1 U24012 ( .A1(n21054), .A2(keyinput_g2), .B1(n21053), .B2(
        keyinput_g119), .ZN(n21052) );
  OAI221_X1 U24013 ( .B1(n21054), .B2(keyinput_g2), .C1(n21053), .C2(
        keyinput_g119), .A(n21052), .ZN(n21058) );
  INV_X1 U24014 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21056) );
  AOI22_X1 U24015 ( .A1(n21273), .A2(keyinput_g62), .B1(keyinput_g38), .B2(
        n21056), .ZN(n21055) );
  OAI221_X1 U24016 ( .B1(n21273), .B2(keyinput_g62), .C1(n21056), .C2(
        keyinput_g38), .A(n21055), .ZN(n21057) );
  OR4_X1 U24017 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21061) );
  NOR4_X1 U24018 ( .A1(n21064), .A2(n21063), .A3(n21062), .A4(n21061), .ZN(
        n21408) );
  OAI22_X1 U24019 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_g122), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .ZN(n21065) );
  AOI221_X1 U24020 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g52), .C2(P1_REIP_REG_31__SCAN_IN), .A(n21065), .ZN(n21072)
         );
  OAI22_X1 U24021 ( .A1(DATAI_6_), .A2(keyinput_g26), .B1(DATAI_18_), .B2(
        keyinput_g14), .ZN(n21066) );
  AOI221_X1 U24022 ( .B1(DATAI_6_), .B2(keyinput_g26), .C1(keyinput_g14), .C2(
        DATAI_18_), .A(n21066), .ZN(n21071) );
  OAI22_X1 U24023 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(keyinput_g71), .B1(
        keyinput_g50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21067) );
  AOI221_X1 U24024 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(keyinput_g71), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g50), .A(n21067), .ZN(
        n21070) );
  OAI22_X1 U24025 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_g72), .B1(
        keyinput_g18), .B2(DATAI_14_), .ZN(n21068) );
  AOI221_X1 U24026 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_g72), .C1(
        DATAI_14_), .C2(keyinput_g18), .A(n21068), .ZN(n21069) );
  NAND4_X1 U24027 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21207) );
  OAI22_X1 U24028 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_g112), .B1(
        keyinput_g68), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n21073) );
  AOI221_X1 U24029 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_g112), .C1(
        P1_REIP_REG_15__SCAN_IN), .C2(keyinput_g68), .A(n21073), .ZN(n21099)
         );
  OAI22_X1 U24030 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g20), .B2(DATAI_12_), .ZN(n21074) );
  AOI221_X1 U24031 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_g76), .C1(
        DATAI_12_), .C2(keyinput_g20), .A(n21074), .ZN(n21077) );
  OAI22_X1 U24032 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        DATAI_15_), .B2(keyinput_g17), .ZN(n21075) );
  AOI221_X1 U24033 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g17), .C2(DATAI_15_), .A(n21075), .ZN(n21076) );
  OAI211_X1 U24034 ( .C1(n21079), .C2(keyinput_g127), .A(n21077), .B(n21076), 
        .ZN(n21078) );
  AOI21_X1 U24035 ( .B1(n21079), .B2(keyinput_g127), .A(n21078), .ZN(n21098)
         );
  AOI22_X1 U24036 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .ZN(n21080) );
  OAI221_X1 U24037 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(
        P1_REIP_REG_4__SCAN_IN), .C2(keyinput_g79), .A(n21080), .ZN(n21087) );
  AOI22_X1 U24038 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .ZN(n21081) );
  OAI221_X1 U24039 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_g57), .A(n21081), .ZN(n21086)
         );
  AOI22_X1 U24040 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_g93), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_g117), .ZN(n21082) );
  OAI221_X1 U24041 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_g117), .A(n21082), .ZN(n21085)
         );
  AOI22_X1 U24042 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_g113), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(keyinput_g97), .ZN(n21083) );
  OAI221_X1 U24043 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_g113), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_g97), .A(n21083), .ZN(n21084) );
  NOR4_X1 U24044 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21097) );
  AOI22_X1 U24045 ( .A1(DATAI_16_), .A2(keyinput_g16), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(keyinput_g77), .ZN(n21088) );
  OAI221_X1 U24046 ( .B1(DATAI_16_), .B2(keyinput_g16), .C1(
        P1_REIP_REG_6__SCAN_IN), .C2(keyinput_g77), .A(n21088), .ZN(n21095) );
  AOI22_X1 U24047 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .ZN(n21089) );
  OAI221_X1 U24048 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(n21089), .ZN(n21094)
         );
  AOI22_X1 U24049 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_g104), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .ZN(n21090) );
  OAI221_X1 U24050 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_g126), .A(n21090), .ZN(n21093)
         );
  AOI22_X1 U24051 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_g64), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput_g98), .ZN(n21091) );
  OAI221_X1 U24052 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_g64), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_g98), .A(n21091), .ZN(n21092) );
  NOR4_X1 U24053 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21096) );
  NAND4_X1 U24054 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21206) );
  AOI22_X1 U24055 ( .A1(n21102), .A2(keyinput_g40), .B1(n21101), .B2(
        keyinput_g12), .ZN(n21100) );
  OAI221_X1 U24056 ( .B1(n21102), .B2(keyinput_g40), .C1(n21101), .C2(
        keyinput_g12), .A(n21100), .ZN(n21112) );
  AOI22_X1 U24057 ( .A1(n21104), .A2(keyinput_g47), .B1(n14306), .B2(
        keyinput_g100), .ZN(n21103) );
  OAI221_X1 U24058 ( .B1(n21104), .B2(keyinput_g47), .C1(n14306), .C2(
        keyinput_g100), .A(n21103), .ZN(n21111) );
  AOI22_X1 U24059 ( .A1(n21384), .A2(keyinput_g56), .B1(n21106), .B2(
        keyinput_g115), .ZN(n21105) );
  OAI221_X1 U24060 ( .B1(n21384), .B2(keyinput_g56), .C1(n21106), .C2(
        keyinput_g115), .A(n21105), .ZN(n21110) );
  INV_X1 U24061 ( .A(DATAI_7_), .ZN(n21212) );
  AOI22_X1 U24062 ( .A1(n21212), .A2(keyinput_g25), .B1(keyinput_g35), .B2(
        n21108), .ZN(n21107) );
  OAI221_X1 U24063 ( .B1(n21212), .B2(keyinput_g25), .C1(n21108), .C2(
        keyinput_g35), .A(n21107), .ZN(n21109) );
  NOR4_X1 U24064 ( .A1(n21112), .A2(n21111), .A3(n21110), .A4(n21109), .ZN(
        n21152) );
  AOI22_X1 U24065 ( .A1(n21220), .A2(keyinput_g55), .B1(n21349), .B2(
        keyinput_g88), .ZN(n21113) );
  OAI221_X1 U24066 ( .B1(n21220), .B2(keyinput_g55), .C1(n21349), .C2(
        keyinput_g88), .A(n21113), .ZN(n21124) );
  INV_X1 U24067 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21115) );
  AOI22_X1 U24068 ( .A1(n21115), .A2(keyinput_g116), .B1(keyinput_g46), .B2(
        n21213), .ZN(n21114) );
  OAI221_X1 U24069 ( .B1(n21115), .B2(keyinput_g116), .C1(n21213), .C2(
        keyinput_g46), .A(n21114), .ZN(n21123) );
  INV_X1 U24070 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n21335) );
  AOI22_X1 U24071 ( .A1(n21335), .A2(keyinput_g102), .B1(keyinput_g34), .B2(
        n21117), .ZN(n21116) );
  OAI221_X1 U24072 ( .B1(n21335), .B2(keyinput_g102), .C1(n21117), .C2(
        keyinput_g34), .A(n21116), .ZN(n21122) );
  AOI22_X1 U24073 ( .A1(n21120), .A2(keyinput_g58), .B1(n21119), .B2(
        keyinput_g66), .ZN(n21118) );
  OAI221_X1 U24074 ( .B1(n21120), .B2(keyinput_g58), .C1(n21119), .C2(
        keyinput_g66), .A(n21118), .ZN(n21121) );
  NOR4_X1 U24075 ( .A1(n21124), .A2(n21123), .A3(n21122), .A4(n21121), .ZN(
        n21151) );
  AOI22_X1 U24076 ( .A1(n21126), .A2(keyinput_g69), .B1(n21334), .B2(
        keyinput_g109), .ZN(n21125) );
  OAI221_X1 U24077 ( .B1(n21126), .B2(keyinput_g69), .C1(n21334), .C2(
        keyinput_g109), .A(n21125), .ZN(n21137) );
  AOI22_X1 U24078 ( .A1(n21129), .A2(keyinput_g27), .B1(n21128), .B2(
        keyinput_g65), .ZN(n21127) );
  OAI221_X1 U24079 ( .B1(n21129), .B2(keyinput_g27), .C1(n21128), .C2(
        keyinput_g65), .A(n21127), .ZN(n21136) );
  AOI22_X1 U24080 ( .A1(n21132), .A2(keyinput_g89), .B1(keyinput_g48), .B2(
        n21131), .ZN(n21130) );
  OAI221_X1 U24081 ( .B1(n21132), .B2(keyinput_g89), .C1(n21131), .C2(
        keyinput_g48), .A(n21130), .ZN(n21135) );
  AOI22_X1 U24082 ( .A1(n21225), .A2(keyinput_g10), .B1(n21353), .B2(
        keyinput_g95), .ZN(n21133) );
  OAI221_X1 U24083 ( .B1(n21225), .B2(keyinput_g10), .C1(n21353), .C2(
        keyinput_g95), .A(n21133), .ZN(n21134) );
  NOR4_X1 U24084 ( .A1(n21137), .A2(n21136), .A3(n21135), .A4(n21134), .ZN(
        n21150) );
  AOI22_X1 U24085 ( .A1(n21229), .A2(keyinput_g92), .B1(keyinput_g75), .B2(
        n21226), .ZN(n21138) );
  OAI221_X1 U24086 ( .B1(n21229), .B2(keyinput_g92), .C1(n21226), .C2(
        keyinput_g75), .A(n21138), .ZN(n21148) );
  AOI22_X1 U24087 ( .A1(n21140), .A2(keyinput_g41), .B1(n21250), .B2(
        keyinput_g107), .ZN(n21139) );
  OAI221_X1 U24088 ( .B1(n21140), .B2(keyinput_g41), .C1(n21250), .C2(
        keyinput_g107), .A(n21139), .ZN(n21147) );
  AOI22_X1 U24089 ( .A1(n21381), .A2(keyinput_g106), .B1(keyinput_g30), .B2(
        n21142), .ZN(n21141) );
  OAI221_X1 U24090 ( .B1(n21381), .B2(keyinput_g106), .C1(n21142), .C2(
        keyinput_g30), .A(n21141), .ZN(n21146) );
  AOI22_X1 U24091 ( .A1(n21219), .A2(keyinput_g74), .B1(keyinput_g6), .B2(
        n21144), .ZN(n21143) );
  OAI221_X1 U24092 ( .B1(n21219), .B2(keyinput_g74), .C1(n21144), .C2(
        keyinput_g6), .A(n21143), .ZN(n21145) );
  NOR4_X1 U24093 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21149) );
  NAND4_X1 U24094 ( .A1(n21152), .A2(n21151), .A3(n21150), .A4(n21149), .ZN(
        n21205) );
  INV_X1 U24095 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21378) );
  AOI22_X1 U24096 ( .A1(n21347), .A2(keyinput_g105), .B1(n21378), .B2(
        keyinput_g103), .ZN(n21153) );
  OAI221_X1 U24097 ( .B1(n21347), .B2(keyinput_g105), .C1(n21378), .C2(
        keyinput_g103), .A(n21153), .ZN(n21163) );
  INV_X1 U24098 ( .A(READY2), .ZN(n21155) );
  AOI22_X1 U24099 ( .A1(n21155), .A2(keyinput_g37), .B1(n21350), .B2(
        keyinput_g11), .ZN(n21154) );
  OAI221_X1 U24100 ( .B1(n21155), .B2(keyinput_g37), .C1(n21350), .C2(
        keyinput_g11), .A(n21154), .ZN(n21162) );
  AOI22_X1 U24101 ( .A1(n21157), .A2(keyinput_g111), .B1(keyinput_g8), .B2(
        n21337), .ZN(n21156) );
  OAI221_X1 U24102 ( .B1(n21157), .B2(keyinput_g111), .C1(n21337), .C2(
        keyinput_g8), .A(n21156), .ZN(n21161) );
  AOI22_X1 U24103 ( .A1(n21228), .A2(keyinput_g91), .B1(n21159), .B2(
        keyinput_g90), .ZN(n21158) );
  OAI221_X1 U24104 ( .B1(n21228), .B2(keyinput_g91), .C1(n21159), .C2(
        keyinput_g90), .A(n21158), .ZN(n21160) );
  NOR4_X1 U24105 ( .A1(n21163), .A2(n21162), .A3(n21161), .A4(n21160), .ZN(
        n21203) );
  AOI22_X1 U24106 ( .A1(n21363), .A2(keyinput_g70), .B1(keyinput_g7), .B2(
        n21165), .ZN(n21164) );
  OAI221_X1 U24107 ( .B1(n21363), .B2(keyinput_g70), .C1(n21165), .C2(
        keyinput_g7), .A(n21164), .ZN(n21175) );
  AOI22_X1 U24108 ( .A1(n21355), .A2(keyinput_g60), .B1(keyinput_g51), .B2(
        n21167), .ZN(n21166) );
  OAI221_X1 U24109 ( .B1(n21355), .B2(keyinput_g60), .C1(n21167), .C2(
        keyinput_g51), .A(n21166), .ZN(n21174) );
  INV_X1 U24110 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21244) );
  AOI22_X1 U24111 ( .A1(n21244), .A2(keyinput_g94), .B1(keyinput_g83), .B2(
        n21169), .ZN(n21168) );
  OAI221_X1 U24112 ( .B1(n21244), .B2(keyinput_g94), .C1(n21169), .C2(
        keyinput_g83), .A(n21168), .ZN(n21173) );
  AOI22_X1 U24113 ( .A1(n21171), .A2(keyinput_g121), .B1(keyinput_g54), .B2(
        n21249), .ZN(n21170) );
  OAI221_X1 U24114 ( .B1(n21171), .B2(keyinput_g121), .C1(n21249), .C2(
        keyinput_g54), .A(n21170), .ZN(n21172) );
  NOR4_X1 U24115 ( .A1(n21175), .A2(n21174), .A3(n21173), .A4(n21172), .ZN(
        n21202) );
  AOI22_X1 U24116 ( .A1(n21254), .A2(keyinput_g33), .B1(n11294), .B2(
        keyinput_g120), .ZN(n21176) );
  OAI221_X1 U24117 ( .B1(n21254), .B2(keyinput_g33), .C1(n11294), .C2(
        keyinput_g120), .A(n21176), .ZN(n21185) );
  AOI22_X1 U24118 ( .A1(n21178), .A2(keyinput_g53), .B1(keyinput_g67), .B2(
        n14637), .ZN(n21177) );
  OAI221_X1 U24119 ( .B1(n21178), .B2(keyinput_g53), .C1(n14637), .C2(
        keyinput_g67), .A(n21177), .ZN(n21184) );
  AOI22_X1 U24120 ( .A1(n10416), .A2(keyinput_g114), .B1(keyinput_g45), .B2(
        n21222), .ZN(n21179) );
  OAI221_X1 U24121 ( .B1(n10416), .B2(keyinput_g114), .C1(n21222), .C2(
        keyinput_g45), .A(n21179), .ZN(n21183) );
  AOI22_X1 U24122 ( .A1(n21364), .A2(keyinput_g73), .B1(n21181), .B2(
        keyinput_g108), .ZN(n21180) );
  OAI221_X1 U24123 ( .B1(n21364), .B2(keyinput_g73), .C1(n21181), .C2(
        keyinput_g108), .A(n21180), .ZN(n21182) );
  NOR4_X1 U24124 ( .A1(n21185), .A2(n21184), .A3(n21183), .A4(n21182), .ZN(
        n21201) );
  AOI22_X1 U24125 ( .A1(n21188), .A2(keyinput_g99), .B1(keyinput_g80), .B2(
        n21187), .ZN(n21186) );
  OAI221_X1 U24126 ( .B1(n21188), .B2(keyinput_g99), .C1(n21187), .C2(
        keyinput_g80), .A(n21186), .ZN(n21199) );
  AOI22_X1 U24127 ( .A1(n21191), .A2(keyinput_g86), .B1(keyinput_g49), .B2(
        n21190), .ZN(n21189) );
  OAI221_X1 U24128 ( .B1(n21191), .B2(keyinput_g86), .C1(n21190), .C2(
        keyinput_g49), .A(n21189), .ZN(n21198) );
  INV_X1 U24129 ( .A(DATAI_11_), .ZN(n21247) );
  AOI22_X1 U24130 ( .A1(n21247), .A2(keyinput_g21), .B1(n10660), .B2(
        keyinput_g118), .ZN(n21192) );
  OAI221_X1 U24131 ( .B1(n21247), .B2(keyinput_g21), .C1(n10660), .C2(
        keyinput_g118), .A(n21192), .ZN(n21197) );
  AOI22_X1 U24132 ( .A1(n21195), .A2(keyinput_g85), .B1(keyinput_g9), .B2(
        n21194), .ZN(n21193) );
  OAI221_X1 U24133 ( .B1(n21195), .B2(keyinput_g85), .C1(n21194), .C2(
        keyinput_g9), .A(n21193), .ZN(n21196) );
  NOR4_X1 U24134 ( .A1(n21199), .A2(n21198), .A3(n21197), .A4(n21196), .ZN(
        n21200) );
  NAND4_X1 U24135 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21204) );
  NOR4_X1 U24136 ( .A1(n21207), .A2(n21206), .A3(n21205), .A4(n21204), .ZN(
        n21407) );
  AOI22_X1 U24137 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_f83), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_f115), .ZN(n21208) );
  OAI221_X1 U24138 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_f83), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_f115), .A(n21208), .ZN(n21217) );
  AOI22_X1 U24139 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21209) );
  OAI221_X1 U24140 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21209), .ZN(n21216)
         );
  AOI22_X1 U24141 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_f121), .ZN(n21210) );
  OAI221_X1 U24142 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_f121), .A(n21210), .ZN(n21215)
         );
  AOI22_X1 U24143 ( .A1(n21213), .A2(keyinput_f46), .B1(n21212), .B2(
        keyinput_f25), .ZN(n21211) );
  OAI221_X1 U24144 ( .B1(n21213), .B2(keyinput_f46), .C1(n21212), .C2(
        keyinput_f25), .A(n21211), .ZN(n21214) );
  NOR4_X1 U24145 ( .A1(n21217), .A2(n21216), .A3(n21215), .A4(n21214), .ZN(
        n21400) );
  AOI22_X1 U24146 ( .A1(n21220), .A2(keyinput_f55), .B1(n21219), .B2(
        keyinput_f74), .ZN(n21218) );
  OAI221_X1 U24147 ( .B1(n21220), .B2(keyinput_f55), .C1(n21219), .C2(
        keyinput_f74), .A(n21218), .ZN(n21233) );
  INV_X1 U24148 ( .A(READY1), .ZN(n21223) );
  AOI22_X1 U24149 ( .A1(n21223), .A2(keyinput_f36), .B1(keyinput_f45), .B2(
        n21222), .ZN(n21221) );
  OAI221_X1 U24150 ( .B1(n21223), .B2(keyinput_f36), .C1(n21222), .C2(
        keyinput_f45), .A(n21221), .ZN(n21232) );
  AOI22_X1 U24151 ( .A1(n21226), .A2(keyinput_f75), .B1(keyinput_f10), .B2(
        n21225), .ZN(n21224) );
  OAI221_X1 U24152 ( .B1(n21226), .B2(keyinput_f75), .C1(n21225), .C2(
        keyinput_f10), .A(n21224), .ZN(n21231) );
  AOI22_X1 U24153 ( .A1(n21229), .A2(keyinput_f92), .B1(n21228), .B2(
        keyinput_f91), .ZN(n21227) );
  OAI221_X1 U24154 ( .B1(n21229), .B2(keyinput_f92), .C1(n21228), .C2(
        keyinput_f91), .A(n21227), .ZN(n21230) );
  NOR4_X1 U24155 ( .A1(n21233), .A2(n21232), .A3(n21231), .A4(n21230), .ZN(
        n21399) );
  OAI22_X1 U24156 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_f76), .B1(
        keyinput_f5), .B2(DATAI_27_), .ZN(n21234) );
  AOI221_X1 U24157 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_f76), .C1(
        DATAI_27_), .C2(keyinput_f5), .A(n21234), .ZN(n21241) );
  OAI22_X1 U24158 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_f84), .B1(
        DATAI_12_), .B2(keyinput_f20), .ZN(n21235) );
  AOI221_X1 U24159 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .C1(
        keyinput_f20), .C2(DATAI_12_), .A(n21235), .ZN(n21240) );
  OAI22_X1 U24160 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .ZN(n21236) );
  AOI221_X1 U24161 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .C1(
        keyinput_f66), .C2(P1_REIP_REG_17__SCAN_IN), .A(n21236), .ZN(n21239)
         );
  OAI22_X1 U24162 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_f87), .B1(
        keyinput_f35), .B2(BS16), .ZN(n21237) );
  AOI221_X1 U24163 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .C1(BS16), 
        .C2(keyinput_f35), .A(n21237), .ZN(n21238) );
  NAND4_X1 U24164 ( .A1(n21241), .A2(n21240), .A3(n21239), .A4(n21238), .ZN(
        n21258) );
  AOI22_X1 U24165 ( .A1(n21244), .A2(keyinput_f94), .B1(keyinput_f113), .B2(
        n21243), .ZN(n21242) );
  OAI221_X1 U24166 ( .B1(n21244), .B2(keyinput_f94), .C1(n21243), .C2(
        keyinput_f113), .A(n21242), .ZN(n21257) );
  AOI22_X1 U24167 ( .A1(n21247), .A2(keyinput_f21), .B1(n21246), .B2(
        keyinput_f63), .ZN(n21245) );
  OAI221_X1 U24168 ( .B1(n21247), .B2(keyinput_f21), .C1(n21246), .C2(
        keyinput_f63), .A(n21245), .ZN(n21256) );
  XOR2_X1 U24169 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_f39), .Z(n21252) );
  AOI22_X1 U24170 ( .A1(n21250), .A2(keyinput_f107), .B1(keyinput_f54), .B2(
        n21249), .ZN(n21248) );
  OAI221_X1 U24171 ( .B1(n21250), .B2(keyinput_f107), .C1(n21249), .C2(
        keyinput_f54), .A(n21248), .ZN(n21251) );
  AOI211_X1 U24172 ( .C1(n21254), .C2(keyinput_f33), .A(n21252), .B(n21251), 
        .ZN(n21253) );
  OAI21_X1 U24173 ( .B1(n21254), .B2(keyinput_f33), .A(n21253), .ZN(n21255) );
  NOR4_X1 U24174 ( .A1(n21258), .A2(n21257), .A3(n21256), .A4(n21255), .ZN(
        n21398) );
  OAI22_X1 U24175 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(keyinput_f0), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21259) );
  AOI221_X1 U24176 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_f0), .A(n21259), .ZN(n21266)
         );
  OAI22_X1 U24177 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f12), .B2(DATAI_20_), .ZN(n21260) );
  AOI221_X1 U24178 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .C1(
        DATAI_20_), .C2(keyinput_f12), .A(n21260), .ZN(n21265) );
  OAI22_X1 U24179 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n21261) );
  AOI221_X1 U24180 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(keyinput_f43), 
        .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n21261), .ZN(n21264) );
  OAI22_X1 U24181 ( .A1(DATAI_10_), .A2(keyinput_f22), .B1(keyinput_f51), .B2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21262) );
  AOI221_X1 U24182 ( .B1(DATAI_10_), .B2(keyinput_f22), .C1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_f51), .A(n21262), .ZN(
        n21263) );
  NAND4_X1 U24183 ( .A1(n21266), .A2(n21265), .A3(n21264), .A4(n21263), .ZN(
        n21396) );
  OAI22_X1 U24184 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(keyinput_f99), .B1(
        keyinput_f108), .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n21267) );
  AOI221_X1 U24185 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(keyinput_f99), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_f108), .A(n21267), .ZN(n21293) );
  OAI22_X1 U24186 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_f112), .B1(
        keyinput_f30), .B2(DATAI_2_), .ZN(n21268) );
  AOI221_X1 U24187 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .C1(
        DATAI_2_), .C2(keyinput_f30), .A(n21268), .ZN(n21271) );
  OAI22_X1 U24188 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_f123), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n21269) );
  AOI221_X1 U24189 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .C1(
        keyinput_f58), .C2(P1_REIP_REG_25__SCAN_IN), .A(n21269), .ZN(n21270)
         );
  OAI211_X1 U24190 ( .C1(n21273), .C2(keyinput_f62), .A(n21271), .B(n21270), 
        .ZN(n21272) );
  AOI21_X1 U24191 ( .B1(n21273), .B2(keyinput_f62), .A(n21272), .ZN(n21292) );
  AOI22_X1 U24192 ( .A1(DATAI_6_), .A2(keyinput_f26), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_f59), .ZN(n21274) );
  OAI221_X1 U24193 ( .B1(DATAI_6_), .B2(keyinput_f26), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_f59), .A(n21274), .ZN(n21281)
         );
  AOI22_X1 U24194 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_f47), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_f127), .ZN(n21275) );
  OAI221_X1 U24195 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_f47), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_f127), .A(n21275), .ZN(n21280)
         );
  AOI22_X1 U24196 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .ZN(n21276) );
  OAI221_X1 U24197 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        P1_EAX_REG_23__SCAN_IN), .C2(keyinput_f124), .A(n21276), .ZN(n21279)
         );
  AOI22_X1 U24198 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_f96), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n21277) );
  OAI221_X1 U24199 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n21277), .ZN(n21278)
         );
  NOR4_X1 U24200 ( .A1(n21281), .A2(n21280), .A3(n21279), .A4(n21278), .ZN(
        n21291) );
  AOI22_X1 U24201 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .ZN(n21282) );
  OAI221_X1 U24202 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_f85), .A(n21282), .ZN(n21289) );
  AOI22_X1 U24203 ( .A1(DATAI_5_), .A2(keyinput_f27), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(keyinput_f72), .ZN(n21283) );
  OAI221_X1 U24204 ( .B1(DATAI_5_), .B2(keyinput_f27), .C1(
        P1_REIP_REG_11__SCAN_IN), .C2(keyinput_f72), .A(n21283), .ZN(n21288)
         );
  AOI22_X1 U24205 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput_f68), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_f125), .ZN(n21284) );
  OAI221_X1 U24206 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput_f68), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_f125), .A(n21284), .ZN(n21287)
         );
  AOI22_X1 U24207 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(keyinput_f90), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .ZN(n21285) );
  OAI221_X1 U24208 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(keyinput_f90), .C1(
        P1_EAX_REG_31__SCAN_IN), .C2(keyinput_f116), .A(n21285), .ZN(n21286)
         );
  NOR4_X1 U24209 ( .A1(n21289), .A2(n21288), .A3(n21287), .A4(n21286), .ZN(
        n21290) );
  NAND4_X1 U24210 ( .A1(n21293), .A2(n21292), .A3(n21291), .A4(n21290), .ZN(
        n21395) );
  AOI22_X1 U24211 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(DATAI_31_), .B2(
        keyinput_f1), .ZN(n21294) );
  OAI221_X1 U24212 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(DATAI_31_), .C2(
        keyinput_f1), .A(n21294), .ZN(n21301) );
  AOI22_X1 U24213 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput_f98), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(keyinput_f122), .ZN(n21295) );
  OAI221_X1 U24214 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput_f98), .C1(
        P1_EAX_REG_25__SCAN_IN), .C2(keyinput_f122), .A(n21295), .ZN(n21300)
         );
  AOI22_X1 U24215 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(DATAI_26_), .B2(
        keyinput_f6), .ZN(n21296) );
  OAI221_X1 U24216 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(DATAI_26_), .C2(
        keyinput_f6), .A(n21296), .ZN(n21299) );
  AOI22_X1 U24217 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput_f81), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .ZN(n21297) );
  OAI221_X1 U24218 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_f81), .C1(
        P1_EBX_REG_4__SCAN_IN), .C2(keyinput_f111), .A(n21297), .ZN(n21298) );
  NOR4_X1 U24219 ( .A1(n21301), .A2(n21300), .A3(n21299), .A4(n21298), .ZN(
        n21329) );
  AOI22_X1 U24220 ( .A1(DATAI_13_), .A2(keyinput_f19), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput_f110), .ZN(n21302) );
  OAI221_X1 U24221 ( .B1(DATAI_13_), .B2(keyinput_f19), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput_f110), .A(n21302), .ZN(n21309) );
  AOI22_X1 U24222 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_14_), .B2(
        keyinput_f18), .ZN(n21303) );
  OAI221_X1 U24223 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_14_), .C2(
        keyinput_f18), .A(n21303), .ZN(n21308) );
  AOI22_X1 U24224 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .ZN(n21304) );
  OAI221_X1 U24225 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_f126), .A(n21304), .ZN(n21307)
         );
  AOI22_X1 U24226 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(
        P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .ZN(n21305) );
  OAI221_X1 U24227 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(
        P1_EBX_REG_26__SCAN_IN), .C2(keyinput_f89), .A(n21305), .ZN(n21306) );
  NOR4_X1 U24228 ( .A1(n21309), .A2(n21308), .A3(n21307), .A4(n21306), .ZN(
        n21328) );
  AOI22_X1 U24229 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(keyinput_f80), .ZN(n21310) );
  OAI221_X1 U24230 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(
        P1_REIP_REG_3__SCAN_IN), .C2(keyinput_f80), .A(n21310), .ZN(n21317) );
  AOI22_X1 U24231 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        DATAI_3_), .B2(keyinput_f29), .ZN(n21311) );
  OAI221_X1 U24232 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        DATAI_3_), .C2(keyinput_f29), .A(n21311), .ZN(n21316) );
  AOI22_X1 U24233 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .ZN(n21312) );
  OAI221_X1 U24234 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_f38), .A(n21312), .ZN(n21315) );
  AOI22_X1 U24235 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput_f86), .ZN(n21313) );
  OAI221_X1 U24236 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput_f86), .A(n21313), .ZN(n21314) );
  NOR4_X1 U24237 ( .A1(n21317), .A2(n21316), .A3(n21315), .A4(n21314), .ZN(
        n21327) );
  AOI22_X1 U24238 ( .A1(DATAI_1_), .A2(keyinput_f31), .B1(DATAI_29_), .B2(
        keyinput_f3), .ZN(n21318) );
  OAI221_X1 U24239 ( .B1(DATAI_1_), .B2(keyinput_f31), .C1(DATAI_29_), .C2(
        keyinput_f3), .A(n21318), .ZN(n21325) );
  AOI22_X1 U24240 ( .A1(READY2), .A2(keyinput_f37), .B1(P1_EAX_REG_28__SCAN_IN), .B2(keyinput_f119), .ZN(n21319) );
  OAI221_X1 U24241 ( .B1(READY2), .B2(keyinput_f37), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n21319), .ZN(n21324)
         );
  AOI22_X1 U24242 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(keyinput_f69), .ZN(n21320) );
  OAI221_X1 U24243 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(keyinput_f69), .A(n21320), .ZN(n21323)
         );
  AOI22_X1 U24244 ( .A1(keyinput_f41), .A2(P1_M_IO_N_REG_SCAN_IN), .B1(
        DATAI_4_), .B2(keyinput_f28), .ZN(n21321) );
  OAI221_X1 U24245 ( .B1(keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .C1(
        DATAI_4_), .C2(keyinput_f28), .A(n21321), .ZN(n21322) );
  NOR4_X1 U24246 ( .A1(n21325), .A2(n21324), .A3(n21323), .A4(n21322), .ZN(
        n21326) );
  NAND4_X1 U24247 ( .A1(n21329), .A2(n21328), .A3(n21327), .A4(n21326), .ZN(
        n21394) );
  INV_X1 U24248 ( .A(keyinput_f50), .ZN(n21331) );
  AOI22_X1 U24249 ( .A1(n21332), .A2(keyinput_f16), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n21331), .ZN(n21330) );
  OAI221_X1 U24250 ( .B1(n21332), .B2(keyinput_f16), .C1(n21331), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n21330), .ZN(n21344) );
  AOI22_X1 U24251 ( .A1(n21335), .A2(keyinput_f102), .B1(keyinput_f109), .B2(
        n21334), .ZN(n21333) );
  OAI221_X1 U24252 ( .B1(n21335), .B2(keyinput_f102), .C1(n21334), .C2(
        keyinput_f109), .A(n21333), .ZN(n21343) );
  AOI22_X1 U24253 ( .A1(n21337), .A2(keyinput_f8), .B1(n10416), .B2(
        keyinput_f114), .ZN(n21336) );
  OAI221_X1 U24254 ( .B1(n21337), .B2(keyinput_f8), .C1(n10416), .C2(
        keyinput_f114), .A(n21336), .ZN(n21342) );
  AOI22_X1 U24255 ( .A1(n21340), .A2(keyinput_f14), .B1(n21339), .B2(
        keyinput_f93), .ZN(n21338) );
  OAI221_X1 U24256 ( .B1(n21340), .B2(keyinput_f14), .C1(n21339), .C2(
        keyinput_f93), .A(n21338), .ZN(n21341) );
  NOR4_X1 U24257 ( .A1(n21344), .A2(n21343), .A3(n21342), .A4(n21341), .ZN(
        n21392) );
  AOI22_X1 U24258 ( .A1(n21347), .A2(keyinput_f105), .B1(n21346), .B2(
        keyinput_f44), .ZN(n21345) );
  OAI221_X1 U24259 ( .B1(n21347), .B2(keyinput_f105), .C1(n21346), .C2(
        keyinput_f44), .A(n21345), .ZN(n21359) );
  AOI22_X1 U24260 ( .A1(n21350), .A2(keyinput_f11), .B1(n21349), .B2(
        keyinput_f88), .ZN(n21348) );
  OAI221_X1 U24261 ( .B1(n21350), .B2(keyinput_f11), .C1(n21349), .C2(
        keyinput_f88), .A(n21348), .ZN(n21358) );
  AOI22_X1 U24262 ( .A1(n21353), .A2(keyinput_f95), .B1(keyinput_f82), .B2(
        n21352), .ZN(n21351) );
  OAI221_X1 U24263 ( .B1(n21353), .B2(keyinput_f95), .C1(n21352), .C2(
        keyinput_f82), .A(n21351), .ZN(n21357) );
  AOI22_X1 U24264 ( .A1(n13564), .A2(keyinput_f77), .B1(keyinput_f60), .B2(
        n21355), .ZN(n21354) );
  OAI221_X1 U24265 ( .B1(n13564), .B2(keyinput_f77), .C1(n21355), .C2(
        keyinput_f60), .A(n21354), .ZN(n21356) );
  NOR4_X1 U24266 ( .A1(n21359), .A2(n21358), .A3(n21357), .A4(n21356), .ZN(
        n21391) );
  INV_X1 U24267 ( .A(keyinput_f48), .ZN(n21361) );
  AOI22_X1 U24268 ( .A1(n14637), .A2(keyinput_f67), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n21361), .ZN(n21360) );
  OAI221_X1 U24269 ( .B1(n14637), .B2(keyinput_f67), .C1(n21361), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21360), .ZN(n21373) );
  AOI22_X1 U24270 ( .A1(n21364), .A2(keyinput_f73), .B1(keyinput_f70), .B2(
        n21363), .ZN(n21362) );
  OAI221_X1 U24271 ( .B1(n21364), .B2(keyinput_f73), .C1(n21363), .C2(
        keyinput_f70), .A(n21362), .ZN(n21372) );
  AOI22_X1 U24272 ( .A1(n14306), .A2(keyinput_f100), .B1(keyinput_f64), .B2(
        n21366), .ZN(n21365) );
  OAI221_X1 U24273 ( .B1(n14306), .B2(keyinput_f100), .C1(n21366), .C2(
        keyinput_f64), .A(n21365), .ZN(n21371) );
  AOI22_X1 U24274 ( .A1(n21369), .A2(keyinput_f4), .B1(n21368), .B2(
        keyinput_f78), .ZN(n21367) );
  OAI221_X1 U24275 ( .B1(n21369), .B2(keyinput_f4), .C1(n21368), .C2(
        keyinput_f78), .A(n21367), .ZN(n21370) );
  NOR4_X1 U24276 ( .A1(n21373), .A2(n21372), .A3(n21371), .A4(n21370), .ZN(
        n21390) );
  AOI22_X1 U24277 ( .A1(n21376), .A2(keyinput_f71), .B1(keyinput_f79), .B2(
        n21375), .ZN(n21374) );
  OAI221_X1 U24278 ( .B1(n21376), .B2(keyinput_f71), .C1(n21375), .C2(
        keyinput_f79), .A(n21374), .ZN(n21388) );
  AOI22_X1 U24279 ( .A1(n21379), .A2(keyinput_f97), .B1(keyinput_f103), .B2(
        n21378), .ZN(n21377) );
  OAI221_X1 U24280 ( .B1(n21379), .B2(keyinput_f97), .C1(n21378), .C2(
        keyinput_f103), .A(n21377), .ZN(n21387) );
  AOI22_X1 U24281 ( .A1(n11294), .A2(keyinput_f120), .B1(keyinput_f106), .B2(
        n21381), .ZN(n21380) );
  OAI221_X1 U24282 ( .B1(n11294), .B2(keyinput_f120), .C1(n21381), .C2(
        keyinput_f106), .A(n21380), .ZN(n21386) );
  INV_X1 U24283 ( .A(keyinput_f49), .ZN(n21383) );
  AOI22_X1 U24284 ( .A1(n21384), .A2(keyinput_f56), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n21383), .ZN(n21382) );
  OAI221_X1 U24285 ( .B1(n21384), .B2(keyinput_f56), .C1(n21383), .C2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .A(n21382), .ZN(n21385) );
  NOR4_X1 U24286 ( .A1(n21388), .A2(n21387), .A3(n21386), .A4(n21385), .ZN(
        n21389) );
  NAND4_X1 U24287 ( .A1(n21392), .A2(n21391), .A3(n21390), .A4(n21389), .ZN(
        n21393) );
  NOR4_X1 U24288 ( .A1(n21396), .A2(n21395), .A3(n21394), .A4(n21393), .ZN(
        n21397) );
  NAND4_X1 U24289 ( .A1(n21400), .A2(n21399), .A3(n21398), .A4(n21397), .ZN(
        n21402) );
  AOI21_X1 U24290 ( .B1(keyinput_f32), .B2(n21402), .A(keyinput_g32), .ZN(
        n21404) );
  INV_X1 U24291 ( .A(keyinput_f32), .ZN(n21401) );
  AOI21_X1 U24292 ( .B1(n21402), .B2(n21401), .A(n21405), .ZN(n21403) );
  AOI22_X1 U24293 ( .A1(n21405), .A2(n21404), .B1(keyinput_g32), .B2(n21403), 
        .ZN(n21406) );
  AOI21_X1 U24294 ( .B1(n21408), .B2(n21407), .A(n21406), .ZN(n21410) );
  AOI22_X1 U24295 ( .A1(n16637), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16639), .ZN(n21409) );
  XNOR2_X1 U24296 ( .A(n21410), .B(n21409), .ZN(U355) );
  AND3_X1 U13680 ( .A1(n10621), .A2(n10622), .A3(n10620), .ZN(n10627) );
  CLKBUF_X1 U11282 ( .A(n10697), .Z(n9839) );
  CLKBUF_X1 U11285 ( .A(n9811), .Z(n9853) );
  CLKBUF_X1 U11332 ( .A(n10668), .Z(n13594) );
  CLKBUF_X1 U11334 ( .A(n11877), .Z(n13277) );
  AND2_X2 U11335 ( .A1(n10616), .A2(n10518), .ZN(n9845) );
  NAND2_X1 U11338 ( .A1(n15128), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15118) );
  CLKBUF_X1 U11599 ( .A(n13137), .Z(n20720) );
  CLKBUF_X1 U11604 ( .A(n16631), .Z(n16634) );
  XOR2_X1 U11654 ( .A(n15042), .B(n15087), .Z(n21411) );
  INV_X1 U11657 ( .A(n12310), .ZN(n9803) );
  CLKBUF_X1 U11677 ( .A(n17644), .Z(n17653) );
endmodule

