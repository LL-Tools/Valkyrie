

module b22_C_gen_AntiSAT_k_256_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6664, n6665, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702;

  INV_X1 U7412 ( .A(P3_STATE_REG_SCAN_IN), .ZN(n10084) );
  CLKBUF_X2 U7413 ( .A(n11026), .Z(n12767) );
  CLKBUF_X2 U7414 ( .A(n9403), .Z(n9560) );
  INV_X1 U7415 ( .A(n8245), .ZN(n8537) );
  NAND3_X1 U7416 ( .A1(n7923), .A2(n7922), .A3(n7000), .ZN(n15315) );
  CLKBUF_X2 U7417 ( .A(n9279), .Z(n9411) );
  NAND2_X1 U7418 ( .A1(n6668), .A2(n6672), .ZN(n7921) );
  NAND2_X2 U7419 ( .A1(n10818), .A2(n6673), .ZN(n12162) );
  AND4_X1 U7420 ( .A1(n10602), .A2(n10601), .A3(n10600), .A4(n10599), .ZN(
        n10888) );
  OR2_X1 U7421 ( .A1(n8068), .A2(n6916), .ZN(n8070) );
  AND2_X1 U7422 ( .A1(n12378), .A2(n14767), .ZN(n12125) );
  AND2_X1 U7423 ( .A1(n10431), .A2(n6934), .ZN(n10189) );
  INV_X1 U7424 ( .A(n10084), .ZN(n6664) );
  INV_X1 U7425 ( .A(n6664), .ZN(n6665) );
  INV_X1 U7426 ( .A(n6664), .ZN(P3_U3151) );
  INV_X1 U7427 ( .A(n9826), .ZN(n9951) );
  INV_X1 U7428 ( .A(n9826), .ZN(n9931) );
  CLKBUF_X3 U7429 ( .A(n11546), .Z(n12770) );
  NOR2_X2 U7430 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n10173) );
  NAND2_X1 U7431 ( .A1(n9580), .A2(n9579), .ZN(n7731) );
  INV_X1 U7432 ( .A(n7731), .ZN(n9729) );
  INV_X1 U7433 ( .A(n8059), .ZN(n7908) );
  INV_X1 U7434 ( .A(n10818), .ZN(n12091) );
  NOR2_X2 U7435 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n10088) );
  INV_X1 U7436 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8910) );
  CLKBUF_X2 U7437 ( .A(n8728), .Z(n8787) );
  INV_X2 U7438 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8478) );
  INV_X1 U7439 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U7440 ( .A1(n8077), .A2(n8082), .ZN(n6869) );
  AND2_X1 U7441 ( .A1(n15226), .A2(n10249), .ZN(n15227) );
  OAI21_X1 U7442 ( .B1(n9525), .B2(n7258), .A(n7256), .ZN(n11599) );
  INV_X2 U7443 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14085) );
  AND2_X1 U7444 ( .A1(n8081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8072) );
  AND2_X2 U7446 ( .A1(n10582), .A2(n14767), .ZN(n10631) );
  AND2_X1 U7447 ( .A1(n14554), .A2(n14428), .ZN(n14537) );
  NAND2_X1 U7448 ( .A1(n14608), .A2(n14422), .ZN(n14424) );
  AND2_X1 U7449 ( .A1(n7322), .A2(n7321), .ZN(n14508) );
  INV_X1 U7450 ( .A(n12194), .ZN(n10570) );
  NAND2_X1 U7451 ( .A1(n10189), .A2(n10191), .ZN(n10187) );
  INV_X1 U7452 ( .A(n10860), .ZN(n12606) );
  NAND2_X1 U7453 ( .A1(n6869), .A2(n7874), .ZN(n10031) );
  OAI21_X1 U7454 ( .B1(n13898), .B2(n9425), .A(n6764), .ZN(n13882) );
  NAND2_X1 U7455 ( .A1(n14200), .A2(n14199), .ZN(n14198) );
  NAND2_X1 U7456 ( .A1(n14424), .A2(n6752), .ZN(n14593) );
  NAND2_X1 U7457 ( .A1(n10067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U7458 ( .A1(n10567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10569) );
  XNOR2_X1 U7459 ( .A(n7778), .B(n10077), .ZN(n7924) );
  AND2_X1 U7460 ( .A1(n6970), .A2(n6968), .ZN(n14481) );
  AND2_X1 U7461 ( .A1(n12378), .A2(n10581), .ZN(n12165) );
  BUF_X1 U7462 ( .A(n12052), .Z(n6673) );
  CLKBUF_X3 U7463 ( .A(n12052), .Z(n6672) );
  OR2_X2 U7464 ( .A1(n8549), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8562) );
  NAND2_X2 U7465 ( .A1(n13558), .A2(n13559), .ZN(n13524) );
  NAND2_X1 U7466 ( .A1(n6869), .A2(n7874), .ZN(n6667) );
  NAND2_X1 U7467 ( .A1(n6869), .A2(n7874), .ZN(n6668) );
  INV_X1 U7468 ( .A(n12165), .ZN(n6669) );
  NOR2_X2 U7469 ( .A1(n15693), .A2(n8888), .ZN(n8889) );
  AND2_X2 U7470 ( .A1(n6858), .A2(n7872), .ZN(n7636) );
  NAND2_X1 U7471 ( .A1(n11430), .A2(n9523), .ZN(n9525) );
  NAND2_X2 U7472 ( .A1(n10202), .A2(n14776), .ZN(n10818) );
  XNOR2_X2 U7473 ( .A(n10194), .B(n10193), .ZN(n10202) );
  OR2_X2 U7474 ( .A1(n13078), .A2(n13091), .ZN(n8661) );
  OAI21_X2 U7475 ( .B1(n11777), .B2(n12251), .A(n11006), .ZN(n11268) );
  OAI21_X2 U7476 ( .B1(n15533), .B2(n7384), .A(n7380), .ZN(n14844) );
  NAND2_X2 U7477 ( .A1(n11491), .A2(n7765), .ZN(n11541) );
  NAND4_X2 U7478 ( .A1(n9272), .A2(n9270), .A3(n9271), .A4(n9273), .ZN(n13673)
         );
  NAND2_X2 U7479 ( .A1(n8072), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n8077) );
  AND3_X1 U7480 ( .A1(n10576), .A2(n12194), .A3(n12189), .ZN(n6670) );
  AND3_X1 U7481 ( .A1(n10576), .A2(n12194), .A3(n12189), .ZN(n15077) );
  NOR2_X2 U7482 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7909) );
  INV_X2 U7483 ( .A(n15366), .ZN(n11094) );
  XNOR2_X2 U7484 ( .A(n10054), .B(n10053), .ZN(n10210) );
  AOI21_X2 U7485 ( .B1(n10255), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15227), .ZN(
        n15246) );
  INV_X1 U7487 ( .A(n10593), .ZN(n12052) );
  OAI21_X2 U7488 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8874), .A(n15696), .ZN(
        n15688) );
  INV_X4 U7489 ( .A(n10683), .ZN(n12990) );
  AOI21_X2 U7490 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10331), .A(n10319), .ZN(
        n10298) );
  NOR2_X2 U7491 ( .A1(n8876), .A2(n15686), .ZN(n8879) );
  AOI21_X2 U7492 ( .B1(n6852), .B2(n6747), .A(n6694), .ZN(n8909) );
  NOR2_X2 U7493 ( .A1(n8909), .A2(n8908), .ZN(n14808) );
  NAND2_X1 U7494 ( .A1(n13525), .A2(n6748), .ZN(n13618) );
  NAND3_X1 U7495 ( .A1(n12867), .A2(n6927), .A3(n13161), .ZN(n12791) );
  OAI22_X1 U7496 ( .A1(n6720), .A2(n12325), .B1(n12327), .B2(n7588), .ZN(
        n12330) );
  AOI21_X1 U7497 ( .B1(n13468), .B2(n9705), .A(n9704), .ZN(n9706) );
  AOI21_X1 U7498 ( .B1(n8782), .B2(n12904), .A(n6813), .ZN(n7711) );
  NAND2_X1 U7499 ( .A1(n8780), .A2(n8779), .ZN(n8782) );
  NAND2_X1 U7500 ( .A1(n13608), .A2(n6997), .ZN(n13481) );
  AND2_X1 U7501 ( .A1(n12681), .A2(n12680), .ZN(n14945) );
  NOR2_X1 U7502 ( .A1(n13705), .A2(n13704), .ZN(n13714) );
  NAND2_X1 U7503 ( .A1(n14508), .A2(n7320), .ZN(n14509) );
  XNOR2_X1 U7504 ( .A(n7333), .B(n13718), .ZN(n13704) );
  OAI211_X1 U7505 ( .C1(n13577), .C2(n9653), .A(n6994), .B(n9658), .ZN(n13635)
         );
  NAND2_X1 U7506 ( .A1(n11962), .A2(n6754), .ZN(n12630) );
  NAND2_X1 U7507 ( .A1(n7905), .A2(n7904), .ZN(n14022) );
  NAND2_X1 U7508 ( .A1(n11781), .A2(n11780), .ZN(n11962) );
  NOR2_X1 U7509 ( .A1(n14805), .A2(n14804), .ZN(n14803) );
  NAND3_X1 U7510 ( .A1(n7675), .A2(n7674), .A3(n11028), .ZN(n11491) );
  AOI21_X1 U7511 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n11106), .A(n11099), .ZN(
        n15262) );
  NAND2_X2 U7513 ( .A1(n12485), .A2(n12486), .ZN(n15540) );
  INV_X1 U7514 ( .A(n11057), .ZN(n10727) );
  CLKBUF_X3 U7515 ( .A(n9826), .Z(n9954) );
  INV_X1 U7516 ( .A(n13671), .ZN(n6907) );
  CLKBUF_X2 U7517 ( .A(P2_U3947), .Z(n6675) );
  XNOR2_X1 U7518 ( .A(n14269), .B(n11397), .ZN(n12220) );
  INV_X2 U7519 ( .A(n6688), .ZN(n9826) );
  INV_X2 U7520 ( .A(n12587), .ZN(n12578) );
  CLKBUF_X2 U7521 ( .A(n9963), .Z(n6676) );
  BUF_X2 U7522 ( .A(n9437), .Z(n9420) );
  CLKBUF_X2 U7523 ( .A(n8254), .Z(n10876) );
  CLKBUF_X2 U7524 ( .A(n9411), .Z(n9496) );
  CLKBUF_X2 U7525 ( .A(n9278), .Z(n9327) );
  CLKBUF_X2 U7526 ( .A(n9753), .Z(n6685) );
  INV_X2 U7527 ( .A(n8224), .ZN(n8516) );
  BUF_X2 U7528 ( .A(n8262), .Z(n12415) );
  INV_X1 U7529 ( .A(n12213), .ZN(n15148) );
  OAI21_X1 U7531 ( .B1(n8674), .B2(n7722), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8198) );
  NAND2_X1 U7532 ( .A1(n7104), .A2(n7101), .ZN(n10779) );
  AND3_X1 U7533 ( .A1(n7669), .A2(n10196), .A3(n7670), .ZN(n7309) );
  INV_X1 U7534 ( .A(n10093), .ZN(n7669) );
  INV_X1 U7535 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8063) );
  OR2_X1 U7537 ( .A1(n12367), .A2(n6808), .ZN(n12369) );
  OR2_X1 U7538 ( .A1(n13373), .A2(n8704), .ZN(n6940) );
  OR2_X1 U7539 ( .A1(n13376), .A2(n8704), .ZN(n7378) );
  AOI21_X1 U7540 ( .B1(n12446), .B2(n12445), .A(n12600), .ZN(n6897) );
  XNOR2_X1 U7541 ( .A(n6874), .B(n10010), .ZN(n13744) );
  NAND2_X1 U7542 ( .A1(n13765), .A2(n13764), .ZN(n13763) );
  AND2_X1 U7543 ( .A1(n7592), .A2(n7590), .ZN(n14680) );
  NAND2_X1 U7544 ( .A1(n13755), .A2(n9495), .ZN(n6874) );
  NAND2_X1 U7545 ( .A1(n8611), .A2(n6941), .ZN(n13084) );
  AND2_X1 U7546 ( .A1(n7035), .A2(n15612), .ZN(n13104) );
  NAND2_X1 U7547 ( .A1(n7712), .A2(n7711), .ZN(n12867) );
  NAND2_X1 U7548 ( .A1(n8216), .A2(n8215), .ZN(n13078) );
  NOR2_X1 U7549 ( .A1(n13804), .A2(n6779), .ZN(n6879) );
  NAND2_X1 U7550 ( .A1(n13142), .A2(n13149), .ZN(n13126) );
  NAND2_X1 U7551 ( .A1(n13822), .A2(n9469), .ZN(n13804) );
  NAND2_X1 U7552 ( .A1(n7680), .A2(n6750), .ZN(n14146) );
  NAND2_X1 U7553 ( .A1(n14231), .A2(n14230), .ZN(n7680) );
  NAND2_X1 U7554 ( .A1(n14503), .A2(n14514), .ZN(n14502) );
  AND2_X1 U7555 ( .A1(n9701), .A2(n9700), .ZN(n13468) );
  NAND2_X1 U7556 ( .A1(n9690), .A2(n6749), .ZN(n13506) );
  NAND2_X1 U7557 ( .A1(n14809), .A2(n14807), .ZN(n14786) );
  NAND2_X1 U7558 ( .A1(n13882), .A2(n9432), .ZN(n9434) );
  OAI21_X1 U7559 ( .B1(n8657), .B2(n7375), .A(n7373), .ZN(n6875) );
  NAND2_X1 U7560 ( .A1(n13481), .A2(n9685), .ZN(n13571) );
  NAND2_X1 U7561 ( .A1(n6876), .A2(n12547), .ZN(n8657) );
  NAND2_X1 U7562 ( .A1(n6974), .A2(n6972), .ZN(n14540) );
  NOR2_X1 U7563 ( .A1(n14945), .A2(n14944), .ZN(n12686) );
  NAND2_X1 U7564 ( .A1(n8180), .A2(n6899), .ZN(n8586) );
  AOI21_X1 U7565 ( .B1(n12377), .B2(n8061), .A(n7880), .ZN(n14050) );
  INV_X1 U7566 ( .A(n12911), .ZN(n6925) );
  OR2_X1 U7567 ( .A1(n11948), .A2(n7149), .ZN(n7145) );
  OR2_X1 U7568 ( .A1(n15299), .A2(n7334), .ZN(n7333) );
  OAI21_X1 U7569 ( .B1(n8545), .B2(n7416), .A(n7414), .ZN(n8178) );
  NAND2_X1 U7570 ( .A1(n8176), .A2(n8175), .ZN(n8545) );
  NAND2_X1 U7571 ( .A1(n6978), .A2(n6977), .ZN(n14735) );
  NAND2_X1 U7572 ( .A1(n8052), .A2(n8051), .ZN(n13986) );
  NAND2_X1 U7573 ( .A1(n11720), .A2(n11719), .ZN(n11913) );
  NAND2_X1 U7574 ( .A1(n6892), .A2(n6891), .ZN(n8176) );
  OR2_X1 U7575 ( .A1(n14887), .A2(n14888), .ZN(n14885) );
  NAND2_X1 U7576 ( .A1(n13635), .A2(n13634), .ZN(n13633) );
  OR2_X1 U7577 ( .A1(n6893), .A2(n6890), .ZN(n6892) );
  OR2_X1 U7578 ( .A1(n11604), .A2(n9358), .ZN(n9360) );
  NAND2_X1 U7579 ( .A1(n7144), .A2(n11474), .ZN(n11674) );
  NAND2_X1 U7580 ( .A1(n13514), .A2(n6757), .ZN(n13577) );
  NAND2_X1 U7581 ( .A1(n8173), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6894) );
  OR2_X1 U7582 ( .A1(n11710), .A2(n11719), .ZN(n6983) );
  NAND2_X1 U7583 ( .A1(n14188), .A2(n12636), .ZN(n14135) );
  OAI21_X1 U7584 ( .B1(n11468), .B2(n7285), .A(n6736), .ZN(n7144) );
  NAND2_X1 U7585 ( .A1(n12630), .A2(n6734), .ZN(n14188) );
  INV_X1 U7586 ( .A(n15026), .ZN(n7519) );
  NAND2_X1 U7587 ( .A1(n8897), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7518) );
  OAI21_X1 U7588 ( .B1(n11644), .B2(n8651), .A(n12498), .ZN(n15533) );
  NAND2_X1 U7589 ( .A1(n6996), .A2(n6995), .ZN(n11618) );
  NAND2_X1 U7590 ( .A1(n8017), .A2(n8016), .ZN(n13959) );
  NAND2_X1 U7591 ( .A1(n11923), .A2(n11922), .ZN(n14416) );
  NAND2_X1 U7592 ( .A1(n11414), .A2(n7728), .ZN(n6996) );
  NAND2_X1 U7593 ( .A1(n8000), .A2(n7999), .ZN(n14889) );
  AOI21_X1 U7594 ( .B1(n13079), .B2(n8619), .A(n8221), .ZN(n13091) );
  OAI21_X1 U7595 ( .B1(n7423), .B2(n6948), .A(n6946), .ZN(n14847) );
  NAND2_X1 U7596 ( .A1(n7004), .A2(n9615), .ZN(n11414) );
  AND2_X1 U7597 ( .A1(n11532), .A2(n15205), .ZN(n11534) );
  OAI211_X1 U7598 ( .C1(n7735), .C2(n6985), .A(n10866), .B(n6984), .ZN(n10864)
         );
  NAND2_X1 U7599 ( .A1(n6935), .A2(n7673), .ZN(n7675) );
  NAND2_X1 U7600 ( .A1(n7975), .A2(n7974), .ZN(n11737) );
  NAND2_X1 U7601 ( .A1(n15262), .A2(n15261), .ZN(n15260) );
  INV_X2 U7602 ( .A(n15623), .ZN(n15625) );
  OAI21_X1 U7603 ( .B1(n7977), .B2(n7064), .A(n7061), .ZN(n7989) );
  NAND2_X1 U7604 ( .A1(n14458), .A2(n14648), .ZN(n15103) );
  NAND2_X1 U7605 ( .A1(n6902), .A2(n8156), .ZN(n8157) );
  NOR2_X1 U7606 ( .A1(n14203), .A2(n15097), .ZN(n14960) );
  INV_X2 U7607 ( .A(n13963), .ZN(n6674) );
  INV_X2 U7608 ( .A(n11545), .ZN(n10604) );
  NAND2_X1 U7609 ( .A1(n15689), .A2(n8881), .ZN(n8884) );
  AND2_X1 U7610 ( .A1(n10925), .A2(n10924), .ZN(n12234) );
  AND2_X1 U7611 ( .A1(n10971), .A2(n10970), .ZN(n15180) );
  XNOR2_X1 U7612 ( .A(n7959), .B(n7958), .ZN(n10993) );
  INV_X1 U7613 ( .A(n6708), .ZN(n11778) );
  OAI22_X1 U7614 ( .A1(n10794), .A2(n10795), .B1(n10772), .B2(n10780), .ZN(
        n11143) );
  NAND2_X1 U7615 ( .A1(n7018), .A2(n8255), .ZN(n10557) );
  CLKBUF_X3 U7616 ( .A(n12240), .Z(n6682) );
  NAND4_X1 U7617 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n13672)
         );
  NAND3_X1 U7618 ( .A1(n8246), .A2(n8247), .A3(n6885), .ZN(n15608) );
  INV_X1 U7619 ( .A(n10888), .ZN(n10887) );
  BUF_X2 U7620 ( .A(n9963), .Z(n6688) );
  NAND4_X1 U7621 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(n9756)
         );
  XNOR2_X1 U7622 ( .A(n8826), .B(n7097), .ZN(n8877) );
  CLKBUF_X3 U7623 ( .A(n9327), .Z(n9559) );
  AND2_X2 U7624 ( .A1(n12606), .A2(n12449), .ZN(n12587) );
  NAND2_X1 U7625 ( .A1(n9503), .A2(n13726), .ZN(n9580) );
  OR2_X1 U7626 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  BUF_X2 U7627 ( .A(n9280), .Z(n9437) );
  OR2_X1 U7628 ( .A1(n7921), .A2(n10594), .ZN(n7913) );
  INV_X2 U7629 ( .A(n7921), .ZN(n8061) );
  NAND2_X1 U7630 ( .A1(n7098), .A2(n8825), .ZN(n8826) );
  BUF_X2 U7631 ( .A(n9281), .Z(n9403) );
  NAND2_X1 U7632 ( .A1(n8208), .A2(n13437), .ZN(n8254) );
  XNOR2_X1 U7633 ( .A(n10192), .B(n10191), .ZN(n12194) );
  NOR2_X1 U7634 ( .A1(n15698), .A2(n15697), .ZN(n8874) );
  INV_X1 U7635 ( .A(n14401), .ZN(n14527) );
  OR2_X1 U7636 ( .A1(n10336), .A2(n10335), .ZN(n7337) );
  XNOR2_X1 U7637 ( .A(n8067), .B(n7869), .ZN(n9753) );
  AND2_X1 U7638 ( .A1(n7520), .A2(n6786), .ZN(n15698) );
  INV_X1 U7639 ( .A(n8122), .ZN(n9993) );
  OR2_X1 U7640 ( .A1(n14792), .A2(n14791), .ZN(n7520) );
  AND2_X1 U7641 ( .A1(n6993), .A2(n8065), .ZN(n7036) );
  CLKBUF_X1 U7642 ( .A(n8635), .Z(n12382) );
  NAND2_X1 U7643 ( .A1(n8066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8067) );
  NOR2_X1 U7644 ( .A1(n15244), .A2(n7338), .ZN(n10336) );
  NOR2_X2 U7645 ( .A1(n12186), .A2(n10577), .ZN(n14401) );
  OR2_X1 U7646 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  NAND2_X1 U7647 ( .A1(n10063), .A2(n10195), .ZN(n14781) );
  INV_X1 U7648 ( .A(n10581), .ZN(n14767) );
  XNOR2_X1 U7649 ( .A(n8198), .B(n8196), .ZN(n8636) );
  XNOR2_X1 U7650 ( .A(n8871), .B(n8870), .ZN(n14792) );
  NAND2_X1 U7651 ( .A1(n7740), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8036) );
  XNOR2_X1 U7652 ( .A(n8206), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U7653 ( .A1(n8064), .A2(n8063), .ZN(n8066) );
  OR3_X1 U7654 ( .A1(n8064), .A2(n14085), .A3(n8063), .ZN(n6993) );
  NAND2_X1 U7655 ( .A1(n13428), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U7656 ( .A(n7557), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10581) );
  AND2_X1 U7657 ( .A1(n8022), .A2(n6802), .ZN(n8064) );
  OR2_X1 U7658 ( .A1(n8205), .A2(n8478), .ZN(n8206) );
  NOR2_X1 U7659 ( .A1(n7681), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U7660 ( .A1(n15700), .A2(n8867), .ZN(n8871) );
  AND3_X1 U7661 ( .A1(n7386), .A2(n8201), .A3(n8476), .ZN(n8205) );
  NAND2_X1 U7662 ( .A1(n7031), .A2(n8132), .ZN(n8249) );
  AND2_X1 U7663 ( .A1(n7387), .A2(n6805), .ZN(n7386) );
  INV_X1 U7664 ( .A(n6859), .ZN(n8013) );
  INV_X1 U7665 ( .A(n10061), .ZN(n7311) );
  NAND2_X1 U7666 ( .A1(n8820), .A2(n7086), .ZN(n8869) );
  AND2_X1 U7667 ( .A1(n7593), .A2(n10062), .ZN(n7308) );
  NOR2_X1 U7668 ( .A1(n7388), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7387) );
  AND3_X1 U7669 ( .A1(n7668), .A2(n7667), .A3(n7669), .ZN(n10431) );
  NAND4_X1 U7670 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10061) );
  AND2_X1 U7671 ( .A1(n7016), .A2(n8358), .ZN(n7217) );
  AND2_X1 U7672 ( .A1(n8136), .A2(n8135), .ZN(n8259) );
  NOR2_X1 U7673 ( .A1(n7672), .A2(n7671), .ZN(n7667) );
  AND2_X1 U7674 ( .A1(n7739), .A2(n7738), .ZN(n7737) );
  AND3_X1 U7675 ( .A1(n7686), .A2(n12177), .A3(n10191), .ZN(n10059) );
  AND2_X1 U7676 ( .A1(n8021), .A2(n8028), .ZN(n7739) );
  NAND2_X1 U7677 ( .A1(n10050), .A2(n7686), .ZN(n7685) );
  AND4_X1 U7678 ( .A1(n8362), .A2(n8428), .A3(n8359), .A4(n8342), .ZN(n7713)
         );
  AND4_X1 U7679 ( .A1(n10048), .A2(n10173), .A3(n10049), .A4(n10043), .ZN(
        n7668) );
  AND2_X1 U7680 ( .A1(n8189), .A2(n8192), .ZN(n7218) );
  AND2_X1 U7681 ( .A1(n7863), .A2(n7865), .ZN(n6987) );
  AND2_X1 U7682 ( .A1(n6991), .A2(n6992), .ZN(n6861) );
  NAND4_X1 U7683 ( .A1(n10046), .A2(n10106), .A3(n10045), .A4(n10044), .ZN(
        n7672) );
  NAND2_X1 U7684 ( .A1(n8103), .A2(n7640), .ZN(n7639) );
  INV_X1 U7685 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10177) );
  INV_X1 U7686 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8114) );
  INV_X1 U7687 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8103) );
  INV_X1 U7688 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8069) );
  INV_X1 U7689 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7990) );
  INV_X1 U7690 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7640) );
  NOR2_X1 U7691 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7867) );
  INV_X1 U7692 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7869) );
  INV_X1 U7693 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8428) );
  INV_X4 U7694 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7695 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n6926) );
  INV_X1 U7696 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13731) );
  INV_X1 U7697 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8362) );
  INV_X1 U7698 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8342) );
  INV_X1 U7699 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8359) );
  INV_X1 U7700 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8190) );
  NOR2_X1 U7701 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8189) );
  NOR2_X1 U7702 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6991) );
  NOR2_X1 U7703 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6992) );
  INV_X1 U7704 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10141) );
  INV_X1 U7705 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8195) );
  INV_X1 U7706 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7724) );
  NOR2_X1 U7707 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n6961) );
  NOR2_X1 U7708 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n6960) );
  INV_X4 U7709 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7710 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10106) );
  INV_X1 U7711 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10043) );
  INV_X1 U7712 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8284) );
  INV_X1 U7713 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10046) );
  INV_X1 U7714 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10049) );
  INV_X1 U7715 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10045) );
  OR2_X1 U7716 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  NOR2_X1 U7717 ( .A1(n10647), .A2(n10648), .ZN(n10646) );
  NAND4_X2 U7718 ( .A1(n6861), .A2(n6988), .A3(n6987), .A4(n6860), .ZN(n6859)
         );
  INV_X1 U7719 ( .A(n10419), .ZN(n10424) );
  NAND2_X2 U7720 ( .A1(n9580), .A2(n9579), .ZN(n6683) );
  NAND2_X1 U7721 ( .A1(n9580), .A2(n9579), .ZN(n6684) );
  NAND4_X2 U7722 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n15587)
         );
  AOI211_X1 U7723 ( .C1(n10298), .C2(n10297), .A(n15298), .B(n10296), .ZN(
        n10307) );
  OAI211_X1 U7724 ( .C1(n7651), .C2(n7646), .A(n7750), .B(n7644), .ZN(n11781)
         );
  AOI22_X2 U7725 ( .A1(n13771), .A2(n13770), .B1(n9555), .B2(n13980), .ZN(
        n13765) );
  AND2_X1 U7726 ( .A1(n12378), .A2(n14767), .ZN(n6677) );
  INV_X4 U7727 ( .A(n6669), .ZN(n6678) );
  OAI222_X1 U7729 ( .A1(n12189), .A2(P1_U3086), .B1(n14775), .B2(n11525), .C1(
        n12062), .C2(n14772), .ZN(P1_U3335) );
  AND2_X1 U7730 ( .A1(n10570), .A2(n12189), .ZN(n12214) );
  AND2_X4 U7731 ( .A1(n10575), .A2(n12214), .ZN(n11545) );
  NOR2_X2 U7732 ( .A1(n13933), .A2(n14031), .ZN(n13915) );
  OR2_X2 U7733 ( .A1(n13953), .A2(n13936), .ZN(n13933) );
  AND2_X1 U7734 ( .A1(n10582), .A2(n14767), .ZN(n6679) );
  AND2_X1 U7735 ( .A1(n10582), .A2(n14767), .ZN(n6680) );
  BUF_X4 U7736 ( .A(n9585), .Z(n6681) );
  NAND2_X1 U7737 ( .A1(n9576), .A2(n13726), .ZN(n9585) );
  AOI21_X2 U7738 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n8896), .A(n14803), .ZN(
        n15027) );
  MUX2_X1 U7739 ( .A(n12189), .B(n10570), .S(n12193), .Z(n12240) );
  NOR2_X2 U7740 ( .A1(n15609), .A2(n10664), .ZN(n10413) );
  XNOR2_X2 U7741 ( .A(n7925), .B(n7924), .ZN(n10892) );
  INV_X1 U7742 ( .A(n8059), .ZN(n6686) );
  NAND2_X2 U7743 ( .A1(n6667), .A2(n10593), .ZN(n8059) );
  NOR2_X2 U7744 ( .A1(n9752), .A2(n9993), .ZN(n9578) );
  OAI21_X2 U7745 ( .B1(n11815), .B2(n9531), .A(n9530), .ZN(n14879) );
  OAI22_X2 U7746 ( .A1(n11788), .A2(n9529), .B1(n9989), .B2(n11795), .ZN(
        n11815) );
  NAND2_X1 U7748 ( .A1(n10461), .A2(n6685), .ZN(n9963) );
  AND2_X1 U7749 ( .A1(n9923), .A2(n9924), .ZN(n7612) );
  NAND2_X1 U7750 ( .A1(n7495), .A2(n7493), .ZN(n14595) );
  AOI21_X1 U7751 ( .B1(n7496), .B2(n7497), .A(n7494), .ZN(n7493) );
  NAND2_X1 U7752 ( .A1(n14732), .A2(n7496), .ZN(n7495) );
  AOI21_X1 U7753 ( .B1(n12923), .B2(n7702), .A(n8793), .ZN(n7701) );
  INV_X1 U7754 ( .A(n13207), .ZN(n6876) );
  INV_X1 U7755 ( .A(n13649), .ZN(n13448) );
  AND2_X1 U7756 ( .A1(n13482), .A2(n9681), .ZN(n6997) );
  NAND2_X1 U7757 ( .A1(n7598), .A2(n12264), .ZN(n7597) );
  INV_X1 U7758 ( .A(n12296), .ZN(n7012) );
  OAI21_X1 U7759 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9883) );
  AND2_X1 U7760 ( .A1(n7609), .A2(n9933), .ZN(n7604) );
  NAND2_X1 U7761 ( .A1(n7608), .A2(n7613), .ZN(n7607) );
  NOR2_X1 U7762 ( .A1(n7254), .A2(n7253), .ZN(n7252) );
  NOR2_X1 U7763 ( .A1(n7807), .A2(n7255), .ZN(n7253) );
  INV_X1 U7764 ( .A(n7546), .ZN(n7254) );
  AND2_X1 U7765 ( .A1(n13986), .A2(n13649), .ZN(n9479) );
  AND2_X1 U7766 ( .A1(n7638), .A2(n7757), .ZN(n6858) );
  NOR2_X1 U7767 ( .A1(n7639), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U7768 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  AOI21_X1 U7769 ( .B1(n7548), .B2(n7813), .A(n7547), .ZN(n7546) );
  INV_X1 U7770 ( .A(n7550), .ZN(n7548) );
  INV_X1 U7771 ( .A(n8011), .ZN(n7547) );
  AND2_X1 U7772 ( .A1(n7294), .A2(n7782), .ZN(n7129) );
  INV_X1 U7773 ( .A(n8767), .ZN(n6924) );
  NAND2_X1 U7774 ( .A1(n12830), .A2(n8778), .ZN(n8780) );
  NAND2_X1 U7775 ( .A1(n12589), .A2(n12584), .ZN(n7034) );
  NOR2_X1 U7776 ( .A1(n13076), .A2(n7434), .ZN(n7433) );
  INV_X1 U7777 ( .A(n8625), .ZN(n7434) );
  INV_X1 U7778 ( .A(n12569), .ZN(n7371) );
  INV_X1 U7779 ( .A(n7370), .ZN(n7369) );
  OAI21_X1 U7780 ( .B1(n8659), .B2(n7371), .A(n12572), .ZN(n7370) );
  OR2_X1 U7781 ( .A1(n13306), .A2(n13090), .ZN(n12579) );
  OR2_X1 U7782 ( .A1(n13179), .A2(n13162), .ZN(n12555) );
  NAND2_X1 U7783 ( .A1(n13217), .A2(n8503), .ZN(n13199) );
  NOR2_X1 U7784 ( .A1(n8479), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7213) );
  NOR2_X1 U7785 ( .A1(n7485), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n6880) );
  AND2_X1 U7786 ( .A1(n8191), .A2(n8190), .ZN(n7016) );
  NOR2_X1 U7787 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8191) );
  NOR2_X1 U7788 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8192) );
  NAND2_X1 U7789 ( .A1(n13827), .A2(n7352), .ZN(n7355) );
  NOR2_X1 U7790 ( .A1(n7353), .A2(n13980), .ZN(n7352) );
  INV_X1 U7791 ( .A(n7354), .ZN(n7353) );
  NOR2_X1 U7792 ( .A1(n13855), .A2(n7278), .ZN(n7277) );
  INV_X1 U7793 ( .A(n9548), .ZN(n7278) );
  AND2_X2 U7794 ( .A1(n10895), .A2(n10575), .ZN(n11546) );
  NAND2_X1 U7795 ( .A1(n14502), .A2(n14446), .ZN(n14484) );
  NAND2_X1 U7796 ( .A1(n14574), .A2(n14440), .ZN(n7516) );
  INV_X1 U7797 ( .A(n7148), .ZN(n7146) );
  OAI21_X1 U7798 ( .B1(n7580), .B2(n7149), .A(n14652), .ZN(n7148) );
  NAND2_X1 U7799 ( .A1(n14735), .A2(n7748), .ZN(n14732) );
  AOI21_X1 U7800 ( .B1(n6709), .B2(n12279), .A(n11932), .ZN(n14433) );
  NAND2_X1 U7801 ( .A1(n7856), .A2(n7855), .ZN(n7879) );
  NAND2_X1 U7802 ( .A1(n7847), .A2(n7846), .ZN(n7884) );
  OAI21_X1 U7803 ( .B1(n8050), .B2(n11728), .A(n7845), .ZN(n7847) );
  NAND2_X1 U7804 ( .A1(n7248), .A2(n10564), .ZN(n7073) );
  AND2_X1 U7805 ( .A1(n7072), .A2(n7075), .ZN(n7071) );
  OR2_X1 U7806 ( .A1(n7248), .A2(n10564), .ZN(n7075) );
  NAND2_X1 U7807 ( .A1(n8033), .A2(n7824), .ZN(n7072) );
  OAI21_X1 U7808 ( .B1(n8027), .B2(n7551), .A(n7820), .ZN(n8034) );
  INV_X1 U7809 ( .A(n8026), .ZN(n7551) );
  XNOR2_X1 U7810 ( .A(n7819), .B(SI_18_), .ZN(n8027) );
  INV_X1 U7811 ( .A(n7671), .ZN(n7670) );
  INV_X1 U7812 ( .A(n7672), .ZN(n7593) );
  NAND2_X1 U7813 ( .A1(n7539), .A2(n7538), .ZN(n7977) );
  AOI21_X1 U7814 ( .B1(n7541), .B2(n7543), .A(n6775), .ZN(n7538) );
  AOI21_X1 U7815 ( .B1(n8882), .B2(n8828), .A(n6849), .ZN(n8830) );
  AND2_X1 U7816 ( .A1(n8829), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6849) );
  AOI21_X1 U7817 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n8841), .A(n8840), .ZN(
        n8901) );
  AOI21_X1 U7818 ( .B1(n7701), .B2(n7703), .A(n7700), .ZN(n7699) );
  INV_X1 U7819 ( .A(n8794), .ZN(n7700) );
  OAI21_X1 U7820 ( .B1(n13425), .B2(n12444), .A(n8723), .ZN(n8728) );
  INV_X1 U7821 ( .A(n13116), .ZN(n13090) );
  OR2_X1 U7822 ( .A1(n10848), .A2(n7715), .ZN(n7718) );
  INV_X1 U7823 ( .A(n8733), .ZN(n7715) );
  NAND2_X1 U7824 ( .A1(n11082), .A2(n6710), .ZN(n7230) );
  OR2_X1 U7825 ( .A1(n11589), .A2(n8746), .ZN(n8748) );
  AND2_X1 U7826 ( .A1(n8387), .A2(n8386), .ZN(n12507) );
  NAND2_X1 U7827 ( .A1(n12791), .A2(n12867), .ZN(n8786) );
  OAI21_X1 U7828 ( .B1(n11859), .B2(n7222), .A(n7219), .ZN(n8756) );
  NAND2_X1 U7829 ( .A1(n7707), .A2(n7223), .ZN(n7222) );
  AND2_X1 U7830 ( .A1(n7704), .A2(n7220), .ZN(n7219) );
  NAND2_X1 U7831 ( .A1(n7707), .A2(n7221), .ZN(n7220) );
  INV_X1 U7832 ( .A(n8243), .ZN(n8619) );
  OR2_X1 U7833 ( .A1(n8243), .A2(n15619), .ZN(n8226) );
  OAI21_X1 U7834 ( .B1(n10796), .B2(n11306), .A(n10776), .ZN(n7478) );
  NAND2_X1 U7835 ( .A1(n11567), .A2(n11568), .ZN(n11896) );
  OR2_X1 U7836 ( .A1(n14819), .A2(n14820), .ZN(n7119) );
  NAND2_X1 U7837 ( .A1(n6943), .A2(n13076), .ZN(n13071) );
  NAND2_X1 U7838 ( .A1(n13084), .A2(n8625), .ZN(n6943) );
  NAND2_X1 U7839 ( .A1(n13089), .A2(n13088), .ZN(n13087) );
  OR2_X1 U7840 ( .A1(n8589), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U7841 ( .A1(n13112), .A2(n8596), .ZN(n13103) );
  NAND2_X1 U7842 ( .A1(n13131), .A2(n8584), .ZN(n13114) );
  NOR2_X1 U7843 ( .A1(n8502), .A2(n7365), .ZN(n7364) );
  INV_X1 U7844 ( .A(n12535), .ZN(n7365) );
  NAND2_X1 U7845 ( .A1(n6878), .A2(n6877), .ZN(n7372) );
  AND2_X1 U7846 ( .A1(n8653), .A2(n12511), .ZN(n6877) );
  OAI21_X1 U7847 ( .B1(n12472), .B2(n6857), .A(n11499), .ZN(n6856) );
  NOR2_X1 U7848 ( .A1(n15551), .A2(n6857), .ZN(n6854) );
  INV_X1 U7849 ( .A(n12447), .ZN(n6857) );
  NAND3_X1 U7850 ( .A1(n10681), .A2(n10693), .A3(n12587), .ZN(n15590) );
  AND3_X1 U7851 ( .A1(n8233), .A2(n8232), .A3(n8231), .ZN(n15606) );
  INV_X1 U7852 ( .A(n12415), .ZN(n8510) );
  INV_X1 U7853 ( .A(n8261), .ZN(n12417) );
  NAND2_X1 U7854 ( .A1(n8680), .A2(n8682), .ZN(n10136) );
  AOI21_X1 U7855 ( .B1(n7411), .B2(n6707), .A(n6839), .ZN(n12408) );
  OR2_X1 U7856 ( .A1(n8613), .A2(n8185), .ZN(n8187) );
  XNOR2_X1 U7857 ( .A(n8197), .B(n8201), .ZN(n8635) );
  OR2_X1 U7858 ( .A1(n8202), .A2(n8478), .ZN(n8197) );
  AND2_X1 U7859 ( .A1(n7386), .A2(n8476), .ZN(n8202) );
  INV_X1 U7860 ( .A(n7394), .ZN(n7393) );
  OAI21_X1 U7861 ( .B1(n8457), .B2(n7395), .A(n8472), .ZN(n7394) );
  OR2_X1 U7862 ( .A1(n8442), .A2(n8441), .ZN(n8444) );
  AND2_X1 U7863 ( .A1(n8147), .A2(n8146), .ZN(n8330) );
  INV_X1 U7864 ( .A(n7404), .ZN(n7403) );
  OAI21_X1 U7865 ( .B1(n8141), .B2(n7405), .A(n8143), .ZN(n7404) );
  NAND2_X1 U7866 ( .A1(n9722), .A2(n9723), .ZN(n9728) );
  XNOR2_X1 U7867 ( .A(n6684), .B(n10727), .ZN(n9599) );
  NAND2_X1 U7868 ( .A1(n9670), .A2(n13545), .ZN(n13548) );
  NAND2_X1 U7869 ( .A1(n13738), .A2(n14050), .ZN(n13737) );
  NAND2_X1 U7870 ( .A1(n13977), .A2(n7751), .ZN(n13757) );
  OR2_X1 U7871 ( .A1(n13456), .A2(n9555), .ZN(n7751) );
  OR2_X1 U7872 ( .A1(n9554), .A2(n7553), .ZN(n7552) );
  AOI21_X1 U7873 ( .B1(n13856), .B2(n7436), .A(n7435), .ZN(n13822) );
  AND3_X1 U7874 ( .A1(n13823), .A2(n6723), .A3(n7437), .ZN(n7435) );
  NAND2_X1 U7875 ( .A1(n13815), .A2(n9553), .ZN(n13797) );
  NOR2_X1 U7876 ( .A1(n13923), .A2(n7453), .ZN(n7452) );
  INV_X1 U7877 ( .A(n9410), .ZN(n7453) );
  NAND2_X1 U7878 ( .A1(n13932), .A2(n13931), .ZN(n13930) );
  NAND2_X1 U7879 ( .A1(n11992), .A2(n7454), .ZN(n13945) );
  AND2_X1 U7880 ( .A1(n13947), .A2(n9392), .ZN(n7454) );
  NAND2_X1 U7881 ( .A1(n10420), .A2(n10419), .ZN(n9287) );
  NAND2_X1 U7882 ( .A1(n7877), .A2(n7876), .ZN(n9982) );
  AOI21_X1 U7883 ( .B1(n7657), .B2(n7660), .A(n7656), .ZN(n7655) );
  INV_X1 U7884 ( .A(n14182), .ZN(n7656) );
  INV_X1 U7885 ( .A(n7657), .ZN(n6932) );
  AND2_X1 U7886 ( .A1(n10626), .A2(n10625), .ZN(n11224) );
  NAND2_X1 U7887 ( .A1(n14433), .A2(n7582), .ZN(n6978) );
  NAND2_X1 U7888 ( .A1(n7143), .A2(n7287), .ZN(n11720) );
  AOI21_X1 U7889 ( .B1(n7289), .B2(n7288), .A(n6768), .ZN(n7287) );
  NAND2_X1 U7890 ( .A1(n11674), .A2(n7289), .ZN(n7143) );
  AOI21_X1 U7891 ( .B1(n7136), .B2(n7135), .A(n7134), .ZN(n11709) );
  AND2_X1 U7892 ( .A1(n15013), .A2(n14137), .ZN(n7134) );
  NAND2_X1 U7893 ( .A1(n11658), .A2(n14260), .ZN(n7135) );
  INV_X1 U7894 ( .A(n11657), .ZN(n7136) );
  XNOR2_X1 U7895 ( .A(n12255), .B(n14263), .ZN(n12105) );
  NAND2_X1 U7896 ( .A1(n12190), .A2(n10202), .ZN(n15102) );
  NOR2_X1 U7897 ( .A1(n14471), .A2(n7173), .ZN(n7172) );
  INV_X1 U7898 ( .A(n7175), .ZN(n7173) );
  AND2_X1 U7899 ( .A1(n7594), .A2(n10193), .ZN(n6981) );
  AND3_X1 U7900 ( .A1(n10048), .A2(n10043), .A3(n10173), .ZN(n7594) );
  XNOR2_X1 U7901 ( .A(n7780), .B(n10074), .ZN(n7933) );
  AND2_X1 U7902 ( .A1(n7234), .A2(n7233), .ZN(n11589) );
  NOR2_X1 U7903 ( .A1(n11591), .A2(n11588), .ZN(n7233) );
  NAND2_X1 U7904 ( .A1(n12253), .A2(n7584), .ZN(n7583) );
  NOR2_X1 U7905 ( .A1(n7192), .A2(n7010), .ZN(n7009) );
  NOR2_X1 U7906 ( .A1(n7598), .A2(n12264), .ZN(n7010) );
  AND2_X1 U7907 ( .A1(n12266), .A2(n7193), .ZN(n7192) );
  INV_X1 U7908 ( .A(n12265), .ZN(n7193) );
  MUX2_X1 U7909 ( .A(n14261), .B(n12638), .S(n6682), .Z(n12265) );
  INV_X1 U7910 ( .A(n9799), .ZN(n7629) );
  NAND2_X1 U7911 ( .A1(n7578), .A2(n12276), .ZN(n7577) );
  NAND2_X1 U7912 ( .A1(n7044), .A2(n12295), .ZN(n12298) );
  NAND2_X1 U7913 ( .A1(n9828), .A2(n6739), .ZN(n7624) );
  AND2_X1 U7914 ( .A1(n12300), .A2(n7565), .ZN(n7564) );
  NAND2_X1 U7915 ( .A1(n7569), .A2(n7566), .ZN(n7565) );
  NAND2_X1 U7916 ( .A1(n7564), .A2(n7567), .ZN(n7563) );
  NOR2_X1 U7917 ( .A1(n7569), .A2(n7568), .ZN(n7567) );
  OAI21_X1 U7918 ( .B1(n12311), .B2(n12310), .A(n12309), .ZN(n7561) );
  NAND2_X1 U7919 ( .A1(n12336), .A2(n7181), .ZN(n7180) );
  NAND2_X1 U7920 ( .A1(n7606), .A2(n7603), .ZN(n7602) );
  INV_X1 U7921 ( .A(n7604), .ZN(n7603) );
  NAND2_X1 U7922 ( .A1(n7604), .A2(n7612), .ZN(n7599) );
  NAND2_X1 U7923 ( .A1(n7605), .A2(n7607), .ZN(n7600) );
  INV_X1 U7924 ( .A(n7808), .ZN(n7255) );
  NOR2_X1 U7925 ( .A1(n9394), .A2(n13540), .ZN(n9393) );
  INV_X1 U7926 ( .A(n7902), .ZN(n7248) );
  OAI21_X1 U7927 ( .B1(n8020), .B2(n7818), .A(n7817), .ZN(n7819) );
  INV_X1 U7928 ( .A(n8018), .ZN(n7816) );
  INV_X1 U7929 ( .A(n7813), .ZN(n7549) );
  NAND2_X1 U7930 ( .A1(n7061), .A2(n7064), .ZN(n7059) );
  NAND2_X1 U7931 ( .A1(n7252), .A2(n7255), .ZN(n7250) );
  AOI21_X1 U7932 ( .B1(n7065), .B2(n7063), .A(n7062), .ZN(n7061) );
  INV_X1 U7933 ( .A(n7805), .ZN(n7062) );
  INV_X1 U7934 ( .A(n7801), .ZN(n7063) );
  AND2_X1 U7935 ( .A1(n7779), .A2(n7781), .ZN(n7082) );
  NAND2_X1 U7936 ( .A1(n11128), .A2(n6741), .ZN(n11129) );
  NAND2_X1 U7937 ( .A1(n15496), .A2(n7121), .ZN(n11133) );
  OR2_X1 U7938 ( .A1(n11160), .A2(n11158), .ZN(n7121) );
  NAND2_X1 U7939 ( .A1(n11380), .A2(n6828), .ZN(n11563) );
  INV_X1 U7940 ( .A(n7433), .ZN(n7430) );
  OR2_X1 U7941 ( .A1(n13165), .A2(n13176), .ZN(n12560) );
  INV_X1 U7942 ( .A(n12551), .ZN(n7375) );
  OR2_X1 U7943 ( .A1(n13228), .A2(n13236), .ZN(n12539) );
  OR2_X1 U7944 ( .A1(n13418), .A2(n12894), .ZN(n12522) );
  NAND2_X1 U7945 ( .A1(n8652), .A2(n12502), .ZN(n7385) );
  INV_X1 U7946 ( .A(n8372), .ZN(n7419) );
  INV_X1 U7947 ( .A(n6715), .ZN(n6947) );
  OR2_X1 U7948 ( .A1(n15608), .A2(n15582), .ZN(n12457) );
  OR2_X1 U7949 ( .A1(n10557), .A2(n11308), .ZN(n12466) );
  NAND2_X1 U7950 ( .A1(n12457), .A2(n12458), .ZN(n12463) );
  OR2_X1 U7951 ( .A1(n15587), .A2(n15606), .ZN(n12455) );
  INV_X1 U7952 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8201) );
  INV_X1 U7953 ( .A(n7722), .ZN(n7720) );
  INV_X1 U7954 ( .A(n7417), .ZN(n7416) );
  AOI21_X1 U7955 ( .B1(n7417), .B2(n7415), .A(n6837), .ZN(n7414) );
  AOI21_X1 U7956 ( .B1(n8544), .B2(n8177), .A(n7418), .ZN(n7417) );
  NAND2_X1 U7957 ( .A1(n7213), .A2(n7212), .ZN(n8633) );
  INV_X1 U7958 ( .A(n8147), .ZN(n6887) );
  INV_X1 U7959 ( .A(n8136), .ZN(n7399) );
  INV_X1 U7960 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7107) );
  INV_X1 U7961 ( .A(n9619), .ZN(n7730) );
  INV_X1 U7962 ( .A(n7729), .ZN(n7728) );
  OAI21_X1 U7963 ( .B1(n11413), .B2(n7730), .A(n13493), .ZN(n7729) );
  AND2_X1 U7964 ( .A1(n9964), .A2(n10013), .ZN(n10015) );
  NAND2_X1 U7965 ( .A1(n14085), .A2(n7331), .ZN(n7330) );
  INV_X1 U7966 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7331) );
  AND2_X1 U7967 ( .A1(n15304), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7334) );
  OR2_X1 U7968 ( .A1(n9955), .A2(n13450), .ZN(n9556) );
  NOR2_X1 U7969 ( .A1(n13931), .A2(n7271), .ZN(n7270) );
  INV_X1 U7970 ( .A(n9536), .ZN(n7271) );
  INV_X1 U7971 ( .A(n13663), .ZN(n9989) );
  INV_X1 U7972 ( .A(n9300), .ZN(n6863) );
  XNOR2_X1 U7973 ( .A(n13672), .B(n15379), .ZN(n9994) );
  NAND2_X1 U7974 ( .A1(n7357), .A2(n7360), .ZN(n13860) );
  INV_X1 U7975 ( .A(n14010), .ZN(n7360) );
  INV_X1 U7976 ( .A(n13873), .ZN(n7357) );
  NAND2_X1 U7977 ( .A1(n6870), .A2(n9351), .ZN(n11604) );
  NOR2_X1 U7978 ( .A1(n8082), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7041) );
  INV_X1 U7979 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6916) );
  INV_X1 U7980 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6915) );
  INV_X1 U7981 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8075) );
  INV_X1 U7982 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8073) );
  INV_X1 U7983 ( .A(n10575), .ZN(n10588) );
  NOR2_X1 U7984 ( .A1(n14661), .A2(n14477), .ZN(n7318) );
  NAND2_X1 U7985 ( .A1(n14484), .A2(n14483), .ZN(n14482) );
  NOR2_X1 U7986 ( .A1(n7514), .A2(n6976), .ZN(n6975) );
  INV_X1 U7987 ( .A(n6800), .ZN(n6976) );
  NAND2_X1 U7988 ( .A1(n7161), .A2(n14426), .ZN(n7160) );
  NAND2_X1 U7989 ( .A1(n12218), .A2(n12215), .ZN(n12100) );
  NAND2_X1 U7990 ( .A1(n12100), .A2(n15085), .ZN(n15086) );
  NAND2_X1 U7991 ( .A1(n14540), .A2(n14442), .ZN(n14541) );
  AOI21_X1 U7992 ( .B1(n14537), .B2(n14544), .A(n6780), .ZN(n14530) );
  NAND2_X1 U7993 ( .A1(n14530), .A2(n14529), .ZN(n14528) );
  NAND2_X1 U7994 ( .A1(n7501), .A2(n14436), .ZN(n7497) );
  NAND2_X1 U7995 ( .A1(n6785), .A2(n14436), .ZN(n7496) );
  NAND2_X1 U7996 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  INV_X1 U7997 ( .A(n7502), .ZN(n7500) );
  AND2_X1 U7998 ( .A1(n14435), .A2(n14434), .ZN(n7502) );
  OAI21_X1 U7999 ( .B1(n15067), .B2(n6753), .A(n7489), .ZN(n6979) );
  NAND2_X1 U8000 ( .A1(n15075), .A2(n11634), .ZN(n7489) );
  OAI21_X1 U8001 ( .B1(n8054), .B2(n8053), .A(n7852), .ZN(n8058) );
  NAND2_X1 U8002 ( .A1(n7844), .A2(n7843), .ZN(n8050) );
  OR2_X1 U8003 ( .A1(n8045), .A2(n8044), .ZN(n7844) );
  INV_X1 U8004 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10047) );
  AND2_X1 U8005 ( .A1(n7809), .A2(n7811), .ZN(n7550) );
  AND2_X1 U8006 ( .A1(n7669), .A2(n7594), .ZN(n7487) );
  NAND2_X1 U8007 ( .A1(n7251), .A2(n7808), .ZN(n7997) );
  NAND2_X1 U8008 ( .A1(n7989), .A2(n7807), .ZN(n7251) );
  OR2_X1 U8009 ( .A1(n10220), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10221) );
  AOI21_X1 U8010 ( .B1(n7788), .B2(n7247), .A(n6778), .ZN(n7246) );
  INV_X1 U8011 ( .A(n7787), .ZN(n7247) );
  NAND2_X1 U8012 ( .A1(n7132), .A2(n7782), .ZN(n7131) );
  NAND2_X1 U8013 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7087), .ZN(n7086) );
  XNOR2_X1 U8014 ( .A(n9000), .B(n7085), .ZN(n8868) );
  NAND2_X1 U8015 ( .A1(n8861), .A2(n8862), .ZN(n7098) );
  NOR2_X1 U8016 ( .A1(n8831), .A2(n8832), .ZN(n8860) );
  NOR2_X1 U8017 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8886), .ZN(n8831) );
  AOI21_X1 U8018 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n8835), .A(n8834), .ZN(
        n8836) );
  NOR2_X1 U8019 ( .A1(n8893), .A2(n8892), .ZN(n8834) );
  INV_X1 U8020 ( .A(n15044), .ZN(n7528) );
  OR2_X1 U8021 ( .A1(n15047), .A2(n7529), .ZN(n7527) );
  INV_X1 U8022 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7526) );
  NOR2_X1 U8023 ( .A1(n8752), .A2(n13274), .ZN(n7708) );
  NAND2_X1 U8024 ( .A1(n7714), .A2(n6755), .ZN(n12830) );
  NAND2_X1 U8025 ( .A1(n12850), .A2(n6760), .ZN(n12857) );
  AOI21_X1 U8026 ( .B1(n8742), .B2(n8741), .A(n7759), .ZN(n8743) );
  NAND2_X1 U8027 ( .A1(n12818), .A2(n8739), .ZN(n8741) );
  NAND2_X1 U8028 ( .A1(n6710), .A2(n11081), .ZN(n7232) );
  NAND2_X1 U8029 ( .A1(n6928), .A2(n7049), .ZN(n8781) );
  INV_X1 U8030 ( .A(n8779), .ZN(n7049) );
  INV_X1 U8031 ( .A(n8780), .ZN(n6928) );
  NAND2_X1 U8032 ( .A1(n10813), .A2(n8707), .ZN(n12444) );
  XNOR2_X1 U8033 ( .A(n12423), .B(n13039), .ZN(n12602) );
  NAND2_X1 U8034 ( .A1(n7021), .A2(n6745), .ZN(n12423) );
  NAND2_X1 U8035 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  AOI21_X1 U8036 ( .B1(n13076), .B2(n7034), .A(n7032), .ZN(n12594) );
  XNOR2_X1 U8037 ( .A(n7407), .B(n13039), .ZN(n12446) );
  INV_X1 U8038 ( .A(n12595), .ZN(n7410) );
  NOR2_X1 U8039 ( .A1(n12442), .A2(n7409), .ZN(n7408) );
  OAI22_X1 U8040 ( .A1(n8243), .A2(n10852), .B1(n10876), .B2(n8268), .ZN(n7363) );
  OR2_X1 U8041 ( .A1(n8245), .A2(n7002), .ZN(n8257) );
  NOR2_X1 U8042 ( .A1(n8516), .A2(n10770), .ZN(n7019) );
  INV_X1 U8043 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8044 ( .A1(n8478), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U8045 ( .A1(n10783), .A2(n10784), .ZN(n11128) );
  XNOR2_X1 U8046 ( .A(n11129), .B(n7476), .ZN(n15444) );
  AOI21_X1 U8047 ( .B1(n7478), .B2(n7477), .A(n6729), .ZN(n11121) );
  INV_X1 U8048 ( .A(n11118), .ZN(n7477) );
  NAND2_X1 U8049 ( .A1(n7115), .A2(n7114), .ZN(n7113) );
  INV_X1 U8050 ( .A(n15450), .ZN(n7114) );
  NAND2_X1 U8051 ( .A1(n15478), .A2(n11132), .ZN(n15498) );
  NAND2_X1 U8052 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  XNOR2_X1 U8053 ( .A(n11133), .B(n11166), .ZN(n15518) );
  AOI21_X1 U8054 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15493), .A(n15484), .ZN(
        n11125) );
  NAND2_X1 U8055 ( .A1(n11135), .A2(n11136), .ZN(n11380) );
  XNOR2_X1 U8056 ( .A(n11563), .B(n11572), .ZN(n11382) );
  AOI21_X1 U8057 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11374), .A(n11373), .ZN(
        n11558) );
  NAND2_X1 U8058 ( .A1(n11896), .A2(n11897), .ZN(n12957) );
  INV_X1 U8059 ( .A(n7108), .ZN(n13002) );
  INV_X1 U8060 ( .A(n7110), .ZN(n7109) );
  AOI21_X1 U8061 ( .B1(n12954), .B2(n12968), .A(n7111), .ZN(n7110) );
  NAND2_X1 U8062 ( .A1(n7119), .A2(n6735), .ZN(n7118) );
  OR2_X1 U8063 ( .A1(n8618), .A2(n8617), .ZN(n13095) );
  INV_X1 U8064 ( .A(n6867), .ZN(n6866) );
  OAI21_X1 U8065 ( .B1(n7367), .B2(n6868), .A(n12580), .ZN(n6867) );
  INV_X1 U8066 ( .A(n12579), .ZN(n6868) );
  OR2_X1 U8067 ( .A1(n8601), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8616) );
  AOI21_X1 U8068 ( .B1(n7369), .B2(n7371), .A(n7368), .ZN(n7367) );
  INV_X1 U8069 ( .A(n12575), .ZN(n7368) );
  NAND2_X1 U8070 ( .A1(n13128), .A2(n12569), .ZN(n13111) );
  OAI21_X1 U8071 ( .B1(n13171), .B2(n6959), .A(n6956), .ZN(n13148) );
  INV_X1 U8072 ( .A(n8556), .ZN(n6959) );
  AND2_X1 U8073 ( .A1(n6957), .A2(n8557), .ZN(n6956) );
  AND3_X1 U8074 ( .A1(n8540), .A2(n8539), .A3(n8538), .ZN(n13162) );
  AND2_X1 U8075 ( .A1(n12560), .A2(n12559), .ZN(n13158) );
  OAI21_X1 U8076 ( .B1(n13199), .B2(n7426), .A(n7424), .ZN(n13173) );
  AOI21_X1 U8077 ( .B1(n7427), .B2(n7425), .A(n6763), .ZN(n7424) );
  INV_X1 U8078 ( .A(n7427), .ZN(n7426) );
  INV_X1 U8079 ( .A(n8522), .ZN(n7425) );
  AND2_X1 U8080 ( .A1(n12555), .A2(n12556), .ZN(n13177) );
  NAND2_X1 U8081 ( .A1(n8657), .A2(n6718), .ZN(n13193) );
  OR2_X1 U8082 ( .A1(n13199), .A2(n13208), .ZN(n13200) );
  AND2_X1 U8083 ( .A1(n12547), .A2(n12548), .ZN(n13208) );
  NAND2_X1 U8084 ( .A1(n7422), .A2(n6698), .ZN(n13217) );
  AOI21_X1 U8085 ( .B1(n6953), .B2(n6955), .A(n6758), .ZN(n6951) );
  NAND2_X1 U8086 ( .A1(n8656), .A2(n12531), .ZN(n13239) );
  NAND2_X1 U8087 ( .A1(n13239), .A2(n13238), .ZN(n13237) );
  AND4_X1 U8088 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n13275)
         );
  AND4_X1 U8089 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(n14863)
         );
  NAND2_X1 U8090 ( .A1(n6783), .A2(n6695), .ZN(n6949) );
  NAND2_X1 U8091 ( .A1(n7423), .A2(n6715), .ZN(n6945) );
  NAND2_X1 U8092 ( .A1(n6965), .A2(n6963), .ZN(n11504) );
  NAND2_X1 U8093 ( .A1(n6966), .A2(n8291), .ZN(n6965) );
  NAND2_X1 U8094 ( .A1(n15569), .A2(n6964), .ZN(n6963) );
  AND2_X1 U8095 ( .A1(n15568), .A2(n8291), .ZN(n6964) );
  NAND2_X1 U8096 ( .A1(n12466), .A2(n12465), .ZN(n11303) );
  NAND2_X1 U8097 ( .A1(n8724), .A2(n12455), .ZN(n15581) );
  NAND2_X1 U8098 ( .A1(n8588), .A2(n8587), .ZN(n13120) );
  OR2_X1 U8099 ( .A1(n12415), .A2(n11597), .ZN(n8587) );
  OR2_X1 U8100 ( .A1(n10309), .A2(n8261), .ZN(n8512) );
  NOR2_X1 U8101 ( .A1(n8188), .A2(n7413), .ZN(n7412) );
  INV_X1 U8102 ( .A(n8186), .ZN(n7413) );
  NAND2_X1 U8103 ( .A1(n6900), .A2(n8182), .ZN(n8598) );
  XNOR2_X1 U8104 ( .A(n8677), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8682) );
  OR2_X1 U8105 ( .A1(n8178), .A2(n11893), .ZN(n8180) );
  NOR2_X1 U8106 ( .A1(n8633), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8630) );
  INV_X1 U8107 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U8108 ( .A1(n6893), .A2(n6894), .ZN(n8523) );
  NAND2_X1 U8109 ( .A1(n7392), .A2(n7390), .ZN(n8492) );
  AOI21_X1 U8110 ( .B1(n7393), .B2(n7395), .A(n7391), .ZN(n7390) );
  INV_X1 U8111 ( .A(n8167), .ZN(n7391) );
  INV_X1 U8112 ( .A(n8165), .ZN(n7395) );
  NAND2_X1 U8113 ( .A1(n8460), .A2(n8165), .ZN(n8473) );
  AND2_X1 U8114 ( .A1(n8167), .A2(n8166), .ZN(n8472) );
  AND2_X1 U8115 ( .A1(n7218), .A2(n8193), .ZN(n7216) );
  NAND2_X1 U8116 ( .A1(n8458), .A2(n8457), .ZN(n8460) );
  AND3_X1 U8117 ( .A1(n7217), .A2(n7218), .A3(n6823), .ZN(n8461) );
  XNOR2_X1 U8118 ( .A(n8157), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8406) );
  NOR2_X1 U8119 ( .A1(n8384), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8399) );
  AND2_X1 U8120 ( .A1(n8141), .A2(n8140), .ZN(n8288) );
  NAND2_X1 U8121 ( .A1(n7107), .A2(n10691), .ZN(n7485) );
  NAND2_X1 U8122 ( .A1(n11414), .A2(n11413), .ZN(n7727) );
  INV_X1 U8123 ( .A(n9578), .ZN(n9579) );
  NAND2_X1 U8124 ( .A1(n7736), .A2(n7735), .ZN(n10705) );
  AOI21_X1 U8125 ( .B1(n7728), .B2(n7730), .A(n7726), .ZN(n7725) );
  INV_X1 U8126 ( .A(n13492), .ZN(n7726) );
  NAND2_X1 U8127 ( .A1(n9992), .A2(n9505), .ZN(n9577) );
  NAND2_X1 U8128 ( .A1(n13596), .A2(n7743), .ZN(n13514) );
  AND2_X1 U8129 ( .A1(n13515), .A2(n9638), .ZN(n7743) );
  NOR2_X1 U8130 ( .A1(n10032), .A2(n10263), .ZN(n13551) );
  OAI21_X1 U8131 ( .B1(n9960), .B2(n7616), .A(n7614), .ZN(n10025) );
  AND2_X1 U8132 ( .A1(n9958), .A2(n9959), .ZN(n7616) );
  NOR2_X1 U8133 ( .A1(n7618), .A2(n7615), .ZN(n7614) );
  NAND2_X1 U8134 ( .A1(n9950), .A2(n6717), .ZN(n9960) );
  INV_X1 U8135 ( .A(n9420), .ZN(n9563) );
  AND2_X1 U8136 ( .A1(n15248), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7338) );
  NOR2_X2 U8137 ( .A1(n7355), .A2(n9955), .ZN(n13759) );
  NOR2_X1 U8138 ( .A1(n6879), .A2(n6777), .ZN(n13775) );
  OR2_X1 U8139 ( .A1(n13799), .A2(n13798), .ZN(n7555) );
  AND2_X1 U8140 ( .A1(n6723), .A2(n13855), .ZN(n7442) );
  NOR2_X1 U8141 ( .A1(n9552), .A2(n13835), .ZN(n7276) );
  AND2_X1 U8142 ( .A1(n7275), .A2(n9551), .ZN(n13838) );
  AOI21_X1 U8143 ( .B1(n9434), .B2(n6904), .A(n6722), .ZN(n13856) );
  NOR2_X1 U8144 ( .A1(n13871), .A2(n6905), .ZN(n6904) );
  INV_X1 U8145 ( .A(n9433), .ZN(n6905) );
  NAND2_X1 U8146 ( .A1(n13856), .A2(n13855), .ZN(n13854) );
  XNOR2_X1 U8147 ( .A(n14010), .B(n9550), .ZN(n13855) );
  NAND2_X1 U8148 ( .A1(n13945), .A2(n9402), .ZN(n13932) );
  OR2_X1 U8149 ( .A1(n13948), .A2(n13947), .ZN(n13950) );
  NAND2_X1 U8150 ( .A1(n8010), .A2(n8009), .ZN(n11993) );
  OR2_X1 U8151 ( .A1(n9378), .A2(n9377), .ZN(n9386) );
  NAND2_X1 U8152 ( .A1(n7996), .A2(n7995), .ZN(n11823) );
  NOR2_X1 U8153 ( .A1(n9368), .A2(n7449), .ZN(n7448) );
  INV_X1 U8154 ( .A(n9359), .ZN(n7449) );
  NAND2_X1 U8155 ( .A1(n7980), .A2(n7979), .ZN(n11607) );
  NAND2_X1 U8156 ( .A1(n6864), .A2(n9317), .ZN(n11233) );
  NAND2_X1 U8157 ( .A1(n11066), .A2(n11069), .ZN(n6864) );
  INV_X1 U8158 ( .A(n15315), .ZN(n6881) );
  NOR2_X1 U8159 ( .A1(n10224), .A2(n9751), .ZN(n9743) );
  INV_X1 U8160 ( .A(n13748), .ZN(n9574) );
  INV_X1 U8161 ( .A(n13972), .ZN(n6912) );
  NAND2_X1 U8162 ( .A1(n8039), .A2(n8038), .ZN(n13907) );
  NAND2_X1 U8163 ( .A1(n8032), .A2(n8031), .ZN(n14031) );
  NAND2_X1 U8164 ( .A1(n8025), .A2(n8024), .ZN(n13936) );
  NAND2_X1 U8165 ( .A1(n10743), .A2(n8123), .ZN(n15398) );
  INV_X1 U8166 ( .A(n7639), .ZN(n7637) );
  XNOR2_X1 U8167 ( .A(n8115), .B(n8114), .ZN(n10035) );
  OAI21_X1 U8168 ( .B1(n8066), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8115) );
  NAND3_X1 U8169 ( .A1(n7864), .A2(n6986), .A3(n15236), .ZN(n6989) );
  INV_X1 U8170 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7864) );
  INV_X1 U8171 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U8172 ( .A1(n7909), .A2(n7863), .ZN(n7927) );
  AOI21_X1 U8173 ( .B1(n11542), .B2(n6834), .A(n7652), .ZN(n7651) );
  INV_X1 U8174 ( .A(n11632), .ZN(n7652) );
  XNOR2_X1 U8175 ( .A(n11027), .B(n11778), .ZN(n11489) );
  NAND2_X1 U8176 ( .A1(n14198), .A2(n6751), .ZN(n14152) );
  AND2_X1 U8177 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  INV_X1 U8178 ( .A(n14124), .ZN(n7660) );
  AND2_X1 U8179 ( .A1(n7658), .A2(n12740), .ZN(n7657) );
  NAND2_X1 U8180 ( .A1(n14124), .A2(n7659), .ZN(n7658) );
  NAND2_X1 U8181 ( .A1(n6834), .A2(n11543), .ZN(n7654) );
  CLKBUF_X1 U8182 ( .A(n7651), .Z(n7024) );
  AND2_X1 U8183 ( .A1(n15149), .A2(n10570), .ZN(n12190) );
  AND2_X1 U8184 ( .A1(n10636), .A2(n11218), .ZN(n10630) );
  NAND2_X1 U8185 ( .A1(n7202), .A2(n7572), .ZN(n12367) );
  NAND2_X1 U8186 ( .A1(n7573), .A2(n12359), .ZN(n7572) );
  OAI21_X1 U8187 ( .B1(n12212), .B2(n12211), .A(n12209), .ZN(n7058) );
  AND4_X1 U8188 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n11777) );
  NOR2_X1 U8189 ( .A1(n12195), .A2(n7317), .ZN(n7316) );
  INV_X1 U8190 ( .A(n7318), .ZN(n7317) );
  NAND2_X1 U8191 ( .A1(n12013), .A2(n12012), .ZN(n14497) );
  AND2_X1 U8192 ( .A1(n14441), .A2(n7511), .ZN(n7138) );
  NAND2_X1 U8193 ( .A1(n7512), .A2(n7516), .ZN(n7511) );
  NAND2_X1 U8194 ( .A1(n7161), .A2(n6714), .ZN(n7512) );
  NAND2_X1 U8195 ( .A1(n14582), .A2(n7513), .ZN(n7510) );
  NAND2_X1 U8196 ( .A1(n14782), .A2(n12116), .ZN(n14572) );
  NOR2_X1 U8197 ( .A1(n14439), .A2(n7168), .ZN(n7167) );
  INV_X1 U8198 ( .A(n14425), .ZN(n7168) );
  OR2_X1 U8199 ( .A1(n7167), .A2(n7166), .ZN(n7165) );
  INV_X1 U8200 ( .A(n14422), .ZN(n14609) );
  AOI21_X1 U8201 ( .B1(n6692), .B2(n7302), .A(n6770), .ZN(n7301) );
  NOR2_X1 U8202 ( .A1(n14419), .A2(n7305), .ZN(n7304) );
  INV_X1 U8203 ( .A(n14418), .ZN(n7305) );
  NOR2_X1 U8204 ( .A1(n14432), .A2(n14652), .ZN(n6977) );
  INV_X1 U8205 ( .A(n15102), .ZN(n14643) );
  NOR2_X1 U8206 ( .A1(n7582), .A2(n7581), .ZN(n7580) );
  INV_X1 U8207 ( .A(n11919), .ZN(n7581) );
  NAND2_X1 U8208 ( .A1(n7146), .A2(n7145), .ZN(n14651) );
  AOI21_X1 U8209 ( .B1(n11709), .B2(n11708), .A(n6773), .ZN(n11710) );
  NAND2_X1 U8210 ( .A1(n11534), .A2(n11658), .ZN(n11672) );
  INV_X1 U8211 ( .A(n11674), .ZN(n7292) );
  INV_X1 U8212 ( .A(n11675), .ZN(n7290) );
  OR2_X1 U8213 ( .A1(n12638), .A2(n14971), .ZN(n7508) );
  NAND2_X1 U8214 ( .A1(n7504), .A2(n11529), .ZN(n7503) );
  XNOR2_X1 U8215 ( .A(n14192), .B(n14262), .ZN(n12106) );
  NAND2_X1 U8216 ( .A1(n12190), .A2(n14283), .ZN(n15097) );
  NAND2_X1 U8217 ( .A1(n12077), .A2(n12076), .ZN(n14721) );
  INV_X1 U8218 ( .A(n15156), .ZN(n15204) );
  NAND2_X1 U8219 ( .A1(n10885), .A2(n11229), .ZN(n15156) );
  NAND2_X1 U8220 ( .A1(n10213), .A2(n10212), .ZN(n10624) );
  INV_X1 U8221 ( .A(n14781), .ZN(n10212) );
  XNOR2_X1 U8222 ( .A(n7879), .B(n7878), .ZN(n12377) );
  AOI21_X1 U8223 ( .B1(n7071), .B2(n7069), .A(n6820), .ZN(n7068) );
  XNOR2_X1 U8224 ( .A(n7888), .B(SI_22_), .ZN(n12053) );
  NAND2_X1 U8225 ( .A1(n7682), .A2(n10568), .ZN(n7681) );
  INV_X1 U8226 ( .A(n7683), .ZN(n7682) );
  XNOR2_X1 U8227 ( .A(n7076), .B(n10564), .ZN(n7903) );
  OAI21_X1 U8228 ( .B1(n7977), .B2(n7976), .A(n7801), .ZN(n7981) );
  NAND2_X1 U8229 ( .A1(n15031), .A2(n7517), .ZN(n7096) );
  OR2_X1 U8230 ( .A1(n15031), .A2(n7517), .ZN(n7090) );
  INV_X1 U8231 ( .A(n8903), .ZN(n7093) );
  NOR2_X1 U8232 ( .A1(n6842), .A2(n6841), .ZN(n8853) );
  AND2_X1 U8233 ( .A1(n8843), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U8234 ( .A1(n8855), .A2(n8856), .ZN(n6842) );
  XNOR2_X1 U8235 ( .A(n8845), .B(n6840), .ZN(n8906) );
  INV_X1 U8236 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n6840) );
  AOI21_X1 U8237 ( .B1(n7699), .B2(n7697), .A(n7696), .ZN(n7695) );
  INV_X1 U8238 ( .A(n7699), .ZN(n7698) );
  NAND2_X1 U8239 ( .A1(n10669), .A2(n8731), .ZN(n10670) );
  AND3_X1 U8240 ( .A1(n8530), .A2(n8529), .A3(n8528), .ZN(n13175) );
  INV_X1 U8241 ( .A(n13375), .ZN(n7039) );
  OR2_X1 U8242 ( .A1(n8261), .A2(n10122), .ZN(n8332) );
  NAND2_X1 U8243 ( .A1(n8727), .A2(n8726), .ZN(n12611) );
  NAND2_X1 U8244 ( .A1(n8534), .A2(n8533), .ZN(n13179) );
  OR2_X1 U8245 ( .A1(n12415), .A2(n10811), .ZN(n8533) );
  OR2_X1 U8246 ( .A1(n8750), .A2(n8749), .ZN(n6930) );
  NAND2_X1 U8247 ( .A1(n6918), .A2(n12843), .ZN(n12846) );
  NAND2_X1 U8248 ( .A1(n12842), .A2(n12844), .ZN(n6918) );
  NAND2_X1 U8249 ( .A1(n13120), .A2(n12943), .ZN(n7226) );
  INV_X1 U8250 ( .A(n12847), .ZN(n7225) );
  NAND2_X1 U8251 ( .A1(n7717), .A2(n7716), .ZN(n11082) );
  NAND2_X1 U8252 ( .A1(n7718), .A2(n6724), .ZN(n7716) );
  NAND2_X1 U8253 ( .A1(n8483), .A2(n8482), .ZN(n13240) );
  OR2_X1 U8254 ( .A1(n10184), .A2(n8261), .ZN(n8483) );
  NAND2_X1 U8255 ( .A1(n8583), .A2(n8582), .ZN(n13314) );
  OR2_X1 U8256 ( .A1(n12415), .A2(n11443), .ZN(n8582) );
  XNOR2_X1 U8257 ( .A(n7215), .B(n8787), .ZN(n10848) );
  XNOR2_X1 U8258 ( .A(n15556), .B(n8734), .ZN(n7215) );
  AND3_X1 U8259 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n11318) );
  OR2_X1 U8260 ( .A1(n8261), .A2(n10120), .ZN(n8302) );
  NAND2_X1 U8261 ( .A1(n8798), .A2(n10659), .ZN(n12931) );
  NAND2_X1 U8262 ( .A1(n12922), .A2(n12923), .ZN(n12921) );
  OAI21_X1 U8263 ( .B1(n12842), .B2(n6921), .A(n6919), .ZN(n12922) );
  AOI21_X1 U8264 ( .B1(n12843), .B2(n6920), .A(n7702), .ZN(n6919) );
  NAND2_X1 U8265 ( .A1(n7420), .A2(n12417), .ZN(n8449) );
  INV_X1 U8266 ( .A(n10160), .ZN(n7420) );
  INV_X1 U8267 ( .A(n13222), .ZN(n13187) );
  INV_X1 U8268 ( .A(n13274), .ZN(n14851) );
  XNOR2_X1 U8269 ( .A(n12957), .B(n12964), .ZN(n11898) );
  XNOR2_X1 U8270 ( .A(n13002), .B(n13007), .ZN(n12982) );
  XNOR2_X1 U8271 ( .A(n7118), .B(n7117), .ZN(n7116) );
  INV_X1 U8272 ( .A(n14838), .ZN(n7117) );
  OAI21_X1 U8273 ( .B1(n14839), .B2(n7469), .A(n7127), .ZN(n7126) );
  NAND2_X1 U8274 ( .A1(n14837), .A2(n7471), .ZN(n7469) );
  AOI21_X1 U8275 ( .B1(n13056), .B2(n15508), .A(n13055), .ZN(n7127) );
  NAND2_X1 U8276 ( .A1(n7474), .A2(n7472), .ZN(n7471) );
  INV_X1 U8277 ( .A(n7118), .ZN(n14839) );
  NOR2_X1 U8278 ( .A1(n15523), .A2(n6835), .ZN(n7468) );
  INV_X1 U8279 ( .A(n7473), .ZN(n7470) );
  XNOR2_X1 U8280 ( .A(n13050), .B(n7124), .ZN(n7123) );
  INV_X1 U8281 ( .A(n13049), .ZN(n7124) );
  NAND2_X1 U8282 ( .A1(n7017), .A2(n13074), .ZN(n13301) );
  NAND2_X1 U8283 ( .A1(n7039), .A2(n7038), .ZN(n7037) );
  AOI21_X1 U8284 ( .B1(n12621), .B2(n12417), .A(n12416), .ZN(n13369) );
  AND2_X1 U8285 ( .A1(n13068), .A2(n15669), .ZN(n8667) );
  AOI21_X1 U8286 ( .B1(n13300), .B2(n15669), .A(n13301), .ZN(n13373) );
  OR2_X1 U8287 ( .A1(n12415), .A2(n11801), .ZN(n8614) );
  NOR2_X1 U8288 ( .A1(n13303), .A2(n7379), .ZN(n13376) );
  AND2_X1 U8289 ( .A1(n13304), .A2(n15662), .ZN(n7379) );
  INV_X1 U8290 ( .A(SI_4_), .ZN(n10074) );
  AND2_X1 U8291 ( .A1(n9727), .A2(n9721), .ZN(n7742) );
  AND2_X1 U8292 ( .A1(n9631), .A2(n9625), .ZN(n7732) );
  NAND2_X1 U8293 ( .A1(n11618), .A2(n9625), .ZN(n11623) );
  AND2_X1 U8294 ( .A1(n13608), .A2(n9681), .ZN(n13483) );
  NAND2_X1 U8295 ( .A1(n8043), .A2(n8042), .ZN(n13996) );
  NOR2_X1 U8296 ( .A1(n6738), .A2(n7462), .ZN(n7461) );
  NOR2_X1 U8297 ( .A1(n10031), .A2(n10282), .ZN(n7462) );
  INV_X1 U8298 ( .A(n15315), .ZN(n10422) );
  XNOR2_X1 U8299 ( .A(n13737), .B(n9982), .ZN(n8071) );
  INV_X1 U8300 ( .A(n14050), .ZN(n13742) );
  INV_X1 U8301 ( .A(n9982), .ZN(n13736) );
  NAND2_X1 U8302 ( .A1(n6873), .A2(n6872), .ZN(n7351) );
  NAND2_X1 U8303 ( .A1(n13744), .A2(n15370), .ZN(n6873) );
  AND2_X1 U8304 ( .A1(n7261), .A2(n7260), .ZN(n6872) );
  INV_X1 U8305 ( .A(n13750), .ZN(n7260) );
  AND2_X1 U8306 ( .A1(n10639), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10214) );
  AOI21_X1 U8307 ( .B1(n7664), .B2(n7666), .A(n6762), .ZN(n7661) );
  NAND2_X1 U8308 ( .A1(n14174), .A2(n7664), .ZN(n7662) );
  NAND2_X1 U8309 ( .A1(n7680), .A2(n12704), .ZN(n14145) );
  NAND2_X1 U8310 ( .A1(n10993), .A2(n12161), .ZN(n7306) );
  NAND2_X1 U8311 ( .A1(n12089), .A2(n12088), .ZN(n14951) );
  INV_X1 U8312 ( .A(n11540), .ZN(n7050) );
  INV_X1 U8313 ( .A(n14261), .ZN(n14971) );
  INV_X1 U8314 ( .A(n15097), .ZN(n14641) );
  XNOR2_X1 U8315 ( .A(n10595), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n14275) );
  AND2_X1 U8316 ( .A1(n10359), .A2(n10358), .ZN(n14400) );
  AND2_X1 U8317 ( .A1(n10359), .A2(n10202), .ZN(n14398) );
  XNOR2_X1 U8318 ( .A(n7241), .B(n14448), .ZN(n14449) );
  AOI21_X1 U8319 ( .B1(n7238), .B2(n7240), .A(n6782), .ZN(n7237) );
  AOI22_X1 U8320 ( .A1(n14470), .A2(n14471), .B1(n14485), .B2(n7172), .ZN(
        n14670) );
  NAND2_X1 U8321 ( .A1(n14485), .A2(n7175), .ZN(n14470) );
  AND2_X1 U8322 ( .A1(n6969), .A2(n6821), .ZN(n6968) );
  NAND2_X1 U8323 ( .A1(n6971), .A2(n14645), .ZN(n6970) );
  NAND2_X1 U8324 ( .A1(n12147), .A2(n12146), .ZN(n14562) );
  NAND2_X1 U8325 ( .A1(n15223), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8326 ( .A1(n15210), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7158) );
  XNOR2_X1 U8327 ( .A(n14430), .B(n14448), .ZN(n14669) );
  NAND2_X1 U8328 ( .A1(n7171), .A2(n7170), .ZN(n14430) );
  OR2_X1 U8329 ( .A1(n7172), .A2(n14429), .ZN(n7170) );
  INV_X1 U8330 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10579) );
  NOR2_X1 U8331 ( .A1(n15694), .A2(n15695), .ZN(n15693) );
  NAND2_X1 U8332 ( .A1(n7525), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U8333 ( .A1(n15043), .A2(n15044), .ZN(n7525) );
  OR2_X1 U8334 ( .A1(n15043), .A2(n15044), .ZN(n7530) );
  NAND2_X1 U8335 ( .A1(n14810), .A2(n15312), .ZN(n14807) );
  OAI21_X1 U8336 ( .B1(n14786), .B2(n14785), .A(n7523), .ZN(n7100) );
  INV_X1 U8337 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U8338 ( .A1(n14786), .A2(n14785), .ZN(n14784) );
  AND2_X1 U8339 ( .A1(n12218), .A2(n6682), .ZN(n7586) );
  OAI21_X1 U8340 ( .B1(n12217), .B2(n12216), .A(n12215), .ZN(n7587) );
  NAND2_X1 U8341 ( .A1(n6794), .A2(n9779), .ZN(n7642) );
  NAND2_X1 U8342 ( .A1(n12252), .A2(n12254), .ZN(n7184) );
  NAND2_X1 U8343 ( .A1(n9788), .A2(n6716), .ZN(n9794) );
  NAND2_X1 U8344 ( .A1(n12267), .A2(n12265), .ZN(n7191) );
  OAI21_X1 U8345 ( .B1(n7596), .B2(n7595), .A(n7009), .ZN(n7190) );
  NAND2_X1 U8346 ( .A1(n12277), .A2(n7576), .ZN(n7575) );
  INV_X1 U8347 ( .A(n12276), .ZN(n7576) );
  NOR2_X1 U8348 ( .A1(n9828), .A2(n6739), .ZN(n7626) );
  NAND2_X1 U8349 ( .A1(n7622), .A2(n6759), .ZN(n9820) );
  INV_X1 U8350 ( .A(n9813), .ZN(n7623) );
  AND2_X1 U8351 ( .A1(n12308), .A2(n7563), .ZN(n7562) );
  NAND2_X1 U8352 ( .A1(n9838), .A2(n6740), .ZN(n7635) );
  MUX2_X1 U8353 ( .A(n14565), .B(n14709), .S(n6682), .Z(n12313) );
  INV_X1 U8354 ( .A(n9888), .ZN(n7620) );
  NOR2_X1 U8355 ( .A1(n9888), .A2(n9891), .ZN(n7621) );
  AND2_X1 U8356 ( .A1(n7588), .A2(n12327), .ZN(n7589) );
  INV_X1 U8357 ( .A(n9912), .ZN(n7631) );
  NAND2_X1 U8358 ( .A1(n7611), .A2(n7610), .ZN(n7609) );
  INV_X1 U8359 ( .A(n9924), .ZN(n7611) );
  INV_X1 U8360 ( .A(n9923), .ZN(n7610) );
  AOI21_X1 U8361 ( .B1(n6726), .B2(n7182), .A(n6689), .ZN(n7178) );
  AND2_X1 U8362 ( .A1(n12338), .A2(n7183), .ZN(n7182) );
  AOI21_X1 U8363 ( .B1(n7976), .B2(n7801), .A(n7066), .ZN(n7065) );
  INV_X1 U8364 ( .A(n7761), .ZN(n7066) );
  AND2_X1 U8365 ( .A1(n13369), .A2(n12947), .ZN(n12441) );
  INV_X1 U8366 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7723) );
  INV_X1 U8367 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8196) );
  INV_X1 U8368 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8194) );
  INV_X1 U8369 ( .A(n8558), .ZN(n7418) );
  INV_X1 U8370 ( .A(n8177), .ZN(n7415) );
  NAND2_X1 U8371 ( .A1(n7601), .A2(n6731), .ZN(n9942) );
  INV_X1 U8372 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8028) );
  INV_X4 U8373 ( .A(n12240), .ZN(n12350) );
  INV_X1 U8374 ( .A(n14417), .ZN(n7149) );
  NAND2_X1 U8375 ( .A1(n7014), .A2(n7013), .ZN(n7307) );
  INV_X1 U8376 ( .A(n7065), .ZN(n7064) );
  INV_X1 U8377 ( .A(n7542), .ZN(n7541) );
  OAI21_X1 U8378 ( .B1(n7793), .B2(n7543), .A(n7797), .ZN(n7542) );
  INV_X1 U8379 ( .A(n7795), .ZN(n7543) );
  AOI21_X1 U8380 ( .B1(n7246), .B2(n7952), .A(n7958), .ZN(n7245) );
  OR2_X1 U8381 ( .A1(n12820), .A2(n11446), .ZN(n8739) );
  NOR2_X1 U8382 ( .A1(n6693), .A2(n11860), .ZN(n7221) );
  AOI21_X1 U8383 ( .B1(n7707), .B2(n8753), .A(n7705), .ZN(n7704) );
  INV_X1 U8384 ( .A(n8755), .ZN(n7705) );
  NOR2_X1 U8385 ( .A1(n12443), .A2(n12419), .ZN(n7022) );
  NAND2_X1 U8386 ( .A1(n12586), .A2(n12587), .ZN(n7033) );
  INV_X1 U8387 ( .A(n12441), .ZN(n12591) );
  NOR2_X1 U8388 ( .A1(n13297), .A2(n12421), .ZN(n12595) );
  NAND2_X1 U8389 ( .A1(n10775), .A2(n10774), .ZN(n10777) );
  NAND2_X1 U8390 ( .A1(n15461), .A2(n7120), .ZN(n11131) );
  OR2_X1 U8391 ( .A1(n11147), .A2(n11145), .ZN(n7120) );
  INV_X1 U8392 ( .A(n12987), .ZN(n7111) );
  NOR2_X1 U8393 ( .A1(n14826), .A2(n13225), .ZN(n7475) );
  NAND2_X1 U8394 ( .A1(n8556), .A2(n6958), .ZN(n6957) );
  INV_X1 U8395 ( .A(n8543), .ZN(n6958) );
  OR2_X1 U8396 ( .A1(n13319), .A2(n13161), .ZN(n12566) );
  AND2_X1 U8397 ( .A1(n13190), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U8398 ( .A1(n13208), .A2(n8522), .ZN(n7428) );
  INV_X1 U8399 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9174) );
  AND2_X1 U8400 ( .A1(n13247), .A2(n6954), .ZN(n6953) );
  OR2_X1 U8401 ( .A1(n13258), .A2(n6955), .ZN(n6954) );
  INV_X1 U8402 ( .A(n8456), .ZN(n6955) );
  OR2_X1 U8403 ( .A1(n8376), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8390) );
  OR2_X1 U8404 ( .A1(n11451), .A2(n11318), .ZN(n12483) );
  NAND2_X1 U8405 ( .A1(n6728), .A2(n15553), .ZN(n6966) );
  NAND2_X1 U8406 ( .A1(n15569), .A2(n15568), .ZN(n6967) );
  NOR2_X1 U8407 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8278) );
  INV_X1 U8408 ( .A(n6894), .ZN(n6890) );
  AND2_X1 U8409 ( .A1(n8288), .A2(n8142), .ZN(n7402) );
  NOR2_X1 U8410 ( .A1(n11200), .A2(n7734), .ZN(n7733) );
  INV_X1 U8411 ( .A(n9610), .ZN(n7734) );
  NAND2_X1 U8412 ( .A1(n13506), .A2(n9696), .ZN(n9701) );
  OR2_X1 U8413 ( .A1(n9965), .A2(n7619), .ZN(n7618) );
  NOR2_X1 U8414 ( .A1(n9959), .A2(n9958), .ZN(n7615) );
  INV_X1 U8415 ( .A(n10010), .ZN(n7537) );
  INV_X1 U8416 ( .A(n9479), .ZN(n7458) );
  OR2_X1 U8417 ( .A1(n9479), .A2(n7459), .ZN(n7457) );
  NOR2_X1 U8418 ( .A1(n13986), .A2(n13811), .ZN(n7354) );
  INV_X1 U8419 ( .A(n7442), .ZN(n7439) );
  NAND2_X1 U8420 ( .A1(n9260), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9450) );
  NOR2_X1 U8421 ( .A1(n13903), .A2(n14022), .ZN(n7359) );
  OR2_X1 U8422 ( .A1(n9418), .A2(n9258), .ZN(n9427) );
  NOR2_X1 U8423 ( .A1(n11823), .A2(n11795), .ZN(n7348) );
  INV_X1 U8424 ( .A(n7448), .ZN(n7444) );
  OR2_X1 U8425 ( .A1(n11236), .A2(n6812), .ZN(n7263) );
  NAND2_X1 U8426 ( .A1(n7361), .A2(n7356), .ZN(n13844) );
  INV_X1 U8427 ( .A(n13860), .ZN(n7356) );
  NOR2_X1 U8428 ( .A1(n11067), .A2(n11208), .ZN(n11234) );
  INV_X1 U8429 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6860) );
  INV_X1 U8430 ( .A(n6989), .ZN(n6988) );
  INV_X1 U8431 ( .A(n12733), .ZN(n7659) );
  INV_X1 U8432 ( .A(n12770), .ZN(n12727) );
  NAND2_X1 U8433 ( .A1(n12360), .A2(n7571), .ZN(n7570) );
  INV_X1 U8434 ( .A(n12359), .ZN(n7571) );
  NAND2_X1 U8435 ( .A1(n7078), .A2(n12350), .ZN(n7077) );
  NAND2_X1 U8436 ( .A1(n14407), .A2(n12176), .ZN(n7078) );
  INV_X1 U8437 ( .A(n14547), .ZN(n7322) );
  OR2_X1 U8438 ( .A1(n14991), .A2(n14951), .ZN(n7328) );
  INV_X1 U8439 ( .A(n7304), .ZN(n7302) );
  NOR2_X1 U8440 ( .A1(n14416), .A2(n11951), .ZN(n7011) );
  INV_X1 U8441 ( .A(n7763), .ZN(n7288) );
  INV_X1 U8442 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U8443 ( .A1(n15107), .A2(n10887), .ZN(n12218) );
  NOR2_X1 U8444 ( .A1(n14647), .A2(n7328), .ZN(n14743) );
  NAND2_X1 U8445 ( .A1(n15107), .A2(n15148), .ZN(n15090) );
  NAND2_X1 U8446 ( .A1(n15077), .A2(n14401), .ZN(n10885) );
  OAI21_X1 U8447 ( .B1(n8041), .B2(n7839), .A(n7838), .ZN(n8045) );
  XNOR2_X1 U8448 ( .A(n7837), .B(SI_24_), .ZN(n8041) );
  INV_X1 U8449 ( .A(n7899), .ZN(n7825) );
  INV_X1 U8450 ( .A(n7824), .ZN(n7069) );
  INV_X1 U8451 ( .A(n7071), .ZN(n7070) );
  NAND2_X1 U8452 ( .A1(n7684), .A2(n7046), .ZN(n7683) );
  INV_X1 U8453 ( .A(n7685), .ZN(n7684) );
  NAND2_X1 U8454 ( .A1(n7060), .A2(n6743), .ZN(n7249) );
  AOI21_X1 U8455 ( .B1(n7546), .B2(n7549), .A(n6776), .ZN(n7544) );
  OAI21_X1 U8456 ( .B1(n10157), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10176) );
  OR2_X1 U8457 ( .A1(n10151), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U8458 ( .A1(n7293), .A2(n7081), .ZN(n7235) );
  NAND2_X1 U8459 ( .A1(n7295), .A2(n7082), .ZN(n7081) );
  OAI21_X1 U8460 ( .B1(n7296), .B2(n7779), .A(n7781), .ZN(n7293) );
  OAI21_X1 U8461 ( .B1(n7299), .B2(n7924), .A(n7933), .ZN(n7298) );
  NAND2_X1 U8462 ( .A1(n7043), .A2(n6756), .ZN(n7772) );
  INV_X1 U8463 ( .A(n7774), .ZN(n7043) );
  INV_X1 U8464 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7281) );
  INV_X1 U8465 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7280) );
  XNOR2_X1 U8466 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n8863) );
  NAND2_X1 U8467 ( .A1(n6853), .A2(n7084), .ZN(n8821) );
  NAND2_X1 U8468 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7085), .ZN(n7084) );
  XNOR2_X1 U8469 ( .A(n8824), .B(n7099), .ZN(n8861) );
  INV_X1 U8470 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9161) );
  AOI21_X1 U8471 ( .B1(n8853), .B2(n8844), .A(n8852), .ZN(n8845) );
  NOR2_X1 U8472 ( .A1(n7697), .A2(n8794), .ZN(n7694) );
  NOR3_X1 U8473 ( .A1(n8794), .A2(n7697), .A3(n12923), .ZN(n7696) );
  INV_X1 U8474 ( .A(n7701), .ZN(n7697) );
  NOR2_X1 U8475 ( .A1(n12782), .A2(n7708), .ZN(n7707) );
  OR2_X1 U8476 ( .A1(n12891), .A2(n8753), .ZN(n7709) );
  NAND2_X1 U8477 ( .A1(n6701), .A2(n12901), .ZN(n6927) );
  NOR2_X1 U8478 ( .A1(n8513), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8526) );
  OAI21_X1 U8479 ( .B1(n6925), .B2(n6924), .A(n6922), .ZN(n7714) );
  NOR2_X1 U8480 ( .A1(n6923), .A2(n6771), .ZN(n6922) );
  NOR2_X1 U8481 ( .A1(n8764), .A2(n6924), .ZN(n6923) );
  AND2_X1 U8482 ( .A1(n8526), .A2(n9174), .ZN(n8535) );
  NAND2_X1 U8483 ( .A1(n8535), .A2(n12834), .ZN(n8549) );
  NOR2_X1 U8484 ( .A1(n8450), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8465) );
  INV_X1 U8485 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9042) );
  XNOR2_X1 U8486 ( .A(n8787), .B(n8734), .ZN(n7214) );
  NAND2_X1 U8487 ( .A1(n8759), .A2(n12948), .ZN(n8760) );
  AND2_X1 U8488 ( .A1(n12844), .A2(n8785), .ZN(n12868) );
  OR2_X1 U8489 ( .A1(n8732), .A2(n15589), .ZN(n8733) );
  INV_X1 U8490 ( .A(n11325), .ZN(n7229) );
  NAND2_X1 U8491 ( .A1(n12417), .A2(n6838), .ZN(n8349) );
  NAND2_X1 U8492 ( .A1(n7690), .A2(n7687), .ZN(n12612) );
  INV_X1 U8493 ( .A(n12611), .ZN(n7687) );
  NAND2_X1 U8494 ( .A1(n8724), .A2(n7691), .ZN(n7690) );
  NAND2_X1 U8495 ( .A1(n7688), .A2(n6937), .ZN(n7691) );
  NAND2_X1 U8496 ( .A1(n6929), .A2(n7689), .ZN(n8727) );
  XNOR2_X1 U8497 ( .A(n7688), .B(n15606), .ZN(n6929) );
  NAND2_X1 U8498 ( .A1(n8484), .A2(n12861), .ZN(n8496) );
  OR2_X1 U8499 ( .A1(n8496), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8513) );
  OR2_X1 U8500 ( .A1(n12578), .A2(n12599), .ZN(n8807) );
  INV_X1 U8501 ( .A(n12844), .ZN(n6920) );
  OAI21_X1 U8502 ( .B1(n10777), .B2(n10780), .A(n10776), .ZN(n10796) );
  NAND2_X1 U8503 ( .A1(n10798), .A2(n10782), .ZN(n10783) );
  NAND2_X1 U8504 ( .A1(n15443), .A2(n11130), .ZN(n15463) );
  NAND2_X1 U8505 ( .A1(n15463), .A2(n15462), .ZN(n15461) );
  OR2_X1 U8506 ( .A1(n15432), .A2(n11122), .ZN(n7115) );
  XNOR2_X1 U8507 ( .A(n11131), .B(n11153), .ZN(n15479) );
  AND2_X1 U8508 ( .A1(n7113), .A2(n7112), .ZN(n11123) );
  NAND2_X1 U8509 ( .A1(n15458), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U8510 ( .A1(n15517), .A2(n11134), .ZN(n11135) );
  NAND2_X1 U8511 ( .A1(n11565), .A2(n11566), .ZN(n11567) );
  AOI21_X1 U8512 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11899), .A(n11894), .ZN(
        n12952) );
  NAND2_X1 U8513 ( .A1(n12984), .A2(n12986), .ZN(n13006) );
  OR2_X1 U8514 ( .A1(n14838), .A2(n13040), .ZN(n7474) );
  NOR2_X1 U8515 ( .A1(n13038), .A2(n7475), .ZN(n7473) );
  AOI21_X1 U8516 ( .B1(n7473), .B2(n14838), .A(n6833), .ZN(n7472) );
  NAND2_X1 U8517 ( .A1(n6719), .A2(n6944), .ZN(n7431) );
  NAND2_X1 U8518 ( .A1(n7430), .A2(n6719), .ZN(n7429) );
  NOR2_X1 U8519 ( .A1(n13088), .A2(n6942), .ZN(n6941) );
  INV_X1 U8520 ( .A(n8610), .ZN(n6942) );
  NAND2_X1 U8521 ( .A1(n8611), .A2(n8610), .ZN(n13086) );
  NAND2_X1 U8522 ( .A1(n13114), .A2(n13113), .ZN(n13112) );
  NAND2_X1 U8523 ( .A1(n13126), .A2(n8659), .ZN(n13128) );
  NOR2_X1 U8524 ( .A1(n8562), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8573) );
  INV_X1 U8525 ( .A(n13148), .ZN(n8570) );
  AND2_X1 U8526 ( .A1(n12566), .A2(n12562), .ZN(n13149) );
  NAND2_X1 U8527 ( .A1(n6875), .A2(n12555), .ZN(n13164) );
  INV_X1 U8528 ( .A(n7374), .ZN(n7373) );
  OAI21_X1 U8529 ( .B1(n6718), .B2(n7375), .A(n12556), .ZN(n7374) );
  AND4_X1 U8530 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n13236)
         );
  AND4_X1 U8531 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n13274)
         );
  AOI21_X1 U8532 ( .B1(n7383), .B2(n7382), .A(n7381), .ZN(n7380) );
  INV_X1 U8533 ( .A(n12502), .ZN(n7382) );
  INV_X1 U8534 ( .A(n12506), .ZN(n7381) );
  INV_X1 U8535 ( .A(n6949), .ZN(n6948) );
  AOI21_X1 U8536 ( .B1(n6947), .B2(n6949), .A(n6784), .ZN(n6946) );
  INV_X1 U8537 ( .A(n12507), .ZN(n14865) );
  OR2_X1 U8538 ( .A1(n8351), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U8539 ( .A1(n7423), .A2(n6713), .ZN(n11765) );
  NOR2_X1 U8540 ( .A1(n8305), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8322) );
  OR2_X1 U8541 ( .A1(n8292), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8305) );
  AND2_X1 U8542 ( .A1(n6967), .A2(n6728), .ZN(n15554) );
  NAND2_X1 U8543 ( .A1(n6967), .A2(n6962), .ZN(n15552) );
  INV_X1 U8544 ( .A(n6966), .ZN(n6962) );
  OR2_X1 U8545 ( .A1(n8261), .A2(n10078), .ZN(n8290) );
  OR2_X1 U8546 ( .A1(n8261), .A2(n10072), .ZN(n8276) );
  AND2_X1 U8547 ( .A1(n11303), .A2(n8253), .ZN(n7001) );
  INV_X1 U8548 ( .A(n12463), .ZN(n15593) );
  NAND2_X1 U8549 ( .A1(n15581), .A2(n15593), .ZN(n15580) );
  NAND2_X1 U8550 ( .A1(n6939), .A2(n12615), .ZN(n6938) );
  NAND2_X1 U8551 ( .A1(n8600), .A2(n8599), .ZN(n13306) );
  OR2_X1 U8552 ( .A1(n12415), .A2(n11728), .ZN(n8599) );
  OR2_X1 U8553 ( .A1(n10170), .A2(n8261), .ZN(n8464) );
  AND2_X1 U8554 ( .A1(n13426), .A2(n10070), .ZN(n10678) );
  OAI21_X1 U8555 ( .B1(n10136), .B2(P3_D_REG_1__SCAN_IN), .A(n8683), .ZN(
        n10652) );
  OAI21_X1 U8556 ( .B1(n8598), .B2(n8183), .A(n8184), .ZN(n8613) );
  OR2_X1 U8557 ( .A1(n8674), .A2(n7721), .ZN(n8672) );
  NAND2_X1 U8558 ( .A1(n8195), .A2(n7724), .ZN(n7721) );
  NAND2_X1 U8559 ( .A1(n8179), .A2(n12375), .ZN(n6899) );
  NAND2_X1 U8560 ( .A1(n8476), .A2(n7387), .ZN(n8674) );
  XNOR2_X1 U8561 ( .A(n8669), .B(n8670), .ZN(n10679) );
  INV_X1 U8562 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8669) );
  OAI21_X1 U8563 ( .B1(n8668), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8670) );
  XNOR2_X1 U8564 ( .A(n8634), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U8565 ( .A1(n6901), .A2(n8170), .ZN(n8505) );
  INV_X1 U8566 ( .A(n7213), .ZN(n8627) );
  OAI21_X1 U8567 ( .B1(n8426), .B2(n8160), .A(n8161), .ZN(n8442) );
  OR2_X1 U8568 ( .A1(n8361), .A2(n8360), .ZN(n8384) );
  AND2_X1 U8569 ( .A1(n8151), .A2(n8150), .ZN(n8364) );
  AOI21_X1 U8570 ( .B1(n8330), .B2(n6888), .A(n6887), .ZN(n6886) );
  INV_X1 U8571 ( .A(n8330), .ZN(n6889) );
  INV_X1 U8572 ( .A(n8145), .ZN(n6888) );
  AND2_X1 U8573 ( .A1(n8149), .A2(n8148), .ZN(n8345) );
  OR2_X1 U8574 ( .A1(n8328), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8343) );
  AOI21_X1 U8575 ( .B1(n8259), .B2(n7397), .A(n7399), .ZN(n7396) );
  XNOR2_X1 U8576 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8229) );
  NAND2_X1 U8577 ( .A1(n9259), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9435) );
  INV_X1 U8578 ( .A(n9427), .ZN(n9259) );
  NAND2_X1 U8579 ( .A1(n13571), .A2(n13570), .ZN(n9690) );
  XNOR2_X1 U8580 ( .A(n6683), .B(n11094), .ZN(n9581) );
  INV_X1 U8581 ( .A(n10024), .ZN(n9984) );
  NAND2_X1 U8582 ( .A1(n7910), .A2(n7329), .ZN(n10254) );
  AND2_X1 U8583 ( .A1(n7332), .A2(n7330), .ZN(n7329) );
  NOR2_X1 U8584 ( .A1(n7982), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n7991) );
  NOR2_X1 U8585 ( .A1(n11843), .A2(n6826), .ZN(n11846) );
  NOR2_X1 U8586 ( .A1(n11846), .A2(n11845), .ZN(n13675) );
  XNOR2_X1 U8587 ( .A(n13676), .B(n13684), .ZN(n15287) );
  NOR2_X1 U8588 ( .A1(n13675), .A2(n7341), .ZN(n13676) );
  AND2_X1 U8589 ( .A1(n13681), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7341) );
  NOR2_X1 U8590 ( .A1(n13702), .A2(n7335), .ZN(n15301) );
  AND2_X1 U8591 ( .A1(n13703), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U8592 ( .A1(n15301), .A2(n15300), .ZN(n15299) );
  INV_X1 U8593 ( .A(n7333), .ZN(n13712) );
  INV_X1 U8594 ( .A(n13551), .ZN(n13447) );
  OR2_X1 U8595 ( .A1(n13763), .A2(n7537), .ZN(n7267) );
  INV_X1 U8596 ( .A(n7265), .ZN(n7264) );
  OAI21_X1 U8597 ( .B1(n7537), .B2(n9556), .A(n14882), .ZN(n7265) );
  NOR2_X1 U8598 ( .A1(n9480), .A2(n13451), .ZN(n13745) );
  AOI21_X1 U8599 ( .B1(n14095), .B2(n8061), .A(n8060), .ZN(n13748) );
  NAND2_X1 U8600 ( .A1(n9556), .A2(n9493), .ZN(n13756) );
  INV_X1 U8601 ( .A(n7355), .ZN(n13778) );
  AND2_X1 U8602 ( .A1(n7555), .A2(n6809), .ZN(n7553) );
  NAND2_X1 U8603 ( .A1(n13827), .A2(n7354), .ZN(n13785) );
  NAND2_X1 U8604 ( .A1(n13827), .A2(n14059), .ZN(n13807) );
  OR2_X1 U8605 ( .A1(n13804), .A2(n7556), .ZN(n7460) );
  NAND2_X1 U8606 ( .A1(n7359), .A2(n7358), .ZN(n13873) );
  INV_X1 U8607 ( .A(n7359), .ZN(n13888) );
  AOI21_X1 U8608 ( .B1(n13947), .B2(n7270), .A(n6781), .ZN(n7268) );
  OR2_X1 U8609 ( .A1(n13952), .A2(n13959), .ZN(n13953) );
  NAND2_X1 U8610 ( .A1(n14890), .A2(n14899), .ZN(n13952) );
  AOI21_X1 U8611 ( .B1(n14879), .B2(n7273), .A(n7272), .ZN(n11983) );
  AND2_X1 U8612 ( .A1(n14889), .A2(n7274), .ZN(n7272) );
  OR2_X1 U8613 ( .A1(n14889), .A2(n7274), .ZN(n7273) );
  NOR2_X2 U8614 ( .A1(n11821), .A2(n14889), .ZN(n14890) );
  OAI21_X1 U8615 ( .B1(n9360), .B2(n7445), .A(n7443), .ZN(n14887) );
  INV_X1 U8616 ( .A(n7446), .ZN(n7445) );
  AOI21_X1 U8617 ( .B1(n7446), .B2(n7444), .A(n6766), .ZN(n7443) );
  NOR2_X1 U8618 ( .A1(n9376), .A2(n7451), .ZN(n7446) );
  INV_X1 U8619 ( .A(n9370), .ZN(n9257) );
  OR2_X1 U8620 ( .A1(n9362), .A2(n9361), .ZN(n9370) );
  NAND2_X1 U8621 ( .A1(n11794), .A2(n14916), .ZN(n11822) );
  OR2_X1 U8622 ( .A1(n9345), .A2(n9255), .ZN(n9352) );
  INV_X1 U8623 ( .A(n7257), .ZN(n7256) );
  OAI21_X1 U8624 ( .B1(n7258), .B2(n9524), .A(n9526), .ZN(n7257) );
  NOR2_X1 U8625 ( .A1(n11519), .A2(n11737), .ZN(n11606) );
  NAND2_X1 U8626 ( .A1(n7345), .A2(n7344), .ZN(n11519) );
  INV_X1 U8627 ( .A(n11435), .ZN(n7345) );
  AND2_X1 U8628 ( .A1(n11234), .A2(n11244), .ZN(n11294) );
  NAND2_X1 U8629 ( .A1(n11294), .A2(n15391), .ZN(n11435) );
  NAND2_X1 U8630 ( .A1(n7263), .A2(n7262), .ZN(n11288) );
  AND2_X1 U8631 ( .A1(n11284), .A2(n6696), .ZN(n7262) );
  NAND2_X1 U8632 ( .A1(n6906), .A2(n6862), .ZN(n6865) );
  NOR2_X1 U8633 ( .A1(n6863), .A2(n9309), .ZN(n6862) );
  OAI21_X1 U8634 ( .B1(n11092), .B2(n11091), .A(n6882), .ZN(n10420) );
  NAND2_X1 U8635 ( .A1(n10380), .A2(n15366), .ZN(n6882) );
  AOI21_X1 U8636 ( .B1(n9738), .B2(n10037), .A(n8116), .ZN(n10459) );
  INV_X1 U8637 ( .A(n13751), .ZN(n7261) );
  NAND2_X1 U8638 ( .A1(n7886), .A2(n7885), .ZN(n13980) );
  INV_X1 U8639 ( .A(n15370), .ZN(n14043) );
  NAND2_X1 U8640 ( .A1(n9360), .A2(n9359), .ZN(n11792) );
  NAND2_X1 U8641 ( .A1(n6917), .A2(n6914), .ZN(n8084) );
  NAND2_X1 U8642 ( .A1(n6916), .A2(n6915), .ZN(n6914) );
  XNOR2_X1 U8643 ( .A(n8076), .B(n8075), .ZN(n10263) );
  NAND2_X1 U8644 ( .A1(n8022), .A2(n7737), .ZN(n7740) );
  INV_X1 U8645 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7940) );
  INV_X1 U8646 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U8647 ( .A1(n6671), .A2(SI_0_), .ZN(n8241) );
  INV_X1 U8648 ( .A(n11636), .ZN(n7646) );
  AND2_X1 U8649 ( .A1(n14239), .A2(n7665), .ZN(n7664) );
  OR2_X1 U8650 ( .A1(n14175), .A2(n7666), .ZN(n7665) );
  INV_X1 U8651 ( .A(n12753), .ZN(n7666) );
  INV_X1 U8652 ( .A(n12138), .ZN(n12148) );
  OR2_X1 U8653 ( .A1(n10985), .A2(n10984), .ZN(n10997) );
  INV_X1 U8654 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10996) );
  XNOR2_X1 U8655 ( .A(n7051), .B(n6708), .ZN(n10607) );
  NAND2_X1 U8656 ( .A1(n11546), .A2(n10603), .ZN(n7052) );
  OR2_X1 U8657 ( .A1(n10997), .A2(n10996), .ZN(n11008) );
  NAND2_X1 U8658 ( .A1(n11545), .A2(n15091), .ZN(n10590) );
  NOR2_X1 U8659 ( .A1(n14169), .A2(n7679), .ZN(n7678) );
  INV_X1 U8660 ( .A(n12652), .ZN(n7679) );
  XNOR2_X1 U8661 ( .A(n11022), .B(n11021), .ZN(n7673) );
  AND2_X1 U8662 ( .A1(n11711), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U8663 ( .A1(n14934), .A2(n7755), .ZN(n12679) );
  OR2_X1 U8664 ( .A1(n12675), .A2(n12674), .ZN(n7755) );
  AND4_X1 U8665 ( .A1(n10977), .A2(n10976), .A3(n10975), .A4(n10974), .ZN(
        n11634) );
  NAND2_X1 U8666 ( .A1(n6680), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10584) );
  OR2_X1 U8667 ( .A1(n10124), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n10140) );
  OR2_X1 U8668 ( .A1(n10493), .A2(n10494), .ZN(n7201) );
  OR2_X1 U8669 ( .A1(n10533), .A2(n10534), .ZN(n7199) );
  OR2_X1 U8670 ( .A1(n10475), .A2(n10476), .ZN(n7197) );
  OR2_X1 U8671 ( .A1(n10506), .A2(n10507), .ZN(n7195) );
  OR2_X1 U8672 ( .A1(n11036), .A2(n11037), .ZN(n7177) );
  XNOR2_X1 U8673 ( .A(n11743), .B(n15056), .ZN(n15052) );
  AND2_X1 U8674 ( .A1(n7177), .A2(n7176), .ZN(n11743) );
  NAND2_X1 U8675 ( .A1(n11742), .A2(n15012), .ZN(n7176) );
  NAND2_X1 U8676 ( .A1(n15052), .A2(n15051), .ZN(n15050) );
  NAND2_X1 U8677 ( .A1(n7047), .A2(n7045), .ZN(n12186) );
  NAND2_X1 U8678 ( .A1(n14760), .A2(n7046), .ZN(n7045) );
  OR2_X1 U8679 ( .A1(n10952), .A2(n7048), .ZN(n7047) );
  NAND2_X1 U8680 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n7048) );
  INV_X1 U8681 ( .A(n7239), .ZN(n7238) );
  OAI21_X1 U8682 ( .B1(n14483), .B2(n7240), .A(n7488), .ZN(n7239) );
  NAND2_X1 U8683 ( .A1(n14673), .A2(n14447), .ZN(n7488) );
  INV_X1 U8684 ( .A(n6712), .ZN(n7240) );
  OR2_X1 U8685 ( .A1(n14497), .A2(n14505), .ZN(n7175) );
  XNOR2_X1 U8686 ( .A(n14467), .B(n14471), .ZN(n6971) );
  NAND2_X1 U8687 ( .A1(n14482), .A2(n6712), .ZN(n14467) );
  OR2_X1 U8688 ( .A1(n14468), .A2(n15097), .ZN(n6969) );
  NAND2_X1 U8689 ( .A1(n14528), .A2(n6746), .ZN(n14515) );
  NAND2_X1 U8690 ( .A1(n14520), .A2(n14444), .ZN(n14503) );
  INV_X1 U8691 ( .A(n14445), .ZN(n14514) );
  NAND2_X1 U8692 ( .A1(n7324), .A2(n7323), .ZN(n14547) );
  INV_X1 U8693 ( .A(n14442), .ZN(n14544) );
  NAND2_X1 U8694 ( .A1(n6973), .A2(n6800), .ZN(n6972) );
  NAND2_X1 U8695 ( .A1(n14582), .A2(n6975), .ZN(n6974) );
  INV_X1 U8696 ( .A(n7138), .ZN(n6973) );
  OAI21_X1 U8697 ( .B1(n14593), .B2(n7162), .A(n7006), .ZN(n14555) );
  INV_X1 U8698 ( .A(n7007), .ZN(n7006) );
  OAI21_X1 U8699 ( .B1(n7165), .B2(n7163), .A(n7160), .ZN(n7007) );
  NAND2_X1 U8700 ( .A1(n14555), .A2(n14427), .ZN(n14554) );
  NAND2_X1 U8701 ( .A1(n7011), .A2(n7325), .ZN(n14614) );
  NOR2_X1 U8702 ( .A1(n14727), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U8703 ( .A1(n14619), .A2(n7327), .ZN(n7326) );
  INV_X1 U8704 ( .A(n7328), .ZN(n7327) );
  NOR3_X1 U8705 ( .A1(n14727), .A2(n14647), .A3(n7328), .ZN(n14631) );
  NOR2_X1 U8706 ( .A1(n12096), .A2(n12095), .ZN(n12121) );
  NAND2_X1 U8707 ( .A1(n14732), .A2(n14434), .ZN(n14626) );
  INV_X1 U8708 ( .A(n12214), .ZN(n10895) );
  OR2_X1 U8709 ( .A1(n11935), .A2(n11934), .ZN(n12096) );
  NAND2_X1 U8710 ( .A1(n11924), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11935) );
  INV_X1 U8711 ( .A(n7011), .ZN(n14647) );
  NOR2_X1 U8712 ( .A1(n14647), .A2(n14951), .ZN(n14742) );
  NAND2_X1 U8713 ( .A1(n6824), .A2(n7312), .ZN(n11951) );
  NAND2_X1 U8714 ( .A1(n7313), .A2(n14258), .ZN(n6982) );
  INV_X1 U8715 ( .A(n12112), .ZN(n11719) );
  NOR2_X1 U8716 ( .A1(n11008), .A2(n11007), .ZN(n11461) );
  NAND2_X1 U8717 ( .A1(n11268), .A2(n6730), .ZN(n7505) );
  NAND2_X1 U8718 ( .A1(n7509), .A2(n7137), .ZN(n7506) );
  NAND2_X1 U8719 ( .A1(n6727), .A2(n12106), .ZN(n7137) );
  NAND2_X1 U8720 ( .A1(n15174), .A2(n14266), .ZN(n7490) );
  NAND2_X1 U8721 ( .A1(n11367), .A2(n7491), .ZN(n6980) );
  NAND2_X1 U8722 ( .A1(n12242), .A2(n12241), .ZN(n7491) );
  NAND2_X1 U8723 ( .A1(n15078), .A2(n15180), .ZN(n15076) );
  AND4_X1 U8724 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n12235) );
  NAND2_X1 U8725 ( .A1(n15086), .A2(n10889), .ZN(n11393) );
  INV_X1 U8726 ( .A(n15091), .ZN(n15096) );
  NAND2_X1 U8727 ( .A1(n11227), .A2(n11226), .ZN(n14458) );
  NAND2_X1 U8728 ( .A1(n12164), .A2(n12163), .ZN(n14661) );
  AOI21_X1 U8729 ( .B1(n14515), .B2(n14445), .A(n7300), .ZN(n14487) );
  AND2_X1 U8730 ( .A1(n14507), .A2(n14524), .ZN(n7300) );
  AND2_X1 U8731 ( .A1(n14599), .A2(n14598), .ZN(n14717) );
  NAND2_X1 U8732 ( .A1(n7492), .A2(n7496), .ZN(n14597) );
  OR2_X1 U8733 ( .A1(n14732), .A2(n7497), .ZN(n7492) );
  NAND2_X1 U8734 ( .A1(n7498), .A2(n7501), .ZN(n14610) );
  NAND2_X1 U8735 ( .A1(n14732), .A2(n7502), .ZN(n7498) );
  XNOR2_X1 U8736 ( .A(n8058), .B(n8057), .ZN(n14095) );
  OAI21_X1 U8737 ( .B1(n7884), .B2(n7849), .A(n7848), .ZN(n8054) );
  XNOR2_X1 U8738 ( .A(n8050), .B(n8049), .ZN(n14105) );
  NAND2_X1 U8739 ( .A1(n7028), .A2(n7027), .ZN(n10067) );
  NOR2_X1 U8740 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7027) );
  INV_X1 U8741 ( .A(n10187), .ZN(n7028) );
  NAND2_X1 U8742 ( .A1(n7067), .A2(n7071), .ZN(n7074) );
  NAND2_X1 U8743 ( .A1(n8034), .A2(n7824), .ZN(n7067) );
  NOR2_X1 U8744 ( .A1(n10055), .A2(n7685), .ZN(n10952) );
  NAND2_X1 U8745 ( .A1(n7545), .A2(n7813), .ZN(n8012) );
  NAND2_X1 U8746 ( .A1(n7997), .A2(n7550), .ZN(n7545) );
  AND2_X1 U8747 ( .A1(n7593), .A2(n7670), .ZN(n7486) );
  NAND2_X1 U8748 ( .A1(n7540), .A2(n7795), .ZN(n7972) );
  NAND2_X1 U8749 ( .A1(n7965), .A2(n7793), .ZN(n7540) );
  OAI21_X1 U8750 ( .B1(n7282), .B2(n7952), .A(n7246), .ZN(n7959) );
  NAND2_X1 U8751 ( .A1(n7282), .A2(n7787), .ZN(n7953) );
  NAND2_X1 U8752 ( .A1(n7669), .A2(n10043), .ZN(n10105) );
  INV_X1 U8753 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10090) );
  AND2_X1 U8754 ( .A1(n7534), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8864) );
  INV_X1 U8755 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7534) );
  XNOR2_X1 U8756 ( .A(n7533), .B(n8863), .ZN(n8866) );
  INV_X1 U8757 ( .A(n8864), .ZN(n7533) );
  XNOR2_X1 U8758 ( .A(n8821), .B(n7083), .ZN(n8873) );
  INV_X1 U8759 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7083) );
  INV_X1 U8760 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U8761 ( .A1(n6850), .A2(n8827), .ZN(n8882) );
  NAND2_X1 U8762 ( .A1(n8877), .A2(n8878), .ZN(n6850) );
  NOR2_X1 U8763 ( .A1(n14793), .A2(n8885), .ZN(n8887) );
  AND2_X1 U8764 ( .A1(n6848), .A2(n6847), .ZN(n8893) );
  NAND2_X1 U8765 ( .A1(n8833), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n6847) );
  OR2_X1 U8766 ( .A1(n8860), .A2(n8859), .ZN(n6848) );
  NAND2_X1 U8767 ( .A1(n6846), .A2(n8838), .ZN(n8858) );
  NAND2_X1 U8768 ( .A1(n8895), .A2(n8837), .ZN(n6846) );
  AND2_X1 U8769 ( .A1(n6845), .A2(n6844), .ZN(n8899) );
  NAND2_X1 U8770 ( .A1(n8839), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n6844) );
  OR2_X1 U8771 ( .A1(n8858), .A2(n8857), .ZN(n6845) );
  OAI22_X1 U8772 ( .A1(n8901), .A2(n8842), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n8900), .ZN(n8855) );
  OR2_X1 U8773 ( .A1(n8261), .A2(n10085), .ZN(n8319) );
  NAND2_X1 U8774 ( .A1(n7709), .A2(n7706), .ZN(n12781) );
  INV_X1 U8775 ( .A(n7708), .ZN(n7706) );
  AND2_X1 U8776 ( .A1(n8580), .A2(n8579), .ZN(n13145) );
  INV_X1 U8777 ( .A(n12791), .ZN(n12870) );
  NAND2_X1 U8778 ( .A1(n12867), .A2(n6927), .ZN(n12792) );
  NAND2_X1 U8779 ( .A1(n7693), .A2(n7699), .ZN(n12816) );
  INV_X2 U8780 ( .A(n8728), .ZN(n7688) );
  INV_X1 U8781 ( .A(n6937), .ZN(n12615) );
  NAND2_X1 U8782 ( .A1(n7714), .A2(n8775), .ZN(n12832) );
  AOI22_X1 U8783 ( .A1(n8757), .A2(n12933), .B1(n8756), .B2(n13275), .ZN(
        n12852) );
  NAND2_X1 U8784 ( .A1(n12852), .A2(n12851), .ZN(n12850) );
  NAND2_X1 U8785 ( .A1(n12850), .A2(n8760), .ZN(n12859) );
  INV_X1 U8786 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U8787 ( .A1(n10670), .A2(n8733), .ZN(n10849) );
  OR2_X1 U8788 ( .A1(n7228), .A2(n7231), .ZN(n11324) );
  INV_X1 U8789 ( .A(n7230), .ZN(n7228) );
  AOI21_X1 U8790 ( .B1(n11859), .B2(n11860), .A(n6693), .ZN(n12891) );
  NAND2_X1 U8791 ( .A1(n8781), .A2(n8782), .ZN(n12903) );
  NAND2_X1 U8792 ( .A1(n8548), .A2(n8547), .ZN(n13165) );
  OR2_X1 U8793 ( .A1(n12415), .A2(n8546), .ZN(n8547) );
  INV_X1 U8794 ( .A(n8749), .ZN(n8747) );
  NAND2_X1 U8795 ( .A1(n10555), .A2(n10556), .ZN(n10669) );
  NAND2_X1 U8796 ( .A1(n12612), .A2(n8727), .ZN(n10555) );
  INV_X1 U8797 ( .A(n12896), .ZN(n12938) );
  NAND2_X1 U8798 ( .A1(n6925), .A2(n8764), .ZN(n12912) );
  INV_X1 U8799 ( .A(n12941), .ZN(n12914) );
  AND2_X1 U8800 ( .A1(n8595), .A2(n8594), .ZN(n13130) );
  AND2_X1 U8801 ( .A1(n8799), .A2(n8801), .ZN(n12936) );
  INV_X1 U8802 ( .A(n12931), .ZN(n12943) );
  AND2_X1 U8803 ( .A1(n10882), .A2(n8212), .ZN(n13072) );
  NAND2_X1 U8804 ( .A1(n8624), .A2(n8623), .ZN(n12928) );
  NAND2_X1 U8805 ( .A1(n8608), .A2(n8607), .ZN(n13116) );
  INV_X1 U8806 ( .A(n13130), .ZN(n12874) );
  INV_X1 U8807 ( .A(n13145), .ZN(n13115) );
  INV_X1 U8808 ( .A(n13175), .ZN(n13204) );
  INV_X1 U8809 ( .A(n7363), .ZN(n7362) );
  OR2_X1 U8810 ( .A1(n8243), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8255) );
  NOR2_X1 U8811 ( .A1(n7020), .A2(n7019), .ZN(n7018) );
  OR2_X1 U8812 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  AOI22_X1 U8813 ( .A1(n8639), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n8224), .B2(
        P3_REG1_REG_2__SCAN_IN), .ZN(n6885) );
  OR2_X1 U8814 ( .A1(n8245), .A2(n8222), .ZN(n8228) );
  OAI21_X1 U8815 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7105), .ZN(n7104) );
  AND2_X1 U8816 ( .A1(n7103), .A2(n7102), .ZN(n7101) );
  AND2_X1 U8817 ( .A1(n7106), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7105) );
  INV_X1 U8818 ( .A(n7478), .ZN(n11119) );
  INV_X1 U8819 ( .A(n15508), .ZN(n15439) );
  XNOR2_X1 U8820 ( .A(n11121), .B(n7476), .ZN(n15433) );
  INV_X1 U8821 ( .A(n7113), .ZN(n15449) );
  INV_X1 U8822 ( .A(n7115), .ZN(n15451) );
  XNOR2_X1 U8823 ( .A(n11123), .B(n11153), .ZN(n15469) );
  OAI21_X1 U8824 ( .B1(n15504), .B2(n7465), .A(n7464), .ZN(n11373) );
  NAND2_X1 U8825 ( .A1(n7466), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U8826 ( .A1(n11126), .A2(n7466), .ZN(n7464) );
  XNOR2_X1 U8827 ( .A(n11558), .B(n11572), .ZN(n11375) );
  NOR2_X1 U8828 ( .A1(n11375), .A2(n8374), .ZN(n11559) );
  OAI21_X1 U8829 ( .B1(n11375), .B2(n7480), .A(n7479), .ZN(n11894) );
  NAND2_X1 U8830 ( .A1(n7481), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7480) );
  NAND2_X1 U8831 ( .A1(n11560), .A2(n7481), .ZN(n7479) );
  INV_X1 U8832 ( .A(n11562), .ZN(n7481) );
  NAND2_X1 U8833 ( .A1(n12959), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U8834 ( .A1(n12962), .A2(n12967), .ZN(n12984) );
  NOR2_X1 U8835 ( .A1(n12953), .A2(n12954), .ZN(n12956) );
  NOR2_X1 U8836 ( .A1(n12956), .A2(n12966), .ZN(n12981) );
  XNOR2_X1 U8837 ( .A(n13006), .B(n13020), .ZN(n12985) );
  NOR2_X1 U8838 ( .A1(n12982), .A2(n12983), .ZN(n13003) );
  NAND2_X1 U8839 ( .A1(n7484), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U8840 ( .A1(n13004), .A2(n7484), .ZN(n7482) );
  INV_X1 U8841 ( .A(n13005), .ZN(n7484) );
  INV_X1 U8842 ( .A(n7119), .ZN(n14821) );
  NAND2_X1 U8843 ( .A1(n7366), .A2(n7367), .ZN(n13100) );
  NAND2_X1 U8844 ( .A1(n13171), .A2(n8543), .ZN(n13159) );
  NAND2_X1 U8845 ( .A1(n13193), .A2(n12551), .ZN(n13178) );
  NAND2_X1 U8846 ( .A1(n8657), .A2(n12548), .ZN(n13191) );
  NAND2_X1 U8847 ( .A1(n8525), .A2(n8524), .ZN(n13332) );
  NAND2_X1 U8848 ( .A1(n13200), .A2(n8522), .ZN(n13185) );
  NAND2_X1 U8849 ( .A1(n13237), .A2(n12535), .ZN(n13214) );
  NAND2_X1 U8850 ( .A1(n7422), .A2(n8490), .ZN(n13219) );
  NAND2_X1 U8851 ( .A1(n8495), .A2(n8494), .ZN(n13228) );
  NAND2_X1 U8852 ( .A1(n13257), .A2(n13258), .ZN(n6952) );
  NAND2_X1 U8853 ( .A1(n7372), .A2(n12425), .ZN(n13277) );
  NAND2_X1 U8854 ( .A1(n8373), .A2(n8372), .ZN(n14860) );
  NAND2_X1 U8855 ( .A1(n6945), .A2(n6949), .ZN(n8373) );
  AND2_X1 U8856 ( .A1(n15623), .A2(n15602), .ZN(n13156) );
  INV_X1 U8857 ( .A(n11762), .ZN(n15577) );
  AND2_X1 U8858 ( .A1(n10566), .A2(n13039), .ZN(n15585) );
  INV_X1 U8859 ( .A(n15576), .ZN(n15618) );
  NAND2_X1 U8860 ( .A1(n15577), .A2(n15583), .ZN(n13289) );
  OAI21_X1 U8861 ( .B1(n13435), .B2(n8261), .A(n7421), .ZN(n13365) );
  OR2_X1 U8862 ( .A1(n12415), .A2(n13431), .ZN(n7421) );
  INV_X1 U8863 ( .A(n13078), .ZN(n13375) );
  NAND2_X1 U8864 ( .A1(n8430), .A2(n8429), .ZN(n13418) );
  NAND2_X1 U8865 ( .A1(n8415), .A2(n8414), .ZN(n13422) );
  OAI22_X1 U8866 ( .A1(n10136), .A2(P3_D_REG_0__SCAN_IN), .B1(n8682), .B2(
        n8681), .ZN(n13425) );
  AND2_X1 U8867 ( .A1(n10679), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13426) );
  INV_X1 U8868 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13429) );
  INV_X1 U8869 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U8870 ( .A1(n12413), .A2(n12412), .ZN(n12621) );
  NAND2_X1 U8871 ( .A1(n8180), .A2(n8179), .ZN(n8581) );
  OAI21_X1 U8872 ( .B1(n8545), .B2(n8544), .A(n8177), .ZN(n8559) );
  XNOR2_X1 U8873 ( .A(n8629), .B(n8628), .ZN(n10860) );
  INV_X1 U8874 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U8875 ( .A(n8632), .B(n8631), .ZN(n10813) );
  OR2_X1 U8876 ( .A1(n8630), .A2(n8478), .ZN(n8632) );
  INV_X1 U8877 ( .A(SI_20_), .ZN(n10564) );
  INV_X1 U8878 ( .A(n8707), .ZN(n10566) );
  INV_X1 U8879 ( .A(SI_19_), .ZN(n10308) );
  NAND2_X1 U8880 ( .A1(n7389), .A2(n7393), .ZN(n8475) );
  OR2_X1 U8881 ( .A1(n8458), .A2(n7395), .ZN(n7389) );
  OR2_X1 U8882 ( .A1(n8481), .A2(n8480), .ZN(n13046) );
  INV_X1 U8883 ( .A(SI_15_), .ZN(n10161) );
  INV_X1 U8884 ( .A(SI_13_), .ZN(n10139) );
  INV_X1 U8885 ( .A(SI_12_), .ZN(n10131) );
  INV_X1 U8886 ( .A(n11574), .ZN(n11899) );
  INV_X1 U8887 ( .A(SI_11_), .ZN(n10116) );
  NAND2_X1 U8888 ( .A1(n8317), .A2(n8145), .ZN(n8331) );
  INV_X1 U8889 ( .A(n11160), .ZN(n15493) );
  INV_X1 U8890 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U8891 ( .A1(n7406), .A2(n8141), .ZN(n8299) );
  NAND2_X1 U8892 ( .A1(n8230), .A2(n8189), .ZN(n8271) );
  NAND2_X1 U8893 ( .A1(n7400), .A2(n8134), .ZN(n8260) );
  NAND2_X1 U8894 ( .A1(n8249), .A2(n8248), .ZN(n7400) );
  OAI211_X1 U8895 ( .C1(P3_IR_REG_31__SCAN_IN), .C2(P3_IR_REG_1__SCAN_IN), .A(
        n7485), .B(n7128), .ZN(n10747) );
  XNOR2_X1 U8896 ( .A(n9732), .B(n9731), .ZN(n9740) );
  XNOR2_X1 U8897 ( .A(n9730), .B(n9729), .ZN(n9731) );
  NAND2_X1 U8898 ( .A1(n13445), .A2(n9728), .ZN(n9732) );
  NAND2_X1 U8899 ( .A1(n7727), .A2(n9619), .ZN(n13491) );
  XNOR2_X1 U8900 ( .A(n9581), .B(n9582), .ZN(n10242) );
  OR2_X1 U8901 ( .A1(n12396), .A2(n6733), .ZN(n10241) );
  AND2_X1 U8902 ( .A1(n13596), .A2(n9638), .ZN(n13516) );
  AND2_X1 U8903 ( .A1(n13633), .A2(n9666), .ZN(n13535) );
  NAND2_X1 U8904 ( .A1(n10705), .A2(n9604), .ZN(n10865) );
  NAND2_X1 U8905 ( .A1(n7736), .A2(n9598), .ZN(n10708) );
  AND2_X1 U8906 ( .A1(n7725), .A2(n9622), .ZN(n6995) );
  AND2_X1 U8907 ( .A1(n9659), .A2(n9647), .ZN(n13579) );
  AND2_X1 U8908 ( .A1(n13514), .A2(n9642), .ZN(n13578) );
  NAND2_X1 U8909 ( .A1(n13598), .A2(n13597), .ZN(n13596) );
  NAND2_X1 U8910 ( .A1(n11624), .A2(n9632), .ZN(n13598) );
  AND2_X1 U8911 ( .A1(n9680), .A2(n9674), .ZN(n7741) );
  NAND2_X1 U8912 ( .A1(n13548), .A2(n9674), .ZN(n13607) );
  NAND2_X1 U8913 ( .A1(n10864), .A2(n9610), .ZN(n11201) );
  NAND2_X1 U8914 ( .A1(n13525), .A2(n9717), .ZN(n13620) );
  NAND2_X1 U8915 ( .A1(n9739), .A2(n13957), .ZN(n13628) );
  INV_X1 U8916 ( .A(n11993), .ZN(n14899) );
  NAND2_X1 U8917 ( .A1(n13577), .A2(n7746), .ZN(n6994) );
  INV_X1 U8918 ( .A(n9956), .ZN(n13647) );
  NAND2_X1 U8919 ( .A1(n9477), .A2(n9476), .ZN(n13649) );
  OR2_X1 U8920 ( .A1(n13789), .A2(n9472), .ZN(n9477) );
  CLKBUF_X1 U8921 ( .A(n13673), .Z(n7040) );
  INV_X1 U8922 ( .A(n7337), .ZN(n10334) );
  NOR2_X1 U8923 ( .A1(n10252), .A2(n10251), .ZN(n10276) );
  AND2_X1 U8924 ( .A1(n7337), .A2(n7336), .ZN(n10252) );
  NAND2_X1 U8925 ( .A1(n10344), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7336) );
  NOR2_X1 U8926 ( .A1(n10281), .A2(n10280), .ZN(n10393) );
  NOR2_X1 U8927 ( .A1(n10296), .A2(n7340), .ZN(n10281) );
  AND2_X1 U8928 ( .A1(n10284), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7340) );
  NOR2_X1 U8929 ( .A1(n10393), .A2(n7339), .ZN(n10396) );
  AND2_X1 U8930 ( .A1(n10397), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U8931 ( .A1(n10396), .A2(n10395), .ZN(n11099) );
  NOR2_X1 U8932 ( .A1(n11104), .A2(n11103), .ZN(n11331) );
  NOR2_X1 U8933 ( .A1(n15273), .A2(n7343), .ZN(n11104) );
  AND2_X1 U8934 ( .A1(n11108), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7343) );
  NOR2_X1 U8935 ( .A1(n11331), .A2(n7342), .ZN(n11335) );
  AND2_X1 U8936 ( .A1(n11332), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U8937 ( .A1(n11335), .A2(n11334), .ZN(n11686) );
  AND2_X1 U8938 ( .A1(n8022), .A2(n8021), .ZN(n8029) );
  NOR2_X1 U8939 ( .A1(n10253), .A2(n14104), .ZN(n15307) );
  NOR2_X1 U8940 ( .A1(n10253), .A2(n10250), .ZN(n15265) );
  NAND2_X1 U8941 ( .A1(n13775), .A2(n13774), .ZN(n13977) );
  NAND2_X1 U8942 ( .A1(n7554), .A2(n7555), .ZN(n13801) );
  NAND2_X1 U8943 ( .A1(n7440), .A2(n7441), .ZN(n13824) );
  NAND2_X1 U8944 ( .A1(n13856), .A2(n7442), .ZN(n7440) );
  AND2_X1 U8945 ( .A1(n13854), .A2(n9449), .ZN(n13836) );
  NAND2_X1 U8946 ( .A1(n7898), .A2(n7897), .ZN(n14010) );
  NAND2_X1 U8947 ( .A1(n9434), .A2(n9433), .ZN(n13872) );
  NAND2_X1 U8948 ( .A1(n13930), .A2(n9410), .ZN(n13922) );
  NAND2_X1 U8949 ( .A1(n13950), .A2(n9536), .ZN(n13927) );
  NAND2_X1 U8950 ( .A1(n11992), .A2(n9392), .ZN(n13943) );
  NAND2_X1 U8951 ( .A1(n7447), .A2(n7450), .ZN(n11819) );
  NAND2_X1 U8952 ( .A1(n9360), .A2(n7448), .ZN(n7447) );
  NAND2_X1 U8953 ( .A1(n6906), .A2(n9300), .ZN(n10834) );
  OR2_X1 U8954 ( .A1(n6674), .A2(n10743), .ZN(n13918) );
  OR2_X1 U8955 ( .A1(n10031), .A2(n10256), .ZN(n7000) );
  INV_X1 U8956 ( .A(n13957), .ZN(n15316) );
  INV_X1 U8957 ( .A(n13966), .ZN(n15320) );
  AOI21_X1 U8958 ( .B1(n13974), .B2(n15370), .A(n6910), .ZN(n6909) );
  NAND2_X1 U8959 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  INV_X1 U8960 ( .A(n13973), .ZN(n6911) );
  INV_X1 U8961 ( .A(n13936), .ZN(n14077) );
  AND2_X2 U8962 ( .A1(n8125), .A2(n10457), .ZN(n15420) );
  AND2_X1 U8963 ( .A1(n10035), .A2(n9734), .ZN(n15362) );
  XNOR2_X1 U8964 ( .A(n8107), .B(n7873), .ZN(n14108) );
  AND2_X1 U8965 ( .A1(n8022), .A2(n6702), .ZN(n8068) );
  INV_X1 U8966 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11196) );
  INV_X1 U8967 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10453) );
  INV_X1 U8968 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10552) );
  INV_X1 U8969 ( .A(n15292), .ZN(n13684) );
  INV_X1 U8970 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10438) );
  INV_X1 U8971 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10219) );
  INV_X1 U8972 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10172) );
  INV_X1 U8973 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10167) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10156) );
  INV_X1 U8975 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U8976 ( .A1(n6990), .A2(n6989), .ZN(n7960) );
  INV_X1 U8977 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10146) );
  INV_X1 U8978 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10132) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10128) );
  INV_X1 U8980 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U8981 ( .A1(n14220), .A2(n12733), .ZN(n14123) );
  NOR2_X1 U8982 ( .A1(n11021), .A2(n11023), .ZN(n11024) );
  INV_X1 U8983 ( .A(n11490), .ZN(n6936) );
  NAND2_X1 U8984 ( .A1(n11962), .A2(n7754), .ZN(n11965) );
  NAND2_X1 U8985 ( .A1(n14198), .A2(n12720), .ZN(n14154) );
  NAND2_X1 U8986 ( .A1(n14977), .A2(n12652), .ZN(n14168) );
  NAND2_X1 U8987 ( .A1(n11662), .A2(n11661), .ZN(n14172) );
  AOI21_X1 U8988 ( .B1(n7655), .B2(n6932), .A(n6761), .ZN(n6931) );
  INV_X1 U8989 ( .A(n7655), .ZN(n6933) );
  NAND2_X1 U8990 ( .A1(n12686), .A2(n14247), .ZN(n14947) );
  AOI21_X1 U8991 ( .B1(n11544), .B2(n11543), .A(n11542), .ZN(n11633) );
  OAI21_X1 U8992 ( .B1(n14220), .B2(n7660), .A(n7657), .ZN(n14181) );
  AND2_X1 U8993 ( .A1(n12630), .A2(n12629), .ZN(n14190) );
  NAND2_X1 U8994 ( .A1(n14146), .A2(n12713), .ZN(n14200) );
  OR2_X1 U8995 ( .A1(n14572), .A2(n15204), .ZN(n14707) );
  INV_X1 U8996 ( .A(n7675), .ZN(n11025) );
  INV_X1 U8997 ( .A(n7673), .ZN(n10824) );
  NAND2_X1 U8998 ( .A1(n7024), .A2(n7649), .ZN(n7648) );
  NAND2_X1 U8999 ( .A1(n7024), .A2(n7654), .ZN(n7647) );
  INV_X1 U9000 ( .A(n7654), .ZN(n7653) );
  AND2_X1 U9001 ( .A1(n14118), .A2(n15156), .ZN(n14981) );
  INV_X1 U9002 ( .A(n14985), .ZN(n14244) );
  NAND2_X1 U9003 ( .A1(n7663), .A2(n12753), .ZN(n14238) );
  NAND2_X1 U9004 ( .A1(n14174), .A2(n14175), .ZN(n7663) );
  NAND4_X1 U9005 ( .A1(n10630), .A2(n10944), .A3(n11224), .A4(n10627), .ZN(
        n14976) );
  INV_X1 U9006 ( .A(n14976), .ZN(n14965) );
  INV_X1 U9007 ( .A(n7058), .ZN(n7057) );
  NAND2_X1 U9008 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  INV_X1 U9009 ( .A(n12374), .ZN(n7055) );
  CLKBUF_X2 U9010 ( .A(P1_U4016), .Z(n14285) );
  NAND2_X1 U9011 ( .A1(n14275), .A2(n14274), .ZN(n14273) );
  NOR2_X1 U9012 ( .A1(n10354), .A2(n10355), .ZN(n10467) );
  NAND2_X1 U9013 ( .A1(n14316), .A2(n7189), .ZN(n10354) );
  OR2_X1 U9014 ( .A1(n10923), .A2(n10353), .ZN(n7189) );
  NOR2_X1 U9015 ( .A1(n10467), .A2(n7188), .ZN(n14333) );
  AND2_X1 U9016 ( .A1(n10468), .A2(n15218), .ZN(n7188) );
  NAND2_X1 U9017 ( .A1(n14333), .A2(n14334), .ZN(n14332) );
  INV_X1 U9018 ( .A(n7201), .ZN(n10492) );
  AND2_X1 U9019 ( .A1(n7201), .A2(n7200), .ZN(n10533) );
  NAND2_X1 U9020 ( .A1(n10495), .A2(n10472), .ZN(n7200) );
  INV_X1 U9021 ( .A(n7199), .ZN(n10532) );
  AND2_X1 U9022 ( .A1(n7199), .A2(n7198), .ZN(n10527) );
  NAND2_X1 U9023 ( .A1(n10535), .A2(n10473), .ZN(n7198) );
  INV_X1 U9024 ( .A(n7197), .ZN(n10505) );
  AND2_X1 U9025 ( .A1(n7197), .A2(n7196), .ZN(n10506) );
  NAND2_X1 U9026 ( .A1(n10512), .A2(n15019), .ZN(n7196) );
  INV_X1 U9027 ( .A(n7195), .ZN(n11035) );
  AND2_X1 U9028 ( .A1(n7195), .A2(n7194), .ZN(n14361) );
  NAND2_X1 U9029 ( .A1(n11041), .A2(n11702), .ZN(n7194) );
  INV_X1 U9030 ( .A(n7177), .ZN(n11741) );
  OAI21_X1 U9031 ( .B1(n14397), .B2(n14396), .A(n7206), .ZN(n7205) );
  AOI21_X1 U9032 ( .B1(n14399), .B2(n14400), .A(n14398), .ZN(n7206) );
  OR2_X1 U9033 ( .A1(n14492), .A2(n14407), .ZN(n7314) );
  AOI21_X1 U9034 ( .B1(n14676), .B2(n15072), .A(n14490), .ZN(n7590) );
  NAND2_X1 U9035 ( .A1(n14491), .A2(n14645), .ZN(n7592) );
  NAND2_X1 U9036 ( .A1(n7510), .A2(n7511), .ZN(n14556) );
  NAND2_X1 U9037 ( .A1(n7164), .A2(n7169), .ZN(n14570) );
  NAND2_X1 U9038 ( .A1(n14593), .A2(n7167), .ZN(n7164) );
  NAND2_X1 U9039 ( .A1(n14582), .A2(n14439), .ZN(n7515) );
  NAND2_X1 U9040 ( .A1(n14593), .A2(n14425), .ZN(n14580) );
  NAND2_X1 U9041 ( .A1(n12064), .A2(n12063), .ZN(n14714) );
  NOR2_X1 U9042 ( .A1(n7560), .A2(n7559), .ZN(n14594) );
  INV_X1 U9043 ( .A(n14423), .ZN(n7559) );
  INV_X1 U9044 ( .A(n14424), .ZN(n7560) );
  NAND2_X1 U9045 ( .A1(n7303), .A2(n14420), .ZN(n14624) );
  NAND2_X1 U9046 ( .A1(n14651), .A2(n7304), .ZN(n7303) );
  NAND2_X1 U9047 ( .A1(n14651), .A2(n14418), .ZN(n14731) );
  AND2_X1 U9048 ( .A1(n6978), .A2(n14431), .ZN(n14640) );
  NAND2_X1 U9049 ( .A1(n7147), .A2(n14417), .ZN(n14653) );
  NAND2_X1 U9050 ( .A1(n11948), .A2(n7580), .ZN(n7147) );
  NAND2_X1 U9051 ( .A1(n11948), .A2(n11919), .ZN(n14414) );
  NAND2_X1 U9052 ( .A1(n7291), .A2(n11675), .ZN(n11676) );
  NAND2_X1 U9053 ( .A1(n7292), .A2(n7763), .ZN(n7291) );
  NAND2_X1 U9054 ( .A1(n11457), .A2(n11456), .ZN(n15013) );
  INV_X1 U9055 ( .A(n12106), .ZN(n7286) );
  AND2_X1 U9056 ( .A1(n7507), .A2(n6727), .ZN(n11475) );
  NAND2_X1 U9057 ( .A1(n11268), .A2(n12105), .ZN(n7507) );
  OR2_X1 U9058 ( .A1(n14458), .A2(n14401), .ZN(n14577) );
  AND2_X1 U9059 ( .A1(n11218), .A2(n11217), .ZN(n15099) );
  INV_X1 U9060 ( .A(n15106), .ZN(n15074) );
  INV_X2 U9061 ( .A(n15103), .ZN(n15112) );
  NAND2_X1 U9062 ( .A1(n14481), .A2(n14675), .ZN(n14748) );
  INV_X1 U9063 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U9064 ( .A1(n14761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7558) );
  XNOR2_X1 U9065 ( .A(n8054), .B(n8053), .ZN(n14769) );
  INV_X1 U9066 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10052) );
  NAND3_X1 U9067 ( .A1(n10051), .A2(n12177), .A3(n10053), .ZN(n7676) );
  XNOR2_X1 U9068 ( .A(n7893), .B(n7892), .ZN(n12144) );
  XNOR2_X1 U9069 ( .A(n7243), .B(n7242), .ZN(n14782) );
  INV_X1 U9070 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7242) );
  NOR2_X1 U9071 ( .A1(n12053), .A2(n6673), .ZN(n7243) );
  INV_X1 U9072 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12074) );
  INV_X1 U9073 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12117) );
  INV_X1 U9074 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10436) );
  INV_X1 U9075 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10550) );
  INV_X1 U9076 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10441) );
  INV_X1 U9077 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10317) );
  INV_X1 U9078 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10179) );
  INV_X1 U9079 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10165) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10158) );
  INV_X1 U9081 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10153) );
  INV_X1 U9082 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10144) );
  INV_X1 U9083 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10134) );
  INV_X1 U9084 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10126) );
  XNOR2_X1 U9085 ( .A(n7934), .B(n7933), .ZN(n10109) );
  NAND2_X1 U9086 ( .A1(n7297), .A2(n7779), .ZN(n7934) );
  XNOR2_X1 U9087 ( .A(n7919), .B(n7920), .ZN(n10822) );
  XNOR2_X1 U9088 ( .A(n7208), .B(n10102), .ZN(n10595) );
  NAND2_X1 U9089 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7208) );
  XNOR2_X1 U9090 ( .A(n8866), .B(n7532), .ZN(n15701) );
  XNOR2_X1 U9091 ( .A(n8884), .B(n7088), .ZN(n14794) );
  NOR2_X1 U9092 ( .A1(n14794), .A2(n14795), .ZN(n14793) );
  XNOR2_X1 U9093 ( .A(n8887), .B(n7524), .ZN(n15694) );
  NOR2_X1 U9094 ( .A1(n8891), .A2(n14796), .ZN(n14801) );
  NOR2_X1 U9095 ( .A1(n8904), .A2(n8903), .ZN(n15034) );
  NOR2_X1 U9096 ( .A1(n7095), .A2(n7094), .ZN(n8904) );
  AND3_X1 U9097 ( .A1(n7518), .A2(n7519), .A3(n7517), .ZN(n7094) );
  NAND2_X1 U9098 ( .A1(n15030), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U9099 ( .A1(n7089), .A2(n7091), .ZN(n15036) );
  NOR2_X1 U9100 ( .A1(n7093), .A2(n7092), .ZN(n7091) );
  INV_X1 U9101 ( .A(n7096), .ZN(n7092) );
  OAI21_X1 U9102 ( .B1(n13378), .B2(n12931), .A(n8816), .ZN(n8817) );
  AOI21_X1 U9103 ( .B1(n7227), .B2(n12924), .A(n7224), .ZN(n12848) );
  NAND2_X1 U9104 ( .A1(n7226), .A2(n7225), .ZN(n7224) );
  NAND2_X1 U9105 ( .A1(n7116), .A2(n14837), .ZN(n14840) );
  NAND2_X1 U9106 ( .A1(n7123), .A2(n15519), .ZN(n7122) );
  INV_X1 U9107 ( .A(n7126), .ZN(n7125) );
  AOI21_X1 U9108 ( .B1(n8700), .B2(n7038), .A(n8702), .ZN(n8703) );
  NAND2_X1 U9109 ( .A1(n6940), .A2(n6705), .ZN(P3_U3487) );
  INV_X1 U9110 ( .A(n7377), .ZN(n7376) );
  OAI22_X1 U9111 ( .A1(n13378), .A2(n13364), .B1(n15685), .B2(n13305), .ZN(
        n7377) );
  OAI21_X1 U9112 ( .B1(n13373), .B2(n15672), .A(n7025), .ZN(P3_U3455) );
  INV_X1 U9113 ( .A(n7026), .ZN(n7025) );
  OAI22_X1 U9114 ( .A1(n13375), .A2(n13423), .B1(n15670), .B2(n13374), .ZN(
        n7026) );
  OAI21_X1 U9115 ( .B1(n13376), .B2(n15672), .A(n7029), .ZN(P3_U3454) );
  AOI21_X1 U9116 ( .B1(n8797), .B2(n8719), .A(n7030), .ZN(n7029) );
  NOR2_X1 U9117 ( .A1(n15670), .A2(n13377), .ZN(n7030) );
  OR2_X1 U9118 ( .A1(n13736), .A2(n14046), .ZN(n7752) );
  AND2_X1 U9119 ( .A1(n9570), .A2(n7456), .ZN(n7455) );
  OR2_X1 U9120 ( .A1(n15431), .A2(n9568), .ZN(n7456) );
  OR2_X1 U9121 ( .A1(n13736), .A2(n14081), .ZN(n7753) );
  AND2_X1 U9122 ( .A1(n9575), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U9123 ( .A1(n7351), .A2(n15420), .ZN(n7259) );
  OR2_X1 U9124 ( .A1(n15420), .A2(n9572), .ZN(n7350) );
  INV_X1 U9125 ( .A(n10214), .ZN(n10069) );
  NAND2_X1 U9126 ( .A1(n7207), .A2(n7203), .ZN(P1_U3262) );
  AOI21_X1 U9127 ( .B1(n7205), .B2(n14401), .A(n7204), .ZN(n7203) );
  OR2_X1 U9128 ( .A1(n14402), .A2(n14401), .ZN(n7207) );
  OAI21_X1 U9129 ( .B1(n15064), .B2(n7766), .A(n14403), .ZN(n7204) );
  NAND2_X1 U9130 ( .A1(n15225), .A2(n15208), .ZN(n7157) );
  OAI21_X1 U9131 ( .B1(n14667), .B2(n15223), .A(n7156), .ZN(n7155) );
  NAND2_X1 U9132 ( .A1(n15212), .A2(n15208), .ZN(n7159) );
  OAI21_X1 U9133 ( .B1(n14667), .B2(n15210), .A(n7158), .ZN(n7154) );
  INV_X1 U9134 ( .A(n7520), .ZN(n14790) );
  INV_X1 U9135 ( .A(n7530), .ZN(n15042) );
  NOR2_X1 U9136 ( .A1(n15048), .A2(n15047), .ZN(n15046) );
  AND2_X1 U9137 ( .A1(n7531), .A2(n7530), .ZN(n15048) );
  NAND2_X1 U9138 ( .A1(n6843), .A2(n14784), .ZN(n14787) );
  OR2_X1 U9139 ( .A1(n14786), .A2(n14785), .ZN(n6843) );
  XNOR2_X1 U9140 ( .A(n7522), .B(n7521), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9141 ( .A(n9250), .B(n8912), .ZN(n7521) );
  NAND2_X1 U9142 ( .A1(n14784), .A2(n7100), .ZN(n7522) );
  AND2_X1 U9143 ( .A1(n12339), .A2(n12341), .ZN(n6689) );
  OR2_X1 U9144 ( .A1(n14416), .A2(n14943), .ZN(n14431) );
  OR2_X1 U9145 ( .A1(n9833), .A2(n9832), .ZN(n6690) );
  OR2_X1 U9146 ( .A1(n9794), .A2(n9793), .ZN(n6691) );
  NOR2_X1 U9147 ( .A1(n14421), .A2(n7568), .ZN(n6692) );
  INV_X1 U9148 ( .A(n11518), .ZN(n7258) );
  NOR2_X1 U9149 ( .A1(n8751), .A2(n14863), .ZN(n6693) );
  INV_X1 U9150 ( .A(n14419), .ZN(n7566) );
  NAND2_X1 U9151 ( .A1(n7306), .A2(n10995), .ZN(n12255) );
  INV_X1 U9152 ( .A(n12255), .ZN(n7013) );
  NAND2_X1 U9153 ( .A1(n14449), .A2(n14645), .ZN(n14668) );
  INV_X1 U9154 ( .A(n14668), .ZN(n7152) );
  AND2_X1 U9155 ( .A1(n15047), .A2(n7529), .ZN(n6694) );
  OR2_X1 U9156 ( .A1(n8370), .A2(n15525), .ZN(n6695) );
  NAND2_X1 U9157 ( .A1(n11244), .A2(n13668), .ZN(n6696) );
  OR2_X1 U9158 ( .A1(n9754), .A2(n13726), .ZN(n6697) );
  AND2_X1 U9159 ( .A1(n8502), .A2(n8490), .ZN(n6698) );
  NOR2_X1 U9160 ( .A1(n8439), .A2(n13276), .ZN(n6699) );
  AND2_X1 U9161 ( .A1(n9549), .A2(n9548), .ZN(n6700) );
  INV_X1 U9162 ( .A(n12338), .ZN(n7181) );
  AND2_X1 U9163 ( .A1(n8782), .A2(n6813), .ZN(n6701) );
  AND2_X1 U9164 ( .A1(n7737), .A2(n8062), .ZN(n6702) );
  AND4_X1 U9165 ( .A1(n7309), .A2(n6981), .A3(n7308), .A4(n7311), .ZN(n6703)
         );
  INV_X1 U9166 ( .A(n11782), .ZN(n12251) );
  AND2_X1 U9167 ( .A1(n10982), .A2(n10981), .ZN(n11782) );
  NAND2_X1 U9168 ( .A1(n12340), .A2(n7579), .ZN(n6704) );
  AND2_X1 U9169 ( .A1(n7037), .A2(n6825), .ZN(n6705) );
  INV_X1 U9170 ( .A(n8797), .ZN(n13378) );
  NAND2_X1 U9171 ( .A1(n8615), .A2(n8614), .ZN(n8797) );
  INV_X1 U9172 ( .A(n6685), .ZN(n9754) );
  XNOR2_X1 U9173 ( .A(n7677), .B(n10052), .ZN(n10209) );
  NAND2_X1 U9174 ( .A1(n11918), .A2(n11917), .ZN(n14938) );
  INV_X1 U9175 ( .A(n14938), .ZN(n7312) );
  AND2_X1 U9176 ( .A1(n9753), .A2(n9752), .ZN(n8090) );
  OR2_X1 U9177 ( .A1(n14770), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6706) );
  AND2_X1 U9178 ( .A1(n12401), .A2(n6706), .ZN(n6707) );
  NAND2_X1 U9179 ( .A1(n10431), .A2(n10433), .ZN(n10055) );
  NAND2_X2 U9180 ( .A1(n8208), .A2(n8207), .ZN(n8243) );
  NAND2_X1 U9181 ( .A1(n15609), .A2(n10447), .ZN(n6937) );
  AND2_X1 U9182 ( .A1(n10896), .A2(n10895), .ZN(n6708) );
  NAND2_X1 U9183 ( .A1(n10681), .A2(n6672), .ZN(n8262) );
  OR2_X1 U9184 ( .A1(n10055), .A2(n7683), .ZN(n10567) );
  AND2_X1 U9185 ( .A1(n6983), .A2(n6982), .ZN(n6709) );
  INV_X1 U9186 ( .A(n7485), .ZN(n8230) );
  AND4_X1 U9187 ( .A1(n12818), .A2(n8738), .A3(n11312), .A4(n8737), .ZN(n6710)
         );
  XNOR2_X1 U9188 ( .A(n9701), .B(n9699), .ZN(n13467) );
  AOI21_X1 U9189 ( .B1(n12377), .B2(n12161), .A(n12160), .ZN(n14660) );
  OR2_X1 U9190 ( .A1(n8674), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n6711) );
  OR2_X1 U9191 ( .A1(n14495), .A2(n14505), .ZN(n6712) );
  NAND2_X1 U9192 ( .A1(n10065), .A2(n10064), .ZN(n10575) );
  NAND2_X1 U9193 ( .A1(n12120), .A2(n12119), .ZN(n14727) );
  AND2_X1 U9194 ( .A1(n8334), .A2(n8321), .ZN(n6713) );
  OR2_X1 U9195 ( .A1(n14709), .A2(n14225), .ZN(n6714) );
  NAND2_X1 U9196 ( .A1(n7080), .A2(n11999), .ZN(n14407) );
  INV_X1 U9197 ( .A(n14407), .ZN(n7319) );
  AND2_X1 U9198 ( .A1(n6695), .A2(n6713), .ZN(n6715) );
  OR2_X1 U9199 ( .A1(n9787), .A2(n9786), .ZN(n6716) );
  OR2_X1 U9200 ( .A1(n9949), .A2(n9948), .ZN(n6717) );
  NOR2_X1 U9201 ( .A1(n14571), .A2(n14562), .ZN(n7324) );
  NAND2_X1 U9202 ( .A1(n11267), .A2(n11266), .ZN(n14192) );
  INV_X1 U9203 ( .A(n10604), .ZN(n12768) );
  INV_X2 U9204 ( .A(n10604), .ZN(n12769) );
  AND2_X1 U9205 ( .A1(n13186), .A2(n12548), .ZN(n6718) );
  NAND2_X1 U9206 ( .A1(n13078), .A2(n10956), .ZN(n6719) );
  OR2_X1 U9207 ( .A1(n12324), .A2(n7589), .ZN(n6720) );
  AND2_X1 U9208 ( .A1(n9592), .A2(n9604), .ZN(n6721) );
  NOR2_X1 U9209 ( .A1(n13877), .A2(n13654), .ZN(n6722) );
  INV_X1 U9210 ( .A(n14420), .ZN(n7568) );
  NAND2_X1 U9211 ( .A1(n8047), .A2(n8046), .ZN(n13811) );
  INV_X1 U9212 ( .A(n15438), .ZN(n7476) );
  OR2_X1 U9213 ( .A1(n13842), .A2(n13652), .ZN(n6723) );
  NAND2_X1 U9214 ( .A1(n7214), .A2(n15556), .ZN(n6724) );
  OR2_X1 U9215 ( .A1(n15044), .A2(n7526), .ZN(n6725) );
  AND2_X1 U9216 ( .A1(n6704), .A2(n7180), .ZN(n6726) );
  NAND2_X1 U9217 ( .A1(n7013), .A2(n14263), .ZN(n6727) );
  NAND2_X1 U9218 ( .A1(n11301), .A2(n8734), .ZN(n6728) );
  INV_X1 U9219 ( .A(n12923), .ZN(n7703) );
  AND2_X1 U9220 ( .A1(n11120), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U9221 ( .A1(n12044), .A2(n12043), .ZN(n14709) );
  NAND2_X1 U9222 ( .A1(n12136), .A2(n12135), .ZN(n14549) );
  INV_X1 U9223 ( .A(n14549), .ZN(n7323) );
  NAND2_X1 U9224 ( .A1(n12031), .A2(n12030), .ZN(n14518) );
  INV_X1 U9225 ( .A(n14518), .ZN(n7321) );
  AND2_X1 U9226 ( .A1(n12105), .A2(n7509), .ZN(n6730) );
  AND3_X1 U9227 ( .A1(n7600), .A2(n9938), .A3(n7599), .ZN(n6731) );
  NAND2_X1 U9228 ( .A1(n13618), .A2(n9721), .ZN(n13443) );
  XNOR2_X1 U9229 ( .A(n8797), .B(n12928), .ZN(n13088) );
  INV_X1 U9230 ( .A(n13088), .ZN(n6944) );
  NAND2_X1 U9231 ( .A1(n12094), .A2(n12093), .ZN(n14991) );
  OR3_X1 U9232 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U9233 ( .A1(n13618), .A2(n7742), .ZN(n13445) );
  AND2_X1 U9234 ( .A1(n6684), .A2(n12400), .ZN(n6733) );
  AND2_X1 U9235 ( .A1(n14189), .A2(n12629), .ZN(n6734) );
  AND2_X1 U9236 ( .A1(n8056), .A2(n8055), .ZN(n14053) );
  INV_X1 U9237 ( .A(n14053), .ZN(n9955) );
  OR2_X1 U9238 ( .A1(n14811), .A2(n13032), .ZN(n6735) );
  AND4_X1 U9239 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n12241) );
  AND2_X1 U9240 ( .A1(n7284), .A2(n12109), .ZN(n6736) );
  AND2_X1 U9241 ( .A1(n7556), .A2(n9553), .ZN(n6737) );
  NOR2_X2 U9242 ( .A1(n8084), .A2(n14084), .ZN(n9264) );
  INV_X1 U9243 ( .A(n9264), .ZN(n14097) );
  NOR2_X1 U9244 ( .A1(n8059), .A2(n10111), .ZN(n6738) );
  AND2_X1 U9245 ( .A1(n9824), .A2(n9823), .ZN(n6739) );
  AND2_X1 U9246 ( .A1(n9836), .A2(n9835), .ZN(n6740) );
  OR2_X1 U9247 ( .A1(n11141), .A2(n15676), .ZN(n6741) );
  OR2_X1 U9248 ( .A1(n10818), .A2(n10595), .ZN(n6742) );
  AND2_X1 U9249 ( .A1(n7252), .A2(n7059), .ZN(n6743) );
  NOR2_X1 U9250 ( .A1(n13003), .A2(n13004), .ZN(n6744) );
  INV_X1 U9251 ( .A(n11795), .ZN(n14916) );
  NAND2_X1 U9252 ( .A1(n7986), .A2(n7985), .ZN(n11795) );
  NOR2_X1 U9253 ( .A1(n11708), .A2(n7290), .ZN(n7289) );
  NOR2_X1 U9254 ( .A1(n12595), .A2(n12422), .ZN(n6745) );
  INV_X1 U9255 ( .A(n14477), .ZN(n14673) );
  NAND2_X1 U9256 ( .A1(n12004), .A2(n12003), .ZN(n14477) );
  OR2_X1 U9257 ( .A1(n7321), .A2(n14538), .ZN(n6746) );
  AND2_X1 U9258 ( .A1(n6926), .A2(n8284), .ZN(n8358) );
  AND2_X1 U9259 ( .A1(n7527), .A2(n6725), .ZN(n6747) );
  AND2_X1 U9260 ( .A1(n9718), .A2(n9717), .ZN(n6748) );
  INV_X1 U9261 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10053) );
  AND2_X1 U9262 ( .A1(n9691), .A2(n9689), .ZN(n6749) );
  AND2_X1 U9263 ( .A1(n12709), .A2(n12704), .ZN(n6750) );
  AND2_X1 U9264 ( .A1(n12722), .A2(n12720), .ZN(n6751) );
  AND2_X1 U9265 ( .A1(n7494), .A2(n14423), .ZN(n6752) );
  INV_X1 U9266 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7532) );
  AND2_X1 U9267 ( .A1(n15180), .A2(n14265), .ZN(n6753) );
  AND2_X1 U9268 ( .A1(n11963), .A2(n7754), .ZN(n6754) );
  AND2_X1 U9269 ( .A1(n8777), .A2(n8775), .ZN(n6755) );
  OR2_X1 U9270 ( .A1(n10083), .A2(SI_1_), .ZN(n6756) );
  AND2_X1 U9271 ( .A1(n13579), .A2(n9642), .ZN(n6757) );
  AND2_X1 U9272 ( .A1(n12849), .A2(n12948), .ZN(n6758) );
  OR2_X1 U9273 ( .A1(n7623), .A2(n9814), .ZN(n6759) );
  INV_X1 U9274 ( .A(n7451), .ZN(n7450) );
  AND2_X1 U9275 ( .A1(n8762), .A2(n8760), .ZN(n6760) );
  AND2_X1 U9276 ( .A1(n12746), .A2(n12745), .ZN(n6761) );
  AND2_X1 U9277 ( .A1(n12760), .A2(n12759), .ZN(n6762) );
  INV_X1 U9278 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10191) );
  INV_X1 U9279 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10568) );
  INV_X1 U9280 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7046) );
  INV_X1 U9281 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7212) );
  AND2_X1 U9282 ( .A1(n13332), .A2(n13204), .ZN(n6763) );
  OR2_X1 U9283 ( .A1(n14072), .A2(n9987), .ZN(n6764) );
  OR2_X1 U9284 ( .A1(n7528), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U9285 ( .A1(n11823), .A2(n13662), .ZN(n6766) );
  AND2_X1 U9286 ( .A1(n7510), .A2(n7138), .ZN(n6767) );
  INV_X1 U9287 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7686) );
  NOR2_X1 U9288 ( .A1(n14172), .A2(n14259), .ZN(n6768) );
  AND2_X1 U9289 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U9290 ( .A1(n14727), .A2(n14957), .ZN(n6770) );
  INV_X1 U9291 ( .A(n7779), .ZN(n7299) );
  INV_X1 U9292 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U9293 ( .A1(n12800), .A2(n8768), .ZN(n6771) );
  INV_X1 U9294 ( .A(n7514), .ZN(n7513) );
  NAND2_X1 U9295 ( .A1(n7516), .A2(n14439), .ZN(n7514) );
  AND2_X1 U9296 ( .A1(n10965), .A2(n10964), .ZN(n15174) );
  AND2_X1 U9297 ( .A1(n15529), .A2(n12507), .ZN(n6772) );
  AND2_X1 U9298 ( .A1(n11707), .A2(n14259), .ZN(n6773) );
  OR2_X1 U9299 ( .A1(n9776), .A2(n9775), .ZN(n6774) );
  AND2_X1 U9300 ( .A1(n7970), .A2(SI_10_), .ZN(n6775) );
  INV_X1 U9301 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10051) );
  AND2_X1 U9302 ( .A1(n8661), .A2(n8660), .ZN(n13076) );
  AND2_X1 U9303 ( .A1(n7815), .A2(n10171), .ZN(n6776) );
  NAND2_X1 U9304 ( .A1(n7457), .A2(n9478), .ZN(n6777) );
  AND2_X1 U9305 ( .A1(n7789), .A2(SI_7_), .ZN(n6778) );
  INV_X1 U9306 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U9307 ( .A1(n7458), .A2(n13799), .ZN(n6779) );
  INV_X1 U9308 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10433) );
  AND2_X1 U9309 ( .A1(n14437), .A2(n12072), .ZN(n14596) );
  INV_X1 U9310 ( .A(n14596), .ZN(n7494) );
  INV_X1 U9311 ( .A(n7384), .ZN(n7383) );
  NAND2_X1 U9312 ( .A1(n14859), .A2(n7385), .ZN(n7384) );
  NAND2_X1 U9313 ( .A1(n10777), .A2(n10780), .ZN(n10776) );
  AND2_X1 U9314 ( .A1(n7323), .A2(n14443), .ZN(n6780) );
  AND2_X1 U9315 ( .A1(n12539), .A2(n12538), .ZN(n13220) );
  INV_X1 U9316 ( .A(n13220), .ZN(n8502) );
  NOR2_X1 U9317 ( .A1(n14077), .A2(n13658), .ZN(n6781) );
  NOR2_X1 U9318 ( .A1(n14673), .A2(n14447), .ZN(n6782) );
  INV_X1 U9319 ( .A(n7606), .ZN(n7605) );
  OAI21_X1 U9320 ( .B1(n7609), .B2(n9933), .A(n9929), .ZN(n7606) );
  NAND2_X1 U9321 ( .A1(n11646), .A2(n15532), .ZN(n6783) );
  OR2_X1 U9322 ( .A1(n6772), .A2(n7419), .ZN(n6784) );
  NAND2_X1 U9323 ( .A1(n12299), .A2(n14435), .ZN(n7501) );
  NAND2_X1 U9324 ( .A1(n14192), .A2(n14138), .ZN(n7509) );
  INV_X1 U9325 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9000) );
  INV_X1 U9326 ( .A(n12336), .ZN(n7183) );
  MUX2_X1 U9327 ( .A(n14504), .B(n14518), .S(n6682), .Z(n12336) );
  INV_X1 U9328 ( .A(n12360), .ZN(n7573) );
  INV_X1 U9329 ( .A(n12277), .ZN(n7578) );
  NAND2_X1 U9330 ( .A1(n7499), .A2(n14609), .ZN(n6785) );
  OR2_X1 U9331 ( .A1(n8871), .A2(n8870), .ZN(n6786) );
  AND2_X1 U9332 ( .A1(n7174), .A2(n14486), .ZN(n6787) );
  AND2_X1 U9333 ( .A1(n7554), .A2(n7553), .ZN(n6788) );
  INV_X1 U9334 ( .A(n14441), .ZN(n14427) );
  OR2_X1 U9335 ( .A1(n6794), .A2(n9779), .ZN(n6789) );
  OR2_X1 U9336 ( .A1(n9799), .A2(n9801), .ZN(n6790) );
  OR2_X1 U9337 ( .A1(n9813), .A2(n9815), .ZN(n6791) );
  AND2_X1 U9338 ( .A1(n7460), .A2(n7459), .ZN(n6792) );
  OR2_X1 U9339 ( .A1(n9838), .A2(n6740), .ZN(n6793) );
  AND2_X1 U9340 ( .A1(n9781), .A2(n9780), .ZN(n6794) );
  AND2_X1 U9341 ( .A1(n7515), .A2(n6714), .ZN(n6795) );
  AND2_X1 U9342 ( .A1(n7074), .A2(n7073), .ZN(n6796) );
  OR2_X1 U9343 ( .A1(n10112), .A2(n8261), .ZN(n6797) );
  INV_X1 U9344 ( .A(n13823), .ZN(n7438) );
  INV_X1 U9345 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14760) );
  AND2_X1 U9346 ( .A1(n6880), .A2(n7713), .ZN(n6798) );
  AND2_X1 U9347 ( .A1(n8654), .A2(n12425), .ZN(n6799) );
  NAND2_X1 U9348 ( .A1(n14562), .A2(n14539), .ZN(n6800) );
  AND2_X1 U9349 ( .A1(n7250), .A2(n7544), .ZN(n6801) );
  AND2_X1 U9350 ( .A1(n6702), .A2(n8069), .ZN(n6802) );
  OR2_X1 U9351 ( .A1(n9912), .A2(n7632), .ZN(n6803) );
  INV_X1 U9352 ( .A(n8142), .ZN(n7405) );
  AND2_X1 U9353 ( .A1(n7537), .A2(n9556), .ZN(n6804) );
  AND2_X1 U9354 ( .A1(n7720), .A2(n8196), .ZN(n6805) );
  OR2_X1 U9355 ( .A1(n7631), .A2(n9913), .ZN(n6806) );
  OR2_X1 U9356 ( .A1(n7629), .A2(n9800), .ZN(n6807) );
  OR2_X1 U9357 ( .A1(n12361), .A2(n12362), .ZN(n6808) );
  INV_X1 U9358 ( .A(n11284), .ZN(n11286) );
  AND2_X1 U9359 ( .A1(n9522), .A2(n9335), .ZN(n11284) );
  NAND2_X1 U9360 ( .A1(n13811), .A2(n9932), .ZN(n6809) );
  INV_X1 U9361 ( .A(n7169), .ZN(n7166) );
  NAND2_X1 U9362 ( .A1(n14438), .A2(n14225), .ZN(n7169) );
  INV_X1 U9363 ( .A(n14429), .ZN(n7174) );
  INV_X1 U9364 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10193) );
  AND2_X1 U9365 ( .A1(n7311), .A2(n10579), .ZN(n6810) );
  AND2_X1 U9366 ( .A1(n8194), .A2(n7212), .ZN(n6811) );
  INV_X1 U9367 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7738) );
  AND2_X1 U9368 ( .A1(n9521), .A2(n11418), .ZN(n6812) );
  INV_X1 U9369 ( .A(n10983), .ZN(n12056) );
  NAND2_X1 U9370 ( .A1(n11706), .A2(n11705), .ZN(n12662) );
  INV_X1 U9371 ( .A(n12662), .ZN(n7313) );
  INV_X1 U9372 ( .A(n15512), .ZN(n11166) );
  OAI21_X1 U9373 ( .B1(n11803), .B2(n12508), .A(n6930), .ZN(n11859) );
  OR2_X1 U9374 ( .A1(n11990), .A2(n11989), .ZN(n11992) );
  NAND2_X1 U9375 ( .A1(n12021), .A2(n12020), .ZN(n14507) );
  INV_X1 U9376 ( .A(n14507), .ZN(n7320) );
  NAND2_X1 U9377 ( .A1(n12912), .A2(n8767), .ZN(n12799) );
  XOR2_X1 U9378 ( .A(n13319), .B(n8787), .Z(n6813) );
  NAND2_X1 U9379 ( .A1(n6878), .A2(n12511), .ZN(n13287) );
  NAND2_X1 U9380 ( .A1(n6952), .A2(n8456), .ZN(n13246) );
  INV_X1 U9381 ( .A(n8756), .ZN(n12932) );
  INV_X1 U9382 ( .A(n8791), .ZN(n7702) );
  NAND2_X1 U9383 ( .A1(n7487), .A2(n7486), .ZN(n6814) );
  NAND2_X1 U9384 ( .A1(n9690), .A2(n9689), .ZN(n13504) );
  NAND2_X1 U9385 ( .A1(n13548), .A2(n7741), .ZN(n13608) );
  NAND2_X1 U9386 ( .A1(n7423), .A2(n8321), .ZN(n11763) );
  NAND2_X1 U9387 ( .A1(n8022), .A2(n7739), .ZN(n8035) );
  NOR2_X1 U9388 ( .A1(n11559), .A2(n11560), .ZN(n6815) );
  AND2_X1 U9389 ( .A1(n8791), .A2(n8790), .ZN(n12843) );
  INV_X1 U9390 ( .A(n12843), .ZN(n6921) );
  AND2_X1 U9391 ( .A1(n7709), .A2(n7707), .ZN(n6816) );
  AND2_X1 U9392 ( .A1(n7291), .A2(n7289), .ZN(n6817) );
  OR2_X1 U9393 ( .A1(n10055), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6818) );
  OR2_X1 U9394 ( .A1(n14053), .A2(n14081), .ZN(n6819) );
  NAND2_X1 U9395 ( .A1(n8555), .A2(n8554), .ZN(n12904) );
  INV_X1 U9396 ( .A(n12904), .ZN(n13176) );
  NAND2_X1 U9397 ( .A1(n7825), .A2(n7073), .ZN(n6820) );
  OR2_X1 U9398 ( .A1(n14469), .A2(n15102), .ZN(n6821) );
  INV_X1 U9399 ( .A(n13161), .ZN(n12873) );
  AND2_X1 U9400 ( .A1(n8568), .A2(n8567), .ZN(n13161) );
  AND2_X1 U9401 ( .A1(n7518), .A2(n7519), .ZN(n6822) );
  AND2_X1 U9402 ( .A1(n7713), .A2(n8230), .ZN(n6823) );
  NAND2_X1 U9403 ( .A1(n10460), .A2(n13957), .ZN(n13963) );
  AND2_X1 U9404 ( .A1(n8013), .A2(n7749), .ZN(n8102) );
  INV_X1 U9405 ( .A(n13364), .ZN(n7038) );
  NAND2_X1 U9406 ( .A1(n7901), .A2(n7900), .ZN(n13877) );
  INV_X1 U9407 ( .A(n13877), .ZN(n7358) );
  NAND2_X1 U9408 ( .A1(n7895), .A2(n7894), .ZN(n13842) );
  INV_X1 U9409 ( .A(n13842), .ZN(n7361) );
  INV_X1 U9410 ( .A(n11989), .ZN(n6913) );
  NOR2_X1 U9411 ( .A1(n11082), .A2(n11081), .ZN(n11080) );
  NAND2_X1 U9412 ( .A1(n8102), .A2(n8103), .ZN(n8099) );
  AND2_X1 U9413 ( .A1(n7015), .A2(n7313), .ZN(n6824) );
  OR2_X1 U9414 ( .A1(n15685), .A2(n13302), .ZN(n6825) );
  NAND2_X1 U9415 ( .A1(n6871), .A2(n9342), .ZN(n11517) );
  OAI21_X1 U9416 ( .B1(n6854), .B2(n6856), .A(n12483), .ZN(n15538) );
  NAND2_X1 U9417 ( .A1(n9525), .A2(n9524), .ZN(n11512) );
  INV_X1 U9418 ( .A(n11255), .ZN(n7014) );
  AND2_X1 U9419 ( .A1(n11849), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6826) );
  NOR2_X1 U9420 ( .A1(n15503), .A2(n11126), .ZN(n6827) );
  NAND2_X1 U9421 ( .A1(n6996), .A2(n7725), .ZN(n11615) );
  INV_X1 U9422 ( .A(n7015), .ZN(n11721) );
  NOR2_X1 U9423 ( .A1(n11672), .A2(n14172), .ZN(n7015) );
  OR2_X1 U9424 ( .A1(n11381), .A2(n11171), .ZN(n6828) );
  INV_X1 U9425 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7088) );
  INV_X1 U9426 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7524) );
  OR2_X1 U9427 ( .A1(n10187), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U9428 ( .A1(n7263), .A2(n6696), .ZN(n6830) );
  AND2_X1 U9429 ( .A1(n15596), .A2(n8253), .ZN(n6831) );
  NAND2_X1 U9430 ( .A1(n8102), .A2(n7637), .ZN(n6832) );
  INV_X1 U9431 ( .A(n10665), .ZN(n12950) );
  INV_X1 U9432 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7097) );
  INV_X1 U9433 ( .A(n15594), .ZN(n15612) );
  AND2_X1 U9434 ( .A1(n10695), .A2(n10694), .ZN(n14837) );
  AND2_X1 U9435 ( .A1(n8795), .A2(n10678), .ZN(n12924) );
  INV_X1 U9436 ( .A(n15431), .ZN(n15429) );
  INV_X1 U9437 ( .A(n10739), .ZN(n13726) );
  INV_X1 U9438 ( .A(n14645), .ZN(n15145) );
  NAND2_X1 U9439 ( .A1(n10629), .A2(n12191), .ZN(n14645) );
  AND2_X1 U9440 ( .A1(n15198), .A2(n15197), .ZN(n15146) );
  NAND2_X1 U9441 ( .A1(n7969), .A2(n7968), .ZN(n15399) );
  INV_X1 U9442 ( .A(n15399), .ZN(n7344) );
  AND2_X1 U9443 ( .A1(n13038), .A2(n7475), .ZN(n6833) );
  OR2_X1 U9444 ( .A1(n11549), .A2(n11548), .ZN(n6834) );
  INV_X1 U9445 ( .A(n6693), .ZN(n7223) );
  INV_X1 U9446 ( .A(n13051), .ZN(n15519) );
  NOR2_X1 U9447 ( .A1(n9752), .A2(n9751), .ZN(n10461) );
  AND2_X1 U9448 ( .A1(n9558), .A2(n9557), .ZN(n13946) );
  INV_X1 U9449 ( .A(n13946), .ZN(n14882) );
  INV_X1 U9450 ( .A(n15587), .ZN(n7689) );
  AND2_X1 U9451 ( .A1(n7472), .A2(n7470), .ZN(n6835) );
  NAND2_X1 U9452 ( .A1(n12455), .A2(n12450), .ZN(n15611) );
  INV_X1 U9453 ( .A(n15611), .ZN(n6939) );
  AND2_X1 U9454 ( .A1(n10670), .A2(n7719), .ZN(n6836) );
  AND2_X1 U9455 ( .A1(n11889), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U9456 ( .A1(n8205), .A2(n8203), .ZN(n13428) );
  NAND2_X1 U9457 ( .A1(n8348), .A2(n8347), .ZN(n6838) );
  AND2_X1 U9458 ( .A1(n14766), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6839) );
  INV_X1 U9459 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7002) );
  INV_X1 U9460 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n8988) );
  INV_X1 U9461 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9033) );
  INV_X1 U9462 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7087) );
  INV_X1 U9463 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7085) );
  INV_X1 U9464 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7099) );
  INV_X1 U9465 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7517) );
  INV_X1 U9466 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7529) );
  INV_X1 U9467 ( .A(n14808), .ZN(n14809) );
  INV_X1 U9468 ( .A(n15043), .ZN(n6851) );
  NAND2_X1 U9469 ( .A1(n6851), .A2(n6765), .ZN(n6852) );
  NAND2_X1 U9470 ( .A1(n8873), .A2(n8872), .ZN(n8822) );
  NAND2_X1 U9471 ( .A1(n8869), .A2(n8868), .ZN(n6853) );
  NAND2_X1 U9472 ( .A1(n6855), .A2(n12447), .ZN(n11500) );
  NAND2_X1 U9473 ( .A1(n15551), .A2(n12472), .ZN(n6855) );
  NAND2_X1 U9474 ( .A1(n7636), .A2(n8013), .ZN(n8081) );
  NAND3_X1 U9475 ( .A1(n6861), .A2(n6988), .A3(n6987), .ZN(n7966) );
  AND2_X1 U9476 ( .A1(n7872), .A2(n7757), .ZN(n7749) );
  NAND2_X1 U9477 ( .A1(n6865), .A2(n9308), .ZN(n11066) );
  OAI21_X2 U9478 ( .B1(n7366), .B2(n6868), .A(n6866), .ZN(n13089) );
  NAND2_X1 U9479 ( .A1(n15580), .A2(n12457), .ZN(n11300) );
  NAND2_X1 U9480 ( .A1(n10413), .A2(n12450), .ZN(n8724) );
  XNOR2_X1 U9481 ( .A(n7907), .B(n7906), .ZN(n10594) );
  XNOR2_X1 U9482 ( .A(n7774), .B(n10117), .ZN(n7907) );
  NAND2_X2 U9483 ( .A1(n7347), .A2(n7346), .ZN(n7774) );
  NAND2_X1 U9484 ( .A1(n11517), .A2(n7258), .ZN(n6870) );
  NAND2_X1 U9485 ( .A1(n11428), .A2(n11429), .ZN(n6871) );
  NAND2_X1 U9486 ( .A1(n14844), .A2(n14845), .ZN(n6878) );
  AND3_X2 U9487 ( .A1(n6798), .A2(n7218), .A3(n7217), .ZN(n8476) );
  XNOR2_X2 U9488 ( .A(n11094), .B(n13674), .ZN(n11092) );
  NAND2_X2 U9489 ( .A1(n6884), .A2(n6883), .ZN(n13674) );
  XNOR2_X2 U9490 ( .A(n13673), .B(n6881), .ZN(n10419) );
  AND2_X1 U9491 ( .A1(n9277), .A2(n9275), .ZN(n6883) );
  AND2_X1 U9492 ( .A1(n9274), .A2(n9276), .ZN(n6884) );
  OAI21_X2 U9493 ( .B1(n8317), .B2(n6889), .A(n6886), .ZN(n8346) );
  NAND2_X1 U9494 ( .A1(n8346), .A2(n8345), .ZN(n8348) );
  OAI21_X1 U9495 ( .B1(n8523), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n6894), .ZN(
        n8532) );
  AOI21_X1 U9496 ( .B1(n6894), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8531), .ZN(
        n6891) );
  OR2_X1 U9497 ( .A1(n8173), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U9498 ( .A1(n6895), .A2(n12607), .ZN(P3_U3296) );
  NAND2_X1 U9499 ( .A1(n6896), .A2(n10677), .ZN(n6895) );
  NAND2_X1 U9500 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  NAND2_X1 U9501 ( .A1(n12602), .A2(n12601), .ZN(n6898) );
  NAND2_X1 U9502 ( .A1(n8586), .A2(n8181), .ZN(n6900) );
  NAND2_X1 U9503 ( .A1(n8505), .A2(n8504), .ZN(n8507) );
  NAND2_X1 U9504 ( .A1(n8492), .A2(n8169), .ZN(n6901) );
  NAND2_X1 U9505 ( .A1(n8129), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U9506 ( .A1(n8406), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U9507 ( .A1(n8397), .A2(n8155), .ZN(n6902) );
  NAND2_X1 U9508 ( .A1(n6903), .A2(n7402), .ZN(n7401) );
  NAND2_X1 U9509 ( .A1(n6903), .A2(n8288), .ZN(n7406) );
  XNOR2_X1 U9510 ( .A(n6903), .B(n8288), .ZN(n10078) );
  NAND2_X1 U9511 ( .A1(n8139), .A2(n8138), .ZN(n6903) );
  NAND4_X1 U9512 ( .A1(n12440), .A2(n13076), .A3(n13102), .A4(n13088), .ZN(
        n7409) );
  NAND2_X1 U9513 ( .A1(n10716), .A2(n10720), .ZN(n6906) );
  XNOR2_X2 U9514 ( .A(n11057), .B(n6907), .ZN(n10720) );
  NAND2_X1 U9515 ( .A1(n6908), .A2(n9292), .ZN(n10716) );
  NAND2_X1 U9516 ( .A1(n10733), .A2(n9994), .ZN(n6908) );
  MUX2_X1 U9517 ( .A(n13975), .B(n6909), .S(n15431), .Z(n13976) );
  MUX2_X1 U9518 ( .A(n14051), .B(n6909), .S(n15420), .Z(n14052) );
  NAND3_X1 U9519 ( .A1(n8083), .A2(P2_IR_REG_29__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n6917) );
  NAND3_X1 U9520 ( .A1(n7636), .A2(n7042), .A3(n7041), .ZN(n8083) );
  INV_X1 U9521 ( .A(n8781), .ZN(n7710) );
  XNOR2_X1 U9522 ( .A(n8748), .B(n8747), .ZN(n11803) );
  OAI21_X2 U9523 ( .B1(n14220), .B2(n6933), .A(n6931), .ZN(n14174) );
  NAND2_X2 U9524 ( .A1(n14249), .A2(n14248), .ZN(n14247) );
  XNOR2_X2 U9525 ( .A(n12679), .B(n12680), .ZN(n14249) );
  INV_X1 U9526 ( .A(n6935), .ZN(n10825) );
  OR2_X2 U9527 ( .A1(n10816), .A2(n10815), .ZN(n6935) );
  XNOR2_X1 U9528 ( .A(n11489), .B(n6936), .ZN(n11028) );
  AND2_X1 U9529 ( .A1(n10576), .A2(n12189), .ZN(n10894) );
  NAND2_X2 U9530 ( .A1(n11546), .A2(n11216), .ZN(n10817) );
  NAND2_X1 U9531 ( .A1(n13133), .A2(n13132), .ZN(n13131) );
  INV_X1 U9532 ( .A(n13173), .ZN(n8542) );
  NAND2_X1 U9533 ( .A1(n6938), .A2(n15591), .ZN(n15613) );
  NAND2_X1 U9534 ( .A1(n6937), .A2(n15611), .ZN(n15591) );
  NAND2_X1 U9535 ( .A1(n14847), .A2(n8404), .ZN(n14848) );
  NAND2_X1 U9536 ( .A1(n6950), .A2(n6951), .ZN(n13233) );
  NAND2_X1 U9537 ( .A1(n13257), .A2(n6953), .ZN(n6950) );
  NAND3_X1 U9538 ( .A1(n6811), .A2(n6961), .A3(n6960), .ZN(n7388) );
  NAND2_X1 U9539 ( .A1(n11504), .A2(n12429), .ZN(n11503) );
  INV_X1 U9540 ( .A(n6979), .ZN(n11249) );
  NAND2_X1 U9541 ( .A1(n6980), .A2(n7490), .ZN(n15067) );
  NAND4_X1 U9542 ( .A1(n6810), .A2(n7309), .A3(n6981), .A4(n7308), .ZN(n14761)
         );
  NAND4_X1 U9543 ( .A1(n7309), .A2(n7308), .A3(n7311), .A4(n7594), .ZN(n10578)
         );
  INV_X1 U9544 ( .A(n6983), .ZN(n11931) );
  INV_X1 U9545 ( .A(n9604), .ZN(n6985) );
  NAND2_X1 U9546 ( .A1(n9593), .A2(n9592), .ZN(n7736) );
  NAND2_X1 U9547 ( .A1(n6721), .A2(n9593), .ZN(n6984) );
  NAND3_X1 U9548 ( .A1(n6991), .A2(n6992), .A3(n7863), .ZN(n6990) );
  NAND3_X1 U9549 ( .A1(n13633), .A2(n13534), .A3(n9666), .ZN(n13533) );
  NAND2_X1 U9550 ( .A1(n8444), .A2(n8163), .ZN(n8458) );
  NAND2_X1 U9551 ( .A1(n7033), .A2(n8661), .ZN(n7032) );
  NAND2_X1 U9552 ( .A1(n8159), .A2(n8158), .ZN(n8426) );
  NAND2_X1 U9553 ( .A1(n14221), .A2(n14222), .ZN(n14220) );
  AOI22_X1 U9554 ( .A1(n14115), .A2(n14116), .B1(n12766), .B2(n12765), .ZN(
        n12775) );
  INV_X1 U9555 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U9556 ( .A1(n10593), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U9557 ( .A1(n14152), .A2(n12725), .ZN(n14221) );
  INV_X1 U9558 ( .A(n7907), .ZN(n7768) );
  NAND2_X1 U9559 ( .A1(n7925), .A2(n7924), .ZN(n7297) );
  NAND2_X1 U9560 ( .A1(n13524), .A2(n13526), .ZN(n13525) );
  AND2_X4 U9561 ( .A1(n6999), .A2(n6998), .ZN(n10593) );
  NAND2_X1 U9562 ( .A1(n7139), .A2(n7766), .ZN(n6998) );
  NAND2_X1 U9563 ( .A1(n7140), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6999) );
  OR2_X1 U9564 ( .A1(n7921), .A2(n10892), .ZN(n7931) );
  AND2_X2 U9565 ( .A1(n11606), .A2(n15410), .ZN(n11794) );
  NAND2_X1 U9566 ( .A1(n10375), .A2(n9591), .ZN(n10408) );
  NAND2_X1 U9567 ( .A1(n11503), .A2(n8304), .ZN(n15541) );
  NAND2_X1 U9568 ( .A1(n13146), .A2(n8571), .ZN(n13133) );
  NAND2_X1 U9569 ( .A1(n8542), .A2(n8541), .ZN(n13171) );
  AOI21_X1 U9570 ( .B1(n13271), .B2(n8440), .A(n6699), .ZN(n13257) );
  NAND2_X1 U9571 ( .A1(n7001), .A2(n15596), .ZN(n11302) );
  NAND2_X1 U9572 ( .A1(n7036), .A2(n8066), .ZN(n9752) );
  INV_X1 U9573 ( .A(n9598), .ZN(n7003) );
  NOR2_X1 U9574 ( .A1(n10707), .A2(n7003), .ZN(n7735) );
  NAND2_X1 U9575 ( .A1(n10864), .A2(n7733), .ZN(n7004) );
  NAND2_X1 U9576 ( .A1(n13755), .A2(n7005), .ZN(n13971) );
  OR2_X1 U9577 ( .A1(n13757), .A2(n13756), .ZN(n7005) );
  NAND2_X1 U9578 ( .A1(n13757), .A2(n13756), .ZN(n13755) );
  NAND2_X1 U9579 ( .A1(n14052), .A2(n6819), .ZN(P2_U3495) );
  INV_X1 U9580 ( .A(n7966), .ZN(n7042) );
  NAND2_X1 U9581 ( .A1(n7150), .A2(n7301), .ZN(n14608) );
  NAND2_X1 U9582 ( .A1(n10979), .A2(n10978), .ZN(n11248) );
  NAND2_X1 U9583 ( .A1(n10922), .A2(n10921), .ZN(n10960) );
  NAND2_X1 U9584 ( .A1(n7142), .A2(n10992), .ZN(n11261) );
  NAND2_X1 U9585 ( .A1(n7141), .A2(n10961), .ZN(n11362) );
  NAND2_X1 U9586 ( .A1(n11618), .A2(n7732), .ZN(n11624) );
  OR2_X1 U9587 ( .A1(n8245), .A2(n8234), .ZN(n8235) );
  NAND2_X1 U9588 ( .A1(n7008), .A2(n12466), .ZN(n15567) );
  NAND2_X1 U9589 ( .A1(n11300), .A2(n12427), .ZN(n7008) );
  NAND2_X1 U9590 ( .A1(n8650), .A2(n12492), .ZN(n11644) );
  NAND2_X1 U9591 ( .A1(n12420), .A2(n12592), .ZN(n7023) );
  INV_X1 U9592 ( .A(n14268), .ZN(n12226) );
  NOR2_X4 U9593 ( .A1(n14497), .A2(n14509), .ZN(n14492) );
  AND2_X1 U9594 ( .A1(n10938), .A2(n12234), .ZN(n11363) );
  NAND2_X1 U9595 ( .A1(n7056), .A2(n7055), .ZN(n7054) );
  AOI21_X1 U9596 ( .B1(n12298), .B2(n12297), .A(n7012), .ZN(n7211) );
  NOR2_X2 U9597 ( .A1(n14192), .A2(n7307), .ZN(n11532) );
  NAND2_X1 U9598 ( .A1(n10240), .A2(n9584), .ZN(n10376) );
  NAND2_X1 U9599 ( .A1(n8252), .A2(n12463), .ZN(n15596) );
  NAND2_X1 U9600 ( .A1(n15541), .A2(n15540), .ZN(n7423) );
  NAND3_X1 U9601 ( .A1(n13071), .A2(n7432), .A3(n15612), .ZN(n7017) );
  NAND2_X1 U9602 ( .A1(n13233), .A2(n13234), .ZN(n7422) );
  NAND2_X1 U9603 ( .A1(n10376), .A2(n10377), .ZN(n10375) );
  NAND2_X1 U9604 ( .A1(n8257), .A2(n8256), .ZN(n7020) );
  NAND2_X1 U9605 ( .A1(n8570), .A2(n8569), .ZN(n13146) );
  OAI21_X1 U9606 ( .B1(n6681), .B2(n12400), .A(n9577), .ZN(n12396) );
  NAND2_X1 U9607 ( .A1(n7053), .A2(n7052), .ZN(n7051) );
  INV_X1 U9608 ( .A(n7351), .ZN(n9571) );
  AOI22_X1 U9609 ( .A1(n12092), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n12091), 
        .B2(n14307), .ZN(n10891) );
  NOR2_X1 U9610 ( .A1(n10646), .A2(n10592), .ZN(n10610) );
  NAND2_X1 U9611 ( .A1(n7378), .A2(n7376), .ZN(P3_U3486) );
  OAI21_X1 U9612 ( .B1(n13094), .B2(n15594), .A(n13093), .ZN(n13303) );
  NAND2_X1 U9613 ( .A1(n14885), .A2(n9384), .ZN(n11990) );
  NAND2_X1 U9614 ( .A1(n7259), .A2(n7349), .ZN(P2_U3496) );
  NAND2_X2 U9615 ( .A1(n14133), .A2(n12648), .ZN(n14977) );
  NOR2_X1 U9616 ( .A1(n10210), .A2(n14781), .ZN(n10064) );
  NAND2_X1 U9617 ( .A1(n10887), .A2(n11545), .ZN(n7053) );
  NAND2_X1 U9618 ( .A1(n7662), .A2(n7661), .ZN(n14115) );
  NAND2_X2 U9619 ( .A1(n13815), .A2(n6737), .ZN(n7554) );
  NAND2_X2 U9620 ( .A1(n7279), .A2(n7276), .ZN(n13815) );
  NAND2_X1 U9621 ( .A1(n9532), .A2(n7747), .ZN(n9535) );
  AND3_X4 U9622 ( .A1(n7931), .A2(n7930), .A3(n7929), .ZN(n15379) );
  NAND2_X1 U9623 ( .A1(n7269), .A2(n7268), .ZN(n13912) );
  NAND2_X1 U9624 ( .A1(n8130), .A2(n8229), .ZN(n7031) );
  XNOR2_X1 U9625 ( .A(n13103), .B(n13102), .ZN(n7035) );
  NAND2_X1 U9626 ( .A1(n14848), .A2(n8405), .ZN(n13284) );
  OAI21_X1 U9627 ( .B1(n9571), .B2(n15429), .A(n7455), .ZN(P2_U3528) );
  NAND2_X1 U9628 ( .A1(n13920), .A2(n9416), .ZN(n13898) );
  OR2_X1 U9629 ( .A1(n10593), .A2(n8131), .ZN(n7347) );
  AND2_X1 U9630 ( .A1(n12257), .A2(n12256), .ZN(n7595) );
  NAND3_X1 U9631 ( .A1(n12294), .A2(n12292), .A3(n12293), .ZN(n7044) );
  NAND3_X1 U9632 ( .A1(n12225), .A2(n12223), .A3(n12224), .ZN(n12232) );
  NAND2_X1 U9633 ( .A1(n7209), .A2(n7562), .ZN(n12311) );
  NAND2_X1 U9634 ( .A1(n7179), .A2(n7178), .ZN(n12344) );
  NAND2_X1 U9635 ( .A1(n7185), .A2(n7184), .ZN(n12258) );
  NAND2_X1 U9636 ( .A1(n7054), .A2(n12373), .ZN(P1_U3242) );
  NAND2_X1 U9637 ( .A1(n7587), .A2(n7586), .ZN(n7585) );
  NAND4_X1 U9638 ( .A1(n7230), .A2(n8743), .A3(n7229), .A4(n7232), .ZN(n7234)
         );
  XNOR2_X2 U9639 ( .A(n11541), .B(n7050), .ZN(n11544) );
  XNOR2_X2 U9640 ( .A(n8204), .B(n13429), .ZN(n12623) );
  NAND2_X1 U9641 ( .A1(n11302), .A2(n8266), .ZN(n15569) );
  NAND4_X1 U9642 ( .A1(n12368), .A2(n12210), .A3(n7057), .A4(n12369), .ZN(
        n7056) );
  NAND2_X1 U9643 ( .A1(n7977), .A2(n7061), .ZN(n7060) );
  OAI21_X1 U9644 ( .B1(n8034), .B2(n7070), .A(n7068), .ZN(n7828) );
  OAI21_X1 U9645 ( .B1(n8034), .B2(n8033), .A(n7824), .ZN(n7076) );
  MUX2_X1 U9646 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n10593), .Z(n7780) );
  NAND2_X1 U9647 ( .A1(n7079), .A2(n7077), .ZN(n12206) );
  OAI21_X1 U9648 ( .B1(n14407), .B2(n12176), .A(n6682), .ZN(n7079) );
  NAND2_X1 U9649 ( .A1(n14083), .A2(n12161), .ZN(n7080) );
  NAND3_X1 U9650 ( .A1(n7519), .A2(n7518), .A3(n15031), .ZN(n15030) );
  NAND3_X1 U9651 ( .A1(n7519), .A2(n7518), .A3(n7090), .ZN(n7089) );
  NAND3_X1 U9652 ( .A1(n7107), .A2(n10691), .A3(P3_IR_REG_2__SCAN_IN), .ZN(
        n7103) );
  AOI21_X1 U9653 ( .B1(n12953), .B2(n12968), .A(n7109), .ZN(n7108) );
  NAND3_X1 U9654 ( .A1(n7125), .A2(n7467), .A3(n7122), .ZN(P3_U3201) );
  NAND3_X1 U9655 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U9656 ( .A1(n7129), .A2(n7925), .ZN(n7130) );
  INV_X1 U9657 ( .A(n7235), .ZN(n7132) );
  NAND3_X1 U9658 ( .A1(n7131), .A2(n7130), .A3(n7784), .ZN(n7948) );
  NAND2_X1 U9659 ( .A1(n7133), .A2(n7235), .ZN(n7944) );
  NAND2_X1 U9660 ( .A1(n7925), .A2(n7294), .ZN(n7133) );
  NAND3_X1 U9661 ( .A1(n13731), .A2(n7280), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7139) );
  NAND3_X1 U9662 ( .A1(n8910), .A2(n7281), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7140) );
  NAND2_X1 U9663 ( .A1(n11362), .A2(n12101), .ZN(n10967) );
  NAND2_X1 U9664 ( .A1(n10960), .A2(n10959), .ZN(n7141) );
  NAND2_X1 U9665 ( .A1(n11261), .A2(n11260), .ZN(n11263) );
  NAND2_X1 U9666 ( .A1(n11248), .A2(n10991), .ZN(n7142) );
  NAND3_X1 U9667 ( .A1(n7146), .A2(n7145), .A3(n6692), .ZN(n7150) );
  OAI21_X1 U9668 ( .B1(n14669), .B2(n7157), .A(n7151), .ZN(P1_U3557) );
  AOI21_X1 U9669 ( .B1(n7152), .B2(n15225), .A(n7155), .ZN(n7151) );
  AOI21_X1 U9670 ( .B1(n7152), .B2(n15212), .A(n7154), .ZN(n7153) );
  OAI21_X1 U9671 ( .B1(n14669), .B2(n7159), .A(n7153), .ZN(P1_U3525) );
  OAI211_X1 U9672 ( .C1(n14593), .C2(n7166), .A(n14569), .B(n7165), .ZN(n14568) );
  INV_X1 U9673 ( .A(n14569), .ZN(n7161) );
  NAND2_X1 U9674 ( .A1(n14426), .A2(n7169), .ZN(n7162) );
  INV_X1 U9675 ( .A(n14426), .ZN(n7163) );
  NAND2_X1 U9676 ( .A1(n14487), .A2(n14486), .ZN(n14485) );
  NAND2_X1 U9677 ( .A1(n14487), .A2(n6787), .ZN(n7171) );
  INV_X2 U9678 ( .A(n10603), .ZN(n15107) );
  NAND2_X2 U9680 ( .A1(n10818), .A2(n10593), .ZN(n11914) );
  NAND2_X1 U9681 ( .A1(n12337), .A2(n6726), .ZN(n7179) );
  OAI211_X1 U9682 ( .C1(n12249), .C2(n12250), .A(n7186), .B(n7583), .ZN(n7185)
         );
  NAND2_X1 U9683 ( .A1(n7187), .A2(n12248), .ZN(n7186) );
  NAND2_X1 U9684 ( .A1(n12249), .A2(n12250), .ZN(n7187) );
  INV_X1 U9685 ( .A(n12270), .ZN(n12273) );
  NAND2_X1 U9686 ( .A1(n7190), .A2(n7191), .ZN(n12270) );
  NAND3_X1 U9687 ( .A1(n12358), .A2(n7570), .A3(n12357), .ZN(n7202) );
  OAI21_X1 U9688 ( .B1(n7211), .B2(n7210), .A(n7564), .ZN(n7209) );
  NOR2_X1 U9689 ( .A1(n12298), .A2(n12297), .ZN(n7210) );
  NAND3_X1 U9690 ( .A1(n6798), .A2(n7216), .A3(n7217), .ZN(n8479) );
  NAND2_X1 U9691 ( .A1(n12845), .A2(n12846), .ZN(n7227) );
  NAND2_X1 U9692 ( .A1(n8743), .A2(n7232), .ZN(n7231) );
  INV_X1 U9693 ( .A(n7234), .ZN(n11323) );
  NAND2_X1 U9694 ( .A1(n14484), .A2(n7238), .ZN(n7236) );
  NAND2_X1 U9695 ( .A1(n7236), .A2(n7237), .ZN(n7241) );
  NAND2_X1 U9696 ( .A1(n7282), .A2(n7246), .ZN(n7244) );
  NAND2_X1 U9697 ( .A1(n7244), .A2(n7245), .ZN(n7792) );
  NAND2_X1 U9698 ( .A1(n7249), .A2(n6801), .ZN(n8020) );
  MUX2_X1 U9699 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n10593), .Z(n7778) );
  NAND2_X1 U9700 ( .A1(n11599), .A2(n11603), .ZN(n9528) );
  NAND2_X1 U9701 ( .A1(n11288), .A2(n9522), .ZN(n11430) );
  NAND2_X1 U9702 ( .A1(n13763), .A2(n6804), .ZN(n7266) );
  NAND3_X1 U9703 ( .A1(n7267), .A2(n7266), .A3(n7264), .ZN(n7536) );
  NAND2_X1 U9704 ( .A1(n13948), .A2(n7270), .ZN(n7269) );
  INV_X1 U9705 ( .A(n13661), .ZN(n7274) );
  NAND2_X1 U9706 ( .A1(n9549), .A2(n7277), .ZN(n7279) );
  CLKBUF_X1 U9707 ( .A(n7279), .Z(n7275) );
  NAND2_X1 U9708 ( .A1(n7948), .A2(n7785), .ZN(n7282) );
  NAND2_X1 U9709 ( .A1(n7283), .A2(n11469), .ZN(n11527) );
  NAND2_X1 U9710 ( .A1(n11468), .A2(n7286), .ZN(n7283) );
  NAND2_X1 U9711 ( .A1(n12106), .A2(n11469), .ZN(n7284) );
  INV_X1 U9712 ( .A(n11469), .ZN(n7285) );
  NAND2_X1 U9713 ( .A1(n11263), .A2(n11262), .ZN(n11468) );
  INV_X1 U9714 ( .A(n7298), .ZN(n7294) );
  INV_X1 U9715 ( .A(n7924), .ZN(n7295) );
  INV_X1 U9716 ( .A(n7933), .ZN(n7296) );
  NAND2_X1 U9717 ( .A1(n12052), .A2(n6769), .ZN(n7915) );
  NAND2_X1 U9718 ( .A1(n7915), .A2(n10574), .ZN(n7906) );
  NAND3_X1 U9719 ( .A1(n15078), .A2(n15180), .A3(n11782), .ZN(n11255) );
  INV_X1 U9720 ( .A(n7307), .ZN(n11278) );
  AND3_X1 U9721 ( .A1(n7593), .A2(n10062), .A3(n7670), .ZN(n7310) );
  NAND3_X1 U9722 ( .A1(n7310), .A2(n7487), .A3(n7311), .ZN(n10195) );
  AND2_X1 U9723 ( .A1(n14492), .A2(n7318), .ZN(n14450) );
  NAND2_X1 U9724 ( .A1(n14492), .A2(n14673), .ZN(n14472) );
  NAND2_X1 U9725 ( .A1(n7316), .A2(n14492), .ZN(n14410) );
  OAI211_X1 U9726 ( .C1(n7316), .C2(n14407), .A(n7315), .B(n7314), .ZN(n14404)
         );
  NAND3_X1 U9727 ( .A1(n7316), .A2(n14492), .A3(n14407), .ZN(n7315) );
  NAND3_X1 U9728 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9729 ( .A1(n11794), .A2(n7348), .ZN(n11821) );
  NAND2_X1 U9730 ( .A1(n12469), .A2(n12470), .ZN(n15568) );
  NAND2_X1 U9731 ( .A1(n15556), .A2(n8734), .ZN(n12470) );
  NAND3_X1 U9732 ( .A1(n8269), .A2(n8270), .A3(n7362), .ZN(n11301) );
  NAND2_X1 U9733 ( .A1(n13237), .A2(n7364), .ZN(n13216) );
  NAND2_X1 U9734 ( .A1(n13126), .A2(n7369), .ZN(n7366) );
  NAND2_X1 U9735 ( .A1(n7372), .A2(n6799), .ZN(n8655) );
  OAI21_X1 U9736 ( .B1(n15533), .B2(n8652), .A(n12502), .ZN(n14858) );
  NAND2_X1 U9737 ( .A1(n8458), .A2(n7393), .ZN(n7392) );
  NAND3_X1 U9738 ( .A1(n8249), .A2(n8248), .A3(n8259), .ZN(n7398) );
  NAND2_X1 U9739 ( .A1(n7398), .A2(n7396), .ZN(n8274) );
  INV_X1 U9740 ( .A(n8134), .ZN(n7397) );
  NAND2_X1 U9741 ( .A1(n7401), .A2(n7403), .ZN(n8315) );
  NAND4_X1 U9742 ( .A1(n7410), .A2(n12591), .A3(n12596), .A4(n7408), .ZN(n7407) );
  NAND2_X1 U9743 ( .A1(n8187), .A2(n7412), .ZN(n7411) );
  NAND2_X1 U9744 ( .A1(n7411), .A2(n6706), .ZN(n12402) );
  NAND2_X1 U9745 ( .A1(n8187), .A2(n8186), .ZN(n8214) );
  NAND2_X1 U9746 ( .A1(n8367), .A2(n8151), .ZN(n8383) );
  NAND2_X1 U9747 ( .A1(n8507), .A2(n8172), .ZN(n8173) );
  NAND2_X1 U9748 ( .A1(n8154), .A2(n8153), .ZN(n8397) );
  OR2_X1 U9749 ( .A1(n8261), .A2(n10081), .ZN(n8251) );
  OAI21_X1 U9750 ( .B1(n13086), .B2(n7431), .A(n7429), .ZN(n8626) );
  NAND2_X1 U9751 ( .A1(n13084), .A2(n7433), .ZN(n7432) );
  NAND2_X1 U9752 ( .A1(n13835), .A2(n9449), .ZN(n7437) );
  NAND2_X1 U9753 ( .A1(n7437), .A2(n6723), .ZN(n7441) );
  NOR2_X1 U9754 ( .A1(n7439), .A2(n7438), .ZN(n7436) );
  NOR2_X1 U9755 ( .A1(n14916), .A2(n9989), .ZN(n7451) );
  NAND2_X1 U9756 ( .A1(n13930), .A2(n7452), .ZN(n13920) );
  INV_X1 U9757 ( .A(n7460), .ZN(n13806) );
  NAND2_X1 U9758 ( .A1(n14059), .A2(n9932), .ZN(n7459) );
  OAI21_X2 U9759 ( .B1(n10109), .B2(n7921), .A(n7461), .ZN(n11057) );
  NAND3_X1 U9760 ( .A1(n7776), .A2(n7463), .A3(n7775), .ZN(n7919) );
  NAND3_X1 U9761 ( .A1(n7770), .A2(SI_2_), .A3(n7771), .ZN(n7463) );
  NOR2_X1 U9762 ( .A1(n15504), .A2(n11165), .ZN(n15503) );
  INV_X1 U9763 ( .A(n11127), .ZN(n7466) );
  XNOR2_X1 U9764 ( .A(n11125), .B(n11166), .ZN(n15504) );
  NAND2_X1 U9765 ( .A1(n14839), .A2(n7468), .ZN(n7467) );
  OAI21_X1 U9766 ( .B1(n12982), .B2(n7483), .A(n7482), .ZN(n13030) );
  OAI211_X2 U9767 ( .C1(n7505), .C2(n12109), .A(n7503), .B(n7508), .ZN(n11657)
         );
  INV_X1 U9768 ( .A(n7506), .ZN(n7504) );
  NAND2_X1 U9769 ( .A1(n11530), .A2(n11529), .ZN(n11528) );
  NAND2_X1 U9770 ( .A1(n7505), .A2(n7506), .ZN(n11530) );
  NAND2_X2 U9771 ( .A1(n7535), .A2(n7777), .ZN(n7925) );
  NAND2_X1 U9772 ( .A1(n7919), .A2(n7920), .ZN(n7535) );
  INV_X1 U9773 ( .A(n7906), .ZN(n7770) );
  NAND2_X1 U9774 ( .A1(n7536), .A2(n9567), .ZN(n13751) );
  NAND2_X1 U9775 ( .A1(n7965), .A2(n7541), .ZN(n7539) );
  INV_X1 U9776 ( .A(n13799), .ZN(n7556) );
  OAI211_X2 U9777 ( .C1(n7554), .C2(n9554), .A(n10006), .B(n7552), .ZN(n13771)
         );
  OR2_X1 U9778 ( .A1(n6703), .A2(n14760), .ZN(n7557) );
  XNOR2_X2 U9779 ( .A(n7558), .B(n10580), .ZN(n12378) );
  NAND2_X1 U9780 ( .A1(n7561), .A2(n12312), .ZN(n12315) );
  INV_X1 U9781 ( .A(n12301), .ZN(n7569) );
  NAND2_X1 U9782 ( .A1(n7574), .A2(n7577), .ZN(n12286) );
  NAND3_X1 U9783 ( .A1(n12275), .A2(n7575), .A3(n12274), .ZN(n7574) );
  INV_X1 U9784 ( .A(n12339), .ZN(n7579) );
  OR2_X2 U9785 ( .A1(n11950), .A2(n12290), .ZN(n11948) );
  INV_X1 U9786 ( .A(n14415), .ZN(n7582) );
  INV_X1 U9787 ( .A(n12252), .ZN(n7584) );
  OAI211_X1 U9788 ( .C1(n6682), .C2(n12219), .A(n7585), .B(n12220), .ZN(n12225) );
  INV_X1 U9789 ( .A(n12326), .ZN(n7588) );
  NAND2_X1 U9790 ( .A1(n14485), .A2(n7591), .ZN(n14676) );
  OR2_X1 U9791 ( .A1(n14487), .A2(n14486), .ZN(n7591) );
  NAND2_X1 U9792 ( .A1(n12262), .A2(n7597), .ZN(n7596) );
  INV_X1 U9793 ( .A(n12263), .ZN(n7598) );
  OAI21_X1 U9794 ( .B1(n9925), .B2(n7607), .A(n7605), .ZN(n9936) );
  OAI21_X1 U9795 ( .B1(n9925), .B2(n7612), .A(n7604), .ZN(n9935) );
  NAND2_X1 U9796 ( .A1(n9925), .A2(n7602), .ZN(n7601) );
  INV_X1 U9797 ( .A(n7612), .ZN(n7608) );
  INV_X1 U9798 ( .A(n9933), .ZN(n7613) );
  NAND2_X1 U9799 ( .A1(n7617), .A2(n7756), .ZN(n10030) );
  NAND2_X1 U9800 ( .A1(n10025), .A2(n9985), .ZN(n7617) );
  INV_X1 U9801 ( .A(n9957), .ZN(n7619) );
  OAI22_X1 U9802 ( .A1(n9889), .A2(n7621), .B1(n7620), .B2(n9890), .ZN(n9896)
         );
  NOR2_X1 U9803 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  NAND3_X1 U9804 ( .A1(n7764), .A2(n9808), .A3(n6791), .ZN(n7622) );
  OAI21_X1 U9805 ( .B1(n7625), .B2(n9822), .A(n7624), .ZN(n9833) );
  OR2_X1 U9806 ( .A1(n9821), .A2(n7626), .ZN(n7625) );
  NAND2_X1 U9807 ( .A1(n7627), .A2(n6807), .ZN(n9807) );
  NAND3_X1 U9808 ( .A1(n7628), .A2(n6691), .A3(n6790), .ZN(n7627) );
  INV_X1 U9809 ( .A(n9795), .ZN(n7628) );
  NAND3_X1 U9810 ( .A1(n9907), .A2(n9906), .A3(n6803), .ZN(n7630) );
  NAND2_X1 U9811 ( .A1(n7630), .A2(n6806), .ZN(n9918) );
  INV_X1 U9812 ( .A(n9913), .ZN(n7632) );
  NAND2_X1 U9813 ( .A1(n7633), .A2(n7635), .ZN(n9843) );
  NAND3_X1 U9814 ( .A1(n7634), .A2(n6690), .A3(n6793), .ZN(n7633) );
  INV_X1 U9815 ( .A(n9834), .ZN(n7634) );
  NAND2_X1 U9816 ( .A1(n7641), .A2(n6789), .ZN(n9787) );
  NAND3_X1 U9817 ( .A1(n7643), .A2(n6774), .A3(n7642), .ZN(n7641) );
  INV_X1 U9818 ( .A(n9774), .ZN(n7643) );
  NAND2_X1 U9819 ( .A1(n11544), .A2(n7645), .ZN(n7644) );
  NOR2_X1 U9820 ( .A1(n7654), .A2(n7646), .ZN(n7645) );
  NAND3_X1 U9821 ( .A1(n7648), .A2(n7647), .A3(n11636), .ZN(n11776) );
  INV_X1 U9822 ( .A(n11544), .ZN(n7649) );
  NAND2_X1 U9823 ( .A1(n7650), .A2(n7024), .ZN(n11637) );
  NAND2_X1 U9824 ( .A1(n11544), .A2(n7653), .ZN(n7650) );
  NAND3_X1 U9825 ( .A1(n10047), .A2(n10141), .A3(n10177), .ZN(n7671) );
  INV_X1 U9826 ( .A(n11024), .ZN(n7674) );
  NOR2_X1 U9827 ( .A1(n11025), .A2(n11024), .ZN(n11029) );
  OAI21_X1 U9828 ( .B1(n10187), .B2(n7676), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7677) );
  NAND2_X1 U9829 ( .A1(n14977), .A2(n7678), .ZN(n14166) );
  NAND2_X1 U9830 ( .A1(n12846), .A2(n7694), .ZN(n7692) );
  NAND2_X1 U9831 ( .A1(n12846), .A2(n7701), .ZN(n7693) );
  OAI211_X1 U9832 ( .C1(n12846), .C2(n7698), .A(n7695), .B(n7692), .ZN(n8796)
         );
  NAND2_X1 U9833 ( .A1(n7710), .A2(n8782), .ZN(n7712) );
  NAND3_X1 U9834 ( .A1(n8781), .A2(n13176), .A3(n8782), .ZN(n12901) );
  NAND3_X1 U9835 ( .A1(n8190), .A2(n8230), .A3(n8189), .ZN(n8361) );
  NAND3_X1 U9836 ( .A1(n10669), .A2(n6724), .A3(n8731), .ZN(n7717) );
  NAND3_X1 U9837 ( .A1(n8195), .A2(n7724), .A3(n7723), .ZN(n7722) );
  XNOR2_X1 U9838 ( .A(n15379), .B(n6684), .ZN(n9594) );
  XNOR2_X1 U9839 ( .A(n6684), .B(n10422), .ZN(n9589) );
  XNOR2_X1 U9840 ( .A(n15386), .B(n6683), .ZN(n9605) );
  XNOR2_X1 U9841 ( .A(n11418), .B(n6684), .ZN(n9618) );
  XNOR2_X1 U9842 ( .A(n11076), .B(n7731), .ZN(n9611) );
  XNOR2_X1 U9843 ( .A(n13498), .B(n6683), .ZN(n9621) );
  XNOR2_X1 U9844 ( .A(n11737), .B(n7731), .ZN(n9626) );
  XNOR2_X1 U9845 ( .A(n11607), .B(n7731), .ZN(n9633) );
  XNOR2_X1 U9846 ( .A(n11795), .B(n7731), .ZN(n9639) );
  XNOR2_X1 U9847 ( .A(n11823), .B(n7731), .ZN(n9643) );
  XNOR2_X1 U9848 ( .A(n13959), .B(n7731), .ZN(n9667) );
  XNOR2_X1 U9849 ( .A(n14889), .B(n7731), .ZN(n9650) );
  XNOR2_X1 U9850 ( .A(n13936), .B(n7731), .ZN(n9671) );
  XNOR2_X1 U9851 ( .A(n11993), .B(n7731), .ZN(n9656) );
  XNOR2_X1 U9852 ( .A(n14031), .B(n7731), .ZN(n9675) );
  XNOR2_X1 U9853 ( .A(n13907), .B(n7731), .ZN(n9682) );
  XNOR2_X1 U9854 ( .A(n14022), .B(n7731), .ZN(n9686) );
  XNOR2_X1 U9855 ( .A(n13811), .B(n7731), .ZN(n9712) );
  XNOR2_X1 U9856 ( .A(n13980), .B(n7731), .ZN(n9722) );
  AOI21_X1 U9857 ( .B1(n11005), .B2(n11004), .A(n11003), .ZN(n11367) );
  NAND2_X2 U9858 ( .A1(n10681), .A2(n10593), .ZN(n8261) );
  INV_X1 U9859 ( .A(n12612), .ZN(n12614) );
  NAND2_X2 U9860 ( .A1(n12623), .A2(n13437), .ZN(n8245) );
  INV_X1 U9861 ( .A(n8207), .ZN(n13437) );
  NAND4_X2 U9862 ( .A1(n8235), .A2(n8237), .A3(n8236), .A4(n8238), .ZN(n15609)
         );
  NAND2_X1 U9863 ( .A1(n6686), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7912) );
  OAI211_X2 U9864 ( .C1(n11914), .C2(n10822), .A(n10821), .B(n10820), .ZN(
        n11397) );
  OR2_X1 U9865 ( .A1(n9920), .A2(n9919), .ZN(n9925) );
  NAND4_X2 U9866 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n15091) );
  AND2_X2 U9867 ( .A1(n12623), .A2(n8207), .ZN(n8224) );
  OAI21_X2 U9868 ( .B1(n10892), .B2(n11914), .A(n10891), .ZN(n12227) );
  INV_X1 U9869 ( .A(n11022), .ZN(n11023) );
  NAND2_X1 U9870 ( .A1(n10607), .A2(n10606), .ZN(n10814) );
  CLKBUF_X1 U9871 ( .A(n9580), .Z(n15412) );
  NAND2_X1 U9872 ( .A1(n8122), .A2(n10739), .ZN(n9751) );
  AND2_X1 U9873 ( .A1(n14053), .A2(n13632), .ZN(n7744) );
  OR2_X1 U9874 ( .A1(n9973), .A2(n9972), .ZN(n7745) );
  OR2_X1 U9875 ( .A1(n15672), .A2(n15605), .ZN(n13423) );
  INV_X1 U9876 ( .A(n13423), .ZN(n8719) );
  AND2_X1 U9877 ( .A1(n8716), .A2(n8715), .ZN(n15672) );
  AND2_X2 U9878 ( .A1(n10658), .A2(n8699), .ZN(n15685) );
  INV_X1 U9879 ( .A(n15685), .ZN(n8704) );
  AND2_X1 U9880 ( .A1(n9649), .A2(n9656), .ZN(n7746) );
  OR2_X1 U9881 ( .A1(n11993), .A2(n9533), .ZN(n7747) );
  AND2_X1 U9882 ( .A1(n14733), .A2(n14734), .ZN(n7748) );
  INV_X1 U9883 ( .A(n12488), .ZN(n8334) );
  OR2_X1 U9884 ( .A1(n11775), .A2(n11774), .ZN(n7750) );
  OR2_X1 U9885 ( .A1(n11961), .A2(n11960), .ZN(n7754) );
  AND2_X1 U9886 ( .A1(n10020), .A2(n10019), .ZN(n7756) );
  AND4_X1 U9887 ( .A1(n7868), .A2(n7867), .A3(n7990), .A4(n7866), .ZN(n7757)
         );
  AND4_X1 U9888 ( .A1(n8471), .A2(n8470), .A3(n8469), .A4(n8468), .ZN(n13260)
         );
  INV_X1 U9889 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12861) );
  AOI21_X1 U9890 ( .B1(n13760), .B2(n9496), .A(n9492), .ZN(n13450) );
  AND2_X1 U9891 ( .A1(n6673), .A2(P2_U3088), .ZN(n14098) );
  INV_X1 U9892 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12834) );
  INV_X1 U9893 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n8878) );
  OR2_X1 U9894 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10684), .ZN(n7758) );
  INV_X1 U9895 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9361) );
  INV_X1 U9896 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8417) );
  INV_X1 U9897 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U9898 ( .A1(n10945), .A2(n10944), .ZN(n15223) );
  INV_X2 U9899 ( .A(n15223), .ZN(n15225) );
  INV_X2 U9900 ( .A(n15210), .ZN(n15212) );
  OR2_X1 U9901 ( .A1(n10032), .A2(n15231), .ZN(n13449) );
  AND2_X1 U9902 ( .A1(n8740), .A2(n12491), .ZN(n7759) );
  INV_X1 U9903 ( .A(n14046), .ZN(n9569) );
  INV_X1 U9904 ( .A(n13630), .ZN(n13632) );
  AND3_X1 U9905 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n7760) );
  AND2_X1 U9906 ( .A1(n7805), .A2(n7804), .ZN(n7761) );
  OR2_X1 U9907 ( .A1(n9963), .A2(n15366), .ZN(n7762) );
  OR2_X1 U9908 ( .A1(n15013), .A2(n14260), .ZN(n7763) );
  INV_X1 U9909 ( .A(n13039), .ZN(n13054) );
  OR2_X1 U9910 ( .A1(n9807), .A2(n9806), .ZN(n7764) );
  OR2_X1 U9911 ( .A1(n11490), .A2(n11489), .ZN(n7765) );
  OAI21_X1 U9912 ( .B1(n12245), .B2(n12244), .A(n12243), .ZN(n12247) );
  MUX2_X1 U9913 ( .A(n14265), .B(n15075), .S(n6682), .Z(n12248) );
  MUX2_X1 U9914 ( .A(n14263), .B(n12255), .S(n6682), .Z(n12256) );
  INV_X1 U9915 ( .A(n9800), .ZN(n9801) );
  MUX2_X1 U9916 ( .A(n14259), .B(n14172), .S(n6682), .Z(n12276) );
  INV_X1 U9917 ( .A(n9862), .ZN(n9855) );
  NAND2_X1 U9918 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  AND2_X1 U9919 ( .A1(n9881), .A2(n9857), .ZN(n9858) );
  MUX2_X1 U9920 ( .A(n14585), .B(n14574), .S(n6682), .Z(n12322) );
  MUX2_X1 U9921 ( .A(n14505), .B(n14497), .S(n6682), .Z(n12342) );
  INV_X1 U9922 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7866) );
  INV_X1 U9923 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7865) );
  INV_X1 U9924 ( .A(n13177), .ZN(n8541) );
  INV_X1 U9925 ( .A(n10017), .ZN(n10018) );
  AND2_X1 U9926 ( .A1(n12441), .A2(n13365), .ZN(n12422) );
  OR2_X1 U9927 ( .A1(n8432), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8450) );
  NOR2_X1 U9928 ( .A1(n8616), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8617) );
  INV_X1 U9929 ( .A(n13149), .ZN(n8569) );
  INV_X1 U9930 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8335) );
  AND2_X1 U9931 ( .A1(n10441), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8160) );
  INV_X1 U9932 ( .A(n13444), .ZN(n9727) );
  INV_X1 U9933 ( .A(n9986), .ZN(n9964) );
  INV_X1 U9934 ( .A(n9441), .ZN(n9260) );
  INV_X1 U9935 ( .A(n13450), .ZN(n9494) );
  INV_X1 U9936 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U9937 ( .A1(n10588), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U9938 ( .A1(n11546), .A2(n12213), .ZN(n10591) );
  INV_X1 U9939 ( .A(n10817), .ZN(n11026) );
  INV_X1 U9940 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11476) );
  OR2_X1 U9941 ( .A1(n14991), .A2(n14942), .ZN(n14434) );
  NAND2_X1 U9942 ( .A1(n7888), .A2(n7831), .ZN(n7836) );
  INV_X1 U9943 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10050) );
  INV_X1 U9944 ( .A(n8758), .ZN(n8759) );
  INV_X1 U9945 ( .A(n8748), .ZN(n8750) );
  INV_X1 U9946 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8277) );
  AND2_X1 U9947 ( .A1(n8617), .A2(n8217), .ZN(n13064) );
  OR2_X1 U9948 ( .A1(n13064), .A2(n8218), .ZN(n13079) );
  NOR2_X1 U9949 ( .A1(n8390), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U9950 ( .A1(n8630), .A2(n8631), .ZN(n8668) );
  AND2_X1 U9951 ( .A1(n8399), .A2(n8398), .ZN(n8408) );
  INV_X1 U9952 ( .A(n13621), .ZN(n9718) );
  INV_X1 U9953 ( .A(n9752), .ZN(n10014) );
  OR2_X1 U9954 ( .A1(n9450), .A2(n13477), .ZN(n9459) );
  NAND2_X1 U9955 ( .A1(n9393), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9418) );
  OR2_X1 U9956 ( .A1(n9470), .A2(n13625), .ZN(n9480) );
  INV_X1 U9957 ( .A(n13447), .ZN(n13622) );
  INV_X1 U9958 ( .A(n10031), .ZN(n8037) );
  AND2_X1 U9959 ( .A1(n14109), .A2(n8106), .ZN(n8108) );
  INV_X1 U9960 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11663) );
  INV_X1 U9961 ( .A(n12633), .ZN(n12634) );
  INV_X1 U9962 ( .A(n14155), .ZN(n12722) );
  INV_X1 U9963 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10929) );
  INV_X1 U9964 ( .A(n11966), .ZN(n11963) );
  AND2_X1 U9965 ( .A1(n14973), .A2(n14974), .ZN(n12648) );
  OR2_X1 U9966 ( .A1(n12123), .A2(n12078), .ZN(n12080) );
  OR2_X1 U9967 ( .A1(n11477), .A2(n11476), .ZN(n11664) );
  INV_X1 U9968 ( .A(n12100), .ZN(n15092) );
  NAND2_X1 U9969 ( .A1(n8058), .A2(n8057), .ZN(n7856) );
  NAND2_X1 U9970 ( .A1(n7821), .A2(n10308), .ZN(n7824) );
  INV_X1 U9971 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8829) );
  NOR2_X1 U9972 ( .A1(n8899), .A2(n8898), .ZN(n8840) );
  OR2_X1 U9973 ( .A1(n12415), .A2(n11054), .ZN(n8560) );
  AND2_X1 U9974 ( .A1(n10671), .A2(n10668), .ZN(n8731) );
  AND2_X1 U9975 ( .A1(n8322), .A2(n12823), .ZN(n8336) );
  OR2_X1 U9976 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  AND2_X1 U9977 ( .A1(n8465), .A2(n9042), .ZN(n8484) );
  NAND2_X1 U9978 ( .A1(n8573), .A2(n8572), .ZN(n8589) );
  OR2_X1 U9979 ( .A1(n8711), .A2(n8710), .ZN(n8810) );
  INV_X1 U9980 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12823) );
  INV_X1 U9981 ( .A(n11564), .ZN(n11572) );
  AND2_X1 U9982 ( .A1(n10690), .A2(n10688), .ZN(n10695) );
  AND2_X1 U9983 ( .A1(n12579), .A2(n12580), .ZN(n13102) );
  AND3_X1 U9984 ( .A1(n8521), .A2(n8520), .A3(n8519), .ZN(n13222) );
  AND4_X1 U9985 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n13249)
         );
  INV_X1 U9986 ( .A(n12894), .ZN(n13286) );
  INV_X1 U9987 ( .A(n10813), .ZN(n12449) );
  AND2_X1 U9988 ( .A1(n8807), .A2(n10651), .ZN(n10655) );
  OR2_X1 U9989 ( .A1(n8262), .A2(n12383), .ZN(n8215) );
  INV_X1 U9990 ( .A(n10681), .ZN(n8509) );
  NAND2_X1 U9991 ( .A1(n8637), .A2(n12587), .ZN(n15588) );
  AND2_X1 U9992 ( .A1(n8708), .A2(n12424), .ZN(n15594) );
  AND2_X1 U9993 ( .A1(n8172), .A2(n8171), .ZN(n8504) );
  AND2_X1 U9994 ( .A1(n8165), .A2(n8164), .ZN(n8457) );
  INV_X1 U9995 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8407) );
  AND2_X1 U9996 ( .A1(n8138), .A2(n8137), .ZN(n8273) );
  INV_X1 U9997 ( .A(n9651), .ZN(n9660) );
  INV_X1 U9998 ( .A(n11622), .ZN(n9631) );
  INV_X1 U9999 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13540) );
  AND2_X1 U10000 ( .A1(n9590), .A2(n9591), .ZN(n10377) );
  NAND2_X1 U10001 ( .A1(n10014), .A2(n9754), .ZN(n10032) );
  AND2_X1 U10002 ( .A1(n9488), .A2(n9481), .ZN(n13779) );
  OR2_X1 U10003 ( .A1(n9435), .A2(n13510), .ZN(n9441) );
  OR2_X1 U10004 ( .A1(n15232), .A2(n14099), .ZN(n10253) );
  INV_X1 U10005 ( .A(n13650), .ZN(n9932) );
  INV_X1 U10006 ( .A(n10004), .ZN(n13871) );
  OR2_X1 U10007 ( .A1(n9386), .A2(n9385), .ZN(n9394) );
  NAND2_X1 U10008 ( .A1(n9528), .A2(n9527), .ZN(n11788) );
  NAND2_X1 U10009 ( .A1(n9743), .A2(n15362), .ZN(n13957) );
  INV_X1 U10010 ( .A(n9576), .ZN(n14001) );
  OR2_X1 U10011 ( .A1(n7993), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8007) );
  INV_X1 U10012 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7863) );
  NOR2_X1 U10013 ( .A1(n11664), .A2(n11663), .ZN(n11711) );
  NAND2_X1 U10014 ( .A1(n12635), .A2(n12634), .ZN(n12636) );
  INV_X1 U10015 ( .A(n12149), .ZN(n12054) );
  OR2_X1 U10016 ( .A1(n14203), .A2(n15102), .ZN(n14969) );
  NOR2_X1 U10017 ( .A1(n12080), .A2(n14202), .ZN(n12066) );
  INV_X1 U10018 ( .A(n10202), .ZN(n14283) );
  INV_X1 U10019 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11007) );
  INV_X1 U10020 ( .A(n11756), .ZN(n12087) );
  AND2_X1 U10021 ( .A1(n14477), .A2(n14447), .ZN(n14429) );
  INV_X1 U10022 ( .A(n14447), .ZN(n14488) );
  INV_X1 U10023 ( .A(n12299), .ZN(n14625) );
  INV_X1 U10024 ( .A(n14260), .ZN(n14137) );
  INV_X1 U10025 ( .A(n14259), .ZN(n14970) );
  AND2_X1 U10026 ( .A1(n10630), .A2(n10640), .ZN(n11226) );
  INV_X1 U10027 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9008) );
  AND2_X1 U10028 ( .A1(n10678), .A2(n15583), .ZN(n10659) );
  AND2_X1 U10029 ( .A1(P3_U3897), .A2(n12382), .ZN(n15508) );
  NAND2_X1 U10030 ( .A1(n8666), .A2(n8695), .ZN(n15599) );
  AND2_X1 U10031 ( .A1(n13216), .A2(n13215), .ZN(n13342) );
  AND2_X1 U10032 ( .A1(n15623), .A2(n14864), .ZN(n15535) );
  INV_X1 U10033 ( .A(n15590), .ZN(n15610) );
  AND2_X2 U10034 ( .A1(n10659), .A2(n15585), .ZN(n15576) );
  NAND2_X1 U10035 ( .A1(n10658), .A2(n10657), .ZN(n10661) );
  INV_X1 U10036 ( .A(n15605), .ZN(n15583) );
  AND4_X1 U10037 ( .A1(n10678), .A2(n8705), .A3(n8710), .A4(n8709), .ZN(n10658) );
  NOR2_X1 U10038 ( .A1(n15670), .A2(n8717), .ZN(n8718) );
  NAND2_X1 U10039 ( .A1(n10860), .A2(n10813), .ZN(n15605) );
  OR2_X1 U10040 ( .A1(n15599), .A2(n15662), .ZN(n15669) );
  AND2_X1 U10041 ( .A1(n10860), .A2(n15585), .ZN(n15662) );
  INV_X1 U10042 ( .A(n13588), .ZN(n13638) );
  AND2_X1 U10043 ( .A1(n10244), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13588) );
  OR2_X1 U10044 ( .A1(n15357), .A2(n10456), .ZN(n9742) );
  AND3_X1 U10045 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n9969) );
  INV_X1 U10046 ( .A(n9496), .ZN(n9472) );
  OR2_X1 U10047 ( .A1(n15232), .A2(n10264), .ZN(n15272) );
  INV_X1 U10048 ( .A(n15265), .ZN(n15298) );
  INV_X1 U10049 ( .A(n15272), .ZN(n15305) );
  INV_X1 U10050 ( .A(n9998), .ZN(n11429) );
  INV_X1 U10051 ( .A(n13961), .ZN(n15319) );
  INV_X1 U10052 ( .A(n13918), .ZN(n15314) );
  NAND2_X1 U10053 ( .A1(n15412), .A2(n15401), .ZN(n15370) );
  NAND2_X1 U10054 ( .A1(n8120), .A2(n8119), .ZN(n10457) );
  INV_X1 U10055 ( .A(n8118), .ZN(n15325) );
  INV_X1 U10056 ( .A(n10457), .ZN(n9735) );
  AND2_X1 U10057 ( .A1(n7994), .A2(n8007), .ZN(n11849) );
  AND2_X1 U10058 ( .A1(n12167), .A2(n12015), .ZN(n14496) );
  INV_X1 U10059 ( .A(n14203), .ZN(n14214) );
  AND4_X1 U10060 ( .A1(n12171), .A2(n12170), .A3(n12169), .A4(n12168), .ZN(
        n14469) );
  AND4_X1 U10061 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n14440) );
  INV_X1 U10062 ( .A(n10356), .ZN(n10359) );
  INV_X1 U10063 ( .A(n14398), .ZN(n15055) );
  INV_X1 U10064 ( .A(n14396), .ZN(n15060) );
  INV_X1 U10065 ( .A(n15099), .ZN(n14648) );
  NAND2_X1 U10066 ( .A1(n15103), .A2(n14990), .ZN(n15106) );
  INV_X1 U10067 ( .A(n14577), .ZN(n15080) );
  XNOR2_X1 U10068 ( .A(n12234), .B(n12235), .ZN(n12231) );
  AND2_X1 U10069 ( .A1(n10897), .A2(n11778), .ZN(n14997) );
  INV_X1 U10070 ( .A(n14623), .ZN(n14654) );
  AND2_X1 U10071 ( .A1(n10623), .A2(n10622), .ZN(n10944) );
  INV_X1 U10072 ( .A(n15146), .ZN(n15208) );
  AND2_X1 U10073 ( .A1(n10575), .A2(n10214), .ZN(n11218) );
  INV_X1 U10074 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10196) );
  AND2_X1 U10075 ( .A1(n10439), .A2(n10316), .ZN(n11704) );
  AND2_X1 U10076 ( .A1(n10690), .A2(n10689), .ZN(n15516) );
  AND3_X1 U10077 ( .A1(n8813), .A2(n8812), .A3(n12608), .ZN(n12896) );
  INV_X1 U10078 ( .A(n12924), .ZN(n12945) );
  INV_X1 U10079 ( .A(n13275), .ZN(n12949) );
  AND2_X2 U10080 ( .A1(n13426), .A2(n10071), .ZN(n10665) );
  MUX2_X1 U10081 ( .A(n10682), .B(n12950), .S(n12603), .Z(n15513) );
  INV_X1 U10082 ( .A(n14837), .ZN(n15523) );
  NAND2_X1 U10083 ( .A1(n15618), .A2(n10661), .ZN(n15623) );
  NAND2_X1 U10084 ( .A1(n15685), .A2(n15583), .ZN(n13364) );
  AOI21_X1 U10085 ( .B1(n8700), .B2(n8719), .A(n8718), .ZN(n8720) );
  INV_X2 U10086 ( .A(n15672), .ZN(n15670) );
  NAND2_X1 U10087 ( .A1(n13426), .A2(n10136), .ZN(n10137) );
  INV_X1 U10088 ( .A(SI_26_), .ZN(n11728) );
  INV_X1 U10089 ( .A(SI_16_), .ZN(n10171) );
  INV_X1 U10090 ( .A(SI_10_), .ZN(n10114) );
  INV_X1 U10091 ( .A(n11147), .ZN(n15458) );
  AND2_X1 U10092 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  OR3_X1 U10093 ( .A1(n15398), .A2(n9742), .A3(n9738), .ZN(n13630) );
  NAND2_X1 U10094 ( .A1(n9487), .A2(n9486), .ZN(n13648) );
  INV_X1 U10095 ( .A(n15307), .ZN(n15279) );
  OR2_X1 U10096 ( .A1(n6674), .A2(n10739), .ZN(n13961) );
  AND2_X1 U10097 ( .A1(n11293), .A2(n11292), .ZN(n15395) );
  OR2_X1 U10098 ( .A1(n6674), .A2(n10732), .ZN(n13966) );
  NAND2_X1 U10099 ( .A1(n15431), .A2(n15398), .ZN(n14046) );
  AND2_X2 U10100 ( .A1(n8125), .A2(n9735), .ZN(n15431) );
  INV_X1 U10101 ( .A(n13811), .ZN(n14059) );
  INV_X1 U10102 ( .A(n13907), .ZN(n14072) );
  AND2_X1 U10103 ( .A1(n15395), .A2(n15394), .ZN(n15427) );
  INV_X1 U10104 ( .A(n15420), .ZN(n15418) );
  INV_X1 U10105 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14107) );
  INV_X1 U10106 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10310) );
  INV_X1 U10107 ( .A(n14118), .ZN(n14241) );
  NAND2_X1 U10108 ( .A1(n11030), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14985) );
  INV_X1 U10109 ( .A(n14440), .ZN(n14585) );
  INV_X1 U10110 ( .A(n11634), .ZN(n14265) );
  OR2_X1 U10111 ( .A1(n10356), .A2(n10597), .ZN(n14396) );
  NAND2_X1 U10112 ( .A1(n10201), .A2(n10199), .ZN(n15064) );
  NAND2_X1 U10113 ( .A1(n15103), .A2(n14997), .ZN(n14623) );
  NAND2_X1 U10114 ( .A1(n10945), .A2(n11225), .ZN(n15210) );
  AND2_X2 U10115 ( .A1(n10624), .A2(n11218), .ZN(n15143) );
  INV_X1 U10116 ( .A(n10576), .ZN(n15149) );
  INV_X1 U10117 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10451) );
  INV_X1 U10118 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10222) );
  INV_X1 U10119 ( .A(n14763), .ZN(n14772) );
  INV_X1 U10120 ( .A(n12950), .ZN(P3_U3897) );
  NOR2_X1 U10121 ( .A1(P2_U3088), .A2(n10042), .ZN(P2_U3947) );
  NOR2_X1 U10122 ( .A1(n10575), .A2(n10069), .ZN(P1_U4016) );
  INV_X1 U10123 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8121) );
  INV_X1 U10124 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10103) );
  INV_X1 U10125 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8131) );
  AND2_X1 U10126 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7767) );
  NAND2_X1 U10127 ( .A1(n10593), .A2(n7767), .ZN(n10574) );
  NAND2_X1 U10128 ( .A1(n7774), .A2(SI_1_), .ZN(n7771) );
  OAI21_X1 U10129 ( .B1(n7768), .B2(n7770), .A(n7771), .ZN(n7769) );
  NAND2_X1 U10130 ( .A1(n7769), .A2(SI_2_), .ZN(n7777) );
  INV_X1 U10131 ( .A(SI_1_), .ZN(n10117) );
  OAI21_X1 U10132 ( .B1(SI_2_), .B2(n10117), .A(n7774), .ZN(n7773) );
  INV_X1 U10133 ( .A(SI_2_), .ZN(n10083) );
  NAND2_X1 U10134 ( .A1(n7773), .A2(n7772), .ZN(n7776) );
  OAI211_X1 U10135 ( .C1(n7774), .C2(SI_1_), .A(n7906), .B(n10083), .ZN(n7775)
         );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6671), .Z(n7920) );
  INV_X1 U10137 ( .A(SI_3_), .ZN(n10077) );
  NAND2_X1 U10138 ( .A1(n7778), .A2(SI_3_), .ZN(n7779) );
  NAND2_X1 U10139 ( .A1(n7780), .A2(SI_4_), .ZN(n7781) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n12052), .Z(n7783) );
  XNOR2_X1 U10141 ( .A(n7783), .B(SI_5_), .ZN(n7943) );
  INV_X1 U10142 ( .A(n7943), .ZN(n7782) );
  NAND2_X1 U10143 ( .A1(n7783), .A2(SI_5_), .ZN(n7784) );
  MUX2_X1 U10144 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6672), .Z(n7786) );
  XNOR2_X1 U10145 ( .A(n7786), .B(SI_6_), .ZN(n7947) );
  INV_X1 U10146 ( .A(n7947), .ZN(n7785) );
  NAND2_X1 U10147 ( .A1(n7786), .A2(SI_6_), .ZN(n7787) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6671), .Z(n7789) );
  XNOR2_X1 U10149 ( .A(n7789), .B(SI_7_), .ZN(n7952) );
  INV_X1 U10150 ( .A(n7952), .ZN(n7788) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6673), .Z(n7790) );
  XNOR2_X1 U10152 ( .A(n7790), .B(SI_8_), .ZN(n7958) );
  NAND2_X1 U10153 ( .A1(n7790), .A2(SI_8_), .ZN(n7791) );
  NAND2_X1 U10154 ( .A1(n7792), .A2(n7791), .ZN(n7965) );
  MUX2_X1 U10155 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6673), .Z(n7794) );
  XNOR2_X1 U10156 ( .A(n7794), .B(SI_9_), .ZN(n7964) );
  INV_X1 U10157 ( .A(n7964), .ZN(n7793) );
  NAND2_X1 U10158 ( .A1(n7794), .A2(SI_9_), .ZN(n7795) );
  MUX2_X1 U10159 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6672), .Z(n7970) );
  INV_X1 U10160 ( .A(n7970), .ZN(n7796) );
  NAND2_X1 U10161 ( .A1(n7796), .A2(n10114), .ZN(n7797) );
  MUX2_X1 U10162 ( .A(n10179), .B(n10172), .S(n6672), .Z(n7798) );
  NAND2_X1 U10163 ( .A1(n7798), .A2(n10116), .ZN(n7801) );
  INV_X1 U10164 ( .A(n7798), .ZN(n7799) );
  NAND2_X1 U10165 ( .A1(n7799), .A2(SI_11_), .ZN(n7800) );
  NAND2_X1 U10166 ( .A1(n7801), .A2(n7800), .ZN(n7976) );
  MUX2_X1 U10167 ( .A(n10222), .B(n10219), .S(n6672), .Z(n7802) );
  NAND2_X1 U10168 ( .A1(n7802), .A2(n10131), .ZN(n7805) );
  INV_X1 U10169 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U10170 ( .A1(n7803), .A2(SI_12_), .ZN(n7804) );
  MUX2_X1 U10171 ( .A(n10317), .B(n10310), .S(n6673), .Z(n7987) );
  INV_X1 U10172 ( .A(n7987), .ZN(n7806) );
  NAND2_X1 U10173 ( .A1(n7806), .A2(SI_13_), .ZN(n7807) );
  NAND2_X1 U10174 ( .A1(n7987), .A2(n10139), .ZN(n7808) );
  MUX2_X1 U10175 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6672), .Z(n7810) );
  NAND2_X1 U10176 ( .A1(n7810), .A2(SI_15_), .ZN(n7811) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6673), .Z(n8002) );
  NAND2_X1 U10178 ( .A1(n8002), .A2(SI_14_), .ZN(n7809) );
  NOR2_X1 U10179 ( .A1(n8002), .A2(SI_14_), .ZN(n7812) );
  INV_X1 U10180 ( .A(n7810), .ZN(n8004) );
  AOI22_X1 U10181 ( .A1(n7812), .A2(n7811), .B1(n10161), .B2(n8004), .ZN(n7813) );
  MUX2_X1 U10182 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n6672), .Z(n7814) );
  XNOR2_X1 U10183 ( .A(n7814), .B(n10171), .ZN(n8011) );
  INV_X1 U10184 ( .A(n7814), .ZN(n7815) );
  MUX2_X1 U10185 ( .A(n10451), .B(n10453), .S(n6672), .Z(n8018) );
  NOR2_X1 U10186 ( .A1(n7816), .A2(SI_17_), .ZN(n7818) );
  NAND2_X1 U10187 ( .A1(n7816), .A2(SI_17_), .ZN(n7817) );
  MUX2_X1 U10188 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6672), .Z(n8026) );
  NAND2_X1 U10189 ( .A1(n7819), .A2(SI_18_), .ZN(n7820) );
  MUX2_X1 U10190 ( .A(n12074), .B(n11196), .S(n6672), .Z(n7821) );
  INV_X1 U10191 ( .A(n7821), .ZN(n7822) );
  NAND2_X1 U10192 ( .A1(n7822), .A2(SI_19_), .ZN(n7823) );
  NAND2_X1 U10193 ( .A1(n7824), .A2(n7823), .ZN(n8033) );
  MUX2_X1 U10194 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6672), .Z(n7902) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6672), .Z(n7826) );
  XNOR2_X1 U10196 ( .A(n7826), .B(SI_21_), .ZN(n7899) );
  NAND2_X1 U10197 ( .A1(n7826), .A2(SI_21_), .ZN(n7827) );
  NAND2_X1 U10198 ( .A1(n7828), .A2(n7827), .ZN(n7888) );
  MUX2_X1 U10199 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6672), .Z(n7896) );
  MUX2_X1 U10200 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6672), .Z(n7891) );
  INV_X1 U10201 ( .A(n7891), .ZN(n7829) );
  INV_X1 U10202 ( .A(SI_23_), .ZN(n11054) );
  NAND2_X1 U10203 ( .A1(n7829), .A2(n11054), .ZN(n7833) );
  OAI21_X1 U10204 ( .B1(SI_22_), .B2(n7896), .A(n7833), .ZN(n7830) );
  INV_X1 U10205 ( .A(n7830), .ZN(n7831) );
  INV_X1 U10206 ( .A(n7896), .ZN(n7832) );
  INV_X1 U10207 ( .A(SI_22_), .ZN(n8546) );
  NOR2_X1 U10208 ( .A1(n7832), .A2(n8546), .ZN(n7834) );
  AOI22_X1 U10209 ( .A1(n7834), .A2(n7833), .B1(n7891), .B2(SI_23_), .ZN(n7835) );
  MUX2_X1 U10210 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6672), .Z(n8040) );
  INV_X1 U10211 ( .A(n8040), .ZN(n7839) );
  NAND2_X1 U10212 ( .A1(n7837), .A2(SI_24_), .ZN(n7838) );
  INV_X1 U10213 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12625) );
  INV_X1 U10214 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14112) );
  MUX2_X1 U10215 ( .A(n12625), .B(n14112), .S(n6673), .Z(n7840) );
  INV_X1 U10216 ( .A(SI_25_), .ZN(n11597) );
  NAND2_X1 U10217 ( .A1(n7840), .A2(n11597), .ZN(n7843) );
  INV_X1 U10218 ( .A(n7840), .ZN(n7841) );
  NAND2_X1 U10219 ( .A1(n7841), .A2(SI_25_), .ZN(n7842) );
  NAND2_X1 U10220 ( .A1(n7843), .A2(n7842), .ZN(n8044) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n6672), .Z(n8048) );
  INV_X1 U10222 ( .A(n8048), .ZN(n7845) );
  NAND2_X1 U10223 ( .A1(n8050), .A2(n11728), .ZN(n7846) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6672), .Z(n7881) );
  NOR2_X1 U10225 ( .A1(n7881), .A2(SI_27_), .ZN(n7849) );
  NAND2_X1 U10226 ( .A1(n7881), .A2(SI_27_), .ZN(n7848) );
  MUX2_X1 U10227 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6673), .Z(n7850) );
  XNOR2_X1 U10228 ( .A(n7850), .B(SI_28_), .ZN(n8053) );
  INV_X1 U10229 ( .A(n7850), .ZN(n7851) );
  INV_X1 U10230 ( .A(SI_28_), .ZN(n12383) );
  NAND2_X1 U10231 ( .A1(n7851), .A2(n12383), .ZN(n7852) );
  MUX2_X1 U10232 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6672), .Z(n7853) );
  INV_X1 U10233 ( .A(SI_29_), .ZN(n13440) );
  XNOR2_X1 U10234 ( .A(n7853), .B(n13440), .ZN(n8057) );
  INV_X1 U10235 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U10236 ( .A1(n7854), .A2(n13440), .ZN(n7855) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6673), .Z(n7857) );
  INV_X1 U10238 ( .A(SI_30_), .ZN(n12414) );
  XNOR2_X1 U10239 ( .A(n7857), .B(n12414), .ZN(n7878) );
  INV_X1 U10240 ( .A(n7878), .ZN(n7859) );
  NAND2_X1 U10241 ( .A1(n7857), .A2(SI_30_), .ZN(n7858) );
  OAI21_X1 U10242 ( .B1(n7879), .B2(n7859), .A(n7858), .ZN(n7862) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6672), .Z(n7860) );
  XNOR2_X1 U10244 ( .A(n7860), .B(SI_31_), .ZN(n7861) );
  XNOR2_X1 U10245 ( .A(n7862), .B(n7861), .ZN(n14083) );
  NOR2_X1 U10246 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n7868) );
  NAND4_X1 U10247 ( .A1(n7869), .A2(n8063), .A3(n8069), .A4(n8062), .ZN(n7871)
         );
  NAND4_X1 U10248 ( .A1(n7738), .A2(n8028), .A3(n8021), .A4(n8114), .ZN(n7870)
         );
  NOR2_X1 U10249 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  NAND2_X1 U10250 ( .A1(n8073), .A2(n8075), .ZN(n8082) );
  NAND3_X1 U10251 ( .A1(n8081), .A2(P2_IR_REG_31__SCAN_IN), .A3(n8075), .ZN(
        n7874) );
  NAND2_X1 U10252 ( .A1(n14083), .A2(n8061), .ZN(n7877) );
  INV_X1 U10253 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7875) );
  OR2_X1 U10254 ( .A1(n8059), .A2(n7875), .ZN(n7876) );
  INV_X1 U10255 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14091) );
  NOR2_X1 U10256 ( .A1(n8059), .A2(n14091), .ZN(n7880) );
  INV_X1 U10257 ( .A(n7881), .ZN(n7882) );
  XNOR2_X1 U10258 ( .A(n7882), .B(SI_27_), .ZN(n7883) );
  XNOR2_X1 U10259 ( .A(n7884), .B(n7883), .ZN(n14102) );
  NAND2_X1 U10260 ( .A1(n14102), .A2(n8061), .ZN(n7886) );
  INV_X1 U10261 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14103) );
  OR2_X1 U10262 ( .A1(n8059), .A2(n14103), .ZN(n7885) );
  INV_X1 U10263 ( .A(n12053), .ZN(n7887) );
  NAND2_X1 U10264 ( .A1(n7887), .A2(n7896), .ZN(n7890) );
  NAND2_X1 U10265 ( .A1(n7888), .A2(SI_22_), .ZN(n7889) );
  NAND2_X1 U10266 ( .A1(n7890), .A2(n7889), .ZN(n7893) );
  XNOR2_X1 U10267 ( .A(n7891), .B(SI_23_), .ZN(n7892) );
  NAND2_X1 U10268 ( .A1(n12144), .A2(n8061), .ZN(n7895) );
  INV_X1 U10269 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11889) );
  OR2_X1 U10270 ( .A1(n8059), .A2(n11889), .ZN(n7894) );
  XNOR2_X1 U10271 ( .A(n12053), .B(n7896), .ZN(n11838) );
  NAND2_X1 U10272 ( .A1(n11838), .A2(n8061), .ZN(n7898) );
  INV_X1 U10273 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11840) );
  OR2_X1 U10274 ( .A1(n8059), .A2(n11840), .ZN(n7897) );
  XNOR2_X1 U10275 ( .A(n6796), .B(n7899), .ZN(n12041) );
  NAND2_X1 U10276 ( .A1(n12041), .A2(n8061), .ZN(n7901) );
  INV_X1 U10277 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12610) );
  OR2_X1 U10278 ( .A1(n8059), .A2(n12610), .ZN(n7900) );
  XNOR2_X1 U10279 ( .A(n7903), .B(n7902), .ZN(n12061) );
  NAND2_X1 U10280 ( .A1(n12061), .A2(n8061), .ZN(n7905) );
  INV_X1 U10281 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11526) );
  OR2_X1 U10282 ( .A1(n8059), .A2(n11526), .ZN(n7904) );
  INV_X1 U10283 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15236) );
  INV_X1 U10284 ( .A(n7909), .ZN(n7910) );
  OR2_X1 U10285 ( .A1(n10031), .A2(n10254), .ZN(n7911) );
  AND3_X2 U10286 ( .A1(n7913), .A2(n7912), .A3(n7911), .ZN(n15366) );
  NAND2_X1 U10287 ( .A1(n8241), .A2(n8129), .ZN(n7914) );
  NAND2_X1 U10288 ( .A1(n7915), .A2(n7914), .ZN(n14113) );
  MUX2_X1 U10289 ( .A(n15236), .B(n14113), .S(n10031), .Z(n12400) );
  NAND2_X1 U10290 ( .A1(n15366), .A2(n12400), .ZN(n11093) );
  NOR2_X1 U10291 ( .A1(n7909), .A2(n14085), .ZN(n7916) );
  MUX2_X1 U10292 ( .A(n14085), .B(n7916), .S(P2_IR_REG_2__SCAN_IN), .Z(n7917)
         );
  INV_X1 U10293 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10294 ( .A1(n7918), .A2(n7927), .ZN(n10256) );
  INV_X1 U10295 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10100) );
  OR2_X1 U10296 ( .A1(n8059), .A2(n10100), .ZN(n7923) );
  OR2_X1 U10297 ( .A1(n7921), .A2(n10822), .ZN(n7922) );
  OR2_X1 U10298 ( .A1(n11093), .A2(n15315), .ZN(n10741) );
  INV_X1 U10299 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10101) );
  OR2_X1 U10300 ( .A1(n8059), .A2(n10101), .ZN(n7930) );
  NAND2_X1 U10301 ( .A1(n7927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  MUX2_X1 U10302 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7926), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7928) );
  OR2_X1 U10303 ( .A1(n7927), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10304 ( .A1(n7928), .A2(n7935), .ZN(n10258) );
  OR2_X1 U10305 ( .A1(n10031), .A2(n10258), .ZN(n7929) );
  INV_X1 U10306 ( .A(n15379), .ZN(n10742) );
  NOR2_X2 U10307 ( .A1(n10741), .A2(n10742), .ZN(n10740) );
  NAND2_X1 U10308 ( .A1(n7935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7932) );
  INV_X1 U10309 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7936) );
  XNOR2_X1 U10310 ( .A(n7932), .B(n7936), .ZN(n10282) );
  NAND2_X1 U10311 ( .A1(n10740), .A2(n10727), .ZN(n10717) );
  INV_X1 U10312 ( .A(n7935), .ZN(n7937) );
  NAND2_X1 U10313 ( .A1(n7937), .A2(n7936), .ZN(n7939) );
  NAND2_X1 U10314 ( .A1(n7939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7938) );
  MUX2_X1 U10315 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7938), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7942) );
  INV_X1 U10316 ( .A(n7939), .ZN(n7941) );
  NAND2_X1 U10317 ( .A1(n7941), .A2(n7940), .ZN(n7954) );
  NAND2_X1 U10318 ( .A1(n7942), .A2(n7954), .ZN(n10283) );
  XNOR2_X1 U10319 ( .A(n7944), .B(n7943), .ZN(n10962) );
  NAND2_X1 U10320 ( .A1(n10962), .A2(n8061), .ZN(n7946) );
  OR2_X1 U10321 ( .A1(n8059), .A2(n10128), .ZN(n7945) );
  OAI211_X1 U10322 ( .C1(n10031), .C2(n10283), .A(n7946), .B(n7945), .ZN(n9791) );
  OR2_X1 U10323 ( .A1(n10717), .A2(n9791), .ZN(n11067) );
  XNOR2_X1 U10324 ( .A(n7948), .B(n7947), .ZN(n10968) );
  NAND2_X1 U10325 ( .A1(n10968), .A2(n8061), .ZN(n7951) );
  NAND2_X1 U10326 ( .A1(n7954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7949) );
  XNOR2_X1 U10327 ( .A(n7949), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U10328 ( .A1(n7908), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8037), .B2(
        n10284), .ZN(n7950) );
  NAND2_X1 U10329 ( .A1(n7951), .A2(n7950), .ZN(n11208) );
  XNOR2_X1 U10330 ( .A(n7953), .B(n7952), .ZN(n10980) );
  NAND2_X1 U10331 ( .A1(n10980), .A2(n8061), .ZN(n7957) );
  OAI21_X1 U10332 ( .B1(n7954), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7955) );
  XNOR2_X1 U10333 ( .A(n7955), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U10334 ( .A1(n7908), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8037), .B2(
        n10397), .ZN(n7956) );
  NAND2_X1 U10335 ( .A1(n7957), .A2(n7956), .ZN(n11418) );
  INV_X1 U10336 ( .A(n11418), .ZN(n11244) );
  NAND2_X1 U10337 ( .A1(n10993), .A2(n8061), .ZN(n7963) );
  OR2_X1 U10338 ( .A1(n7960), .A2(n6916), .ZN(n7961) );
  XNOR2_X1 U10339 ( .A(n7961), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U10340 ( .A1(n7908), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8037), .B2(
        n11106), .ZN(n7962) );
  NAND2_X1 U10341 ( .A1(n7963), .A2(n7962), .ZN(n13498) );
  INV_X1 U10342 ( .A(n13498), .ZN(n15391) );
  XNOR2_X1 U10343 ( .A(n7965), .B(n7964), .ZN(n11264) );
  NAND2_X1 U10344 ( .A1(n11264), .A2(n8061), .ZN(n7969) );
  NAND2_X1 U10345 ( .A1(n7966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7967) );
  XNOR2_X1 U10346 ( .A(n7967), .B(P2_IR_REG_9__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U10347 ( .A1(n7908), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8037), .B2(
        n15267), .ZN(n7968) );
  XNOR2_X1 U10348 ( .A(n7970), .B(SI_10_), .ZN(n7971) );
  XNOR2_X1 U10349 ( .A(n7972), .B(n7971), .ZN(n11470) );
  NAND2_X1 U10350 ( .A1(n11470), .A2(n8061), .ZN(n7975) );
  NAND2_X1 U10351 ( .A1(n6859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7973) );
  XNOR2_X1 U10352 ( .A(n7973), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U10353 ( .A1(n7908), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8037), 
        .B2(n11108), .ZN(n7974) );
  XNOR2_X1 U10354 ( .A(n7977), .B(n7976), .ZN(n11454) );
  NAND2_X1 U10355 ( .A1(n11454), .A2(n8061), .ZN(n7980) );
  OR2_X1 U10356 ( .A1(n6859), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10357 ( .A1(n7982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7978) );
  XNOR2_X1 U10358 ( .A(n7978), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U10359 ( .A1(n7908), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8037), 
        .B2(n11332), .ZN(n7979) );
  INV_X1 U10360 ( .A(n11607), .ZN(n15410) );
  XNOR2_X1 U10361 ( .A(n7981), .B(n7761), .ZN(n11659) );
  NAND2_X1 U10362 ( .A1(n11659), .A2(n8061), .ZN(n7986) );
  INV_X1 U10363 ( .A(n7991), .ZN(n7983) );
  NAND2_X1 U10364 ( .A1(n7983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7984) );
  XNOR2_X1 U10365 ( .A(n7984), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U10366 ( .A1(n7908), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8037), 
        .B2(n11687), .ZN(n7985) );
  XNOR2_X1 U10367 ( .A(n7987), .B(SI_13_), .ZN(n7988) );
  XNOR2_X1 U10368 ( .A(n7989), .B(n7988), .ZN(n11703) );
  NAND2_X1 U10369 ( .A1(n11703), .A2(n8061), .ZN(n7996) );
  NAND2_X1 U10370 ( .A1(n7991), .A2(n7990), .ZN(n7993) );
  NAND2_X1 U10371 ( .A1(n7993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7992) );
  MUX2_X1 U10372 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7992), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7994) );
  AOI22_X1 U10373 ( .A1(n7908), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8037), 
        .B2(n11849), .ZN(n7995) );
  INV_X1 U10374 ( .A(SI_14_), .ZN(n10148) );
  XNOR2_X1 U10375 ( .A(n7997), .B(n10148), .ZN(n8003) );
  XNOR2_X1 U10376 ( .A(n8003), .B(n8002), .ZN(n11915) );
  NAND2_X1 U10377 ( .A1(n11915), .A2(n8061), .ZN(n8000) );
  NAND2_X1 U10378 ( .A1(n8007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7998) );
  XNOR2_X1 U10379 ( .A(n7998), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U10380 ( .A1(n7908), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8037), 
        .B2(n13681), .ZN(n7999) );
  INV_X1 U10381 ( .A(n7997), .ZN(n8001) );
  OAI22_X1 U10382 ( .A1(n8003), .A2(n8002), .B1(n8001), .B2(SI_14_), .ZN(n8006) );
  XNOR2_X1 U10383 ( .A(n8004), .B(SI_15_), .ZN(n8005) );
  XNOR2_X1 U10384 ( .A(n8006), .B(n8005), .ZN(n11920) );
  NAND2_X1 U10385 ( .A1(n11920), .A2(n8061), .ZN(n8010) );
  OAI21_X1 U10386 ( .B1(n8007), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8008) );
  XNOR2_X1 U10387 ( .A(n8008), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U10388 ( .A1(n7908), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8037), 
        .B2(n15292), .ZN(n8009) );
  XNOR2_X1 U10389 ( .A(n8012), .B(n8011), .ZN(n12086) );
  NAND2_X1 U10390 ( .A1(n12086), .A2(n8061), .ZN(n8017) );
  AND2_X2 U10391 ( .A1(n8013), .A2(n7757), .ZN(n8022) );
  INV_X1 U10392 ( .A(n8022), .ZN(n8014) );
  NAND2_X1 U10393 ( .A1(n8014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U10394 ( .A(n8015), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U10395 ( .A1(n7908), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8037), 
        .B2(n13703), .ZN(n8016) );
  XNOR2_X1 U10396 ( .A(n8018), .B(SI_17_), .ZN(n8019) );
  XNOR2_X1 U10397 ( .A(n8020), .B(n8019), .ZN(n12090) );
  NAND2_X1 U10398 ( .A1(n12090), .A2(n8061), .ZN(n8025) );
  OR2_X1 U10399 ( .A1(n8029), .A2(n6916), .ZN(n8023) );
  XNOR2_X1 U10400 ( .A(n8023), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U10401 ( .A1(n7908), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8037), 
        .B2(n15304), .ZN(n8024) );
  XNOR2_X1 U10402 ( .A(n8027), .B(n8026), .ZN(n12115) );
  NAND2_X1 U10403 ( .A1(n12115), .A2(n8061), .ZN(n8032) );
  NAND2_X1 U10404 ( .A1(n8035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8030) );
  XNOR2_X1 U10405 ( .A(n8030), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13718) );
  AOI22_X1 U10406 ( .A1(n7908), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8037), 
        .B2(n13718), .ZN(n8031) );
  XNOR2_X1 U10407 ( .A(n8034), .B(n8033), .ZN(n12073) );
  NAND2_X1 U10408 ( .A1(n12073), .A2(n8061), .ZN(n8039) );
  XNOR2_X2 U10409 ( .A(n8036), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U10410 ( .A1(n7908), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8037), 
        .B2(n10739), .ZN(n8038) );
  NAND2_X1 U10411 ( .A1(n13915), .A2(n14072), .ZN(n13903) );
  XNOR2_X1 U10412 ( .A(n8041), .B(n8040), .ZN(n12134) );
  NAND2_X1 U10413 ( .A1(n12134), .A2(n8061), .ZN(n8043) );
  INV_X1 U10414 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11893) );
  OR2_X1 U10415 ( .A1(n8059), .A2(n11893), .ZN(n8042) );
  NOR2_X4 U10416 ( .A1(n13844), .A2(n13996), .ZN(n13827) );
  XNOR2_X1 U10417 ( .A(n8045), .B(n8044), .ZN(n12624) );
  NAND2_X1 U10418 ( .A1(n12624), .A2(n8061), .ZN(n8047) );
  OR2_X1 U10419 ( .A1(n8059), .A2(n14112), .ZN(n8046) );
  XNOR2_X1 U10420 ( .A(n8048), .B(n11728), .ZN(n8049) );
  NAND2_X1 U10421 ( .A1(n14105), .A2(n8061), .ZN(n8052) );
  OR2_X1 U10422 ( .A1(n8059), .A2(n14107), .ZN(n8051) );
  NAND2_X1 U10423 ( .A1(n14769), .A2(n8061), .ZN(n8056) );
  INV_X1 U10424 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14101) );
  OR2_X1 U10425 ( .A1(n8059), .A2(n14101), .ZN(n8055) );
  INV_X1 U10426 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14096) );
  NOR2_X1 U10427 ( .A1(n8059), .A2(n14096), .ZN(n8060) );
  AND2_X2 U10428 ( .A1(n13759), .A2(n13748), .ZN(n13738) );
  INV_X1 U10429 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10430 ( .A1(n6916), .A2(n8063), .ZN(n8065) );
  XNOR2_X2 U10431 ( .A(n8070), .B(n8069), .ZN(n8122) );
  AND2_X2 U10432 ( .A1(n8090), .A2(n8122), .ZN(n9576) );
  NOR2_X2 U10433 ( .A1(n8071), .A2(n14001), .ZN(n13732) );
  INV_X1 U10434 ( .A(n8072), .ZN(n8074) );
  NAND2_X1 U10435 ( .A1(n8074), .A2(n8073), .ZN(n8078) );
  NAND2_X1 U10436 ( .A1(n8078), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8076) );
  INV_X1 U10437 ( .A(n10263), .ZN(n15231) );
  INV_X2 U10438 ( .A(n13449), .ZN(n13610) );
  NAND2_X1 U10439 ( .A1(n8078), .A2(n8077), .ZN(n14104) );
  INV_X1 U10440 ( .A(P2_B_REG_SCAN_IN), .ZN(n8079) );
  OR2_X1 U10441 ( .A1(n14104), .A2(n8079), .ZN(n8080) );
  NAND2_X1 U10442 ( .A1(n13610), .A2(n8080), .ZN(n9565) );
  NOR2_X2 U10443 ( .A1(n8083), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8085) );
  BUF_X1 U10444 ( .A(n8085), .Z(n14084) );
  OR2_X2 U10445 ( .A1(n8085), .A2(n14085), .ZN(n8086) );
  XNOR2_X2 U10446 ( .A(n8086), .B(P2_IR_REG_30__SCAN_IN), .ZN(n14090) );
  NOR2_X2 U10447 ( .A1(n14097), .A2(n14090), .ZN(n9278) );
  NAND2_X1 U10448 ( .A1(n9559), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8089) );
  AND2_X2 U10449 ( .A1(n14097), .A2(n14090), .ZN(n9280) );
  NAND2_X1 U10450 ( .A1(n9420), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8088) );
  NOR2_X2 U10451 ( .A1(n14090), .A2(n9264), .ZN(n9281) );
  NAND2_X1 U10452 ( .A1(n9560), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8087) );
  NOR2_X1 U10453 ( .A1(n9565), .A2(n9969), .ZN(n13733) );
  NOR2_X1 U10454 ( .A1(n13732), .A2(n13733), .ZN(n8126) );
  INV_X1 U10455 ( .A(n8090), .ZN(n10224) );
  NOR4_X1 U10456 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8094) );
  NOR4_X1 U10457 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8093) );
  NOR4_X1 U10458 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8092) );
  NOR4_X1 U10459 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8091) );
  NAND4_X1 U10460 ( .A1(n8094), .A2(n8093), .A3(n8092), .A4(n8091), .ZN(n8110)
         );
  NOR2_X1 U10461 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8098) );
  NOR4_X1 U10462 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8097) );
  NOR4_X1 U10463 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8096) );
  NOR4_X1 U10464 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8095) );
  NAND4_X1 U10465 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(n8109)
         );
  NAND2_X1 U10466 ( .A1(n8099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8100) );
  MUX2_X1 U10467 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8100), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8101) );
  NAND2_X1 U10468 ( .A1(n8101), .A2(n6832), .ZN(n14109) );
  OR2_X1 U10469 ( .A1(n8102), .A2(n6916), .ZN(n8104) );
  MUX2_X1 U10470 ( .A(n8104), .B(P2_IR_REG_31__SCAN_IN), .S(n8103), .Z(n8105)
         );
  NAND2_X1 U10471 ( .A1(n8105), .A2(n8099), .ZN(n11892) );
  XNOR2_X1 U10472 ( .A(n11892), .B(P2_B_REG_SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10473 ( .A1(n6832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8107) );
  OR2_X1 U10474 ( .A1(n8108), .A2(n14108), .ZN(n8118) );
  OAI21_X1 U10475 ( .B1(n8110), .B2(n8109), .A(n15325), .ZN(n9736) );
  OR2_X1 U10476 ( .A1(n8118), .A2(P2_D_REG_1__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10477 ( .A1(n14108), .A2(n14109), .ZN(n8111) );
  NAND2_X1 U10478 ( .A1(n8112), .A2(n8111), .ZN(n15361) );
  NAND3_X1 U10479 ( .A1(n9736), .A2(n15361), .A3(P2_STATE_REG_SCAN_IN), .ZN(
        n8113) );
  NOR2_X1 U10480 ( .A1(n9743), .A2(n8113), .ZN(n8117) );
  INV_X1 U10481 ( .A(n10032), .ZN(n9738) );
  NAND2_X1 U10482 ( .A1(n8122), .A2(n13726), .ZN(n10037) );
  NOR3_X1 U10483 ( .A1(n14108), .A2(n11892), .A3(n14109), .ZN(n10034) );
  INV_X1 U10484 ( .A(n10034), .ZN(n9733) );
  NAND2_X1 U10485 ( .A1(n10035), .A2(n9733), .ZN(n8116) );
  AND2_X1 U10486 ( .A1(n8117), .A2(n10459), .ZN(n8125) );
  OR2_X1 U10487 ( .A1(n8118), .A2(P2_D_REG_0__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10488 ( .A1(n14108), .A2(n11892), .ZN(n8119) );
  MUX2_X1 U10489 ( .A(n8121), .B(n8126), .S(n15431), .Z(n8124) );
  NAND2_X1 U10490 ( .A1(n8090), .A2(n9993), .ZN(n10743) );
  NAND2_X1 U10491 ( .A1(n8090), .A2(n10739), .ZN(n8123) );
  NAND2_X1 U10492 ( .A1(n8124), .A2(n7752), .ZN(P2_U3530) );
  INV_X1 U10493 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8127) );
  MUX2_X1 U10494 ( .A(n8127), .B(n8126), .S(n15420), .Z(n8128) );
  NAND2_X1 U10495 ( .A1(n15420), .A2(n15398), .ZN(n14081) );
  NAND2_X1 U10496 ( .A1(n8128), .A2(n7753), .ZN(P2_U3498) );
  INV_X1 U10497 ( .A(n8240), .ZN(n8130) );
  NAND2_X1 U10498 ( .A1(n8131), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U10499 ( .A1(n10100), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8134) );
  INV_X1 U10500 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U10501 ( .A1(n10819), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8133) );
  AND2_X1 U10502 ( .A1(n8134), .A2(n8133), .ZN(n8248) );
  NAND2_X1 U10503 ( .A1(n10101), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8136) );
  INV_X1 U10504 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U10505 ( .A1(n10096), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U10506 ( .A1(n10111), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8138) );
  INV_X1 U10507 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U10508 ( .A1(n10110), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10509 ( .A1(n8274), .A2(n8273), .ZN(n8139) );
  NAND2_X1 U10510 ( .A1(n10128), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10511 ( .A1(n10126), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10512 ( .A1(n10134), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10513 ( .A1(n10132), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10514 ( .A1(n10144), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10515 ( .A1(n10146), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10516 ( .A1(n8145), .A2(n8144), .ZN(n8314) );
  NAND2_X1 U10517 ( .A1(n10153), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10518 ( .A1(n10150), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10519 ( .A1(n10158), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U10520 ( .A1(n10156), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10521 ( .A1(n8348), .A2(n8149), .ZN(n8365) );
  NAND2_X1 U10522 ( .A1(n10165), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10523 ( .A1(n10167), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10524 ( .A1(n8365), .A2(n8364), .ZN(n8367) );
  NAND2_X1 U10525 ( .A1(n10172), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10526 ( .A1(n8383), .A2(n8152), .ZN(n8154) );
  NAND2_X1 U10527 ( .A1(n10179), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8153) );
  XNOR2_X1 U10528 ( .A(n10219), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8396) );
  INV_X1 U10529 ( .A(n8396), .ZN(n8155) );
  NAND2_X1 U10530 ( .A1(n10222), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U10531 ( .A1(n8157), .A2(n10317), .ZN(n8158) );
  NAND2_X1 U10532 ( .A1(n10438), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10533 ( .A1(n10550), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10534 ( .A1(n10552), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10535 ( .A1(n8163), .A2(n8162), .ZN(n8441) );
  NAND2_X1 U10536 ( .A1(n10436), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8165) );
  INV_X1 U10537 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U10538 ( .A1(n10430), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10539 ( .A1(n10451), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10540 ( .A1(n10453), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10541 ( .A1(n12117), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8170) );
  INV_X1 U10542 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U10543 ( .A1(n10950), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10544 ( .A1(n8170), .A2(n8168), .ZN(n8491) );
  INV_X1 U10545 ( .A(n8491), .ZN(n8169) );
  NAND2_X1 U10546 ( .A1(n12074), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10547 ( .A1(n11196), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8171) );
  INV_X1 U10548 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U10549 ( .A1(n12042), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10550 ( .A1(n12610), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10551 ( .A1(n8175), .A2(n8174), .ZN(n8531) );
  XNOR2_X1 U10552 ( .A(n11840), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10553 ( .A1(n11840), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8177) );
  XNOR2_X1 U10554 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8558) );
  NAND2_X1 U10555 ( .A1(n8178), .A2(n11893), .ZN(n8179) );
  NAND2_X1 U10556 ( .A1(n14112), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10557 ( .A1(n12625), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8182) );
  NOR2_X1 U10558 ( .A1(n14107), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10559 ( .A1(n14107), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8184) );
  AND2_X1 U10560 ( .A1(n14103), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8185) );
  INV_X1 U10561 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14773) );
  NAND2_X1 U10562 ( .A1(n14773), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8186) );
  NOR2_X1 U10563 ( .A1(n14101), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8188) );
  INV_X1 U10564 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14770) );
  XNOR2_X1 U10565 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12401) );
  XNOR2_X1 U10566 ( .A(n12402), .B(n12401), .ZN(n13436) );
  NAND2_X4 U10567 ( .A1(n8635), .A2(n8636), .ZN(n10681) );
  NAND2_X1 U10568 ( .A1(n13436), .A2(n12417), .ZN(n8200) );
  OR2_X1 U10569 ( .A1(n12415), .A2(n13440), .ZN(n8199) );
  NAND2_X1 U10570 ( .A1(n8200), .A2(n8199), .ZN(n8700) );
  NAND2_X1 U10571 ( .A1(n8278), .A2(n8277), .ZN(n8292) );
  NAND2_X1 U10572 ( .A1(n8336), .A2(n8335), .ZN(n8351) );
  NAND2_X1 U10573 ( .A1(n8418), .A2(n8417), .ZN(n8432) );
  INV_X1 U10574 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8572) );
  INV_X1 U10575 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8217) );
  INV_X1 U10576 ( .A(n12623), .ZN(n8208) );
  NAND2_X1 U10577 ( .A1(n13064), .A2(n8619), .ZN(n10882) );
  INV_X1 U10578 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8701) );
  INV_X2 U10579 ( .A(n8254), .ZN(n8639) );
  NAND2_X1 U10580 ( .A1(n8639), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10581 ( .A1(n8537), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8209) );
  OAI211_X1 U10582 ( .C1(n8701), .C2(n8516), .A(n8210), .B(n8209), .ZN(n8211)
         );
  INV_X1 U10583 ( .A(n8211), .ZN(n8212) );
  OR2_X1 U10584 ( .A1(n8700), .A2(n13072), .ZN(n12592) );
  NAND2_X1 U10585 ( .A1(n8700), .A2(n13072), .ZN(n12588) );
  NAND2_X1 U10586 ( .A1(n12592), .A2(n12588), .ZN(n12442) );
  XNOR2_X1 U10587 ( .A(n14101), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8213) );
  XNOR2_X1 U10588 ( .A(n8214), .B(n8213), .ZN(n12379) );
  NAND2_X1 U10589 ( .A1(n12379), .A2(n12417), .ZN(n8216) );
  NOR2_X1 U10590 ( .A1(n8617), .A2(n8217), .ZN(n8218) );
  INV_X1 U10591 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13374) );
  NAND2_X1 U10592 ( .A1(n8224), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10593 ( .A1(n8639), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8219) );
  OAI211_X1 U10594 ( .C1(n13374), .C2(n8245), .A(n8220), .B(n8219), .ZN(n8221)
         );
  INV_X1 U10595 ( .A(n13091), .ZN(n10956) );
  INV_X1 U10596 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8222) );
  INV_X1 U10597 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8223) );
  OR2_X1 U10598 ( .A1(n8254), .A2(n8223), .ZN(n8227) );
  INV_X1 U10599 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15619) );
  NAND2_X1 U10600 ( .A1(n8224), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8225) );
  OR2_X1 U10601 ( .A1(n8262), .A2(n10117), .ZN(n8233) );
  XNOR2_X1 U10602 ( .A(n8229), .B(n8240), .ZN(n10118) );
  OR2_X1 U10603 ( .A1(n8261), .A2(n10118), .ZN(n8232) );
  OR2_X1 U10604 ( .A1(n10681), .A2(n10747), .ZN(n8231) );
  NAND2_X1 U10605 ( .A1(n15587), .A2(n15606), .ZN(n12450) );
  NAND2_X1 U10606 ( .A1(n8639), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8238) );
  INV_X1 U10607 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10700) );
  OR2_X1 U10608 ( .A1(n8516), .A2(n10700), .ZN(n8237) );
  INV_X1 U10609 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11184) );
  OR2_X1 U10610 ( .A1(n8243), .A2(n11184), .ZN(n8236) );
  INV_X1 U10611 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8234) );
  INV_X1 U10612 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U10613 ( .A1(n10571), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8239) );
  AND2_X1 U10614 ( .A1(n8240), .A2(n8239), .ZN(n8242) );
  OAI21_X1 U10615 ( .B1(n6672), .B2(n8242), .A(n8241), .ZN(n13442) );
  MUX2_X1 U10616 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13442), .S(n10681), .Z(n10447) );
  INV_X1 U10617 ( .A(n15606), .ZN(n8725) );
  OR2_X1 U10618 ( .A1(n15587), .A2(n8725), .ZN(n15592) );
  NAND2_X1 U10619 ( .A1(n15591), .A2(n15592), .ZN(n8252) );
  INV_X1 U10620 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10750) );
  INV_X1 U10621 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15586) );
  OR2_X1 U10622 ( .A1(n8243), .A2(n15586), .ZN(n8247) );
  INV_X1 U10623 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U10624 ( .A(n8249), .B(n8248), .ZN(n10081) );
  OR2_X1 U10625 ( .A1(n8262), .A2(SI_2_), .ZN(n8250) );
  OAI211_X1 U10626 ( .C1(n10779), .C2(n10681), .A(n8251), .B(n8250), .ZN(
        n15582) );
  NAND2_X1 U10627 ( .A1(n15608), .A2(n15582), .ZN(n12458) );
  INV_X1 U10628 ( .A(n15608), .ZN(n10673) );
  NAND2_X1 U10629 ( .A1(n10673), .A2(n15582), .ZN(n8253) );
  INV_X1 U10630 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11306) );
  OR2_X1 U10631 ( .A1(n8254), .A2(n11306), .ZN(n8256) );
  INV_X1 U10632 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U10633 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6732), .ZN(n8258) );
  XNOR2_X1 U10634 ( .A(n8258), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10805) );
  XNOR2_X1 U10635 ( .A(n8260), .B(n8259), .ZN(n10075) );
  OR2_X1 U10636 ( .A1(n8261), .A2(n10075), .ZN(n8264) );
  OR2_X1 U10637 ( .A1(n8262), .A2(SI_3_), .ZN(n8263) );
  OAI211_X1 U10638 ( .C1(n10805), .C2(n10681), .A(n8264), .B(n8263), .ZN(
        n11308) );
  NAND2_X1 U10639 ( .A1(n10557), .A2(n11308), .ZN(n12465) );
  INV_X1 U10640 ( .A(n11308), .ZN(n8265) );
  NAND2_X1 U10641 ( .A1(n10557), .A2(n8265), .ZN(n8266) );
  NAND2_X1 U10642 ( .A1(n8537), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8270) );
  OR2_X1 U10643 ( .A1(n8516), .A2(n15676), .ZN(n8269) );
  AND2_X1 U10644 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8267) );
  NOR2_X1 U10645 ( .A1(n8278), .A2(n8267), .ZN(n10852) );
  INV_X1 U10646 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10647 ( .A1(n8271), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8272) );
  XNOR2_X1 U10648 ( .A(n8272), .B(n8190), .ZN(n11120) );
  INV_X1 U10649 ( .A(n11120), .ZN(n11141) );
  XNOR2_X1 U10650 ( .A(n8274), .B(n8273), .ZN(n10072) );
  OR2_X1 U10651 ( .A1(n8262), .A2(SI_4_), .ZN(n8275) );
  OAI211_X1 U10652 ( .C1(n11141), .C2(n10681), .A(n8276), .B(n8275), .ZN(
        n15574) );
  NAND2_X1 U10653 ( .A1(n11301), .A2(n15574), .ZN(n12469) );
  INV_X1 U10654 ( .A(n15574), .ZN(n8734) );
  NAND2_X1 U10655 ( .A1(n8537), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8283) );
  INV_X1 U10656 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15678) );
  OR2_X1 U10657 ( .A1(n8516), .A2(n15678), .ZN(n8282) );
  OR2_X1 U10658 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  AND2_X1 U10659 ( .A1(n8292), .A2(n8279), .ZN(n11084) );
  OR2_X1 U10660 ( .A1(n8243), .A2(n11084), .ZN(n8281) );
  INV_X1 U10661 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15564) );
  OR2_X1 U10662 ( .A1(n10876), .A2(n15564), .ZN(n8280) );
  NAND4_X1 U10663 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n11505) );
  NOR2_X1 U10664 ( .A1(n8361), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8311) );
  INV_X1 U10665 ( .A(n8311), .ZN(n8287) );
  NAND2_X1 U10666 ( .A1(n8361), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8285) );
  MUX2_X1 U10667 ( .A(n8285), .B(P3_IR_REG_31__SCAN_IN), .S(n8284), .Z(n8286)
         );
  NAND2_X1 U10668 ( .A1(n8287), .A2(n8286), .ZN(n15438) );
  OR2_X1 U10669 ( .A1(n12415), .A2(SI_5_), .ZN(n8289) );
  OAI211_X1 U10670 ( .C1(n7476), .C2(n10681), .A(n8290), .B(n8289), .ZN(n15561) );
  OR2_X1 U10671 ( .A1(n11505), .A2(n15561), .ZN(n12447) );
  NAND2_X1 U10672 ( .A1(n11505), .A2(n15561), .ZN(n12474) );
  NAND2_X1 U10673 ( .A1(n12447), .A2(n12474), .ZN(n15553) );
  INV_X1 U10674 ( .A(n15553), .ZN(n12472) );
  INV_X1 U10675 ( .A(n11505), .ZN(n15570) );
  NAND2_X1 U10676 ( .A1(n15570), .A2(n15561), .ZN(n8291) );
  NAND2_X1 U10677 ( .A1(n8537), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8297) );
  INV_X1 U10678 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11145) );
  OR2_X1 U10679 ( .A1(n8516), .A2(n11145), .ZN(n8296) );
  INV_X1 U10680 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11146) );
  OR2_X1 U10681 ( .A1(n10876), .A2(n11146), .ZN(n8295) );
  NAND2_X1 U10682 ( .A1(n8292), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8293) );
  AND2_X1 U10683 ( .A1(n8305), .A2(n8293), .ZN(n11502) );
  OR2_X1 U10684 ( .A1(n8243), .A2(n11502), .ZN(n8294) );
  NAND4_X1 U10685 ( .A1(n8297), .A2(n8296), .A3(n8295), .A4(n8294), .ZN(n11451) );
  INV_X1 U10686 ( .A(SI_6_), .ZN(n10119) );
  OR2_X1 U10687 ( .A1(n8262), .A2(n10119), .ZN(n8303) );
  XNOR2_X1 U10688 ( .A(n10132), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8298) );
  XNOR2_X1 U10689 ( .A(n8299), .B(n8298), .ZN(n10120) );
  OR2_X1 U10690 ( .A1(n8311), .A2(n8478), .ZN(n8300) );
  XNOR2_X1 U10691 ( .A(n8300), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11147) );
  OR2_X1 U10692 ( .A1(n10681), .A2(n15458), .ZN(n8301) );
  NAND2_X1 U10693 ( .A1(n11451), .A2(n11318), .ZN(n12479) );
  NAND2_X1 U10694 ( .A1(n12483), .A2(n12479), .ZN(n12429) );
  INV_X1 U10695 ( .A(n11318), .ZN(n11501) );
  NAND2_X1 U10696 ( .A1(n11451), .A2(n11501), .ZN(n8304) );
  NAND2_X1 U10697 ( .A1(n8537), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8310) );
  INV_X1 U10698 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11151) );
  OR2_X1 U10699 ( .A1(n8516), .A2(n11151), .ZN(n8309) );
  AND2_X1 U10700 ( .A1(n8305), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8306) );
  NOR2_X1 U10701 ( .A1(n8322), .A2(n8306), .ZN(n15547) );
  OR2_X1 U10702 ( .A1(n8243), .A2(n15547), .ZN(n8308) );
  INV_X1 U10703 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11152) );
  OR2_X1 U10704 ( .A1(n10876), .A2(n11152), .ZN(n8307) );
  NAND4_X1 U10705 ( .A1(n8310), .A2(n8309), .A3(n8308), .A4(n8307), .ZN(n12951) );
  NAND2_X1 U10706 ( .A1(n8311), .A2(n8359), .ZN(n8328) );
  NAND2_X1 U10707 ( .A1(n8328), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8313) );
  XNOR2_X1 U10708 ( .A(n8313), .B(n8312), .ZN(n15475) );
  INV_X1 U10709 ( .A(n15475), .ZN(n11153) );
  NAND2_X1 U10710 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  AND2_X1 U10711 ( .A1(n8317), .A2(n8316), .ZN(n10085) );
  OR2_X1 U10712 ( .A1(n12415), .A2(SI_7_), .ZN(n8318) );
  OAI211_X1 U10713 ( .C1(n11153), .C2(n10681), .A(n8319), .B(n8318), .ZN(
        n15546) );
  OR2_X1 U10714 ( .A1(n12951), .A2(n15546), .ZN(n12485) );
  NAND2_X1 U10715 ( .A1(n12951), .A2(n15546), .ZN(n12486) );
  INV_X1 U10716 ( .A(n15546), .ZN(n8320) );
  NAND2_X1 U10717 ( .A1(n12951), .A2(n8320), .ZN(n8321) );
  NAND2_X1 U10718 ( .A1(n8537), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8327) );
  INV_X1 U10719 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11159) );
  OR2_X1 U10720 ( .A1(n10876), .A2(n11159), .ZN(n8326) );
  INV_X1 U10721 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11158) );
  OR2_X1 U10722 ( .A1(n8516), .A2(n11158), .ZN(n8325) );
  NOR2_X1 U10723 ( .A1(n8322), .A2(n12823), .ZN(n8323) );
  OR2_X1 U10724 ( .A1(n8336), .A2(n8323), .ZN(n12825) );
  INV_X1 U10725 ( .A(n12825), .ZN(n11761) );
  OR2_X1 U10726 ( .A1(n8243), .A2(n11761), .ZN(n8324) );
  NAND4_X1 U10727 ( .A1(n8327), .A2(n8326), .A3(n8325), .A4(n8324), .ZN(n12491) );
  NAND2_X1 U10728 ( .A1(n8343), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8329) );
  XNOR2_X1 U10729 ( .A(n8329), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11160) );
  INV_X1 U10730 ( .A(SI_8_), .ZN(n10121) );
  OR2_X1 U10731 ( .A1(n8262), .A2(n10121), .ZN(n8333) );
  XNOR2_X1 U10732 ( .A(n8331), .B(n8330), .ZN(n10122) );
  OAI211_X1 U10733 ( .C1(n10681), .C2(n15493), .A(n8333), .B(n8332), .ZN(
        n12824) );
  XNOR2_X1 U10734 ( .A(n12491), .B(n12824), .ZN(n12488) );
  NAND2_X1 U10735 ( .A1(n8537), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8341) );
  INV_X1 U10736 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11165) );
  OR2_X1 U10737 ( .A1(n10876), .A2(n11165), .ZN(n8340) );
  INV_X1 U10738 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11164) );
  OR2_X1 U10739 ( .A1(n8516), .A2(n11164), .ZN(n8339) );
  OR2_X1 U10740 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  AND2_X1 U10741 ( .A1(n8351), .A2(n8337), .ZN(n11327) );
  OR2_X1 U10742 ( .A1(n8243), .A2(n11327), .ZN(n8338) );
  NAND4_X1 U10743 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), .ZN(n15528) );
  OAI21_X1 U10744 ( .B1(n8343), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8344) );
  XNOR2_X1 U10745 ( .A(n8342), .B(n8344), .ZN(n15512) );
  OR2_X1 U10746 ( .A1(n12415), .A2(SI_9_), .ZN(n8350) );
  OR2_X1 U10747 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  OAI211_X1 U10748 ( .C1(n11166), .C2(n10681), .A(n8350), .B(n8349), .ZN(
        n11651) );
  OR2_X1 U10749 ( .A1(n15528), .A2(n11651), .ZN(n12497) );
  NAND2_X1 U10750 ( .A1(n15528), .A2(n11651), .ZN(n12498) );
  NAND2_X1 U10751 ( .A1(n12497), .A2(n12498), .ZN(n12430) );
  OR2_X1 U10752 ( .A1(n12491), .A2(n12824), .ZN(n11645) );
  AND2_X1 U10753 ( .A1(n12430), .A2(n11645), .ZN(n11646) );
  NAND2_X1 U10754 ( .A1(n8537), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8357) );
  INV_X1 U10755 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11171) );
  OR2_X1 U10756 ( .A1(n8516), .A2(n11171), .ZN(n8356) );
  NAND2_X1 U10757 ( .A1(n8351), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10758 ( .A1(n8376), .A2(n8352), .ZN(n15531) );
  INV_X1 U10759 ( .A(n15531), .ZN(n8353) );
  OR2_X1 U10760 ( .A1(n8243), .A2(n8353), .ZN(n8355) );
  INV_X1 U10761 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11172) );
  OR2_X1 U10762 ( .A1(n10876), .A2(n11172), .ZN(n8354) );
  NAND4_X1 U10763 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n11807) );
  NAND3_X1 U10764 ( .A1(n8358), .A2(n8359), .A3(n8342), .ZN(n8360) );
  NAND2_X1 U10765 ( .A1(n8384), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U10766 ( .A(n8363), .B(n8362), .ZN(n11374) );
  INV_X1 U10767 ( .A(n11374), .ZN(n11381) );
  OR2_X1 U10768 ( .A1(n12415), .A2(SI_10_), .ZN(n8368) );
  OR2_X1 U10769 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  AND2_X1 U10770 ( .A1(n8367), .A2(n8366), .ZN(n10112) );
  OAI211_X1 U10771 ( .C1(n11381), .C2(n10681), .A(n8368), .B(n6797), .ZN(
        n15534) );
  OR2_X1 U10772 ( .A1(n11807), .A2(n15534), .ZN(n12502) );
  NAND2_X1 U10773 ( .A1(n11807), .A2(n15534), .ZN(n12501) );
  NAND2_X1 U10774 ( .A1(n12502), .A2(n12501), .ZN(n15532) );
  INV_X1 U10775 ( .A(n15532), .ZN(n8370) );
  INV_X1 U10776 ( .A(n11651), .ZN(n8369) );
  NAND2_X1 U10777 ( .A1(n15528), .A2(n8369), .ZN(n15525) );
  INV_X1 U10778 ( .A(n15534), .ZN(n8371) );
  NAND2_X1 U10779 ( .A1(n11807), .A2(n8371), .ZN(n8372) );
  NAND2_X1 U10780 ( .A1(n8537), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8381) );
  INV_X1 U10781 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8374) );
  OR2_X1 U10782 ( .A1(n10876), .A2(n8374), .ZN(n8380) );
  INV_X1 U10783 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8375) );
  OR2_X1 U10784 ( .A1(n8516), .A2(n8375), .ZN(n8379) );
  NAND2_X1 U10785 ( .A1(n8376), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8377) );
  AND2_X1 U10786 ( .A1(n8390), .A2(n8377), .ZN(n11806) );
  OR2_X1 U10787 ( .A1(n8243), .A2(n11806), .ZN(n8378) );
  NAND4_X1 U10788 ( .A1(n8381), .A2(n8380), .A3(n8379), .A4(n8378), .ZN(n15529) );
  XNOR2_X1 U10789 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8382) );
  XNOR2_X1 U10790 ( .A(n8383), .B(n8382), .ZN(n10115) );
  NAND2_X1 U10791 ( .A1(n10115), .A2(n12417), .ZN(n8387) );
  NOR2_X1 U10792 ( .A1(n8399), .A2(n8478), .ZN(n8385) );
  XNOR2_X1 U10793 ( .A(n8385), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U10794 ( .A1(n8510), .A2(n10116), .B1(n8509), .B2(n11564), .ZN(
        n8386) );
  NAND2_X1 U10795 ( .A1(n8537), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8395) );
  INV_X1 U10796 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n8388) );
  OR2_X1 U10797 ( .A1(n10876), .A2(n8388), .ZN(n8394) );
  INV_X1 U10798 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8389) );
  OR2_X1 U10799 ( .A1(n8516), .A2(n8389), .ZN(n8393) );
  AND2_X1 U10800 ( .A1(n8390), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8391) );
  NOR2_X1 U10801 ( .A1(n8418), .A2(n8391), .ZN(n11863) );
  OR2_X1 U10802 ( .A1(n8243), .A2(n11863), .ZN(n8392) );
  XNOR2_X1 U10803 ( .A(n8397), .B(n8396), .ZN(n10129) );
  NAND2_X1 U10804 ( .A1(n10129), .A2(n12417), .ZN(n8402) );
  INV_X1 U10805 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8398) );
  NOR2_X1 U10806 ( .A1(n8408), .A2(n8478), .ZN(n8400) );
  XNOR2_X1 U10807 ( .A(n8400), .B(n8407), .ZN(n11574) );
  AOI22_X1 U10808 ( .A1(n8510), .A2(SI_12_), .B1(n8509), .B2(n11574), .ZN(
        n8401) );
  NAND2_X1 U10809 ( .A1(n8402), .A2(n8401), .ZN(n14854) );
  NAND2_X1 U10810 ( .A1(n14863), .A2(n14854), .ZN(n12511) );
  INV_X1 U10811 ( .A(n14854), .ZN(n8403) );
  INV_X1 U10812 ( .A(n14863), .ZN(n11805) );
  NAND2_X1 U10813 ( .A1(n8403), .A2(n11805), .ZN(n12512) );
  NAND2_X1 U10814 ( .A1(n12511), .A2(n12512), .ZN(n14849) );
  INV_X1 U10815 ( .A(n15529), .ZN(n12508) );
  NAND2_X1 U10816 ( .A1(n12508), .A2(n14865), .ZN(n14846) );
  AND2_X1 U10817 ( .A1(n14849), .A2(n14846), .ZN(n8404) );
  NAND2_X1 U10818 ( .A1(n14854), .A2(n11805), .ZN(n8405) );
  XNOR2_X1 U10819 ( .A(n8406), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U10820 ( .A1(n10138), .A2(n12417), .ZN(n8415) );
  AND2_X1 U10821 ( .A1(n8408), .A2(n8407), .ZN(n8412) );
  INV_X1 U10822 ( .A(n8412), .ZN(n8409) );
  NAND2_X1 U10823 ( .A1(n8409), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8410) );
  INV_X1 U10824 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8411) );
  MUX2_X1 U10825 ( .A(n8410), .B(P3_IR_REG_31__SCAN_IN), .S(n8411), .Z(n8413)
         );
  NAND2_X1 U10826 ( .A1(n8412), .A2(n8411), .ZN(n8445) );
  NAND2_X1 U10827 ( .A1(n8413), .A2(n8445), .ZN(n12958) );
  AOI22_X1 U10828 ( .A1(n8510), .A2(n10139), .B1(n8509), .B2(n12958), .ZN(
        n8414) );
  NAND2_X1 U10829 ( .A1(n8537), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8423) );
  INV_X1 U10830 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13291) );
  OR2_X1 U10831 ( .A1(n10876), .A2(n13291), .ZN(n8422) );
  INV_X1 U10832 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8416) );
  OR2_X1 U10833 ( .A1(n8516), .A2(n8416), .ZN(n8421) );
  OR2_X1 U10834 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  AND2_X1 U10835 ( .A1(n8419), .A2(n8432), .ZN(n13290) );
  OR2_X1 U10836 ( .A1(n8243), .A2(n13290), .ZN(n8420) );
  NAND2_X1 U10837 ( .A1(n13422), .A2(n13274), .ZN(n8424) );
  NAND2_X1 U10838 ( .A1(n13284), .A2(n8424), .ZN(n13271) );
  OR2_X1 U10839 ( .A1(n13422), .A2(n13274), .ZN(n13270) );
  XNOR2_X1 U10840 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8425) );
  XNOR2_X1 U10841 ( .A(n8426), .B(n8425), .ZN(n10147) );
  NAND2_X1 U10842 ( .A1(n10147), .A2(n12417), .ZN(n8430) );
  NAND2_X1 U10843 ( .A1(n8445), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8427) );
  XNOR2_X1 U10844 ( .A(n8428), .B(n8427), .ZN(n12976) );
  AOI22_X1 U10845 ( .A1(n8510), .A2(n10148), .B1(n8509), .B2(n12976), .ZN(
        n8429) );
  NAND2_X1 U10846 ( .A1(n8224), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8437) );
  INV_X1 U10847 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8431) );
  OR2_X1 U10848 ( .A1(n10876), .A2(n8431), .ZN(n8436) );
  NAND2_X1 U10849 ( .A1(n8432), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8433) );
  AND2_X1 U10850 ( .A1(n8450), .A2(n8433), .ZN(n12784) );
  OR2_X1 U10851 ( .A1(n8243), .A2(n12784), .ZN(n8435) );
  INV_X1 U10852 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13416) );
  OR2_X1 U10853 ( .A1(n8245), .A2(n13416), .ZN(n8434) );
  NAND4_X1 U10854 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n12894) );
  OR2_X1 U10855 ( .A1(n13418), .A2(n13286), .ZN(n8438) );
  AND2_X1 U10856 ( .A1(n13270), .A2(n8438), .ZN(n8440) );
  INV_X1 U10857 ( .A(n8438), .ZN(n8439) );
  NAND2_X1 U10858 ( .A1(n13418), .A2(n12894), .ZN(n12525) );
  NAND2_X1 U10859 ( .A1(n12522), .A2(n12525), .ZN(n13276) );
  NAND2_X1 U10860 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  NAND2_X1 U10861 ( .A1(n8444), .A2(n8443), .ZN(n10160) );
  OAI21_X1 U10862 ( .B1(n8445), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8447) );
  INV_X1 U10863 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8446) );
  XNOR2_X1 U10864 ( .A(n8447), .B(n8446), .ZN(n13007) );
  INV_X1 U10865 ( .A(n13007), .ZN(n13020) );
  AOI22_X1 U10866 ( .A1(n8510), .A2(SI_15_), .B1(n8509), .B2(n13020), .ZN(
        n8448) );
  NAND2_X1 U10867 ( .A1(n8449), .A2(n8448), .ZN(n13264) );
  NAND2_X1 U10868 ( .A1(n8224), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8455) );
  INV_X1 U10869 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12983) );
  OR2_X1 U10870 ( .A1(n10876), .A2(n12983), .ZN(n8454) );
  AND2_X1 U10871 ( .A1(n8450), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8451) );
  NOR2_X1 U10872 ( .A1(n8465), .A2(n8451), .ZN(n12937) );
  OR2_X1 U10873 ( .A1(n8243), .A2(n12937), .ZN(n8453) );
  INV_X1 U10874 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13412) );
  OR2_X1 U10875 ( .A1(n8245), .A2(n13412), .ZN(n8452) );
  OR2_X1 U10876 ( .A1(n13264), .A2(n13275), .ZN(n12524) );
  NAND2_X1 U10877 ( .A1(n13264), .A2(n13275), .ZN(n12530) );
  NAND2_X1 U10878 ( .A1(n12524), .A2(n12530), .ZN(n13258) );
  NAND2_X1 U10879 ( .A1(n13264), .A2(n12949), .ZN(n8456) );
  OR2_X1 U10880 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  NAND2_X1 U10881 ( .A1(n8460), .A2(n8459), .ZN(n10170) );
  OR2_X1 U10882 ( .A1(n8461), .A2(n8478), .ZN(n8462) );
  XNOR2_X1 U10883 ( .A(n8462), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U10884 ( .A1(n8510), .A2(SI_16_), .B1(n8509), .B2(n13045), .ZN(
        n8463) );
  NAND2_X1 U10885 ( .A1(n8464), .A2(n8463), .ZN(n12849) );
  NAND2_X1 U10886 ( .A1(n8537), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8471) );
  INV_X1 U10887 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13351) );
  OR2_X1 U10888 ( .A1(n8516), .A2(n13351), .ZN(n8470) );
  INV_X1 U10889 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13022) );
  OR2_X1 U10890 ( .A1(n10876), .A2(n13022), .ZN(n8469) );
  NOR2_X1 U10891 ( .A1(n8465), .A2(n9042), .ZN(n8466) );
  OR2_X1 U10892 ( .A1(n8484), .A2(n8466), .ZN(n13252) );
  INV_X1 U10893 ( .A(n13252), .ZN(n8467) );
  OR2_X1 U10894 ( .A1(n8243), .A2(n8467), .ZN(n8468) );
  OR2_X1 U10895 ( .A1(n12849), .A2(n13260), .ZN(n12532) );
  NAND2_X1 U10896 ( .A1(n12849), .A2(n13260), .ZN(n12531) );
  NAND2_X1 U10897 ( .A1(n12532), .A2(n12531), .ZN(n13247) );
  INV_X1 U10898 ( .A(n13260), .ZN(n12948) );
  OR2_X1 U10899 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  NAND2_X1 U10900 ( .A1(n8475), .A2(n8474), .ZN(n10184) );
  NOR2_X1 U10901 ( .A1(n8476), .A2(n8478), .ZN(n8477) );
  MUX2_X1 U10902 ( .A(n8478), .B(n8477), .S(P3_IR_REG_17__SCAN_IN), .Z(n8481)
         );
  INV_X1 U10903 ( .A(n8479), .ZN(n8480) );
  INV_X1 U10904 ( .A(n13046), .ZN(n14811) );
  AOI22_X1 U10905 ( .A1(n8510), .A2(SI_17_), .B1(n8509), .B2(n14811), .ZN(
        n8482) );
  OR2_X1 U10906 ( .A1(n8484), .A2(n12861), .ZN(n8485) );
  NAND2_X1 U10907 ( .A1(n8496), .A2(n8485), .ZN(n13241) );
  NAND2_X1 U10908 ( .A1(n8619), .A2(n13241), .ZN(n8489) );
  INV_X1 U10909 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13347) );
  OR2_X1 U10910 ( .A1(n8516), .A2(n13347), .ZN(n8488) );
  INV_X1 U10911 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14820) );
  OR2_X1 U10912 ( .A1(n10876), .A2(n14820), .ZN(n8487) );
  INV_X1 U10913 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13404) );
  OR2_X1 U10914 ( .A1(n8245), .A2(n13404), .ZN(n8486) );
  OR2_X1 U10915 ( .A1(n13240), .A2(n13249), .ZN(n12540) );
  NAND2_X1 U10916 ( .A1(n13240), .A2(n13249), .ZN(n12535) );
  NAND2_X1 U10917 ( .A1(n12540), .A2(n12535), .ZN(n13234) );
  INV_X1 U10918 ( .A(n13249), .ZN(n12915) );
  NAND2_X1 U10919 ( .A1(n13240), .A2(n12915), .ZN(n8490) );
  XNOR2_X1 U10920 ( .A(n8492), .B(n8491), .ZN(n10273) );
  NAND2_X1 U10921 ( .A1(n10273), .A2(n12417), .ZN(n8495) );
  NAND2_X1 U10922 ( .A1(n8479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10923 ( .A(n8493), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14826) );
  AOI22_X1 U10924 ( .A1(n8510), .A2(SI_18_), .B1(n8509), .B2(n14826), .ZN(
        n8494) );
  NAND2_X1 U10925 ( .A1(n8496), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U10926 ( .A1(n8513), .A2(n8497), .ZN(n13223) );
  NAND2_X1 U10927 ( .A1(n8619), .A2(n13223), .ZN(n8501) );
  INV_X1 U10928 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13343) );
  OR2_X1 U10929 ( .A1(n8516), .A2(n13343), .ZN(n8500) );
  INV_X1 U10930 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13225) );
  OR2_X1 U10931 ( .A1(n10876), .A2(n13225), .ZN(n8499) );
  INV_X1 U10932 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13400) );
  OR2_X1 U10933 ( .A1(n8245), .A2(n13400), .ZN(n8498) );
  NAND2_X1 U10934 ( .A1(n13228), .A2(n13236), .ZN(n12538) );
  INV_X1 U10935 ( .A(n13236), .ZN(n13203) );
  OR2_X1 U10936 ( .A1(n13228), .A2(n13203), .ZN(n8503) );
  OR2_X1 U10937 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  NAND2_X1 U10938 ( .A1(n8507), .A2(n8506), .ZN(n10309) );
  NAND2_X1 U10939 ( .A1(n8627), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8508) );
  XNOR2_X2 U10940 ( .A(n8508), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U10941 ( .A1(n8510), .A2(SI_19_), .B1(n13039), .B2(n8509), .ZN(
        n8511) );
  NAND2_X1 U10942 ( .A1(n8512), .A2(n8511), .ZN(n12798) );
  AND2_X1 U10943 ( .A1(n8513), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8514) );
  OR2_X1 U10944 ( .A1(n8514), .A2(n8526), .ZN(n13209) );
  NAND2_X1 U10945 ( .A1(n13209), .A2(n8619), .ZN(n8521) );
  INV_X1 U10946 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n8515) );
  OR2_X1 U10947 ( .A1(n10876), .A2(n8515), .ZN(n8518) );
  INV_X1 U10948 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13339) );
  OR2_X1 U10949 ( .A1(n8516), .A2(n13339), .ZN(n8517) );
  AND2_X1 U10950 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  NAND2_X1 U10951 ( .A1(n8537), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8519) );
  OR2_X1 U10952 ( .A1(n12798), .A2(n13222), .ZN(n12547) );
  NAND2_X1 U10953 ( .A1(n12798), .A2(n13222), .ZN(n12548) );
  NAND2_X1 U10954 ( .A1(n12798), .A2(n13187), .ZN(n8522) );
  INV_X1 U10955 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12062) );
  XNOR2_X1 U10956 ( .A(n8523), .B(n12062), .ZN(n10563) );
  NAND2_X1 U10957 ( .A1(n10563), .A2(n12417), .ZN(n8525) );
  OR2_X1 U10958 ( .A1(n12415), .A2(n10564), .ZN(n8524) );
  NOR2_X1 U10959 ( .A1(n8526), .A2(n9174), .ZN(n8527) );
  OR2_X1 U10960 ( .A1(n8535), .A2(n8527), .ZN(n13194) );
  NAND2_X1 U10961 ( .A1(n13194), .A2(n8619), .ZN(n8530) );
  AOI22_X1 U10962 ( .A1(n8639), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n8224), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U10963 ( .A1(n8537), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8528) );
  XNOR2_X1 U10964 ( .A(n13332), .B(n13175), .ZN(n13190) );
  XNOR2_X1 U10965 ( .A(n8532), .B(n8531), .ZN(n10810) );
  NAND2_X1 U10966 ( .A1(n10810), .A2(n12417), .ZN(n8534) );
  INV_X1 U10967 ( .A(SI_21_), .ZN(n10811) );
  OR2_X1 U10968 ( .A1(n8535), .A2(n12834), .ZN(n8536) );
  NAND2_X1 U10969 ( .A1(n8549), .A2(n8536), .ZN(n13180) );
  NAND2_X1 U10970 ( .A1(n13180), .A2(n8619), .ZN(n8540) );
  AOI22_X1 U10971 ( .A1(n8639), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n8224), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10972 ( .A1(n8537), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10973 ( .A1(n13179), .A2(n13162), .ZN(n12556) );
  INV_X1 U10974 ( .A(n13162), .ZN(n13188) );
  OR2_X1 U10975 ( .A1(n13179), .A2(n13188), .ZN(n8543) );
  XNOR2_X1 U10976 ( .A(n8545), .B(n8544), .ZN(n10862) );
  NAND2_X1 U10977 ( .A1(n10862), .A2(n12417), .ZN(n8548) );
  NAND2_X1 U10978 ( .A1(n8549), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10979 ( .A1(n8562), .A2(n8550), .ZN(n13166) );
  NAND2_X1 U10980 ( .A1(n13166), .A2(n8619), .ZN(n8555) );
  INV_X1 U10981 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U10982 ( .A1(n8639), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10983 ( .A1(n8224), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8551) );
  OAI211_X1 U10984 ( .C1(n13387), .C2(n8245), .A(n8552), .B(n8551), .ZN(n8553)
         );
  INV_X1 U10985 ( .A(n8553), .ZN(n8554) );
  NAND2_X1 U10986 ( .A1(n13165), .A2(n12904), .ZN(n8556) );
  OR2_X1 U10987 ( .A1(n13165), .A2(n12904), .ZN(n8557) );
  XNOR2_X1 U10988 ( .A(n8559), .B(n8558), .ZN(n11052) );
  NAND2_X1 U10989 ( .A1(n11052), .A2(n12417), .ZN(n8561) );
  NAND2_X2 U10990 ( .A1(n8561), .A2(n8560), .ZN(n13319) );
  XNOR2_X1 U10991 ( .A(n8562), .B(P3_REG3_REG_23__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U10992 ( .A1(n13152), .A2(n8619), .ZN(n8568) );
  INV_X1 U10993 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10994 ( .A1(n8639), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U10995 ( .A1(n8224), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8563) );
  OAI211_X1 U10996 ( .C1(n8565), .C2(n8245), .A(n8564), .B(n8563), .ZN(n8566)
         );
  INV_X1 U10997 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U10998 ( .A1(n13319), .A2(n13161), .ZN(n12562) );
  NAND2_X1 U10999 ( .A1(n13319), .A2(n12873), .ZN(n8571) );
  OR2_X1 U11000 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  NAND2_X1 U11001 ( .A1(n8589), .A2(n8574), .ZN(n13137) );
  NAND2_X1 U11002 ( .A1(n13137), .A2(n8619), .ZN(n8580) );
  INV_X1 U11003 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11004 ( .A1(n8639), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U11005 ( .A1(n8224), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8575) );
  OAI211_X1 U11006 ( .C1(n8577), .C2(n8245), .A(n8576), .B(n8575), .ZN(n8578)
         );
  INV_X1 U11007 ( .A(n8578), .ZN(n8579) );
  INV_X1 U11008 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12375) );
  XNOR2_X1 U11009 ( .A(n8581), .B(n12375), .ZN(n11442) );
  NAND2_X1 U11010 ( .A1(n11442), .A2(n12417), .ZN(n8583) );
  INV_X1 U11011 ( .A(SI_24_), .ZN(n11443) );
  OR2_X1 U11012 ( .A1(n13145), .A2(n13314), .ZN(n12567) );
  NAND2_X1 U11013 ( .A1(n13314), .A2(n13145), .ZN(n12569) );
  NAND2_X1 U11014 ( .A1(n12567), .A2(n12569), .ZN(n13132) );
  NAND2_X1 U11015 ( .A1(n13314), .A2(n13115), .ZN(n8584) );
  XNOR2_X1 U11016 ( .A(n14112), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U11017 ( .A(n8586), .B(n8585), .ZN(n11595) );
  NAND2_X1 U11018 ( .A1(n11595), .A2(n12417), .ZN(n8588) );
  NAND2_X1 U11019 ( .A1(n8589), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U11020 ( .A1(n8601), .A2(n8590), .ZN(n13121) );
  NAND2_X1 U11021 ( .A1(n13121), .A2(n8619), .ZN(n8595) );
  INV_X1 U11022 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U11023 ( .A1(n8639), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11024 ( .A1(n8224), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8591) );
  OAI211_X1 U11025 ( .C1(n13381), .C2(n8245), .A(n8592), .B(n8591), .ZN(n8593)
         );
  INV_X1 U11026 ( .A(n8593), .ZN(n8594) );
  OR2_X1 U11027 ( .A1(n13120), .A2(n13130), .ZN(n12574) );
  NAND2_X1 U11028 ( .A1(n13120), .A2(n13130), .ZN(n12575) );
  NAND2_X1 U11029 ( .A1(n12574), .A2(n12575), .ZN(n13113) );
  NAND2_X1 U11030 ( .A1(n13120), .A2(n12874), .ZN(n8596) );
  XNOR2_X1 U11031 ( .A(n14107), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8597) );
  XNOR2_X1 U11032 ( .A(n8598), .B(n8597), .ZN(n11726) );
  NAND2_X1 U11033 ( .A1(n11726), .A2(n12417), .ZN(n8600) );
  NAND2_X1 U11034 ( .A1(n8601), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11035 ( .A1(n8616), .A2(n8602), .ZN(n13106) );
  NAND2_X1 U11036 ( .A1(n13106), .A2(n8619), .ZN(n8608) );
  INV_X1 U11037 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11038 ( .A1(n8224), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11039 ( .A1(n8639), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8603) );
  OAI211_X1 U11040 ( .C1(n8605), .C2(n8245), .A(n8604), .B(n8603), .ZN(n8606)
         );
  INV_X1 U11041 ( .A(n8606), .ZN(n8607) );
  OR2_X1 U11042 ( .A1(n13306), .A2(n13116), .ZN(n8609) );
  NAND2_X1 U11043 ( .A1(n13103), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U11044 ( .A1(n13306), .A2(n13116), .ZN(n8610) );
  XNOR2_X1 U11045 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8612) );
  XNOR2_X1 U11046 ( .A(n8613), .B(n8612), .ZN(n11800) );
  NAND2_X1 U11047 ( .A1(n11800), .A2(n12417), .ZN(n8615) );
  INV_X1 U11048 ( .A(SI_27_), .ZN(n11801) );
  AND2_X1 U11049 ( .A1(n8616), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11050 ( .A1(n13095), .A2(n8619), .ZN(n8624) );
  INV_X1 U11051 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U11052 ( .A1(n8639), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11053 ( .A1(n8224), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U11054 ( .C1(n13377), .C2(n8245), .A(n8621), .B(n8620), .ZN(n8622)
         );
  INV_X1 U11055 ( .A(n8622), .ZN(n8623) );
  OR2_X1 U11056 ( .A1(n8797), .A2(n12928), .ZN(n8625) );
  NAND2_X1 U11057 ( .A1(n13078), .A2(n13091), .ZN(n8660) );
  XOR2_X1 U11058 ( .A(n12442), .B(n8626), .Z(n8647) );
  NAND2_X1 U11059 ( .A1(n8668), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11060 ( .A1(n12606), .A2(n13039), .ZN(n8708) );
  NAND2_X1 U11061 ( .A1(n8633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U11062 ( .A1(n12449), .A2(n8707), .ZN(n12424) );
  INV_X1 U11063 ( .A(n12382), .ZN(n12603) );
  INV_X1 U11064 ( .A(n8636), .ZN(n10683) );
  NAND2_X1 U11065 ( .A1(n12603), .A2(n10683), .ZN(n10693) );
  NAND2_X1 U11066 ( .A1(n10681), .A2(n10693), .ZN(n8637) );
  AND2_X1 U11067 ( .A1(n12603), .A2(P3_B_REG_SCAN_IN), .ZN(n8638) );
  OR2_X1 U11068 ( .A1(n15588), .A2(n8638), .ZN(n13057) );
  INV_X1 U11069 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11070 ( .A1(n8639), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11071 ( .A1(n8224), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8640) );
  OAI211_X1 U11072 ( .C1(n8642), .C2(n8245), .A(n8641), .B(n8640), .ZN(n8643)
         );
  INV_X1 U11073 ( .A(n8643), .ZN(n8644) );
  AND2_X1 U11074 ( .A1(n10882), .A2(n8644), .ZN(n12418) );
  OAI22_X1 U11075 ( .A1(n13091), .A2(n15590), .B1(n13057), .B2(n12418), .ZN(
        n8645) );
  INV_X1 U11076 ( .A(n8645), .ZN(n8646) );
  OAI21_X1 U11077 ( .B1(n8647), .B2(n15594), .A(n8646), .ZN(n13063) );
  INV_X1 U11078 ( .A(n10447), .ZN(n10664) );
  INV_X1 U11079 ( .A(n11303), .ZN(n12427) );
  INV_X1 U11080 ( .A(n15568), .ZN(n15566) );
  NAND2_X1 U11081 ( .A1(n15567), .A2(n15566), .ZN(n8648) );
  NAND2_X1 U11082 ( .A1(n8648), .A2(n12470), .ZN(n15551) );
  INV_X1 U11083 ( .A(n12429), .ZN(n11499) );
  INV_X1 U11084 ( .A(n15540), .ZN(n15539) );
  NAND2_X1 U11085 ( .A1(n15538), .A2(n15539), .ZN(n8649) );
  NAND2_X1 U11086 ( .A1(n8649), .A2(n12485), .ZN(n11760) );
  NAND2_X1 U11087 ( .A1(n11760), .A2(n12488), .ZN(n8650) );
  INV_X1 U11088 ( .A(n12491), .ZN(n15542) );
  NAND2_X1 U11089 ( .A1(n15542), .A2(n12824), .ZN(n12492) );
  INV_X1 U11090 ( .A(n12497), .ZN(n8651) );
  INV_X1 U11091 ( .A(n12501), .ZN(n8652) );
  XNOR2_X1 U11092 ( .A(n15529), .B(n12507), .ZN(n14859) );
  OR2_X1 U11093 ( .A1(n15529), .A2(n14865), .ZN(n12506) );
  INV_X1 U11094 ( .A(n14849), .ZN(n14845) );
  NOR2_X1 U11095 ( .A1(n13422), .A2(n14851), .ZN(n12517) );
  INV_X1 U11096 ( .A(n12517), .ZN(n8653) );
  NAND2_X1 U11097 ( .A1(n13422), .A2(n14851), .ZN(n12425) );
  INV_X1 U11098 ( .A(n13276), .ZN(n8654) );
  NAND2_X1 U11099 ( .A1(n8655), .A2(n12522), .ZN(n13263) );
  INV_X1 U11100 ( .A(n13258), .ZN(n13262) );
  NAND2_X1 U11101 ( .A1(n13263), .A2(n13262), .ZN(n13261) );
  NAND2_X1 U11102 ( .A1(n13261), .A2(n12530), .ZN(n13251) );
  INV_X1 U11103 ( .A(n13247), .ZN(n13250) );
  NAND2_X1 U11104 ( .A1(n13251), .A2(n13250), .ZN(n8656) );
  INV_X1 U11105 ( .A(n13234), .ZN(n13238) );
  NAND2_X1 U11106 ( .A1(n13216), .A2(n12539), .ZN(n13207) );
  OR2_X1 U11107 ( .A1(n13332), .A2(n13175), .ZN(n12551) );
  NAND2_X1 U11108 ( .A1(n13165), .A2(n13176), .ZN(n12559) );
  NAND2_X1 U11109 ( .A1(n13164), .A2(n12559), .ZN(n8658) );
  NAND2_X1 U11110 ( .A1(n8658), .A2(n12560), .ZN(n13142) );
  INV_X1 U11111 ( .A(n12566), .ZN(n13127) );
  NOR2_X1 U11112 ( .A1(n13132), .A2(n13127), .ZN(n8659) );
  INV_X1 U11113 ( .A(n13113), .ZN(n12572) );
  NAND2_X1 U11114 ( .A1(n13306), .A2(n13090), .ZN(n12580) );
  INV_X1 U11115 ( .A(n12928), .ZN(n13101) );
  NAND2_X1 U11116 ( .A1(n8797), .A2(n13101), .ZN(n13075) );
  AND2_X1 U11117 ( .A1(n8660), .A2(n13075), .ZN(n12586) );
  INV_X1 U11118 ( .A(n8661), .ZN(n12585) );
  AOI21_X2 U11119 ( .B1(n13087), .B2(n12586), .A(n12585), .ZN(n12420) );
  XOR2_X1 U11120 ( .A(n12442), .B(n12420), .Z(n13068) );
  OAI21_X1 U11121 ( .B1(n10860), .B2(n8707), .A(n13039), .ZN(n8662) );
  NAND2_X1 U11122 ( .A1(n8662), .A2(n10813), .ZN(n8664) );
  OAI21_X1 U11123 ( .B1(n8707), .B2(n12449), .A(n10860), .ZN(n8663) );
  NAND2_X1 U11124 ( .A1(n8664), .A2(n8663), .ZN(n8802) );
  NAND2_X1 U11125 ( .A1(n8802), .A2(n15605), .ZN(n10443) );
  NAND2_X1 U11126 ( .A1(n10566), .A2(n13054), .ZN(n8696) );
  OR2_X1 U11127 ( .A1(n10443), .A2(n8696), .ZN(n8666) );
  AND2_X1 U11128 ( .A1(n8707), .A2(n13054), .ZN(n8665) );
  NAND2_X1 U11129 ( .A1(n12606), .A2(n8665), .ZN(n8695) );
  NOR2_X1 U11130 ( .A1(n13063), .A2(n8667), .ZN(n8721) );
  NAND2_X1 U11131 ( .A1(n6711), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8671) );
  MUX2_X1 U11132 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8671), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8673) );
  NAND2_X1 U11133 ( .A1(n8673), .A2(n8672), .ZN(n11598) );
  NAND2_X1 U11134 ( .A1(n8674), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8675) );
  MUX2_X1 U11135 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8675), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8676) );
  NAND2_X1 U11136 ( .A1(n8676), .A2(n6711), .ZN(n11445) );
  NOR2_X1 U11137 ( .A1(n11598), .A2(n11445), .ZN(n8678) );
  NAND2_X1 U11138 ( .A1(n8672), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11139 ( .A1(n8678), .A2(n8682), .ZN(n10070) );
  XNOR2_X1 U11140 ( .A(n11445), .B(P3_B_REG_SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11141 ( .A1(n8679), .A2(n11598), .ZN(n8680) );
  INV_X1 U11142 ( .A(n11445), .ZN(n8681) );
  INV_X1 U11143 ( .A(n8682), .ZN(n11729) );
  NAND2_X1 U11144 ( .A1(n11729), .A2(n11598), .ZN(n8683) );
  OR2_X1 U11145 ( .A1(n13425), .A2(n10652), .ZN(n8705) );
  NAND2_X1 U11146 ( .A1(n13425), .A2(n10652), .ZN(n8710) );
  NOR2_X1 U11147 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8687) );
  NOR4_X1 U11148 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8686) );
  NOR4_X1 U11149 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8685) );
  NOR4_X1 U11150 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8684) );
  NAND4_X1 U11151 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n8694)
         );
  NOR4_X1 U11152 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8691) );
  NOR4_X1 U11153 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8690) );
  NOR4_X1 U11154 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8689) );
  NOR4_X1 U11155 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8688) );
  NAND4_X1 U11156 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n8693)
         );
  INV_X1 U11157 ( .A(n10136), .ZN(n8692) );
  OAI21_X1 U11158 ( .B1(n8694), .B2(n8693), .A(n8692), .ZN(n8709) );
  INV_X1 U11159 ( .A(n8696), .ZN(n12599) );
  NAND2_X1 U11160 ( .A1(n12578), .A2(n8695), .ZN(n10651) );
  OAI22_X1 U11161 ( .A1(n15605), .A2(n8707), .B1(n13039), .B2(n10860), .ZN(
        n8697) );
  AOI21_X1 U11162 ( .B1(n8697), .B2(n8696), .A(n12587), .ZN(n8698) );
  MUX2_X1 U11163 ( .A(n10655), .B(n8698), .S(n10652), .Z(n8699) );
  INV_X1 U11164 ( .A(n8700), .ZN(n13066) );
  NOR2_X1 U11165 ( .A1(n15685), .A2(n8701), .ZN(n8702) );
  OAI21_X1 U11166 ( .B1(n8721), .B2(n8704), .A(n8703), .ZN(P3_U3488) );
  INV_X1 U11167 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U11168 ( .A1(n8706), .A2(n8709), .ZN(n8803) );
  OR2_X1 U11169 ( .A1(n8708), .A2(n12444), .ZN(n8804) );
  INV_X1 U11170 ( .A(n8709), .ZN(n8711) );
  INV_X1 U11171 ( .A(n8802), .ZN(n8712) );
  OAI22_X1 U11172 ( .A1(n8803), .A2(n8804), .B1(n8810), .B2(n8712), .ZN(n8713)
         );
  NAND2_X1 U11173 ( .A1(n8713), .A2(n10678), .ZN(n8716) );
  NAND2_X1 U11174 ( .A1(n10678), .A2(n12599), .ZN(n8800) );
  NOR2_X1 U11175 ( .A1(n8800), .A2(n12578), .ZN(n8811) );
  INV_X1 U11176 ( .A(n8803), .ZN(n8714) );
  NAND2_X1 U11177 ( .A1(n8811), .A2(n8714), .ZN(n8715) );
  INV_X1 U11178 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8717) );
  OAI21_X1 U11179 ( .B1(n8721), .B2(n15672), .A(n8720), .ZN(P3_U3456) );
  NAND2_X1 U11180 ( .A1(n10813), .A2(n13039), .ZN(n8722) );
  NAND2_X1 U11181 ( .A1(n8722), .A2(n10566), .ZN(n8723) );
  XNOR2_X1 U11182 ( .A(n8797), .B(n7688), .ZN(n12810) );
  NOR2_X1 U11183 ( .A1(n12810), .A2(n12928), .ZN(n12806) );
  AOI21_X1 U11184 ( .B1(n12810), .B2(n12928), .A(n12806), .ZN(n8794) );
  XNOR2_X1 U11185 ( .A(n13165), .B(n8787), .ZN(n8779) );
  XNOR2_X1 U11186 ( .A(n13240), .B(n8787), .ZN(n8761) );
  INV_X1 U11187 ( .A(n8761), .ZN(n8763) );
  NAND3_X1 U11188 ( .A1(n15587), .A2(n7688), .A3(n8725), .ZN(n8726) );
  XNOR2_X1 U11189 ( .A(n15582), .B(n8728), .ZN(n8729) );
  XNOR2_X1 U11190 ( .A(n10673), .B(n8729), .ZN(n10556) );
  XNOR2_X1 U11191 ( .A(n11308), .B(n7688), .ZN(n8732) );
  XNOR2_X1 U11192 ( .A(n8732), .B(n10557), .ZN(n10671) );
  INV_X1 U11193 ( .A(n8729), .ZN(n8730) );
  NAND2_X1 U11194 ( .A1(n10673), .A2(n8730), .ZN(n10668) );
  INV_X1 U11195 ( .A(n10557), .ZN(n15589) );
  INV_X1 U11196 ( .A(n11301), .ZN(n15556) );
  XNOR2_X1 U11197 ( .A(n15561), .B(n8787), .ZN(n8735) );
  XNOR2_X1 U11198 ( .A(n8735), .B(n11505), .ZN(n11081) );
  XNOR2_X1 U11199 ( .A(n15540), .B(n7688), .ZN(n12818) );
  XNOR2_X1 U11200 ( .A(n12824), .B(n7688), .ZN(n8740) );
  XNOR2_X1 U11201 ( .A(n8740), .B(n12491), .ZN(n12820) );
  INV_X1 U11202 ( .A(n12820), .ZN(n8738) );
  OR2_X1 U11203 ( .A1(n11505), .A2(n8735), .ZN(n11312) );
  INV_X1 U11204 ( .A(n11451), .ZN(n15555) );
  XNOR2_X1 U11205 ( .A(n11318), .B(n8787), .ZN(n11314) );
  INV_X1 U11206 ( .A(n11314), .ZN(n8736) );
  NAND2_X1 U11207 ( .A1(n15555), .A2(n8736), .ZN(n8737) );
  INV_X1 U11208 ( .A(n12951), .ZN(n11319) );
  INV_X1 U11209 ( .A(n12818), .ZN(n11448) );
  OAI21_X1 U11210 ( .B1(n11319), .B2(n12820), .A(n11448), .ZN(n8742) );
  NAND2_X1 U11211 ( .A1(n11314), .A2(n11451), .ZN(n11446) );
  XNOR2_X1 U11212 ( .A(n11651), .B(n8787), .ZN(n8744) );
  XNOR2_X1 U11213 ( .A(n8744), .B(n15528), .ZN(n11325) );
  NOR2_X1 U11214 ( .A1(n8744), .A2(n15528), .ZN(n11588) );
  XNOR2_X1 U11215 ( .A(n15534), .B(n8787), .ZN(n8745) );
  XNOR2_X1 U11216 ( .A(n8745), .B(n11807), .ZN(n11591) );
  AND2_X1 U11217 ( .A1(n8745), .A2(n11807), .ZN(n8746) );
  XNOR2_X1 U11218 ( .A(n12507), .B(n8787), .ZN(n8749) );
  XNOR2_X1 U11219 ( .A(n14854), .B(n8787), .ZN(n8751) );
  NAND2_X1 U11220 ( .A1(n8751), .A2(n14863), .ZN(n11860) );
  XNOR2_X1 U11221 ( .A(n13422), .B(n8787), .ZN(n12889) );
  NOR2_X1 U11222 ( .A1(n12889), .A2(n14851), .ZN(n8753) );
  INV_X1 U11223 ( .A(n12889), .ZN(n8752) );
  XNOR2_X1 U11224 ( .A(n13418), .B(n7688), .ZN(n8754) );
  NAND2_X1 U11225 ( .A1(n8754), .A2(n13286), .ZN(n8755) );
  OAI21_X1 U11226 ( .B1(n8754), .B2(n13286), .A(n8755), .ZN(n12782) );
  NAND2_X1 U11227 ( .A1(n12932), .A2(n12949), .ZN(n8757) );
  XNOR2_X1 U11228 ( .A(n13264), .B(n8787), .ZN(n12933) );
  XNOR2_X1 U11229 ( .A(n12849), .B(n8787), .ZN(n8758) );
  XNOR2_X1 U11230 ( .A(n8758), .B(n12948), .ZN(n12851) );
  XNOR2_X1 U11231 ( .A(n8761), .B(n13249), .ZN(n12860) );
  INV_X1 U11232 ( .A(n12860), .ZN(n8762) );
  OAI21_X1 U11233 ( .B1(n8763), .B2(n12915), .A(n12857), .ZN(n12911) );
  XNOR2_X1 U11234 ( .A(n13228), .B(n8787), .ZN(n8765) );
  XNOR2_X1 U11235 ( .A(n8765), .B(n13236), .ZN(n12910) );
  INV_X1 U11236 ( .A(n12910), .ZN(n8764) );
  INV_X1 U11237 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11238 ( .A1(n8766), .A2(n13203), .ZN(n8767) );
  XNOR2_X1 U11239 ( .A(n12798), .B(n8787), .ZN(n8769) );
  XNOR2_X1 U11240 ( .A(n8769), .B(n13187), .ZN(n12800) );
  XNOR2_X1 U11241 ( .A(n13332), .B(n8787), .ZN(n12881) );
  NAND2_X1 U11242 ( .A1(n12881), .A2(n13175), .ZN(n8768) );
  INV_X1 U11243 ( .A(n8768), .ZN(n8774) );
  INV_X1 U11244 ( .A(n8769), .ZN(n8770) );
  NAND2_X1 U11245 ( .A1(n8770), .A2(n13187), .ZN(n12879) );
  INV_X1 U11246 ( .A(n12881), .ZN(n8771) );
  NAND2_X1 U11247 ( .A1(n8771), .A2(n13204), .ZN(n8772) );
  AND2_X1 U11248 ( .A1(n12879), .A2(n8772), .ZN(n8773) );
  XNOR2_X1 U11249 ( .A(n13179), .B(n8787), .ZN(n8776) );
  NAND2_X1 U11250 ( .A1(n8776), .A2(n13162), .ZN(n8778) );
  OAI21_X1 U11251 ( .B1(n8776), .B2(n13162), .A(n8778), .ZN(n12833) );
  INV_X1 U11252 ( .A(n12833), .ZN(n8777) );
  XNOR2_X1 U11253 ( .A(n13314), .B(n8787), .ZN(n8783) );
  NAND2_X1 U11254 ( .A1(n8783), .A2(n13145), .ZN(n12844) );
  INV_X1 U11255 ( .A(n8783), .ZN(n8784) );
  NAND2_X1 U11256 ( .A1(n8784), .A2(n13115), .ZN(n8785) );
  NAND2_X1 U11257 ( .A1(n8786), .A2(n12868), .ZN(n12842) );
  XNOR2_X1 U11258 ( .A(n13120), .B(n8787), .ZN(n8788) );
  NAND2_X1 U11259 ( .A1(n8788), .A2(n13130), .ZN(n8791) );
  INV_X1 U11260 ( .A(n8788), .ZN(n8789) );
  NAND2_X1 U11261 ( .A1(n8789), .A2(n12874), .ZN(n8790) );
  XNOR2_X1 U11262 ( .A(n13306), .B(n7688), .ZN(n8792) );
  NOR2_X1 U11263 ( .A1(n8792), .A2(n13116), .ZN(n8793) );
  AOI21_X1 U11264 ( .B1(n8792), .B2(n13116), .A(n8793), .ZN(n12923) );
  OAI22_X1 U11265 ( .A1(n8803), .A2(n10443), .B1(n8810), .B2(n8804), .ZN(n8795) );
  NAND2_X1 U11266 ( .A1(n8796), .A2(n12924), .ZN(n8819) );
  INV_X1 U11267 ( .A(n15585), .ZN(n15617) );
  NAND2_X1 U11268 ( .A1(n8803), .A2(n15617), .ZN(n8798) );
  NOR2_X1 U11269 ( .A1(n8800), .A2(n15588), .ZN(n8799) );
  INV_X1 U11270 ( .A(n8810), .ZN(n8801) );
  NOR2_X1 U11271 ( .A1(n8800), .A2(n15590), .ZN(n12604) );
  NAND2_X1 U11272 ( .A1(n12604), .A2(n8801), .ZN(n12941) );
  NAND2_X1 U11273 ( .A1(n8803), .A2(n8802), .ZN(n8808) );
  INV_X1 U11274 ( .A(n8804), .ZN(n8805) );
  NAND2_X1 U11275 ( .A1(n8810), .A2(n8805), .ZN(n8806) );
  NAND4_X1 U11276 ( .A1(n8808), .A2(n10070), .A3(n8807), .A4(n8806), .ZN(n8809) );
  NAND2_X1 U11277 ( .A1(n8809), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11278 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  OR2_X1 U11279 ( .A1(n10679), .A2(P3_U3151), .ZN(n12608) );
  AOI22_X1 U11280 ( .A1(n13095), .A2(n12938), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(n6665), .ZN(n8814) );
  OAI21_X1 U11281 ( .B1(n13090), .B2(n12941), .A(n8814), .ZN(n8815) );
  AOI21_X1 U11282 ( .B1(n10956), .B2(n12936), .A(n8815), .ZN(n8816) );
  INV_X1 U11283 ( .A(n8817), .ZN(n8818) );
  NAND2_X1 U11284 ( .A1(n8819), .A2(n8818), .ZN(P3_U3154) );
  INV_X1 U11285 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8843) );
  XOR2_X1 U11286 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n8856) );
  INV_X1 U11287 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8841) );
  INV_X1 U11288 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8839) );
  INV_X1 U11289 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n8835) );
  INV_X1 U11290 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U11291 ( .A1(n8864), .A2(n8863), .ZN(n8820) );
  NAND2_X1 U11292 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U11293 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U11294 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8824), .ZN(n8825) );
  NAND2_X1 U11295 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8826), .ZN(n8827) );
  NAND2_X1 U11296 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9008), .ZN(n8828) );
  NOR2_X1 U11297 ( .A1(n8830), .A2(n9161), .ZN(n8832) );
  XNOR2_X1 U11298 ( .A(n9161), .B(n8830), .ZN(n8886) );
  INV_X1 U11299 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9227) );
  XNOR2_X1 U11300 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9227), .ZN(n8859) );
  XNOR2_X1 U11301 ( .A(n8835), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11302 ( .A1(n8836), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n8838) );
  XOR2_X1 U11303 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8836), .Z(n8895) );
  INV_X1 U11304 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11305 ( .A(n8839), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n8857) );
  XNOR2_X1 U11306 ( .A(n8841), .B(P3_ADDR_REG_12__SCAN_IN), .ZN(n8898) );
  INV_X1 U11307 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8900) );
  AND2_X1 U11308 ( .A1(n8900), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n8842) );
  INV_X1 U11309 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U11310 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12993), .ZN(n8844) );
  NOR2_X1 U11311 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12993), .ZN(n8852) );
  NAND2_X1 U11312 ( .A1(n8845), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8847) );
  INV_X1 U11313 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U11314 ( .A1(n8906), .A2(n13013), .ZN(n8846) );
  NAND2_X1 U11315 ( .A1(n8847), .A2(n8846), .ZN(n8848) );
  NOR2_X1 U11316 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8848), .ZN(n8851) );
  INV_X1 U11317 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n8849) );
  XNOR2_X1 U11318 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8848), .ZN(n8907) );
  NOR2_X1 U11319 ( .A1(n8849), .A2(n8907), .ZN(n8850) );
  NOR2_X1 U11320 ( .A1(n8851), .A2(n8850), .ZN(n8914) );
  XOR2_X1 U11321 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n8913) );
  XOR2_X1 U11322 ( .A(n8914), .B(n8913), .Z(n14785) );
  AOI21_X1 U11323 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n12993), .A(n8852), .ZN(
        n8854) );
  XOR2_X1 U11324 ( .A(n8854), .B(n8853), .Z(n15044) );
  XNOR2_X1 U11325 ( .A(n8856), .B(n8855), .ZN(n15040) );
  XOR2_X1 U11326 ( .A(n8858), .B(n8857), .Z(n15028) );
  XOR2_X1 U11327 ( .A(n8860), .B(n8859), .Z(n8890) );
  XNOR2_X1 U11328 ( .A(n8862), .B(n8861), .ZN(n8875) );
  AND2_X1 U11329 ( .A1(n8875), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n8876) );
  NOR2_X1 U11330 ( .A1(n8866), .A2(n7532), .ZN(n8867) );
  AOI21_X1 U11331 ( .B1(n9033), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n8864), .ZN(
        n8865) );
  INV_X1 U11332 ( .A(n8865), .ZN(n15692) );
  NAND2_X1 U11333 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15692), .ZN(n15702) );
  NOR2_X1 U11334 ( .A1(n15702), .A2(n15701), .ZN(n15700) );
  XOR2_X1 U11335 ( .A(n8869), .B(n8868), .Z(n8870) );
  INV_X1 U11336 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14791) );
  XOR2_X1 U11337 ( .A(n8873), .B(n8872), .Z(n15697) );
  NAND2_X1 U11338 ( .A1(n15698), .A2(n15697), .ZN(n15696) );
  XNOR2_X1 U11339 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8875), .ZN(n15687) );
  NOR2_X1 U11340 ( .A1(n15688), .A2(n15687), .ZN(n15686) );
  XOR2_X1 U11341 ( .A(n8878), .B(n8877), .Z(n8880) );
  NAND2_X1 U11342 ( .A1(n8879), .A2(n8880), .ZN(n8881) );
  XOR2_X1 U11343 ( .A(n8880), .B(n8879), .Z(n15691) );
  INV_X1 U11344 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15690) );
  NAND2_X1 U11345 ( .A1(n15691), .A2(n15690), .ZN(n15689) );
  NOR2_X1 U11346 ( .A1(n8884), .A2(n7088), .ZN(n8885) );
  XOR2_X1 U11347 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9008), .Z(n8883) );
  XOR2_X1 U11348 ( .A(n8883), .B(n8882), .Z(n14795) );
  NOR2_X1 U11349 ( .A1(n8887), .A2(n7524), .ZN(n8888) );
  XOR2_X1 U11350 ( .A(n8886), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n15695) );
  NOR2_X1 U11351 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  XNOR2_X1 U11352 ( .A(n8890), .B(n8889), .ZN(n14798) );
  INV_X1 U11353 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14797) );
  NOR2_X1 U11354 ( .A1(n14798), .A2(n14797), .ZN(n14796) );
  XOR2_X1 U11355 ( .A(n8893), .B(n8892), .Z(n14800) );
  NAND2_X1 U11356 ( .A1(n14801), .A2(n14800), .ZN(n8894) );
  NOR2_X1 U11357 ( .A1(n14801), .A2(n14800), .ZN(n14799) );
  AOI21_X2 U11358 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n8894), .A(n14799), .ZN(
        n14805) );
  XOR2_X1 U11359 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n8895), .Z(n14804) );
  NAND2_X1 U11360 ( .A1(n14805), .A2(n14804), .ZN(n8896) );
  NAND2_X1 U11361 ( .A1(n15028), .A2(n15027), .ZN(n8897) );
  NOR2_X1 U11362 ( .A1(n15028), .A2(n15027), .ZN(n15026) );
  XOR2_X1 U11363 ( .A(n8899), .B(n8898), .Z(n15031) );
  XOR2_X1 U11364 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(n8900), .Z(n8902) );
  XOR2_X1 U11365 ( .A(n8902), .B(n8901), .Z(n8903) );
  INV_X1 U11366 ( .A(n15034), .ZN(n15035) );
  INV_X1 U11367 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15037) );
  NAND2_X1 U11368 ( .A1(n15037), .A2(n15036), .ZN(n15033) );
  NAND2_X1 U11369 ( .A1(n15035), .A2(n15033), .ZN(n15039) );
  NOR2_X1 U11370 ( .A1(n15040), .A2(n15039), .ZN(n8905) );
  NAND2_X1 U11371 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  OAI21_X2 U11372 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n8905), .A(n15038), .ZN(
        n15043) );
  XOR2_X1 U11373 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n8906), .Z(n15047) );
  XOR2_X1 U11374 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8907), .Z(n8908) );
  INV_X1 U11375 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U11376 ( .A1(n8909), .A2(n8908), .ZN(n14810) );
  XNOR2_X1 U11377 ( .A(n8910), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11378 ( .A(n8911), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8912) );
  INV_X1 U11379 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n8916) );
  NOR2_X1 U11380 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  AOI21_X1 U11381 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n8916), .A(n8915), .ZN(
        n9249) );
  OAI22_X1 U11382 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g122), .B2(P1_IR_REG_15__SCAN_IN), .ZN(n8917) );
  AOI221_X1 U11383 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_g122), .A(n8917), .ZN(n8924) );
  OAI22_X1 U11384 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        SI_16_), .B2(keyinput_g16), .ZN(n8918) );
  AOI221_X1 U11385 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        keyinput_g16), .C2(SI_16_), .A(n8918), .ZN(n8923) );
  OAI22_X1 U11386 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g124), .B1(
        P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n8919) );
  AOI221_X1 U11387 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g93), .C2(P3_DATAO_REG_3__SCAN_IN), .A(n8919), .ZN(n8922) );
  OAI22_X1 U11388 ( .A1(SI_12_), .A2(keyinput_g20), .B1(keyinput_g85), .B2(
        P3_DATAO_REG_11__SCAN_IN), .ZN(n8920) );
  AOI221_X1 U11389 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P3_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n8920), .ZN(n8921) );
  NAND4_X1 U11390 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n8952)
         );
  OAI22_X1 U11391 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P3_ADDR_REG_3__SCAN_IN), 
        .B2(keyinput_g100), .ZN(n8925) );
  AOI221_X1 U11392 ( .B1(SI_29_), .B2(keyinput_g3), .C1(keyinput_g100), .C2(
        P3_ADDR_REG_3__SCAN_IN), .A(n8925), .ZN(n8932) );
  OAI22_X1 U11393 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g67), .B2(
        P3_DATAO_REG_29__SCAN_IN), .ZN(n8926) );
  AOI221_X1 U11394 ( .B1(SI_25_), .B2(keyinput_g7), .C1(
        P3_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n8926), .ZN(n8931) );
  OAI22_X1 U11395 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .ZN(n8927) );
  AOI221_X1 U11396 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g66), .C2(P3_DATAO_REG_30__SCAN_IN), .A(n8927), .ZN(n8930) );
  OAI22_X1 U11397 ( .A1(SI_26_), .A2(keyinput_g6), .B1(P1_IR_REG_11__SCAN_IN), 
        .B2(keyinput_g118), .ZN(n8928) );
  AOI221_X1 U11398 ( .B1(SI_26_), .B2(keyinput_g6), .C1(keyinput_g118), .C2(
        P1_IR_REG_11__SCAN_IN), .A(n8928), .ZN(n8929) );
  NAND4_X1 U11399 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n8951)
         );
  OAI22_X1 U11400 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g123), .B1(
        keyinput_g91), .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n8933) );
  AOI221_X1 U11401 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g123), .C1(
        P3_DATAO_REG_5__SCAN_IN), .C2(keyinput_g91), .A(n8933), .ZN(n8940) );
  OAI22_X1 U11402 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(
        P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .ZN(n8934) );
  AOI221_X1 U11403 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        keyinput_g89), .C2(P3_DATAO_REG_7__SCAN_IN), .A(n8934), .ZN(n8939) );
  OAI22_X1 U11404 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P1_IR_REG_2__SCAN_IN), 
        .B2(keyinput_g109), .ZN(n8935) );
  AOI221_X1 U11405 ( .B1(SI_8_), .B2(keyinput_g24), .C1(keyinput_g109), .C2(
        P1_IR_REG_2__SCAN_IN), .A(n8935), .ZN(n8938) );
  OAI22_X1 U11406 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g88), .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n8936) );
  AOI221_X1 U11407 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P3_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n8936), .ZN(n8937) );
  NAND4_X1 U11408 ( .A1(n8940), .A2(n8939), .A3(n8938), .A4(n8937), .ZN(n8950)
         );
  OAI22_X1 U11409 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_g107), .ZN(n8941) );
  AOI221_X1 U11410 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g107), .C2(P1_IR_REG_0__SCAN_IN), .A(n8941), .ZN(n8948) );
  OAI22_X1 U11411 ( .A1(SI_27_), .A2(keyinput_g5), .B1(keyinput_g12), .B2(
        SI_20_), .ZN(n8942) );
  AOI221_X1 U11412 ( .B1(SI_27_), .B2(keyinput_g5), .C1(SI_20_), .C2(
        keyinput_g12), .A(n8942), .ZN(n8947) );
  OAI22_X1 U11413 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n8943) );
  AOI221_X1 U11414 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        keyinput_g41), .C2(P3_REG3_REG_19__SCAN_IN), .A(n8943), .ZN(n8946) );
  OAI22_X1 U11415 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g114), .ZN(n8944) );
  AOI221_X1 U11416 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        keyinput_g114), .C2(P1_IR_REG_7__SCAN_IN), .A(n8944), .ZN(n8945) );
  NAND4_X1 U11417 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(n8949)
         );
  NOR4_X1 U11418 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n8949), .ZN(n9247)
         );
  OAI22_X1 U11419 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_g101), .B1(
        P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_g96), .ZN(n8953) );
  AOI221_X1 U11420 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_g101), .C1(
        keyinput_g96), .C2(P3_DATAO_REG_0__SCAN_IN), .A(n8953), .ZN(n8960) );
  OAI22_X1 U11421 ( .A1(SI_7_), .A2(keyinput_g25), .B1(
        P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .ZN(n8954) );
  AOI221_X1 U11422 ( .B1(SI_7_), .B2(keyinput_g25), .C1(keyinput_g80), .C2(
        P3_DATAO_REG_16__SCAN_IN), .A(n8954), .ZN(n8959) );
  OAI22_X1 U11423 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n8955) );
  AOI221_X1 U11424 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        keyinput_g75), .C2(P3_DATAO_REG_21__SCAN_IN), .A(n8955), .ZN(n8958) );
  OAI22_X1 U11425 ( .A1(SI_15_), .A2(keyinput_g17), .B1(
        P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .ZN(n8956) );
  AOI221_X1 U11426 ( .B1(SI_15_), .B2(keyinput_g17), .C1(keyinput_g94), .C2(
        P3_DATAO_REG_2__SCAN_IN), .A(n8956), .ZN(n8957) );
  NAND4_X1 U11427 ( .A1(n8960), .A2(n8959), .A3(n8958), .A4(n8957), .ZN(n9076)
         );
  OAI22_X1 U11428 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g126), .B1(
        keyinput_g127), .B2(P1_IR_REG_20__SCAN_IN), .ZN(n8961) );
  AOI221_X1 U11429 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n8961), .ZN(n8986) );
  INV_X1 U11430 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10235) );
  OAI22_X1 U11431 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g120), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .ZN(n8962) );
  AOI221_X1 U11432 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g120), .C1(
        keyinput_g70), .C2(P3_DATAO_REG_26__SCAN_IN), .A(n8962), .ZN(n8965) );
  OAI22_X1 U11433 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        keyinput_g83), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n8963) );
  AOI221_X1 U11434 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P3_DATAO_REG_13__SCAN_IN), .C2(keyinput_g83), .A(n8963), .ZN(n8964) );
  OAI211_X1 U11435 ( .C1(n10235), .C2(keyinput_g77), .A(n8965), .B(n8964), 
        .ZN(n8966) );
  AOI21_X1 U11436 ( .B1(n10235), .B2(keyinput_g77), .A(n8966), .ZN(n8985) );
  AOI22_X1 U11437 ( .A1(P3_DATAO_REG_18__SCAN_IN), .A2(keyinput_g78), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_g105), .ZN(n8967) );
  OAI221_X1 U11438 ( .B1(P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .C1(
        P3_ADDR_REG_8__SCAN_IN), .C2(keyinput_g105), .A(n8967), .ZN(n8974) );
  AOI22_X1 U11439 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .ZN(n8968) );
  OAI221_X1 U11440 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P3_ADDR_REG_7__SCAN_IN), .C2(keyinput_g104), .A(n8968), .ZN(n8973) );
  AOI22_X1 U11441 ( .A1(P3_DATAO_REG_6__SCAN_IN), .A2(keyinput_g90), .B1(SI_0_), .B2(keyinput_g32), .ZN(n8969) );
  OAI221_X1 U11442 ( .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .C1(
        SI_0_), .C2(keyinput_g32), .A(n8969), .ZN(n8972) );
  AOI22_X1 U11443 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g110), .B1(SI_31_), 
        .B2(keyinput_g1), .ZN(n8970) );
  OAI221_X1 U11444 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g110), .C1(SI_31_), .C2(keyinput_g1), .A(n8970), .ZN(n8971) );
  NOR4_X1 U11445 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(n8984)
         );
  AOI22_X1 U11446 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n8975) );
  OAI221_X1 U11447 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_22_), .C2(
        keyinput_g10), .A(n8975), .ZN(n8982) );
  AOI22_X1 U11448 ( .A1(SI_21_), .A2(keyinput_g11), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n8976) );
  OAI221_X1 U11449 ( .B1(SI_21_), .B2(keyinput_g11), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n8976), .ZN(n8981) );
  AOI22_X1 U11450 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_18_), .B2(keyinput_g14), .ZN(n8977) );
  OAI221_X1 U11451 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        SI_18_), .C2(keyinput_g14), .A(n8977), .ZN(n8980) );
  AOI22_X1 U11452 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_1_), .B2(
        keyinput_g31), .ZN(n8978) );
  OAI221_X1 U11453 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_1_), .C2(
        keyinput_g31), .A(n8978), .ZN(n8979) );
  NOR4_X1 U11454 ( .A1(n8982), .A2(n8981), .A3(n8980), .A4(n8979), .ZN(n8983)
         );
  NAND4_X1 U11455 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .ZN(n9075)
         );
  INV_X1 U11456 ( .A(SI_17_), .ZN(n10185) );
  AOI22_X1 U11457 ( .A1(n10185), .A2(keyinput_g15), .B1(n15586), .B2(
        keyinput_g59), .ZN(n8987) );
  OAI221_X1 U11458 ( .B1(n10185), .B2(keyinput_g15), .C1(n15586), .C2(
        keyinput_g59), .A(n8987), .ZN(n8996) );
  XOR2_X1 U11459 ( .A(n8988), .B(keyinput_g98), .Z(n8992) );
  XNOR2_X1 U11460 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g113), .ZN(n8991) );
  XNOR2_X1 U11461 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n8990) );
  XNOR2_X1 U11462 ( .A(SI_5_), .B(keyinput_g27), .ZN(n8989) );
  NAND4_X1 U11463 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(n8989), .ZN(n8995)
         );
  XNOR2_X1 U11464 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_g81), .ZN(n8994)
         );
  XNOR2_X1 U11465 ( .A(keyinput_g56), .B(n8417), .ZN(n8993) );
  NOR4_X1 U11466 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n9029)
         );
  INV_X1 U11467 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U11468 ( .A1(n11443), .A2(keyinput_g8), .B1(n12935), .B2(
        keyinput_g63), .ZN(n8997) );
  OAI221_X1 U11469 ( .B1(n11443), .B2(keyinput_g8), .C1(n12935), .C2(
        keyinput_g63), .A(n8997), .ZN(n9006) );
  INV_X1 U11470 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9162) );
  AOI22_X1 U11471 ( .A1(n9162), .A2(keyinput_g62), .B1(keyinput_g102), .B2(
        n7097), .ZN(n8998) );
  OAI221_X1 U11472 ( .B1(n9162), .B2(keyinput_g62), .C1(n7097), .C2(
        keyinput_g102), .A(n8998), .ZN(n9005) );
  INV_X1 U11473 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U11474 ( .A1(n10884), .A2(keyinput_g65), .B1(n6665), .B2(
        keyinput_g34), .ZN(n8999) );
  OAI221_X1 U11475 ( .B1(n10884), .B2(keyinput_g65), .C1(n6665), .C2(
        keyinput_g34), .A(n8999), .ZN(n9004) );
  XOR2_X1 U11476 ( .A(n9000), .B(keyinput_g99), .Z(n9002) );
  XNOR2_X1 U11477 ( .A(SI_3_), .B(keyinput_g29), .ZN(n9001) );
  NAND2_X1 U11478 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  NOR4_X1 U11479 ( .A1(n9006), .A2(n9005), .A3(n9004), .A4(n9003), .ZN(n9028)
         );
  AOI22_X1 U11480 ( .A1(n10116), .A2(keyinput_g21), .B1(keyinput_g103), .B2(
        n9008), .ZN(n9007) );
  OAI221_X1 U11481 ( .B1(n10116), .B2(keyinput_g21), .C1(n9008), .C2(
        keyinput_g103), .A(n9007), .ZN(n9012) );
  INV_X1 U11482 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n10169) );
  INV_X1 U11483 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9177) );
  AOI22_X1 U11484 ( .A1(n10169), .A2(keyinput_g82), .B1(n9177), .B2(
        keyinput_g38), .ZN(n9009) );
  OAI221_X1 U11485 ( .B1(n10169), .B2(keyinput_g82), .C1(n9177), .C2(
        keyinput_g38), .A(n9009), .ZN(n9011) );
  XOR2_X1 U11486 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g125), .Z(n9010) );
  OR3_X1 U11487 ( .A1(n9012), .A2(n9011), .A3(n9010), .ZN(n9016) );
  INV_X1 U11488 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11489 ( .A1(n10239), .A2(keyinput_g76), .B1(n12414), .B2(
        keyinput_g2), .ZN(n9013) );
  OAI221_X1 U11490 ( .B1(n10239), .B2(keyinput_g76), .C1(n12414), .C2(
        keyinput_g2), .A(n9013), .ZN(n9015) );
  INV_X1 U11491 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n10958) );
  XNOR2_X1 U11492 ( .A(n10958), .B(keyinput_g68), .ZN(n9014) );
  NOR3_X1 U11493 ( .A1(n9016), .A2(n9015), .A3(n9014), .ZN(n9027) );
  INV_X1 U11494 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n10233) );
  INV_X1 U11495 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U11496 ( .A1(n10233), .A2(keyinput_g87), .B1(keyinput_g95), .B2(
        n10392), .ZN(n9017) );
  OAI221_X1 U11497 ( .B1(n10233), .B2(keyinput_g87), .C1(n10392), .C2(
        keyinput_g95), .A(n9017), .ZN(n9025) );
  INV_X1 U11498 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9164) );
  AOI22_X1 U11499 ( .A1(n10046), .A2(keyinput_g119), .B1(n9164), .B2(
        keyinput_g60), .ZN(n9018) );
  OAI221_X1 U11500 ( .B1(n10046), .B2(keyinput_g119), .C1(n9164), .C2(
        keyinput_g60), .A(n9018), .ZN(n9024) );
  INV_X1 U11501 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n10548) );
  XNOR2_X1 U11502 ( .A(n10548), .B(keyinput_g71), .ZN(n9023) );
  XNOR2_X1 U11503 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n9021) );
  XNOR2_X1 U11504 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9020) );
  XNOR2_X1 U11505 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g117), .ZN(n9019)
         );
  NAND3_X1 U11506 ( .A1(n9021), .A2(n9020), .A3(n9019), .ZN(n9022) );
  NOR4_X1 U11507 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n9026)
         );
  NAND4_X1 U11508 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(n9074)
         );
  INV_X1 U11509 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n10418) );
  INV_X1 U11510 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9031) );
  AOI22_X1 U11511 ( .A1(n10418), .A2(keyinput_g72), .B1(n9031), .B2(
        keyinput_g0), .ZN(n9030) );
  OAI221_X1 U11512 ( .B1(n10418), .B2(keyinput_g72), .C1(n9031), .C2(
        keyinput_g0), .A(n9030), .ZN(n9040) );
  INV_X1 U11513 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U11514 ( .A1(n10181), .A2(keyinput_g92), .B1(n9033), .B2(
        keyinput_g97), .ZN(n9032) );
  OAI221_X1 U11515 ( .B1(n10181), .B2(keyinput_g92), .C1(n9033), .C2(
        keyinput_g97), .A(n9032), .ZN(n9039) );
  INV_X1 U11516 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U11517 ( .A1(n10809), .A2(keyinput_g69), .B1(n12823), .B2(
        keyinput_g43), .ZN(n9034) );
  OAI221_X1 U11518 ( .B1(n10809), .B2(keyinput_g69), .C1(n12823), .C2(
        keyinput_g43), .A(n9034), .ZN(n9038) );
  XNOR2_X1 U11519 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n9036) );
  XNOR2_X1 U11520 ( .A(SI_28_), .B(keyinput_g4), .ZN(n9035) );
  NAND2_X1 U11521 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NOR4_X1 U11522 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(n9072)
         );
  INV_X1 U11523 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U11524 ( .A1(n9042), .A2(keyinput_g48), .B1(keyinput_g84), .B2(
        n10272), .ZN(n9041) );
  OAI221_X1 U11525 ( .B1(n9042), .B2(keyinput_g48), .C1(n10272), .C2(
        keyinput_g84), .A(n9041), .ZN(n9051) );
  INV_X1 U11526 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U11527 ( .A1(n10374), .A2(keyinput_g73), .B1(n8277), .B2(
        keyinput_g49), .ZN(n9043) );
  OAI221_X1 U11528 ( .B1(n10374), .B2(keyinput_g73), .C1(n8277), .C2(
        keyinput_g49), .A(n9043), .ZN(n9050) );
  INV_X1 U11529 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9045) );
  AOI22_X1 U11530 ( .A1(n10308), .A2(keyinput_g13), .B1(keyinput_g106), .B2(
        n9045), .ZN(n9044) );
  OAI221_X1 U11531 ( .B1(n10308), .B2(keyinput_g13), .C1(n9045), .C2(
        keyinput_g106), .A(n9044), .ZN(n9049) );
  XNOR2_X1 U11532 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n9047)
         );
  XNOR2_X1 U11533 ( .A(SI_6_), .B(keyinput_g26), .ZN(n9046) );
  NAND2_X1 U11534 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  NOR4_X1 U11535 ( .A1(n9051), .A2(n9050), .A3(n9049), .A4(n9048), .ZN(n9071)
         );
  AOI22_X1 U11536 ( .A1(n12861), .A2(keyinput_g50), .B1(keyinput_g19), .B2(
        n10139), .ZN(n9052) );
  OAI221_X1 U11537 ( .B1(n12861), .B2(keyinput_g50), .C1(n10139), .C2(
        keyinput_g19), .A(n9052), .ZN(n9060) );
  INV_X2 U11538 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11539 ( .A1(n9174), .A2(keyinput_g55), .B1(keyinput_g121), .B2(
        n10044), .ZN(n9053) );
  OAI221_X1 U11540 ( .B1(n9174), .B2(keyinput_g55), .C1(n10044), .C2(
        keyinput_g121), .A(n9053), .ZN(n9059) );
  XOR2_X1 U11541 ( .A(n12834), .B(keyinput_g45), .Z(n9057) );
  XNOR2_X1 U11542 ( .A(SI_14_), .B(keyinput_g18), .ZN(n9056) );
  XNOR2_X1 U11543 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g112), .ZN(n9055) );
  XNOR2_X1 U11544 ( .A(SI_9_), .B(keyinput_g23), .ZN(n9054) );
  NAND4_X1 U11545 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9058)
         );
  NOR3_X1 U11546 ( .A1(n9060), .A2(n9059), .A3(n9058), .ZN(n9070) );
  INV_X1 U11547 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11317) );
  INV_X1 U11548 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U11549 ( .A1(n11317), .A2(keyinput_g61), .B1(keyinput_g116), .B2(
        n10162), .ZN(n9061) );
  OAI221_X1 U11550 ( .B1(n11317), .B2(keyinput_g61), .C1(n10162), .C2(
        keyinput_g116), .A(n9061), .ZN(n9068) );
  INV_X1 U11551 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11384) );
  INV_X1 U11552 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U11553 ( .A1(n11384), .A2(keyinput_g58), .B1(keyinput_g74), .B2(
        n10237), .ZN(n9062) );
  OAI221_X1 U11554 ( .B1(n11384), .B2(keyinput_g58), .C1(n10237), .C2(
        keyinput_g74), .A(n9062), .ZN(n9067) );
  INV_X1 U11555 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9183) );
  AOI22_X1 U11556 ( .A1(n11054), .A2(keyinput_g9), .B1(n9183), .B2(
        keyinput_g47), .ZN(n9063) );
  OAI221_X1 U11557 ( .B1(n11054), .B2(keyinput_g9), .C1(n9183), .C2(
        keyinput_g47), .A(n9063), .ZN(n9066) );
  INV_X1 U11558 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11309) );
  INV_X1 U11559 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U11560 ( .A1(n11309), .A2(keyinput_g40), .B1(n11137), .B2(
        keyinput_g39), .ZN(n9064) );
  OAI221_X1 U11561 ( .B1(n11309), .B2(keyinput_g40), .C1(n11137), .C2(
        keyinput_g39), .A(n9064), .ZN(n9065) );
  NOR4_X1 U11562 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(n9069)
         );
  NAND4_X1 U11563 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n9073)
         );
  NOR4_X1 U11564 ( .A1(n9076), .A2(n9075), .A3(n9074), .A4(n9073), .ZN(n9246)
         );
  XOR2_X1 U11565 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g115), .Z(n9245) );
  XNOR2_X1 U11566 ( .A(n10235), .B(keyinput_f77), .ZN(n9083) );
  AOI22_X1 U11567 ( .A1(SI_0_), .A2(keyinput_f32), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n9077) );
  OAI221_X1 U11568 ( .B1(SI_0_), .B2(keyinput_f32), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n9077), .ZN(n9082) );
  AOI22_X1 U11569 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f113), .B1(SI_14_), 
        .B2(keyinput_f18), .ZN(n9078) );
  OAI221_X1 U11570 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .C1(SI_14_), .C2(keyinput_f18), .A(n9078), .ZN(n9081) );
  AOI22_X1 U11571 ( .A1(keyinput_f92), .A2(P3_DATAO_REG_4__SCAN_IN), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f126), .ZN(n9079) );
  OAI221_X1 U11572 ( .B1(keyinput_f92), .B2(P3_DATAO_REG_4__SCAN_IN), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n9079), .ZN(n9080) );
  NOR4_X1 U11573 ( .A1(n9083), .A2(n9082), .A3(n9081), .A4(n9080), .ZN(n9111)
         );
  AOI22_X1 U11574 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_B_REG_SCAN_IN), .B2(
        keyinput_f64), .ZN(n9084) );
  OAI221_X1 U11575 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P3_B_REG_SCAN_IN), 
        .C2(keyinput_f64), .A(n9084), .ZN(n9091) );
  AOI22_X1 U11576 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_f103), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n9085) );
  OAI221_X1 U11577 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_f103), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n9085), .ZN(n9090) );
  AOI22_X1 U11578 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_f100), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n9086) );
  OAI221_X1 U11579 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_f100), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n9086), .ZN(n9089) );
  AOI22_X1 U11580 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f112), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f124), .ZN(n9087) );
  OAI221_X1 U11581 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f124), .A(n9087), .ZN(n9088) );
  NOR4_X1 U11582 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), .ZN(n9110)
         );
  AOI22_X1 U11583 ( .A1(keyinput_f68), .A2(P3_DATAO_REG_28__SCAN_IN), .B1(
        keyinput_f78), .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n9092) );
  OAI221_X1 U11584 ( .B1(keyinput_f68), .B2(P3_DATAO_REG_28__SCAN_IN), .C1(
        keyinput_f78), .C2(P3_DATAO_REG_18__SCAN_IN), .A(n9092), .ZN(n9099) );
  AOI22_X1 U11585 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n9093) );
  OAI221_X1 U11586 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_27_), .C2(
        keyinput_f5), .A(n9093), .ZN(n9098) );
  AOI22_X1 U11587 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n9094) );
  OAI221_X1 U11588 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n9094), .ZN(n9097) );
  AOI22_X1 U11589 ( .A1(SI_26_), .A2(keyinput_f6), .B1(SI_9_), .B2(
        keyinput_f23), .ZN(n9095) );
  OAI221_X1 U11590 ( .B1(SI_26_), .B2(keyinput_f6), .C1(SI_9_), .C2(
        keyinput_f23), .A(n9095), .ZN(n9096) );
  NOR4_X1 U11591 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), .ZN(n9109)
         );
  AOI22_X1 U11592 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_13_), .B2(keyinput_f19), .ZN(n9100) );
  OAI221_X1 U11593 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_13_), .C2(keyinput_f19), .A(n9100), .ZN(n9107) );
  AOI22_X1 U11594 ( .A1(keyinput_f66), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n9101) );
  OAI221_X1 U11595 ( .B1(keyinput_f66), .B2(P3_DATAO_REG_30__SCAN_IN), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n9101), .ZN(n9106) );
  AOI22_X1 U11596 ( .A1(keyinput_f33), .A2(P3_RD_REG_SCAN_IN), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f117), .ZN(n9102) );
  OAI221_X1 U11597 ( .B1(keyinput_f33), .B2(P3_RD_REG_SCAN_IN), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_f117), .A(n9102), .ZN(n9105) );
  AOI22_X1 U11598 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n9103) );
  OAI221_X1 U11599 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9103), .ZN(n9104) );
  NOR4_X1 U11600 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9108)
         );
  NAND4_X1 U11601 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n9241)
         );
  AOI22_X1 U11602 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n9112) );
  OAI221_X1 U11603 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n9112), .ZN(n9119) );
  AOI22_X1 U11604 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f119), .ZN(n9113) );
  OAI221_X1 U11605 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f119), .A(n9113), .ZN(n9118) );
  AOI22_X1 U11606 ( .A1(keyinput_f81), .A2(P3_DATAO_REG_15__SCAN_IN), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .ZN(n9114) );
  OAI221_X1 U11607 ( .B1(keyinput_f81), .B2(P3_DATAO_REG_15__SCAN_IN), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f123), .A(n9114), .ZN(n9117) );
  AOI22_X1 U11608 ( .A1(SI_21_), .A2(keyinput_f11), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n9115) );
  OAI221_X1 U11609 ( .B1(SI_21_), .B2(keyinput_f11), .C1(SI_23_), .C2(
        keyinput_f9), .A(n9115), .ZN(n9116) );
  NOR4_X1 U11610 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(n9147)
         );
  AOI22_X1 U11611 ( .A1(SI_17_), .A2(keyinput_f15), .B1(SI_22_), .B2(
        keyinput_f10), .ZN(n9120) );
  OAI221_X1 U11612 ( .B1(SI_17_), .B2(keyinput_f15), .C1(SI_22_), .C2(
        keyinput_f10), .A(n9120), .ZN(n9127) );
  AOI22_X1 U11613 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_f101), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_f111), .ZN(n9121) );
  OAI221_X1 U11614 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f111), .A(n9121), .ZN(n9126) );
  AOI22_X1 U11615 ( .A1(keyinput_f89), .A2(P3_DATAO_REG_7__SCAN_IN), .B1(
        P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_f98), .ZN(n9122) );
  OAI221_X1 U11616 ( .B1(keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .C1(
        P3_ADDR_REG_1__SCAN_IN), .C2(keyinput_f98), .A(n9122), .ZN(n9125) );
  AOI22_X1 U11617 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f114), .B1(SI_18_), 
        .B2(keyinput_f14), .ZN(n9123) );
  OAI221_X1 U11618 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f114), .C1(SI_18_), .C2(keyinput_f14), .A(n9123), .ZN(n9124) );
  NOR4_X1 U11619 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n9146)
         );
  AOI22_X1 U11620 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(SI_6_), 
        .B2(keyinput_f26), .ZN(n9128) );
  OAI221_X1 U11621 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(SI_6_), .C2(keyinput_f26), .A(n9128), .ZN(n9135) );
  AOI22_X1 U11622 ( .A1(keyinput_f83), .A2(P3_DATAO_REG_13__SCAN_IN), .B1(
        P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_f99), .ZN(n9129) );
  OAI221_X1 U11623 ( .B1(keyinput_f83), .B2(P3_DATAO_REG_13__SCAN_IN), .C1(
        P3_ADDR_REG_2__SCAN_IN), .C2(keyinput_f99), .A(n9129), .ZN(n9134) );
  AOI22_X1 U11624 ( .A1(keyinput_f80), .A2(P3_DATAO_REG_16__SCAN_IN), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9130) );
  OAI221_X1 U11625 ( .B1(keyinput_f80), .B2(P3_DATAO_REG_16__SCAN_IN), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9130), .ZN(n9133) );
  AOI22_X1 U11626 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(SI_20_), 
        .B2(keyinput_f12), .ZN(n9131) );
  OAI221_X1 U11627 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(SI_20_), .C2(keyinput_f12), .A(n9131), .ZN(n9132) );
  NOR4_X1 U11628 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n9145)
         );
  AOI22_X1 U11629 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_8_), .B2(
        keyinput_f24), .ZN(n9136) );
  OAI221_X1 U11630 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_8_), .C2(
        keyinput_f24), .A(n9136), .ZN(n9143) );
  AOI22_X1 U11631 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n9137) );
  OAI221_X1 U11632 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n9137), .ZN(n9142) );
  AOI22_X1 U11633 ( .A1(keyinput_f75), .A2(P3_DATAO_REG_21__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n9138) );
  OAI221_X1 U11634 ( .B1(keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n9138), .ZN(n9141) );
  AOI22_X1 U11635 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n9139) );
  OAI221_X1 U11636 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n9139), .ZN(n9140) );
  NOR4_X1 U11637 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), .ZN(n9144)
         );
  NAND4_X1 U11638 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(n9240)
         );
  AOI22_X1 U11639 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_f122), .B1(SI_25_), .B2(keyinput_f7), .ZN(n9148) );
  OAI221_X1 U11640 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_f122), .C1(
        SI_25_), .C2(keyinput_f7), .A(n9148), .ZN(n9149) );
  INV_X1 U11641 ( .A(n9149), .ZN(n9159) );
  AOI22_X1 U11642 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(keyinput_f97), .B1(SI_28_), .B2(keyinput_f4), .ZN(n9150) );
  OAI221_X1 U11643 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_f97), .C1(
        SI_28_), .C2(keyinput_f4), .A(n9150), .ZN(n9151) );
  INV_X1 U11644 ( .A(n9151), .ZN(n9158) );
  XNOR2_X1 U11645 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f109), .ZN(n9154) );
  XNOR2_X1 U11646 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f107), .ZN(n9153) );
  XNOR2_X1 U11647 ( .A(keyinput_f56), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n9152)
         );
  AND3_X1 U11648 ( .A1(n9154), .A2(n9153), .A3(n9152), .ZN(n9157) );
  INV_X1 U11649 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10390) );
  INV_X1 U11650 ( .A(keyinput_f94), .ZN(n9155) );
  XNOR2_X1 U11651 ( .A(n10390), .B(n9155), .ZN(n9156) );
  AND4_X1 U11652 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n9195)
         );
  AOI22_X1 U11653 ( .A1(n9162), .A2(keyinput_f62), .B1(keyinput_f104), .B2(
        n9161), .ZN(n9160) );
  OAI221_X1 U11654 ( .B1(n9162), .B2(keyinput_f62), .C1(n9161), .C2(
        keyinput_f104), .A(n9160), .ZN(n9171) );
  AOI22_X1 U11655 ( .A1(n10239), .A2(keyinput_f76), .B1(n9164), .B2(
        keyinput_f60), .ZN(n9163) );
  OAI221_X1 U11656 ( .B1(n10239), .B2(keyinput_f76), .C1(n9164), .C2(
        keyinput_f60), .A(n9163), .ZN(n9170) );
  INV_X1 U11657 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U11658 ( .A1(n11184), .A2(keyinput_f54), .B1(n11569), .B2(
        keyinput_f46), .ZN(n9165) );
  OAI221_X1 U11659 ( .B1(n11184), .B2(keyinput_f54), .C1(n11569), .C2(
        keyinput_f46), .A(n9165), .ZN(n9169) );
  XNOR2_X1 U11660 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f110), .ZN(n9167) );
  XNOR2_X1 U11661 ( .A(SI_3_), .B(keyinput_f29), .ZN(n9166) );
  NAND2_X1 U11662 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  NOR4_X1 U11663 ( .A1(n9171), .A2(n9170), .A3(n9169), .A4(n9168), .ZN(n9194)
         );
  INV_X1 U11664 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U11665 ( .A1(n10308), .A2(keyinput_f13), .B1(keyinput_f93), .B2(
        n10388), .ZN(n9172) );
  OAI221_X1 U11666 ( .B1(n10308), .B2(keyinput_f13), .C1(n10388), .C2(
        keyinput_f93), .A(n9172), .ZN(n9181) );
  INV_X1 U11667 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U11668 ( .A1(n9174), .A2(keyinput_f55), .B1(keyinput_f85), .B2(
        n10386), .ZN(n9173) );
  OAI221_X1 U11669 ( .B1(n9174), .B2(keyinput_f55), .C1(n10386), .C2(
        keyinput_f85), .A(n9173), .ZN(n9180) );
  INV_X1 U11670 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10314) );
  INV_X1 U11671 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U11672 ( .A1(n10314), .A2(keyinput_f120), .B1(keyinput_f90), .B2(
        n10231), .ZN(n9175) );
  OAI221_X1 U11673 ( .B1(n10314), .B2(keyinput_f120), .C1(n10231), .C2(
        keyinput_f90), .A(n9175), .ZN(n9179) );
  AOI22_X1 U11674 ( .A1(n10044), .A2(keyinput_f121), .B1(n9177), .B2(
        keyinput_f38), .ZN(n9176) );
  OAI221_X1 U11675 ( .B1(n10044), .B2(keyinput_f121), .C1(n9177), .C2(
        keyinput_f38), .A(n9176), .ZN(n9178) );
  NOR4_X1 U11676 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n9193)
         );
  INV_X1 U11677 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U11678 ( .A1(n9183), .A2(keyinput_f47), .B1(keyinput_f96), .B2(
        n10384), .ZN(n9182) );
  OAI221_X1 U11679 ( .B1(n9183), .B2(keyinput_f47), .C1(n10384), .C2(
        keyinput_f96), .A(n9182), .ZN(n9191) );
  AOI22_X1 U11680 ( .A1(n10162), .A2(keyinput_f116), .B1(keyinput_f74), .B2(
        n10237), .ZN(n9184) );
  OAI221_X1 U11681 ( .B1(n10162), .B2(keyinput_f116), .C1(n10237), .C2(
        keyinput_f74), .A(n9184), .ZN(n9190) );
  AOI22_X1 U11682 ( .A1(n10374), .A2(keyinput_f73), .B1(n7097), .B2(
        keyinput_f102), .ZN(n9185) );
  OAI221_X1 U11683 ( .B1(n10374), .B2(keyinput_f73), .C1(n7097), .C2(
        keyinput_f102), .A(n9185), .ZN(n9189) );
  XNOR2_X1 U11684 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_f39), .ZN(n9187)
         );
  XNOR2_X1 U11685 ( .A(SI_2_), .B(keyinput_f30), .ZN(n9186) );
  NAND2_X1 U11686 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  NOR4_X1 U11687 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n9192)
         );
  NAND4_X1 U11688 ( .A1(n9195), .A2(n9194), .A3(n9193), .A4(n9192), .ZN(n9239)
         );
  INV_X1 U11689 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U11690 ( .A1(n10884), .A2(keyinput_f65), .B1(keyinput_f70), .B2(
        n10667), .ZN(n9196) );
  OAI221_X1 U11691 ( .B1(n10884), .B2(keyinput_f65), .C1(n10667), .C2(
        keyinput_f70), .A(n9196), .ZN(n9200) );
  XNOR2_X1 U11692 ( .A(n10233), .B(keyinput_f87), .ZN(n9199) );
  XNOR2_X1 U11693 ( .A(n10074), .B(keyinput_f28), .ZN(n9198) );
  XOR2_X1 U11694 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f125), .Z(n9197) );
  OR4_X1 U11695 ( .A1(n9200), .A2(n9199), .A3(n9198), .A4(n9197), .ZN(n9204)
         );
  INV_X1 U11696 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11697 ( .A1(n10131), .A2(keyinput_f20), .B1(keyinput_f79), .B2(
        n10208), .ZN(n9201) );
  OAI221_X1 U11698 ( .B1(n10131), .B2(keyinput_f20), .C1(n10208), .C2(
        keyinput_f79), .A(n9201), .ZN(n9203) );
  INV_X1 U11699 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10183) );
  XNOR2_X1 U11700 ( .A(n10183), .B(keyinput_f91), .ZN(n9202) );
  NOR3_X1 U11701 ( .A1(n9204), .A2(n9203), .A3(n9202), .ZN(n9237) );
  AOI22_X1 U11702 ( .A1(n10114), .A2(keyinput_f22), .B1(keyinput_f17), .B2(
        n10161), .ZN(n9205) );
  OAI221_X1 U11703 ( .B1(n10114), .B2(keyinput_f22), .C1(n10161), .C2(
        keyinput_f17), .A(n9205), .ZN(n9208) );
  INV_X1 U11704 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n10858) );
  XNOR2_X1 U11705 ( .A(n10858), .B(keyinput_f67), .ZN(n9207) );
  XOR2_X1 U11706 ( .A(SI_7_), .B(keyinput_f25), .Z(n9206) );
  OR3_X1 U11707 ( .A1(n9208), .A2(n9207), .A3(n9206), .ZN(n9214) );
  INV_X1 U11708 ( .A(keyinput_f0), .ZN(n9210) );
  AOI22_X1 U11709 ( .A1(n10392), .A2(keyinput_f95), .B1(P3_WR_REG_SCAN_IN), 
        .B2(n9210), .ZN(n9209) );
  OAI221_X1 U11710 ( .B1(n10392), .B2(keyinput_f95), .C1(n9210), .C2(
        P3_WR_REG_SCAN_IN), .A(n9209), .ZN(n9213) );
  AOI22_X1 U11711 ( .A1(n10548), .A2(keyinput_f71), .B1(n11443), .B2(
        keyinput_f8), .ZN(n9211) );
  OAI221_X1 U11712 ( .B1(n10548), .B2(keyinput_f71), .C1(n11443), .C2(
        keyinput_f8), .A(n9211), .ZN(n9212) );
  NOR3_X1 U11713 ( .A1(n9214), .A2(n9213), .A3(n9212), .ZN(n9236) );
  INV_X1 U11714 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U11715 ( .A1(n10809), .A2(keyinput_f69), .B1(n12783), .B2(
        keyinput_f37), .ZN(n9215) );
  OAI221_X1 U11716 ( .B1(n10809), .B2(keyinput_f69), .C1(n12783), .C2(
        keyinput_f37), .A(n9215), .ZN(n9218) );
  XNOR2_X1 U11717 ( .A(n10418), .B(keyinput_f72), .ZN(n9217) );
  XOR2_X1 U11718 ( .A(SI_1_), .B(keyinput_f31), .Z(n9216) );
  OR3_X1 U11719 ( .A1(n9218), .A2(n9217), .A3(n9216), .ZN(n9223) );
  AOI22_X1 U11720 ( .A1(n10272), .A2(keyinput_f84), .B1(n8277), .B2(
        keyinput_f49), .ZN(n9219) );
  OAI221_X1 U11721 ( .B1(n10272), .B2(keyinput_f84), .C1(n8277), .C2(
        keyinput_f49), .A(n9219), .ZN(n9222) );
  INV_X1 U11722 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U11723 ( .A1(n13440), .A2(keyinput_f3), .B1(keyinput_f88), .B2(
        n10270), .ZN(n9220) );
  OAI221_X1 U11724 ( .B1(n13440), .B2(keyinput_f3), .C1(n10270), .C2(
        keyinput_f88), .A(n9220), .ZN(n9221) );
  NOR3_X1 U11725 ( .A1(n9223), .A2(n9222), .A3(n9221), .ZN(n9235) );
  AOI22_X1 U11726 ( .A1(n11317), .A2(keyinput_f61), .B1(keyinput_f16), .B2(
        n10171), .ZN(n9224) );
  OAI221_X1 U11727 ( .B1(n11317), .B2(keyinput_f61), .C1(n10171), .C2(
        keyinput_f16), .A(n9224), .ZN(n9233) );
  INV_X1 U11728 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U11729 ( .A1(n10229), .A2(keyinput_f86), .B1(n8217), .B2(
        keyinput_f42), .ZN(n9225) );
  OAI221_X1 U11730 ( .B1(n10229), .B2(keyinput_f86), .C1(n8217), .C2(
        keyinput_f42), .A(n9225), .ZN(n9232) );
  AOI22_X1 U11731 ( .A1(n15586), .A2(keyinput_f59), .B1(keyinput_f105), .B2(
        n9227), .ZN(n9226) );
  OAI221_X1 U11732 ( .B1(n15586), .B2(keyinput_f59), .C1(n9227), .C2(
        keyinput_f105), .A(n9226), .ZN(n9231) );
  INV_X1 U11733 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9229) );
  AOI22_X1 U11734 ( .A1(n9229), .A2(keyinput_f36), .B1(keyinput_f82), .B2(
        n10169), .ZN(n9228) );
  OAI221_X1 U11735 ( .B1(n9229), .B2(keyinput_f36), .C1(n10169), .C2(
        keyinput_f82), .A(n9228), .ZN(n9230) );
  NOR4_X1 U11736 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n9234)
         );
  NAND4_X1 U11737 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(n9238)
         );
  NOR4_X1 U11738 ( .A1(n9241), .A2(n9240), .A3(n9239), .A4(n9238), .ZN(n9243)
         );
  XOR2_X1 U11739 ( .A(keyinput_g115), .B(keyinput_f115), .Z(n9242) );
  NOR2_X1 U11740 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  AOI211_X1 U11741 ( .C1(n9247), .C2(n9246), .A(n9245), .B(n9244), .ZN(n9248)
         );
  XNOR2_X1 U11742 ( .A(n9249), .B(n9248), .ZN(n9250) );
  INV_X1 U11743 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U11744 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9302) );
  INV_X1 U11745 ( .A(n9302), .ZN(n9251) );
  NAND2_X1 U11746 ( .A1(n9251), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9311) );
  INV_X1 U11747 ( .A(n9311), .ZN(n9252) );
  NAND2_X1 U11748 ( .A1(n9252), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9319) );
  INV_X1 U11749 ( .A(n9319), .ZN(n9253) );
  NAND2_X1 U11750 ( .A1(n9253), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9329) );
  INV_X1 U11751 ( .A(n9329), .ZN(n9254) );
  NAND2_X1 U11752 ( .A1(n9254), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U11753 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n9255) );
  INV_X1 U11754 ( .A(n9352), .ZN(n9256) );
  NAND2_X1 U11755 ( .A1(n9256), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11756 ( .A1(n9257), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9378) );
  INV_X1 U11757 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9377) );
  INV_X1 U11758 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11759 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9258) );
  INV_X1 U11760 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13510) );
  INV_X1 U11761 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13477) );
  INV_X1 U11762 ( .A(n9459), .ZN(n9261) );
  NAND2_X1 U11763 ( .A1(n9261), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9461) );
  INV_X1 U11764 ( .A(n9461), .ZN(n9262) );
  NAND2_X1 U11765 ( .A1(n9262), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9470) );
  INV_X1 U11766 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U11767 ( .A1(n9461), .A2(n13529), .ZN(n9263) );
  NAND2_X1 U11768 ( .A1(n9470), .A2(n9263), .ZN(n13809) );
  AND2_X2 U11769 ( .A1(n9264), .A2(n14090), .ZN(n9279) );
  OR2_X1 U11770 ( .A1(n13809), .A2(n9472), .ZN(n9269) );
  INV_X1 U11771 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U11772 ( .A1(n9559), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11773 ( .A1(n9560), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9265) );
  OAI211_X1 U11774 ( .C1(n13808), .C2(n9563), .A(n9266), .B(n9265), .ZN(n9267)
         );
  INV_X1 U11775 ( .A(n9267), .ZN(n9268) );
  NAND2_X1 U11776 ( .A1(n9269), .A2(n9268), .ZN(n13650) );
  NAND2_X1 U11777 ( .A1(n9403), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11778 ( .A1(n9411), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11779 ( .A1(n9327), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11780 ( .A1(n9437), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11781 ( .A1(n9281), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11782 ( .A1(n9279), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11783 ( .A1(n9278), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11784 ( .A1(n9280), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11785 ( .A1(n9278), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11786 ( .A1(n9279), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11787 ( .A1(n9280), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11788 ( .A1(n9281), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9282) );
  INV_X1 U11789 ( .A(n12400), .ZN(n9992) );
  NAND2_X1 U11790 ( .A1(n9756), .A2(n9992), .ZN(n9991) );
  INV_X1 U11791 ( .A(n9991), .ZN(n11091) );
  INV_X1 U11792 ( .A(n13673), .ZN(n10409) );
  NAND2_X1 U11793 ( .A1(n10409), .A2(n10422), .ZN(n9286) );
  NAND2_X1 U11794 ( .A1(n9287), .A2(n9286), .ZN(n10733) );
  INV_X1 U11795 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11796 ( .A1(n9411), .A2(n9294), .ZN(n9291) );
  NAND2_X1 U11797 ( .A1(n9403), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11798 ( .A1(n9327), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U11799 ( .A1(n9437), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9288) );
  INV_X1 U11800 ( .A(n13672), .ZN(n10379) );
  NAND2_X1 U11801 ( .A1(n10379), .A2(n15379), .ZN(n9292) );
  NAND2_X1 U11802 ( .A1(n9403), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9299) );
  INV_X1 U11803 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11804 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  AND2_X1 U11805 ( .A1(n9295), .A2(n9302), .ZN(n11056) );
  NAND2_X1 U11806 ( .A1(n9411), .A2(n11056), .ZN(n9298) );
  NAND2_X1 U11807 ( .A1(n9327), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11808 ( .A1(n9437), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9296) );
  NAND4_X1 U11809 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n13671) );
  NAND2_X1 U11810 ( .A1(n6907), .A2(n10727), .ZN(n9300) );
  NAND2_X1 U11811 ( .A1(n9559), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11812 ( .A1(n9403), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9306) );
  INV_X1 U11813 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U11814 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  AND2_X1 U11815 ( .A1(n9311), .A2(n9303), .ZN(n10867) );
  NAND2_X1 U11816 ( .A1(n9496), .A2(n10867), .ZN(n9305) );
  NAND2_X1 U11817 ( .A1(n9420), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9304) );
  NAND4_X1 U11818 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n13670) );
  NOR2_X1 U11819 ( .A1(n13670), .A2(n9791), .ZN(n9309) );
  NAND2_X1 U11820 ( .A1(n13670), .A2(n9791), .ZN(n9308) );
  NAND2_X1 U11821 ( .A1(n9327), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U11822 ( .A1(n9560), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9315) );
  INV_X1 U11823 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11824 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  AND2_X1 U11825 ( .A1(n9319), .A2(n9312), .ZN(n11207) );
  NAND2_X1 U11826 ( .A1(n9496), .A2(n11207), .ZN(n9314) );
  NAND2_X1 U11827 ( .A1(n9420), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9313) );
  NAND4_X1 U11828 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n13669) );
  XNOR2_X1 U11829 ( .A(n13669), .B(n11208), .ZN(n11065) );
  INV_X1 U11830 ( .A(n11065), .ZN(n11069) );
  NAND2_X1 U11831 ( .A1(n13669), .A2(n11208), .ZN(n9317) );
  NAND2_X1 U11832 ( .A1(n9403), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9324) );
  INV_X1 U11833 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11834 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  AND2_X1 U11835 ( .A1(n9329), .A2(n9320), .ZN(n11409) );
  NAND2_X1 U11836 ( .A1(n9411), .A2(n11409), .ZN(n9323) );
  NAND2_X1 U11837 ( .A1(n9327), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11838 ( .A1(n9420), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9321) );
  NAND4_X1 U11839 ( .A1(n9324), .A2(n9323), .A3(n9322), .A4(n9321), .ZN(n13668) );
  INV_X1 U11840 ( .A(n13668), .ZN(n9521) );
  XNOR2_X1 U11841 ( .A(n9521), .B(n11418), .ZN(n11237) );
  NAND2_X1 U11842 ( .A1(n11233), .A2(n11237), .ZN(n9326) );
  NAND2_X1 U11843 ( .A1(n11418), .A2(n13668), .ZN(n9325) );
  NAND2_X1 U11844 ( .A1(n9326), .A2(n9325), .ZN(n11285) );
  NAND2_X1 U11845 ( .A1(n9327), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11846 ( .A1(n9403), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9333) );
  INV_X1 U11847 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11848 ( .A1(n9329), .A2(n9328), .ZN(n9330) );
  AND2_X1 U11849 ( .A1(n9345), .A2(n9330), .ZN(n13497) );
  NAND2_X1 U11850 ( .A1(n9496), .A2(n13497), .ZN(n9332) );
  NAND2_X1 U11851 ( .A1(n9420), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9331) );
  NAND4_X1 U11852 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n13667) );
  INV_X1 U11853 ( .A(n13667), .ZN(n9812) );
  NAND2_X1 U11854 ( .A1(n13498), .A2(n9812), .ZN(n9522) );
  OR2_X1 U11855 ( .A1(n13498), .A2(n9812), .ZN(n9335) );
  NAND2_X1 U11856 ( .A1(n11285), .A2(n11286), .ZN(n9337) );
  NAND2_X1 U11857 ( .A1(n13498), .A2(n13667), .ZN(n9336) );
  NAND2_X1 U11858 ( .A1(n9337), .A2(n9336), .ZN(n11428) );
  NAND2_X1 U11859 ( .A1(n9559), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11860 ( .A1(n9403), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9340) );
  XNOR2_X1 U11861 ( .A(n9345), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n11612) );
  NAND2_X1 U11862 ( .A1(n9411), .A2(n11612), .ZN(n9339) );
  NAND2_X1 U11863 ( .A1(n9420), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9338) );
  NAND4_X1 U11864 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n13666) );
  XNOR2_X1 U11865 ( .A(n15399), .B(n13666), .ZN(n9998) );
  NAND2_X1 U11866 ( .A1(n15399), .A2(n13666), .ZN(n9342) );
  NAND2_X1 U11867 ( .A1(n9559), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U11868 ( .A1(n9560), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9349) );
  INV_X1 U11869 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9344) );
  INV_X1 U11870 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9343) );
  OAI21_X1 U11871 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9346) );
  AND2_X1 U11872 ( .A1(n9346), .A2(n9352), .ZN(n11626) );
  NAND2_X1 U11873 ( .A1(n9496), .A2(n11626), .ZN(n9348) );
  NAND2_X1 U11874 ( .A1(n9437), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9347) );
  NAND4_X1 U11875 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n13665) );
  XNOR2_X1 U11876 ( .A(n11737), .B(n13665), .ZN(n11518) );
  NAND2_X1 U11877 ( .A1(n11737), .A2(n13665), .ZN(n9351) );
  NAND2_X1 U11878 ( .A1(n9559), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11879 ( .A1(n9560), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9356) );
  INV_X1 U11880 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U11881 ( .A1(n9352), .A2(n13600), .ZN(n9353) );
  AND2_X1 U11882 ( .A1(n9362), .A2(n9353), .ZN(n13599) );
  NAND2_X1 U11883 ( .A1(n9496), .A2(n13599), .ZN(n9355) );
  NAND2_X1 U11884 ( .A1(n9420), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9354) );
  NAND4_X1 U11885 ( .A1(n9357), .A2(n9356), .A3(n9355), .A4(n9354), .ZN(n13664) );
  AND2_X1 U11886 ( .A1(n11607), .A2(n13664), .ZN(n9358) );
  OR2_X1 U11887 ( .A1(n11607), .A2(n13664), .ZN(n9359) );
  NAND2_X1 U11888 ( .A1(n9559), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11889 ( .A1(n9403), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U11890 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  AND2_X1 U11891 ( .A1(n9370), .A2(n9363), .ZN(n13518) );
  NAND2_X1 U11892 ( .A1(n9496), .A2(n13518), .ZN(n9365) );
  NAND2_X1 U11893 ( .A1(n9437), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9364) );
  NAND4_X1 U11894 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n13663) );
  NOR2_X1 U11895 ( .A1(n11795), .A2(n13663), .ZN(n9368) );
  NAND2_X1 U11896 ( .A1(n9560), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9375) );
  INV_X1 U11897 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11898 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  AND2_X1 U11899 ( .A1(n9378), .A2(n9371), .ZN(n13580) );
  NAND2_X1 U11900 ( .A1(n9411), .A2(n13580), .ZN(n9374) );
  NAND2_X1 U11901 ( .A1(n9559), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11902 ( .A1(n9420), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9372) );
  NAND4_X1 U11903 ( .A1(n9375), .A2(n9374), .A3(n9373), .A4(n9372), .ZN(n13662) );
  AND2_X1 U11904 ( .A1(n11823), .A2(n13662), .ZN(n9376) );
  NAND2_X1 U11905 ( .A1(n9559), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11906 ( .A1(n9403), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11907 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  AND2_X1 U11908 ( .A1(n9386), .A2(n9379), .ZN(n14884) );
  NAND2_X1 U11909 ( .A1(n9496), .A2(n14884), .ZN(n9381) );
  NAND2_X1 U11910 ( .A1(n9420), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9380) );
  NAND4_X1 U11911 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9380), .ZN(n13661) );
  XNOR2_X1 U11912 ( .A(n14889), .B(n13661), .ZN(n14888) );
  NAND2_X1 U11913 ( .A1(n14889), .A2(n13661), .ZN(n9384) );
  NAND2_X1 U11914 ( .A1(n9559), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U11915 ( .A1(n9403), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11916 ( .A1(n9386), .A2(n9385), .ZN(n9387) );
  AND2_X1 U11917 ( .A1(n9394), .A2(n9387), .ZN(n13636) );
  NAND2_X1 U11918 ( .A1(n9411), .A2(n13636), .ZN(n9389) );
  NAND2_X1 U11919 ( .A1(n9420), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9388) );
  NAND4_X1 U11920 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n13660) );
  XNOR2_X1 U11921 ( .A(n11993), .B(n13660), .ZN(n11989) );
  OR2_X1 U11922 ( .A1(n11993), .A2(n13660), .ZN(n9392) );
  NAND2_X1 U11923 ( .A1(n9559), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U11924 ( .A1(n9560), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9398) );
  INV_X1 U11925 ( .A(n9393), .ZN(n9404) );
  NAND2_X1 U11926 ( .A1(n9394), .A2(n13540), .ZN(n9395) );
  AND2_X1 U11927 ( .A1(n9404), .A2(n9395), .ZN(n13539) );
  NAND2_X1 U11928 ( .A1(n9496), .A2(n13539), .ZN(n9397) );
  NAND2_X1 U11929 ( .A1(n9420), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9396) );
  NAND4_X1 U11930 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n13659) );
  INV_X1 U11931 ( .A(n13659), .ZN(n9400) );
  OR2_X1 U11932 ( .A1(n13959), .A2(n9400), .ZN(n9536) );
  NAND2_X1 U11933 ( .A1(n13959), .A2(n9400), .ZN(n9401) );
  NAND2_X1 U11934 ( .A1(n9536), .A2(n9401), .ZN(n13947) );
  INV_X1 U11935 ( .A(n13947), .ZN(n13942) );
  NAND2_X1 U11936 ( .A1(n13959), .A2(n13659), .ZN(n9402) );
  NAND2_X1 U11937 ( .A1(n9559), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U11938 ( .A1(n9403), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9408) );
  INV_X1 U11939 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U11940 ( .A1(n9404), .A2(n15297), .ZN(n9405) );
  AND2_X1 U11941 ( .A1(n9418), .A2(n9405), .ZN(n13935) );
  NAND2_X1 U11942 ( .A1(n9411), .A2(n13935), .ZN(n9407) );
  NAND2_X1 U11943 ( .A1(n9420), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9406) );
  NAND4_X1 U11944 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n13658) );
  INV_X1 U11945 ( .A(n13658), .ZN(n9872) );
  XNOR2_X1 U11946 ( .A(n13936), .B(n9872), .ZN(n13931) );
  NAND2_X1 U11947 ( .A1(n13936), .A2(n13658), .ZN(n9410) );
  NAND2_X1 U11948 ( .A1(n9559), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9415) );
  XNOR2_X1 U11949 ( .A(n9418), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U11950 ( .A1(n13916), .A2(n9411), .ZN(n9414) );
  NAND2_X1 U11951 ( .A1(n9560), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11952 ( .A1(n9437), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9412) );
  NAND4_X1 U11953 ( .A1(n9415), .A2(n9414), .A3(n9413), .A4(n9412), .ZN(n13657) );
  XNOR2_X1 U11954 ( .A(n14031), .B(n13657), .ZN(n13923) );
  OR2_X1 U11955 ( .A1(n14031), .A2(n13657), .ZN(n9416) );
  INV_X1 U11956 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13613) );
  INV_X1 U11957 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9417) );
  OAI21_X1 U11958 ( .B1(n9418), .B2(n13613), .A(n9417), .ZN(n9419) );
  AND2_X1 U11959 ( .A1(n9419), .A2(n9427), .ZN(n13487) );
  NAND2_X1 U11960 ( .A1(n13487), .A2(n9496), .ZN(n9424) );
  NAND2_X1 U11961 ( .A1(n9559), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11962 ( .A1(n9560), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11963 ( .A1(n9420), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9421) );
  NAND4_X1 U11964 ( .A1(n9424), .A2(n9423), .A3(n9422), .A4(n9421), .ZN(n13656) );
  NOR2_X1 U11965 ( .A1(n13907), .A2(n13656), .ZN(n9425) );
  INV_X1 U11966 ( .A(n13656), .ZN(n9987) );
  INV_X1 U11967 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9431) );
  INV_X1 U11968 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11969 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U11970 ( .A1(n9435), .A2(n9428), .ZN(n13891) );
  OR2_X1 U11971 ( .A1(n13891), .A2(n9472), .ZN(n9430) );
  AOI22_X1 U11972 ( .A1(n9559), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n9560), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n9429) );
  OAI211_X1 U11973 ( .C1(n9563), .C2(n9431), .A(n9430), .B(n9429), .ZN(n13655)
         );
  OR2_X1 U11974 ( .A1(n14022), .A2(n13655), .ZN(n9432) );
  NAND2_X1 U11975 ( .A1(n14022), .A2(n13655), .ZN(n9433) );
  NAND2_X1 U11976 ( .A1(n9435), .A2(n13510), .ZN(n9436) );
  NAND2_X1 U11977 ( .A1(n9441), .A2(n9436), .ZN(n13875) );
  AOI22_X1 U11978 ( .A1(n9559), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n9560), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11979 ( .A1(n9437), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9438) );
  OAI211_X1 U11980 ( .C1(n13875), .C2(n9472), .A(n9439), .B(n9438), .ZN(n13654) );
  INV_X1 U11981 ( .A(n13654), .ZN(n9547) );
  XNOR2_X1 U11982 ( .A(n13877), .B(n9547), .ZN(n10004) );
  INV_X1 U11983 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11984 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  NAND2_X1 U11985 ( .A1(n9450), .A2(n9442), .ZN(n13858) );
  OR2_X1 U11986 ( .A1(n13858), .A2(n9472), .ZN(n9448) );
  INV_X1 U11987 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11988 ( .A1(n9559), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11989 ( .A1(n9560), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9443) );
  OAI211_X1 U11990 ( .C1(n9445), .C2(n9563), .A(n9444), .B(n9443), .ZN(n9446)
         );
  INV_X1 U11991 ( .A(n9446), .ZN(n9447) );
  NAND2_X1 U11992 ( .A1(n9448), .A2(n9447), .ZN(n13653) );
  INV_X1 U11993 ( .A(n13653), .ZN(n9550) );
  NAND2_X1 U11994 ( .A1(n14010), .A2(n13653), .ZN(n9449) );
  NAND2_X1 U11995 ( .A1(n9450), .A2(n13477), .ZN(n9451) );
  AND2_X1 U11996 ( .A1(n9459), .A2(n9451), .ZN(n13476) );
  NAND2_X1 U11997 ( .A1(n13476), .A2(n9496), .ZN(n9457) );
  INV_X1 U11998 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U11999 ( .A1(n9559), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U12000 ( .A1(n9560), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9452) );
  OAI211_X1 U12001 ( .C1(n9454), .C2(n9563), .A(n9453), .B(n9452), .ZN(n9455)
         );
  INV_X1 U12002 ( .A(n9455), .ZN(n9456) );
  NAND2_X1 U12003 ( .A1(n9457), .A2(n9456), .ZN(n13652) );
  INV_X1 U12004 ( .A(n13652), .ZN(n9697) );
  XNOR2_X1 U12005 ( .A(n13842), .B(n9697), .ZN(n13835) );
  INV_X1 U12006 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U12007 ( .A1(n9459), .A2(n9458), .ZN(n9460) );
  NAND2_X1 U12008 ( .A1(n9461), .A2(n9460), .ZN(n13565) );
  OR2_X1 U12009 ( .A1(n13565), .A2(n9472), .ZN(n9467) );
  INV_X1 U12010 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U12011 ( .A1(n9559), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U12012 ( .A1(n9560), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U12013 ( .C1(n9464), .C2(n9563), .A(n9463), .B(n9462), .ZN(n9465)
         );
  INV_X1 U12014 ( .A(n9465), .ZN(n9466) );
  NAND2_X1 U12015 ( .A1(n9467), .A2(n9466), .ZN(n13651) );
  INV_X1 U12016 ( .A(n13651), .ZN(n9928) );
  NAND2_X1 U12017 ( .A1(n13996), .A2(n9928), .ZN(n13798) );
  OR2_X1 U12018 ( .A1(n13996), .A2(n9928), .ZN(n9468) );
  NAND2_X1 U12019 ( .A1(n13798), .A2(n9468), .ZN(n13823) );
  NAND2_X1 U12020 ( .A1(n13996), .A2(n13651), .ZN(n9469) );
  XNOR2_X1 U12021 ( .A(n13811), .B(n9932), .ZN(n13799) );
  INV_X1 U12022 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U12023 ( .A1(n9470), .A2(n13625), .ZN(n9471) );
  NAND2_X1 U12024 ( .A1(n9480), .A2(n9471), .ZN(n13789) );
  INV_X1 U12025 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U12026 ( .A1(n9559), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U12027 ( .A1(n9560), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9473) );
  OAI211_X1 U12028 ( .C1(n13788), .C2(n9563), .A(n9474), .B(n9473), .ZN(n9475)
         );
  INV_X1 U12029 ( .A(n9475), .ZN(n9476) );
  INV_X1 U12030 ( .A(n13986), .ZN(n13787) );
  NAND2_X1 U12031 ( .A1(n13787), .A2(n13448), .ZN(n9478) );
  INV_X1 U12032 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13451) );
  INV_X1 U12033 ( .A(n13745), .ZN(n9488) );
  NAND2_X1 U12034 ( .A1(n9480), .A2(n13451), .ZN(n9481) );
  NAND2_X1 U12035 ( .A1(n13779), .A2(n9496), .ZN(n9487) );
  INV_X1 U12036 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U12037 ( .A1(n9559), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U12038 ( .A1(n9560), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9482) );
  OAI211_X1 U12039 ( .C1(n9484), .C2(n9563), .A(n9483), .B(n9482), .ZN(n9485)
         );
  INV_X1 U12040 ( .A(n9485), .ZN(n9486) );
  XNOR2_X1 U12041 ( .A(n13980), .B(n13648), .ZN(n13770) );
  INV_X1 U12042 ( .A(n13770), .ZN(n13774) );
  INV_X1 U12043 ( .A(n13980), .ZN(n13456) );
  INV_X1 U12044 ( .A(n13648), .ZN(n9555) );
  XNOR2_X1 U12045 ( .A(n9488), .B(P2_REG3_REG_28__SCAN_IN), .ZN(n13760) );
  INV_X1 U12046 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U12047 ( .A1(n9559), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U12048 ( .A1(n9560), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9489) );
  OAI211_X1 U12049 ( .C1(n9491), .C2(n9563), .A(n9490), .B(n9489), .ZN(n9492)
         );
  NAND2_X1 U12050 ( .A1(n9955), .A2(n13450), .ZN(n9493) );
  NAND2_X1 U12051 ( .A1(n9955), .A2(n9494), .ZN(n9495) );
  NAND3_X1 U12052 ( .A1(n13745), .A2(n9496), .A3(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9502) );
  INV_X1 U12053 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U12054 ( .A1(n9559), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U12055 ( .A1(n9560), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9497) );
  OAI211_X1 U12056 ( .C1(n9499), .C2(n9563), .A(n9498), .B(n9497), .ZN(n9500)
         );
  INV_X1 U12057 ( .A(n9500), .ZN(n9501) );
  AND2_X1 U12058 ( .A1(n9502), .A2(n9501), .ZN(n9956) );
  XNOR2_X1 U12059 ( .A(n9574), .B(n13647), .ZN(n10010) );
  XNOR2_X1 U12060 ( .A(n9578), .B(n6685), .ZN(n9503) );
  OR2_X1 U12061 ( .A1(n9754), .A2(n9751), .ZN(n15401) );
  INV_X1 U12062 ( .A(n13759), .ZN(n9504) );
  AOI211_X1 U12063 ( .C1(n9574), .C2(n9504), .A(n14001), .B(n13738), .ZN(
        n13750) );
  INV_X1 U12064 ( .A(n9756), .ZN(n9505) );
  INV_X1 U12065 ( .A(n9577), .ZN(n11088) );
  NAND2_X1 U12066 ( .A1(n11088), .A2(n11092), .ZN(n9507) );
  INV_X1 U12067 ( .A(n13674), .ZN(n10380) );
  NAND2_X1 U12068 ( .A1(n10380), .A2(n11094), .ZN(n9506) );
  NAND2_X1 U12069 ( .A1(n9507), .A2(n9506), .ZN(n10423) );
  NAND2_X1 U12070 ( .A1(n10423), .A2(n10424), .ZN(n9509) );
  NAND2_X1 U12071 ( .A1(n10409), .A2(n15315), .ZN(n9508) );
  NAND2_X1 U12072 ( .A1(n9509), .A2(n9508), .ZN(n10734) );
  INV_X1 U12073 ( .A(n9994), .ZN(n10735) );
  NAND2_X1 U12074 ( .A1(n10734), .A2(n10735), .ZN(n9511) );
  NAND2_X1 U12075 ( .A1(n10379), .A2(n10742), .ZN(n9510) );
  NAND2_X1 U12076 ( .A1(n9511), .A2(n9510), .ZN(n10719) );
  INV_X1 U12077 ( .A(n10720), .ZN(n9512) );
  NAND2_X1 U12078 ( .A1(n10719), .A2(n9512), .ZN(n9514) );
  NAND2_X1 U12079 ( .A1(n6907), .A2(n11057), .ZN(n9513) );
  NAND2_X1 U12080 ( .A1(n9514), .A2(n9513), .ZN(n10835) );
  XNOR2_X1 U12081 ( .A(n13670), .B(n9791), .ZN(n10836) );
  NAND2_X1 U12082 ( .A1(n10835), .A2(n10836), .ZN(n9517) );
  INV_X1 U12083 ( .A(n13670), .ZN(n9515) );
  NAND2_X1 U12084 ( .A1(n9515), .A2(n9791), .ZN(n9516) );
  NAND2_X1 U12085 ( .A1(n9517), .A2(n9516), .ZN(n11068) );
  NAND2_X1 U12086 ( .A1(n11068), .A2(n11065), .ZN(n9520) );
  INV_X1 U12087 ( .A(n13669), .ZN(n9518) );
  NAND2_X1 U12088 ( .A1(n9518), .A2(n11208), .ZN(n9519) );
  NAND2_X1 U12089 ( .A1(n9520), .A2(n9519), .ZN(n11236) );
  INV_X1 U12090 ( .A(n13666), .ZN(n11514) );
  OR2_X1 U12091 ( .A1(n15399), .A2(n11514), .ZN(n9523) );
  NAND2_X1 U12092 ( .A1(n15399), .A2(n11514), .ZN(n9524) );
  INV_X1 U12093 ( .A(n13665), .ZN(n9827) );
  NAND2_X1 U12094 ( .A1(n11737), .A2(n9827), .ZN(n9526) );
  XNOR2_X1 U12095 ( .A(n11607), .B(n13664), .ZN(n11603) );
  INV_X1 U12096 ( .A(n13664), .ZN(n11513) );
  NAND2_X1 U12097 ( .A1(n11607), .A2(n11513), .ZN(n9527) );
  AND2_X1 U12098 ( .A1(n11795), .A2(n9989), .ZN(n9529) );
  INV_X1 U12099 ( .A(n13662), .ZN(n9990) );
  NOR2_X1 U12100 ( .A1(n11823), .A2(n9990), .ZN(n9531) );
  NAND2_X1 U12101 ( .A1(n11823), .A2(n9990), .ZN(n9530) );
  INV_X1 U12102 ( .A(n11983), .ZN(n9532) );
  INV_X1 U12103 ( .A(n13660), .ZN(n9533) );
  NAND2_X1 U12104 ( .A1(n11993), .A2(n9533), .ZN(n9534) );
  NAND2_X1 U12105 ( .A1(n9535), .A2(n9534), .ZN(n13948) );
  INV_X1 U12106 ( .A(n13657), .ZN(n9887) );
  AND2_X1 U12107 ( .A1(n14031), .A2(n9887), .ZN(n9537) );
  OR2_X1 U12108 ( .A1(n13912), .A2(n9537), .ZN(n9539) );
  OR2_X1 U12109 ( .A1(n14031), .A2(n9887), .ZN(n9538) );
  NAND2_X1 U12110 ( .A1(n9539), .A2(n9538), .ZN(n13900) );
  NAND2_X1 U12111 ( .A1(n13907), .A2(n9987), .ZN(n9540) );
  NAND2_X1 U12112 ( .A1(n13900), .A2(n9540), .ZN(n9542) );
  OR2_X1 U12113 ( .A1(n13907), .A2(n9987), .ZN(n9541) );
  NAND2_X1 U12114 ( .A1(n9542), .A2(n9541), .ZN(n13866) );
  INV_X1 U12115 ( .A(n13655), .ZN(n9543) );
  NAND2_X1 U12116 ( .A1(n14022), .A2(n9543), .ZN(n13867) );
  NAND2_X1 U12117 ( .A1(n13866), .A2(n13867), .ZN(n9544) );
  OR2_X1 U12118 ( .A1(n14022), .A2(n9543), .ZN(n9988) );
  NAND2_X1 U12119 ( .A1(n9544), .A2(n9988), .ZN(n9546) );
  NAND2_X1 U12120 ( .A1(n13877), .A2(n9547), .ZN(n9545) );
  NAND2_X1 U12121 ( .A1(n9546), .A2(n9545), .ZN(n9549) );
  OR2_X1 U12122 ( .A1(n13877), .A2(n9547), .ZN(n9548) );
  NAND2_X1 U12123 ( .A1(n14010), .A2(n9550), .ZN(n9551) );
  INV_X1 U12124 ( .A(n9551), .ZN(n9552) );
  INV_X1 U12125 ( .A(n13835), .ZN(n13837) );
  NOR2_X1 U12126 ( .A1(n13842), .A2(n9697), .ZN(n13816) );
  NOR2_X1 U12127 ( .A1(n13823), .A2(n13816), .ZN(n9553) );
  OR2_X1 U12128 ( .A1(n13986), .A2(n13448), .ZN(n10007) );
  INV_X1 U12129 ( .A(n10007), .ZN(n9554) );
  NAND2_X1 U12130 ( .A1(n13986), .A2(n13448), .ZN(n10006) );
  INV_X1 U12131 ( .A(n13756), .ZN(n13764) );
  NAND2_X1 U12132 ( .A1(n10014), .A2(n9993), .ZN(n9558) );
  NAND2_X1 U12133 ( .A1(n9754), .A2(n10739), .ZN(n9557) );
  INV_X1 U12134 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U12135 ( .A1(n9559), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U12136 ( .A1(n9560), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9561) );
  OAI211_X1 U12137 ( .C1(n9563), .C2(n13739), .A(n9562), .B(n9561), .ZN(n13646) );
  INV_X1 U12138 ( .A(n13646), .ZN(n9564) );
  OAI22_X1 U12139 ( .A1(n13450), .A2(n13447), .B1(n9565), .B2(n9564), .ZN(
        n9566) );
  INV_X1 U12140 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U12141 ( .A1(n9574), .A2(n9569), .ZN(n9570) );
  INV_X1 U12142 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9572) );
  INV_X1 U12143 ( .A(n14081), .ZN(n9573) );
  NAND2_X1 U12144 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  NAND2_X1 U12145 ( .A1(n6681), .A2(n13674), .ZN(n9582) );
  NAND2_X1 U12146 ( .A1(n10241), .A2(n10242), .ZN(n10240) );
  INV_X1 U12147 ( .A(n9581), .ZN(n9583) );
  NAND2_X1 U12148 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  INV_X1 U12149 ( .A(n9589), .ZN(n9587) );
  NAND2_X1 U12150 ( .A1(n6681), .A2(n13673), .ZN(n9588) );
  INV_X1 U12151 ( .A(n9588), .ZN(n9586) );
  NAND2_X1 U12152 ( .A1(n9587), .A2(n9586), .ZN(n9590) );
  NAND2_X1 U12153 ( .A1(n9589), .A2(n9588), .ZN(n9591) );
  INV_X1 U12154 ( .A(n10408), .ZN(n9593) );
  NAND2_X1 U12155 ( .A1(n6681), .A2(n13672), .ZN(n9595) );
  XNOR2_X1 U12156 ( .A(n9594), .B(n9595), .ZN(n10407) );
  INV_X1 U12157 ( .A(n10407), .ZN(n9592) );
  INV_X1 U12158 ( .A(n9594), .ZN(n9597) );
  INV_X1 U12159 ( .A(n9595), .ZN(n9596) );
  NAND2_X1 U12160 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  NAND2_X1 U12161 ( .A1(n6681), .A2(n13671), .ZN(n9600) );
  NAND2_X1 U12162 ( .A1(n9599), .A2(n9600), .ZN(n9604) );
  INV_X1 U12163 ( .A(n9599), .ZN(n9602) );
  INV_X1 U12164 ( .A(n9600), .ZN(n9601) );
  NAND2_X1 U12165 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NAND2_X1 U12166 ( .A1(n9604), .A2(n9603), .ZN(n10707) );
  INV_X1 U12167 ( .A(n9791), .ZN(n15386) );
  NAND2_X1 U12168 ( .A1(n6681), .A2(n13670), .ZN(n9606) );
  NAND2_X1 U12169 ( .A1(n9605), .A2(n9606), .ZN(n9610) );
  INV_X1 U12170 ( .A(n9605), .ZN(n9608) );
  INV_X1 U12171 ( .A(n9606), .ZN(n9607) );
  NAND2_X1 U12172 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  AND2_X1 U12173 ( .A1(n9610), .A2(n9609), .ZN(n10866) );
  INV_X1 U12174 ( .A(n11208), .ZN(n11076) );
  NAND2_X1 U12175 ( .A1(n6681), .A2(n13669), .ZN(n9612) );
  XNOR2_X1 U12176 ( .A(n9611), .B(n9612), .ZN(n11200) );
  INV_X1 U12177 ( .A(n9611), .ZN(n9614) );
  INV_X1 U12178 ( .A(n9612), .ZN(n9613) );
  NAND2_X1 U12179 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  NAND2_X1 U12180 ( .A1(n6681), .A2(n13668), .ZN(n9616) );
  XNOR2_X1 U12181 ( .A(n9618), .B(n9616), .ZN(n11413) );
  INV_X1 U12182 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12183 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AND2_X1 U12184 ( .A1(n6681), .A2(n13667), .ZN(n9620) );
  OR2_X1 U12185 ( .A1(n9621), .A2(n9620), .ZN(n13493) );
  NAND2_X1 U12186 ( .A1(n9621), .A2(n9620), .ZN(n13492) );
  XNOR2_X1 U12187 ( .A(n15399), .B(n9729), .ZN(n9624) );
  NAND2_X1 U12188 ( .A1(n6681), .A2(n13666), .ZN(n9623) );
  XNOR2_X1 U12189 ( .A(n9624), .B(n9623), .ZN(n11616) );
  INV_X1 U12190 ( .A(n11616), .ZN(n9622) );
  NAND2_X1 U12191 ( .A1(n9624), .A2(n9623), .ZN(n9625) );
  AND2_X1 U12192 ( .A1(n6681), .A2(n13665), .ZN(n9627) );
  NAND2_X1 U12193 ( .A1(n9626), .A2(n9627), .ZN(n9632) );
  INV_X1 U12194 ( .A(n9626), .ZN(n9629) );
  INV_X1 U12195 ( .A(n9627), .ZN(n9628) );
  NAND2_X1 U12196 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  NAND2_X1 U12197 ( .A1(n9632), .A2(n9630), .ZN(n11622) );
  AND2_X1 U12198 ( .A1(n6681), .A2(n13664), .ZN(n9634) );
  NAND2_X1 U12199 ( .A1(n9633), .A2(n9634), .ZN(n9638) );
  INV_X1 U12200 ( .A(n9633), .ZN(n9636) );
  INV_X1 U12201 ( .A(n9634), .ZN(n9635) );
  NAND2_X1 U12202 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  AND2_X1 U12203 ( .A1(n9638), .A2(n9637), .ZN(n13597) );
  NAND2_X1 U12204 ( .A1(n6681), .A2(n13663), .ZN(n9640) );
  XNOR2_X1 U12205 ( .A(n9639), .B(n9640), .ZN(n13515) );
  INV_X1 U12206 ( .A(n9639), .ZN(n9641) );
  NAND2_X1 U12207 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  AND2_X1 U12208 ( .A1(n6681), .A2(n13662), .ZN(n9644) );
  NAND2_X1 U12209 ( .A1(n9643), .A2(n9644), .ZN(n9659) );
  INV_X1 U12210 ( .A(n9643), .ZN(n9646) );
  INV_X1 U12211 ( .A(n9644), .ZN(n9645) );
  NAND2_X1 U12212 ( .A1(n9646), .A2(n9645), .ZN(n9647) );
  AND2_X1 U12213 ( .A1(n6681), .A2(n13661), .ZN(n9651) );
  INV_X1 U12214 ( .A(n9659), .ZN(n9648) );
  AOI21_X1 U12215 ( .B1(n9650), .B2(n9651), .A(n9648), .ZN(n9649) );
  INV_X1 U12216 ( .A(n9656), .ZN(n9652) );
  INV_X1 U12217 ( .A(n9650), .ZN(n9661) );
  NAND2_X1 U12218 ( .A1(n9661), .A2(n9660), .ZN(n9655) );
  NAND2_X1 U12219 ( .A1(n9652), .A2(n9655), .ZN(n9653) );
  AND2_X1 U12220 ( .A1(n9659), .A2(n9660), .ZN(n9654) );
  OAI22_X1 U12221 ( .A1(n9661), .A2(n9654), .B1(n9659), .B2(n9660), .ZN(n9657)
         );
  NAND2_X1 U12222 ( .A1(n9656), .A2(n9655), .ZN(n9664) );
  OAI21_X1 U12223 ( .B1(n9657), .B2(n9656), .A(n9664), .ZN(n9658) );
  AND2_X1 U12224 ( .A1(n6681), .A2(n13660), .ZN(n13634) );
  NAND2_X1 U12225 ( .A1(n13577), .A2(n9659), .ZN(n13459) );
  INV_X1 U12226 ( .A(n13459), .ZN(n9663) );
  XNOR2_X1 U12227 ( .A(n9661), .B(n9660), .ZN(n13460) );
  INV_X1 U12228 ( .A(n13460), .ZN(n9662) );
  NAND2_X1 U12229 ( .A1(n9663), .A2(n9662), .ZN(n13457) );
  INV_X1 U12230 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U12231 ( .A1(n13457), .A2(n9665), .ZN(n9666) );
  NAND2_X1 U12232 ( .A1(n6681), .A2(n13659), .ZN(n9668) );
  XNOR2_X1 U12233 ( .A(n9667), .B(n9668), .ZN(n13534) );
  INV_X1 U12234 ( .A(n9667), .ZN(n9669) );
  NAND2_X1 U12235 ( .A1(n9669), .A2(n9668), .ZN(n13544) );
  NAND2_X1 U12236 ( .A1(n13533), .A2(n13544), .ZN(n9670) );
  NAND2_X1 U12237 ( .A1(n6681), .A2(n13658), .ZN(n9672) );
  XNOR2_X1 U12238 ( .A(n9671), .B(n9672), .ZN(n13545) );
  INV_X1 U12239 ( .A(n9671), .ZN(n9673) );
  NAND2_X1 U12240 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  AND2_X1 U12241 ( .A1(n6681), .A2(n13657), .ZN(n9676) );
  NAND2_X1 U12242 ( .A1(n9675), .A2(n9676), .ZN(n9681) );
  INV_X1 U12243 ( .A(n9675), .ZN(n9678) );
  INV_X1 U12244 ( .A(n9676), .ZN(n9677) );
  NAND2_X1 U12245 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  NAND2_X1 U12246 ( .A1(n9681), .A2(n9679), .ZN(n13606) );
  INV_X1 U12247 ( .A(n13606), .ZN(n9680) );
  NAND2_X1 U12248 ( .A1(n6681), .A2(n13656), .ZN(n9683) );
  XNOR2_X1 U12249 ( .A(n9682), .B(n9683), .ZN(n13482) );
  INV_X1 U12250 ( .A(n9682), .ZN(n9684) );
  NAND2_X1 U12251 ( .A1(n9684), .A2(n9683), .ZN(n9685) );
  NAND2_X1 U12252 ( .A1(n6681), .A2(n13655), .ZN(n9687) );
  XNOR2_X1 U12253 ( .A(n9686), .B(n9687), .ZN(n13570) );
  INV_X1 U12254 ( .A(n9686), .ZN(n9688) );
  NAND2_X1 U12255 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  XNOR2_X1 U12256 ( .A(n13877), .B(n9729), .ZN(n9692) );
  NAND2_X1 U12257 ( .A1(n13654), .A2(n6681), .ZN(n9693) );
  XNOR2_X1 U12258 ( .A(n9692), .B(n9693), .ZN(n13505) );
  INV_X1 U12259 ( .A(n13505), .ZN(n9691) );
  INV_X1 U12260 ( .A(n9692), .ZN(n9695) );
  INV_X1 U12261 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U12262 ( .A1(n9695), .A2(n9694), .ZN(n9696) );
  XNOR2_X1 U12263 ( .A(n14010), .B(n9729), .ZN(n9699) );
  XNOR2_X1 U12264 ( .A(n13842), .B(n9729), .ZN(n13469) );
  NAND2_X1 U12265 ( .A1(n13653), .A2(n6681), .ZN(n13591) );
  AOI21_X1 U12266 ( .B1(n13469), .B2(n9697), .A(n13591), .ZN(n9698) );
  NAND2_X1 U12267 ( .A1(n13467), .A2(n9698), .ZN(n9707) );
  INV_X1 U12268 ( .A(n9699), .ZN(n9700) );
  AND2_X1 U12269 ( .A1(n13652), .A2(n6681), .ZN(n9702) );
  INV_X1 U12270 ( .A(n9702), .ZN(n13473) );
  NAND2_X1 U12271 ( .A1(n13469), .A2(n13473), .ZN(n9705) );
  INV_X1 U12272 ( .A(n13469), .ZN(n9703) );
  AND2_X1 U12273 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  NAND2_X1 U12274 ( .A1(n9707), .A2(n9706), .ZN(n13561) );
  XNOR2_X1 U12275 ( .A(n13996), .B(n9729), .ZN(n9708) );
  NAND2_X1 U12276 ( .A1(n13651), .A2(n6681), .ZN(n9709) );
  NAND2_X1 U12277 ( .A1(n9708), .A2(n9709), .ZN(n13563) );
  NAND2_X1 U12278 ( .A1(n13561), .A2(n13563), .ZN(n13558) );
  INV_X1 U12279 ( .A(n9708), .ZN(n9711) );
  INV_X1 U12280 ( .A(n9709), .ZN(n9710) );
  NAND2_X1 U12281 ( .A1(n9711), .A2(n9710), .ZN(n13559) );
  AND2_X1 U12282 ( .A1(n13650), .A2(n6681), .ZN(n9713) );
  NAND2_X1 U12283 ( .A1(n9712), .A2(n9713), .ZN(n9717) );
  INV_X1 U12284 ( .A(n9712), .ZN(n9715) );
  INV_X1 U12285 ( .A(n9713), .ZN(n9714) );
  NAND2_X1 U12286 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  AND2_X1 U12287 ( .A1(n9717), .A2(n9716), .ZN(n13526) );
  XNOR2_X1 U12288 ( .A(n13986), .B(n9729), .ZN(n9720) );
  NAND2_X1 U12289 ( .A1(n13649), .A2(n6681), .ZN(n9719) );
  XNOR2_X1 U12290 ( .A(n9720), .B(n9719), .ZN(n13621) );
  NAND2_X1 U12291 ( .A1(n9720), .A2(n9719), .ZN(n9721) );
  AND2_X1 U12292 ( .A1(n13648), .A2(n6681), .ZN(n9723) );
  INV_X1 U12293 ( .A(n9722), .ZN(n9725) );
  INV_X1 U12294 ( .A(n9723), .ZN(n9724) );
  NAND2_X1 U12295 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  NAND2_X1 U12296 ( .A1(n9728), .A2(n9726), .ZN(n13444) );
  INV_X1 U12297 ( .A(n6681), .ZN(n12395) );
  OR2_X1 U12298 ( .A1(n13450), .A2(n12395), .ZN(n9730) );
  AND2_X1 U12299 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9733), .ZN(n9734) );
  NAND2_X1 U12300 ( .A1(n15362), .A2(n9735), .ZN(n15357) );
  INV_X1 U12301 ( .A(n15361), .ZN(n9737) );
  NAND2_X1 U12302 ( .A1(n9737), .A2(n9736), .ZN(n10456) );
  OR2_X1 U12303 ( .A1(n9742), .A2(n10743), .ZN(n9739) );
  AOI21_X1 U12304 ( .B1(n9740), .B2(n13632), .A(n13628), .ZN(n9750) );
  INV_X1 U12305 ( .A(n9740), .ZN(n9741) );
  NAND2_X1 U12306 ( .A1(n9741), .A2(n7744), .ZN(n9749) );
  AOI22_X1 U12307 ( .A1(n13647), .A2(n13610), .B1(n13648), .B2(n13622), .ZN(
        n13766) );
  OR2_X1 U12308 ( .A1(n9742), .A2(n10037), .ZN(n13624) );
  OR2_X1 U12309 ( .A1(n13766), .A2(n13624), .ZN(n9747) );
  INV_X1 U12310 ( .A(n9743), .ZN(n9744) );
  OAI21_X1 U12311 ( .B1(n10456), .B2(n10457), .A(n9744), .ZN(n9745) );
  NAND2_X1 U12312 ( .A1(n10459), .A2(n9745), .ZN(n10244) );
  AOI22_X1 U12313 ( .A1(n13760), .A2(n13588), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9746) );
  OAI211_X1 U12314 ( .C1(n9750), .C2(n14053), .A(n9749), .B(n9748), .ZN(
        P2_U3192) );
  NAND2_X1 U12315 ( .A1(n9756), .A2(n12400), .ZN(n12394) );
  NAND2_X1 U12316 ( .A1(n9963), .A2(n9992), .ZN(n9755) );
  NAND2_X1 U12317 ( .A1(n9578), .A2(n6697), .ZN(n9757) );
  NAND3_X1 U12318 ( .A1(n12394), .A2(n9755), .A3(n9757), .ZN(n9759) );
  OAI211_X1 U12319 ( .C1(n9757), .C2(n12400), .A(n6676), .B(n9756), .ZN(n9758)
         );
  NAND2_X1 U12320 ( .A1(n9759), .A2(n9758), .ZN(n9765) );
  NAND2_X1 U12321 ( .A1(n13674), .A2(n6676), .ZN(n9760) );
  NAND2_X1 U12322 ( .A1(n7762), .A2(n9760), .ZN(n9766) );
  NAND2_X1 U12323 ( .A1(n9765), .A2(n9766), .ZN(n9764) );
  NAND2_X1 U12324 ( .A1(n9826), .A2(n13674), .ZN(n9762) );
  NAND2_X1 U12325 ( .A1(n6688), .A2(n11094), .ZN(n9761) );
  NAND2_X1 U12326 ( .A1(n9762), .A2(n9761), .ZN(n9763) );
  NAND2_X1 U12327 ( .A1(n9764), .A2(n9763), .ZN(n9770) );
  INV_X1 U12328 ( .A(n9765), .ZN(n9768) );
  INV_X1 U12329 ( .A(n9766), .ZN(n9767) );
  NAND2_X1 U12330 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  NAND2_X1 U12331 ( .A1(n9770), .A2(n9769), .ZN(n9776) );
  NAND2_X1 U12332 ( .A1(n9826), .A2(n7040), .ZN(n9772) );
  NAND2_X1 U12333 ( .A1(n6688), .A2(n15315), .ZN(n9771) );
  NAND2_X1 U12334 ( .A1(n9772), .A2(n9771), .ZN(n9775) );
  AOI22_X1 U12335 ( .A1(n9826), .A2(n15315), .B1(n6688), .B2(n7040), .ZN(n9773) );
  AOI21_X1 U12336 ( .B1(n9776), .B2(n9775), .A(n9773), .ZN(n9774) );
  NAND2_X1 U12337 ( .A1(n13672), .A2(n6676), .ZN(n9778) );
  OR2_X1 U12338 ( .A1(n6676), .A2(n15379), .ZN(n9777) );
  NAND2_X1 U12339 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  NAND2_X1 U12340 ( .A1(n9826), .A2(n13672), .ZN(n9781) );
  NAND2_X1 U12341 ( .A1(n6688), .A2(n10742), .ZN(n9780) );
  NAND2_X1 U12342 ( .A1(n9826), .A2(n13671), .ZN(n9783) );
  NAND2_X1 U12343 ( .A1(n9931), .A2(n11057), .ZN(n9782) );
  NAND2_X1 U12344 ( .A1(n9783), .A2(n9782), .ZN(n9786) );
  AOI22_X1 U12345 ( .A1(n9826), .A2(n11057), .B1(n9951), .B2(n13671), .ZN(
        n9784) );
  AOI21_X1 U12346 ( .B1(n9787), .B2(n9786), .A(n9784), .ZN(n9785) );
  INV_X1 U12347 ( .A(n9785), .ZN(n9788) );
  NAND2_X1 U12348 ( .A1(n13670), .A2(n9931), .ZN(n9790) );
  OR2_X1 U12349 ( .A1(n9951), .A2(n15386), .ZN(n9789) );
  NAND2_X1 U12350 ( .A1(n9790), .A2(n9789), .ZN(n9793) );
  AOI22_X1 U12351 ( .A1(n9826), .A2(n13670), .B1(n9951), .B2(n9791), .ZN(n9792) );
  AOI21_X1 U12352 ( .B1(n9794), .B2(n9793), .A(n9792), .ZN(n9795) );
  NAND2_X1 U12353 ( .A1(n9826), .A2(n13669), .ZN(n9797) );
  NAND2_X1 U12354 ( .A1(n9931), .A2(n11208), .ZN(n9796) );
  NAND2_X1 U12355 ( .A1(n9797), .A2(n9796), .ZN(n9800) );
  NAND2_X1 U12356 ( .A1(n13669), .A2(n9931), .ZN(n9798) );
  OAI21_X1 U12357 ( .B1(n11076), .B2(n9931), .A(n9798), .ZN(n9799) );
  NAND2_X1 U12358 ( .A1(n11418), .A2(n9954), .ZN(n9803) );
  NAND2_X1 U12359 ( .A1(n13668), .A2(n9931), .ZN(n9802) );
  NAND2_X1 U12360 ( .A1(n9803), .A2(n9802), .ZN(n9806) );
  AOI22_X1 U12361 ( .A1(n11418), .A2(n9951), .B1(n9954), .B2(n13668), .ZN(
        n9804) );
  AOI21_X1 U12362 ( .B1(n9807), .B2(n9806), .A(n9804), .ZN(n9805) );
  INV_X1 U12363 ( .A(n9805), .ZN(n9808) );
  NAND2_X1 U12364 ( .A1(n13498), .A2(n9951), .ZN(n9810) );
  NAND2_X1 U12365 ( .A1(n9826), .A2(n13667), .ZN(n9809) );
  NAND2_X1 U12366 ( .A1(n9810), .A2(n9809), .ZN(n9814) );
  NAND2_X1 U12367 ( .A1(n13498), .A2(n9826), .ZN(n9811) );
  OAI21_X1 U12368 ( .B1(n9812), .B2(n9826), .A(n9811), .ZN(n9813) );
  INV_X1 U12369 ( .A(n9814), .ZN(n9815) );
  NAND2_X1 U12370 ( .A1(n15399), .A2(n9954), .ZN(n9817) );
  NAND2_X1 U12371 ( .A1(n13666), .A2(n9951), .ZN(n9816) );
  NAND2_X1 U12372 ( .A1(n9817), .A2(n9816), .ZN(n9819) );
  AOI22_X1 U12373 ( .A1(n15399), .A2(n9931), .B1(n9954), .B2(n13666), .ZN(
        n9818) );
  AOI21_X1 U12374 ( .B1(n9820), .B2(n9819), .A(n9818), .ZN(n9822) );
  NOR2_X1 U12375 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  NAND2_X1 U12376 ( .A1(n11737), .A2(n9931), .ZN(n9824) );
  NAND2_X1 U12377 ( .A1(n9954), .A2(n13665), .ZN(n9823) );
  NAND2_X1 U12378 ( .A1(n11737), .A2(n9954), .ZN(n9825) );
  OAI21_X1 U12379 ( .B1(n9827), .B2(n9954), .A(n9825), .ZN(n9828) );
  NAND2_X1 U12380 ( .A1(n11607), .A2(n9954), .ZN(n9830) );
  NAND2_X1 U12381 ( .A1(n13664), .A2(n9951), .ZN(n9829) );
  NAND2_X1 U12382 ( .A1(n9830), .A2(n9829), .ZN(n9832) );
  AOI22_X1 U12383 ( .A1(n11607), .A2(n9931), .B1(n9954), .B2(n13664), .ZN(
        n9831) );
  AOI21_X1 U12384 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9834) );
  NAND2_X1 U12385 ( .A1(n11795), .A2(n9931), .ZN(n9836) );
  NAND2_X1 U12386 ( .A1(n9954), .A2(n13663), .ZN(n9835) );
  NAND2_X1 U12387 ( .A1(n11795), .A2(n9954), .ZN(n9837) );
  OAI21_X1 U12388 ( .B1(n9989), .B2(n9954), .A(n9837), .ZN(n9838) );
  NAND2_X1 U12389 ( .A1(n11823), .A2(n9954), .ZN(n9840) );
  NAND2_X1 U12390 ( .A1(n13662), .A2(n9951), .ZN(n9839) );
  NAND2_X1 U12391 ( .A1(n9840), .A2(n9839), .ZN(n9842) );
  AOI22_X1 U12392 ( .A1(n11823), .A2(n9931), .B1(n9954), .B2(n13662), .ZN(
        n9841) );
  AOI21_X1 U12393 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9860) );
  NOR2_X1 U12394 ( .A1(n9843), .A2(n9842), .ZN(n9859) );
  AND2_X1 U12395 ( .A1(n13658), .A2(n9954), .ZN(n9844) );
  AOI21_X1 U12396 ( .B1(n13936), .B2(n9931), .A(n9844), .ZN(n9878) );
  OR2_X1 U12397 ( .A1(n13936), .A2(n13658), .ZN(n9873) );
  AND2_X1 U12398 ( .A1(n13659), .A2(n9954), .ZN(n9845) );
  AOI21_X1 U12399 ( .B1(n13959), .B2(n9931), .A(n9845), .ZN(n9864) );
  NAND2_X1 U12400 ( .A1(n13959), .A2(n9954), .ZN(n9847) );
  NAND2_X1 U12401 ( .A1(n13659), .A2(n9951), .ZN(n9846) );
  NAND2_X1 U12402 ( .A1(n9847), .A2(n9846), .ZN(n9863) );
  AOI22_X1 U12403 ( .A1(n9878), .A2(n9873), .B1(n9864), .B2(n9863), .ZN(n9867)
         );
  AND2_X1 U12404 ( .A1(n13660), .A2(n9954), .ZN(n9848) );
  AOI21_X1 U12405 ( .B1(n11993), .B2(n9951), .A(n9848), .ZN(n9869) );
  NAND2_X1 U12406 ( .A1(n11993), .A2(n9954), .ZN(n9850) );
  NAND2_X1 U12407 ( .A1(n13660), .A2(n9951), .ZN(n9849) );
  NAND2_X1 U12408 ( .A1(n9850), .A2(n9849), .ZN(n9868) );
  NAND2_X1 U12409 ( .A1(n9869), .A2(n9868), .ZN(n9851) );
  AND2_X1 U12410 ( .A1(n9867), .A2(n9851), .ZN(n9881) );
  NAND2_X1 U12411 ( .A1(n14889), .A2(n9931), .ZN(n9853) );
  NAND2_X1 U12412 ( .A1(n9954), .A2(n13661), .ZN(n9852) );
  NAND2_X1 U12413 ( .A1(n9853), .A2(n9852), .ZN(n9861) );
  INV_X1 U12414 ( .A(n9861), .ZN(n9856) );
  AND2_X1 U12415 ( .A1(n13661), .A2(n9951), .ZN(n9854) );
  AOI21_X1 U12416 ( .B1(n14889), .B2(n9954), .A(n9854), .ZN(n9862) );
  AND2_X1 U12417 ( .A1(n9862), .A2(n9861), .ZN(n9880) );
  INV_X1 U12418 ( .A(n9863), .ZN(n9866) );
  INV_X1 U12419 ( .A(n9864), .ZN(n9865) );
  NAND2_X1 U12420 ( .A1(n9866), .A2(n9865), .ZN(n9877) );
  INV_X1 U12421 ( .A(n9867), .ZN(n9870) );
  OR3_X1 U12422 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n9876) );
  NAND2_X1 U12423 ( .A1(n13936), .A2(n9954), .ZN(n9871) );
  OAI21_X1 U12424 ( .B1(n9872), .B2(n9954), .A(n9871), .ZN(n9874) );
  MUX2_X1 U12425 ( .A(n9877), .B(n9874), .S(n9873), .Z(n9875) );
  OAI211_X1 U12426 ( .C1(n9878), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9879)
         );
  AOI21_X1 U12427 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9882) );
  NAND2_X1 U12428 ( .A1(n9883), .A2(n9882), .ZN(n9889) );
  NAND2_X1 U12429 ( .A1(n14031), .A2(n9951), .ZN(n9885) );
  NAND2_X1 U12430 ( .A1(n9954), .A2(n13657), .ZN(n9884) );
  NAND2_X1 U12431 ( .A1(n9885), .A2(n9884), .ZN(n9890) );
  NAND2_X1 U12432 ( .A1(n14031), .A2(n9954), .ZN(n9886) );
  OAI21_X1 U12433 ( .B1(n9887), .B2(n9954), .A(n9886), .ZN(n9888) );
  INV_X1 U12434 ( .A(n9890), .ZN(n9891) );
  NAND2_X1 U12435 ( .A1(n13907), .A2(n9954), .ZN(n9893) );
  NAND2_X1 U12436 ( .A1(n13656), .A2(n9931), .ZN(n9892) );
  NAND2_X1 U12437 ( .A1(n9893), .A2(n9892), .ZN(n9895) );
  AOI22_X1 U12438 ( .A1(n13907), .A2(n9951), .B1(n9954), .B2(n13656), .ZN(
        n9894) );
  AOI21_X1 U12439 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9898) );
  OR2_X1 U12440 ( .A1(n9898), .A2(n9897), .ZN(n9904) );
  NAND2_X1 U12441 ( .A1(n14022), .A2(n9951), .ZN(n9900) );
  NAND2_X1 U12442 ( .A1(n13655), .A2(n9954), .ZN(n9899) );
  NAND2_X1 U12443 ( .A1(n9900), .A2(n9899), .ZN(n9903) );
  AOI22_X1 U12444 ( .A1(n14022), .A2(n9954), .B1(n13655), .B2(n9931), .ZN(
        n9901) );
  AOI21_X1 U12445 ( .B1(n9904), .B2(n9903), .A(n9901), .ZN(n9902) );
  INV_X1 U12446 ( .A(n9902), .ZN(n9907) );
  NOR2_X1 U12447 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  INV_X1 U12448 ( .A(n9905), .ZN(n9906) );
  NAND2_X1 U12449 ( .A1(n13877), .A2(n9954), .ZN(n9909) );
  NAND2_X1 U12450 ( .A1(n13654), .A2(n9951), .ZN(n9908) );
  NAND2_X1 U12451 ( .A1(n9909), .A2(n9908), .ZN(n9913) );
  NAND2_X1 U12452 ( .A1(n13877), .A2(n9931), .ZN(n9911) );
  NAND2_X1 U12453 ( .A1(n13654), .A2(n9954), .ZN(n9910) );
  NAND2_X1 U12454 ( .A1(n9911), .A2(n9910), .ZN(n9912) );
  NAND2_X1 U12455 ( .A1(n14010), .A2(n6676), .ZN(n9915) );
  NAND2_X1 U12456 ( .A1(n13653), .A2(n9954), .ZN(n9914) );
  NAND2_X1 U12457 ( .A1(n9915), .A2(n9914), .ZN(n9917) );
  AOI22_X1 U12458 ( .A1(n14010), .A2(n9954), .B1(n13653), .B2(n9951), .ZN(
        n9916) );
  AOI21_X1 U12459 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9920) );
  NOR2_X1 U12460 ( .A1(n9918), .A2(n9917), .ZN(n9919) );
  NAND2_X1 U12461 ( .A1(n13842), .A2(n9954), .ZN(n9922) );
  NAND2_X1 U12462 ( .A1(n13652), .A2(n9951), .ZN(n9921) );
  NAND2_X1 U12463 ( .A1(n9922), .A2(n9921), .ZN(n9924) );
  AOI22_X1 U12464 ( .A1(n13842), .A2(n9931), .B1(n9954), .B2(n13652), .ZN(
        n9923) );
  AND2_X1 U12465 ( .A1(n13651), .A2(n9954), .ZN(n9926) );
  AOI21_X1 U12466 ( .B1(n13996), .B2(n6688), .A(n9926), .ZN(n9933) );
  NAND2_X1 U12467 ( .A1(n13996), .A2(n9954), .ZN(n9927) );
  OAI21_X1 U12468 ( .B1(n9928), .B2(n9954), .A(n9927), .ZN(n9929) );
  NAND2_X1 U12469 ( .A1(n13811), .A2(n6688), .ZN(n9930) );
  OAI21_X1 U12470 ( .B1(n9932), .B2(n6688), .A(n9930), .ZN(n9937) );
  NAND3_X1 U12471 ( .A1(n9936), .A2(n9937), .A3(n9935), .ZN(n9943) );
  AND2_X1 U12472 ( .A1(n13650), .A2(n6688), .ZN(n9934) );
  AOI21_X1 U12473 ( .B1(n13811), .B2(n9954), .A(n9934), .ZN(n9938) );
  INV_X1 U12474 ( .A(n9937), .ZN(n9940) );
  INV_X1 U12475 ( .A(n9938), .ZN(n9939) );
  OR2_X1 U12476 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  NAND3_X1 U12477 ( .A1(n9943), .A2(n9942), .A3(n9941), .ZN(n9949) );
  NAND2_X1 U12478 ( .A1(n13986), .A2(n6676), .ZN(n9945) );
  NAND2_X1 U12479 ( .A1(n13649), .A2(n9954), .ZN(n9944) );
  NAND2_X1 U12480 ( .A1(n9945), .A2(n9944), .ZN(n9948) );
  AOI22_X1 U12481 ( .A1(n13986), .A2(n9954), .B1(n13649), .B2(n6688), .ZN(
        n9946) );
  AOI21_X1 U12482 ( .B1(n9949), .B2(n9948), .A(n9946), .ZN(n9947) );
  INV_X1 U12483 ( .A(n9947), .ZN(n9950) );
  NAND2_X1 U12484 ( .A1(n13980), .A2(n9954), .ZN(n9953) );
  NAND2_X1 U12485 ( .A1(n13648), .A2(n6688), .ZN(n9952) );
  NAND2_X1 U12486 ( .A1(n9953), .A2(n9952), .ZN(n9959) );
  AOI22_X1 U12487 ( .A1(n9955), .A2(n9954), .B1(n9494), .B2(n6676), .ZN(n9967)
         );
  OAI22_X1 U12488 ( .A1(n14053), .A2(n9954), .B1(n13450), .B2(n6688), .ZN(
        n9966) );
  OAI22_X1 U12489 ( .A1(n13748), .A2(n6676), .B1(n9956), .B2(n9954), .ZN(n9970) );
  AOI22_X1 U12490 ( .A1(n9574), .A2(n6688), .B1(n9954), .B2(n13647), .ZN(n9971) );
  NOR2_X1 U12491 ( .A1(n9970), .A2(n9971), .ZN(n9968) );
  AOI21_X1 U12492 ( .B1(n9967), .B2(n9966), .A(n9968), .ZN(n9957) );
  AOI22_X1 U12493 ( .A1(n13980), .A2(n6676), .B1(n9954), .B2(n13648), .ZN(
        n9958) );
  NOR2_X1 U12494 ( .A1(n9954), .A2(n9969), .ZN(n9979) );
  OAI211_X1 U12495 ( .C1(n6685), .C2(n9993), .A(n10014), .B(n10037), .ZN(n9961) );
  OAI21_X1 U12496 ( .B1(n9979), .B2(n9961), .A(n13646), .ZN(n9962) );
  OAI21_X1 U12497 ( .B1(n14050), .B2(n6676), .A(n9962), .ZN(n9973) );
  AOI22_X1 U12498 ( .A1(n13742), .A2(n6676), .B1(n9954), .B2(n13646), .ZN(
        n9972) );
  XNOR2_X1 U12499 ( .A(n9982), .B(n9969), .ZN(n9986) );
  NAND2_X1 U12500 ( .A1(n7745), .A2(n9964), .ZN(n9965) );
  NOR4_X1 U12501 ( .A1(n9986), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9978)
         );
  INV_X1 U12502 ( .A(n9969), .ZN(n13645) );
  NAND2_X1 U12503 ( .A1(n9954), .A2(n13645), .ZN(n9976) );
  MUX2_X1 U12504 ( .A(n13645), .B(n9954), .S(n9982), .Z(n9975) );
  AOI22_X1 U12505 ( .A1(n9973), .A2(n9972), .B1(n9971), .B2(n9970), .ZN(n9974)
         );
  AOI21_X1 U12506 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9977) );
  OAI21_X1 U12507 ( .B1(n9978), .B2(n9977), .A(n7745), .ZN(n10024) );
  INV_X1 U12508 ( .A(n9979), .ZN(n9981) );
  NAND2_X1 U12509 ( .A1(n9982), .A2(n9954), .ZN(n9980) );
  OAI211_X1 U12510 ( .C1(n9982), .C2(n13645), .A(n9981), .B(n9980), .ZN(n10023) );
  INV_X1 U12511 ( .A(n10023), .ZN(n9983) );
  NOR2_X1 U12512 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  XNOR2_X1 U12513 ( .A(n13742), .B(n13646), .ZN(n10012) );
  XNOR2_X1 U12514 ( .A(n13907), .B(n9987), .ZN(n13899) );
  NAND2_X1 U12515 ( .A1(n9988), .A2(n13867), .ZN(n13885) );
  XNOR2_X1 U12516 ( .A(n11795), .B(n9989), .ZN(n11793) );
  XNOR2_X1 U12517 ( .A(n11823), .B(n9990), .ZN(n11820) );
  OAI21_X1 U12518 ( .B1(n9756), .B2(n9992), .A(n9991), .ZN(n10225) );
  NAND4_X1 U12519 ( .A1(n10424), .A2(n11092), .A3(n9993), .A4(n10225), .ZN(
        n9995) );
  NOR3_X1 U12520 ( .A1(n9995), .A2(n10720), .A3(n9994), .ZN(n9996) );
  NAND4_X1 U12521 ( .A1(n9996), .A2(n11284), .A3(n10836), .A4(n11065), .ZN(
        n9997) );
  NOR2_X1 U12522 ( .A1(n9997), .A2(n11237), .ZN(n9999) );
  NAND4_X1 U12523 ( .A1(n11603), .A2(n9999), .A3(n11518), .A4(n9998), .ZN(
        n10000) );
  OR4_X1 U12524 ( .A1(n13947), .A2(n11793), .A3(n11820), .A4(n10000), .ZN(
        n10001) );
  NOR2_X1 U12525 ( .A1(n13931), .A2(n10001), .ZN(n10002) );
  NAND4_X1 U12526 ( .A1(n13923), .A2(n10002), .A3(n11989), .A4(n14888), .ZN(
        n10003) );
  OR4_X1 U12527 ( .A1(n10004), .A2(n13899), .A3(n13885), .A4(n10003), .ZN(
        n10005) );
  OR3_X1 U12528 ( .A1(n13823), .A2(n13855), .A3(n10005), .ZN(n10008) );
  NAND2_X1 U12529 ( .A1(n10007), .A2(n10006), .ZN(n13792) );
  OR4_X1 U12530 ( .A1(n10008), .A2(n13799), .A3(n13835), .A4(n13792), .ZN(
        n10009) );
  NOR2_X1 U12531 ( .A1(n13756), .A2(n10009), .ZN(n10011) );
  AND4_X1 U12532 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n13770), .ZN(
        n10013) );
  AOI21_X1 U12533 ( .B1(n10015), .B2(n10739), .A(n10014), .ZN(n10027) );
  INV_X1 U12534 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U12535 ( .A1(n10016), .A2(n13726), .ZN(n10026) );
  NAND2_X1 U12536 ( .A1(n10027), .A2(n10026), .ZN(n10020) );
  MUX2_X1 U12537 ( .A(n9752), .B(n6685), .S(n8122), .Z(n10017) );
  NAND2_X1 U12538 ( .A1(n10018), .A2(n10739), .ZN(n10019) );
  OAI21_X1 U12539 ( .B1(n9752), .B2(n10739), .A(n10037), .ZN(n10021) );
  AOI21_X1 U12540 ( .B1(n9578), .B2(n6685), .A(n10021), .ZN(n10022) );
  NAND2_X1 U12541 ( .A1(n10025), .A2(n7760), .ZN(n10029) );
  AND3_X1 U12542 ( .A1(n10027), .A2(n9751), .A3(n10026), .ZN(n10028) );
  AOI21_X1 U12543 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10041) );
  OR2_X1 U12544 ( .A1(n10035), .A2(P2_U3088), .ZN(n11887) );
  INV_X1 U12545 ( .A(n10035), .ZN(n10033) );
  OAI21_X1 U12546 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10036) );
  NAND2_X1 U12547 ( .A1(n10035), .A2(n10034), .ZN(n10042) );
  AND2_X1 U12548 ( .A1(n10036), .A2(n10042), .ZN(n15232) );
  AND2_X1 U12549 ( .A1(n15232), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15289) );
  INV_X1 U12550 ( .A(n15289), .ZN(n15313) );
  NOR4_X1 U12551 ( .A1(n15313), .A2(n10263), .A3(n10037), .A4(n14104), .ZN(
        n10039) );
  OAI21_X1 U12552 ( .B1(n11887), .B2(n9754), .A(P2_B_REG_SCAN_IN), .ZN(n10038)
         );
  OR2_X1 U12553 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  OAI21_X1 U12554 ( .B1(n10041), .B2(n11887), .A(n10040), .ZN(P2_U3328) );
  NAND2_X1 U12555 ( .A1(n10088), .A2(n10090), .ZN(n10093) );
  NOR2_X1 U12556 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n10048) );
  INV_X1 U12557 ( .A(n10209), .ZN(n10065) );
  NOR2_X1 U12558 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n10058) );
  NOR2_X1 U12559 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n10057) );
  NOR2_X1 U12560 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n10056) );
  OAI21_X1 U12561 ( .B1(n10055), .B2(n10061), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10060) );
  MUX2_X1 U12562 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10060), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10063) );
  NOR3_X1 U12563 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U12564 ( .A1(n6829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10066) );
  MUX2_X1 U12565 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10066), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n10068) );
  NAND2_X1 U12566 ( .A1(n10068), .A2(n10067), .ZN(n10639) );
  INV_X1 U12567 ( .A(n10070), .ZN(n10071) );
  NAND2_X1 U12568 ( .A1(n6672), .A2(P3_U3151), .ZN(n13430) );
  NAND2_X1 U12569 ( .A1(n10593), .A2(n6665), .ZN(n12381) );
  INV_X1 U12570 ( .A(n10072), .ZN(n10073) );
  OAI222_X1 U12571 ( .A1(P3_U3151), .A2(n11120), .B1(n13430), .B2(n10074), 
        .C1(n12381), .C2(n10073), .ZN(P3_U3291) );
  INV_X1 U12572 ( .A(n10805), .ZN(n10780) );
  INV_X1 U12573 ( .A(n10075), .ZN(n10076) );
  OAI222_X1 U12574 ( .A1(n6665), .A2(n10780), .B1(n13430), .B2(n10077), .C1(
        n12381), .C2(n10076), .ZN(P3_U3292) );
  INV_X1 U12575 ( .A(SI_5_), .ZN(n10080) );
  INV_X1 U12576 ( .A(n10078), .ZN(n10079) );
  OAI222_X1 U12577 ( .A1(n6665), .A2(n15438), .B1(n13430), .B2(n10080), .C1(
        n12381), .C2(n10079), .ZN(P3_U3290) );
  INV_X1 U12578 ( .A(n10779), .ZN(n10773) );
  INV_X1 U12579 ( .A(n10081), .ZN(n10082) );
  OAI222_X1 U12580 ( .A1(n6665), .A2(n10773), .B1(n13430), .B2(n10083), .C1(
        n12381), .C2(n10082), .ZN(P3_U3293) );
  INV_X1 U12581 ( .A(SI_7_), .ZN(n10087) );
  INV_X1 U12582 ( .A(n10085), .ZN(n10086) );
  OAI222_X1 U12583 ( .A1(P3_U3151), .A2(n15475), .B1(n13430), .B2(n10087), 
        .C1(n12381), .C2(n10086), .ZN(P3_U3288) );
  INV_X1 U12584 ( .A(n10088), .ZN(n10089) );
  NAND2_X1 U12585 ( .A1(n10089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U12586 ( .A(n10091), .B(n10090), .ZN(n14288) );
  NAND2_X1 U12587 ( .A1(n10593), .A2(P1_U3086), .ZN(n14775) );
  NAND2_X1 U12588 ( .A1(n6673), .A2(P1_U3086), .ZN(n14777) );
  OAI222_X1 U12589 ( .A1(n14288), .A2(P1_U3086), .B1(n14775), .B2(n10822), 
        .C1(n10819), .C2(n14777), .ZN(P1_U3353) );
  NAND2_X1 U12590 ( .A1(n10093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10094) );
  MUX2_X1 U12591 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10094), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n10095) );
  AND2_X1 U12592 ( .A1(n10105), .A2(n10095), .ZN(n14307) );
  INV_X1 U12593 ( .A(n14307), .ZN(n10097) );
  OAI222_X1 U12594 ( .A1(n10097), .A2(P1_U3086), .B1(n14775), .B2(n10892), 
        .C1(n10096), .C2(n14777), .ZN(P1_U3352) );
  INV_X1 U12595 ( .A(SI_9_), .ZN(n10098) );
  OAI222_X1 U12596 ( .A1(n6665), .A2(n15512), .B1(n13430), .B2(n10098), .C1(
        n12381), .C2(n6838), .ZN(P3_U3286) );
  NOR2_X1 U12597 ( .A1(n6672), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14088) );
  NAND2_X1 U12598 ( .A1(n14088), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n10099) );
  INV_X1 U12599 ( .A(n10254), .ZN(n10255) );
  NAND2_X1 U12600 ( .A1(n10255), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15230) );
  OAI211_X1 U12601 ( .C1(n10594), .C2(n14111), .A(n10099), .B(n15230), .ZN(
        P2_U3326) );
  INV_X2 U12602 ( .A(n14088), .ZN(n14106) );
  INV_X2 U12603 ( .A(n14098), .ZN(n14111) );
  OAI222_X1 U12604 ( .A1(n14106), .A2(n10100), .B1(n14111), .B2(n10822), .C1(
        P2_U3088), .C2(n10256), .ZN(P2_U3325) );
  OAI222_X1 U12605 ( .A1(n14106), .A2(n10101), .B1(n14111), .B2(n10892), .C1(
        P2_U3088), .C2(n10258), .ZN(P2_U3324) );
  INV_X1 U12606 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10102) );
  INV_X1 U12607 ( .A(n14775), .ZN(n11890) );
  INV_X1 U12608 ( .A(n11890), .ZN(n14780) );
  INV_X1 U12609 ( .A(n14777), .ZN(n14763) );
  OAI222_X1 U12610 ( .A1(n10595), .A2(P1_U3086), .B1(n14780), .B2(n10594), 
        .C1(n10103), .C2(n14772), .ZN(P1_U3354) );
  NAND2_X1 U12611 ( .A1(n10105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10104) );
  MUX2_X1 U12612 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10104), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n10108) );
  INV_X1 U12613 ( .A(n10105), .ZN(n10107) );
  NAND2_X1 U12614 ( .A1(n10107), .A2(n10106), .ZN(n10124) );
  NAND2_X1 U12615 ( .A1(n10108), .A2(n10124), .ZN(n10923) );
  OAI222_X1 U12616 ( .A1(n10923), .A2(P1_U3086), .B1(n14775), .B2(n10109), 
        .C1(n10110), .C2(n14777), .ZN(P1_U3351) );
  OAI222_X1 U12617 ( .A1(n14106), .A2(n10111), .B1(n14111), .B2(n10109), .C1(
        P2_U3088), .C2(n10282), .ZN(P2_U3323) );
  INV_X1 U12618 ( .A(n10112), .ZN(n10113) );
  OAI222_X1 U12619 ( .A1(P3_U3151), .A2(n11374), .B1(n13430), .B2(n10114), 
        .C1(n12381), .C2(n10113), .ZN(P3_U3285) );
  OAI222_X1 U12620 ( .A1(n6665), .A2(n11564), .B1(n13430), .B2(n10116), .C1(
        n12381), .C2(n10115), .ZN(P3_U3284) );
  INV_X1 U12621 ( .A(n12381), .ZN(n11051) );
  INV_X1 U12622 ( .A(n11051), .ZN(n13439) );
  CLKBUF_X1 U12623 ( .A(n13430), .Z(n13441) );
  OAI222_X1 U12624 ( .A1(n13439), .A2(n10118), .B1(n13441), .B2(n10117), .C1(
        P3_U3151), .C2(n10747), .ZN(P3_U3294) );
  OAI222_X1 U12625 ( .A1(P3_U3151), .A2(n15458), .B1(n13439), .B2(n10120), 
        .C1(n10119), .C2(n13441), .ZN(P3_U3289) );
  OAI222_X1 U12626 ( .A1(n15493), .A2(n6665), .B1(n13439), .B2(n10122), .C1(
        n10121), .C2(n13441), .ZN(P3_U3287) );
  NAND2_X1 U12627 ( .A1(n10124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U12628 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10123), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n10125) );
  AND2_X1 U12629 ( .A1(n10125), .A2(n10140), .ZN(n10963) );
  INV_X1 U12630 ( .A(n10963), .ZN(n10468) );
  INV_X1 U12631 ( .A(n10962), .ZN(n10127) );
  OAI222_X1 U12632 ( .A1(n10468), .A2(P1_U3086), .B1(n14775), .B2(n10127), 
        .C1(n10126), .C2(n14777), .ZN(P1_U3350) );
  OAI222_X1 U12633 ( .A1(n14106), .A2(n10128), .B1(n14111), .B2(n10127), .C1(
        P2_U3088), .C2(n10283), .ZN(P2_U3322) );
  INV_X1 U12634 ( .A(n10129), .ZN(n10130) );
  OAI222_X1 U12635 ( .A1(P3_U3151), .A2(n11899), .B1(n13430), .B2(n10131), 
        .C1(n12381), .C2(n10130), .ZN(P3_U3283) );
  INV_X1 U12636 ( .A(n10968), .ZN(n10135) );
  INV_X1 U12637 ( .A(n10284), .ZN(n10304) );
  OAI222_X1 U12638 ( .A1(n14106), .A2(n10132), .B1(n14111), .B2(n10135), .C1(
        P2_U3088), .C2(n10304), .ZN(P2_U3321) );
  NAND2_X1 U12639 ( .A1(n10140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10133) );
  XNOR2_X1 U12640 ( .A(n10133), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10969) );
  INV_X1 U12641 ( .A(n10969), .ZN(n14329) );
  OAI222_X1 U12642 ( .A1(n14329), .A2(P1_U3086), .B1(n14775), .B2(n10135), 
        .C1(n10134), .C2(n14777), .ZN(P1_U3349) );
  AND2_X1 U12643 ( .A1(n10137), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12644 ( .A1(n10137), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12645 ( .A1(n10137), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12646 ( .A1(n10137), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12647 ( .A1(n10137), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12648 ( .A1(n10137), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12649 ( .A1(n10137), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12650 ( .A1(n10137), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12651 ( .A1(n10137), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12652 ( .A1(n10137), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12653 ( .A1(n10137), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12654 ( .A1(n10137), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12655 ( .A1(n10137), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12656 ( .A1(n10137), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12657 ( .A1(n10137), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12658 ( .A1(n10137), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12659 ( .A1(n10137), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12660 ( .A1(n10137), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12661 ( .A1(n10137), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12662 ( .A1(n10137), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12663 ( .A1(n10137), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12664 ( .A1(n10137), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12665 ( .A1(n10137), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12666 ( .A1(n10137), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12667 ( .A1(n10137), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12668 ( .A1(n10137), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12669 ( .A1(n10137), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12670 ( .A1(n10137), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12671 ( .A1(n10137), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12672 ( .A1(n10137), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  OAI222_X1 U12673 ( .A1(n6665), .A2(n12958), .B1(n13430), .B2(n10139), .C1(
        n12381), .C2(n10138), .ZN(P3_U3282) );
  INV_X1 U12674 ( .A(n10140), .ZN(n10142) );
  NAND2_X1 U12675 ( .A1(n10142), .A2(n10141), .ZN(n10151) );
  NAND2_X1 U12676 ( .A1(n10151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10143) );
  XNOR2_X1 U12677 ( .A(n10143), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14350) );
  INV_X1 U12678 ( .A(n14350), .ZN(n10470) );
  INV_X1 U12679 ( .A(n10980), .ZN(n10145) );
  OAI222_X1 U12680 ( .A1(n10470), .A2(P1_U3086), .B1(n14775), .B2(n10145), 
        .C1(n10144), .C2(n14777), .ZN(P1_U3348) );
  INV_X1 U12681 ( .A(n10397), .ZN(n10292) );
  OAI222_X1 U12682 ( .A1(n14106), .A2(n10146), .B1(n14111), .B2(n10145), .C1(
        P2_U3088), .C2(n10292), .ZN(P2_U3320) );
  OAI222_X1 U12683 ( .A1(P3_U3151), .A2(n12976), .B1(n13430), .B2(n10148), 
        .C1(n12381), .C2(n10147), .ZN(P3_U3281) );
  INV_X1 U12684 ( .A(n10993), .ZN(n10154) );
  INV_X1 U12685 ( .A(n11106), .ZN(n10149) );
  OAI222_X1 U12686 ( .A1(n14106), .A2(n10150), .B1(n14111), .B2(n10154), .C1(
        P2_U3088), .C2(n10149), .ZN(P2_U3319) );
  NAND2_X1 U12687 ( .A1(n10157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10152) );
  XNOR2_X1 U12688 ( .A(n10152), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10994) );
  INV_X1 U12689 ( .A(n10994), .ZN(n10495) );
  OAI222_X1 U12690 ( .A1(n10495), .A2(P1_U3086), .B1(n14775), .B2(n10154), 
        .C1(n10153), .C2(n14777), .ZN(P1_U3347) );
  INV_X1 U12691 ( .A(n11264), .ZN(n10159) );
  INV_X1 U12692 ( .A(n15267), .ZN(n10155) );
  OAI222_X1 U12693 ( .A1(n14106), .A2(n10156), .B1(n14111), .B2(n10159), .C1(
        P2_U3088), .C2(n10155), .ZN(P2_U3318) );
  XNOR2_X1 U12694 ( .A(n10176), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11265) );
  INV_X1 U12695 ( .A(n11265), .ZN(n10535) );
  OAI222_X1 U12696 ( .A1(n10535), .A2(P1_U3086), .B1(n14775), .B2(n10159), 
        .C1(n10158), .C2(n14777), .ZN(P1_U3346) );
  OAI222_X1 U12697 ( .A1(n6665), .A2(n13007), .B1(n13441), .B2(n10161), .C1(
        n13439), .C2(n10160), .ZN(P3_U3280) );
  NAND2_X1 U12698 ( .A1(n10176), .A2(n10162), .ZN(n10163) );
  NAND2_X1 U12699 ( .A1(n10163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10164) );
  XNOR2_X1 U12700 ( .A(n10164), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11471) );
  INV_X1 U12701 ( .A(n11471), .ZN(n10522) );
  INV_X1 U12702 ( .A(n11470), .ZN(n10166) );
  OAI222_X1 U12703 ( .A1(n10522), .A2(P1_U3086), .B1(n14780), .B2(n10166), 
        .C1(n10165), .C2(n14777), .ZN(P1_U3345) );
  INV_X1 U12704 ( .A(n11108), .ZN(n15271) );
  OAI222_X1 U12705 ( .A1(n14106), .A2(n10167), .B1(n14111), .B2(n10166), .C1(
        P2_U3088), .C2(n15271), .ZN(P2_U3317) );
  NAND2_X1 U12706 ( .A1(n12894), .A2(n10665), .ZN(n10168) );
  OAI21_X1 U12707 ( .B1(n10665), .B2(n10169), .A(n10168), .ZN(P3_U3505) );
  INV_X1 U12708 ( .A(n13045), .ZN(n13031) );
  OAI222_X1 U12709 ( .A1(n13441), .A2(n10171), .B1(n13439), .B2(n10170), .C1(
        n13031), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12710 ( .A(n11454), .ZN(n10178) );
  INV_X1 U12711 ( .A(n11332), .ZN(n11338) );
  OAI222_X1 U12712 ( .A1(n14106), .A2(n10172), .B1(n14111), .B2(n10178), .C1(
        P2_U3088), .C2(n11338), .ZN(P2_U3316) );
  INV_X1 U12713 ( .A(n10173), .ZN(n10174) );
  NAND2_X1 U12714 ( .A1(n10174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U12715 ( .A1(n10176), .A2(n10175), .ZN(n10220) );
  XNOR2_X1 U12716 ( .A(n10220), .B(n10177), .ZN(n11455) );
  INV_X1 U12717 ( .A(n11455), .ZN(n10512) );
  OAI222_X1 U12718 ( .A1(n14777), .A2(n10179), .B1(n14780), .B2(n10178), .C1(
        P1_U3086), .C2(n10512), .ZN(P1_U3344) );
  NAND2_X1 U12719 ( .A1(n11301), .A2(n10665), .ZN(n10180) );
  OAI21_X1 U12720 ( .B1(n10665), .B2(n10181), .A(n10180), .ZN(P3_U3495) );
  NAND2_X1 U12721 ( .A1(n11505), .A2(n10665), .ZN(n10182) );
  OAI21_X1 U12722 ( .B1(n10665), .B2(n10183), .A(n10182), .ZN(P3_U3496) );
  OAI222_X1 U12723 ( .A1(P3_U3151), .A2(n13046), .B1(n13441), .B2(n10185), 
        .C1(n12381), .C2(n10184), .ZN(P3_U3278) );
  INV_X1 U12724 ( .A(n11218), .ZN(n10186) );
  OR2_X1 U12725 ( .A1(n10639), .A2(P1_U3086), .ZN(n12374) );
  NAND2_X1 U12726 ( .A1(n10186), .A2(n12374), .ZN(n10201) );
  NAND2_X1 U12727 ( .A1(n10187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10188) );
  XNOR2_X1 U12728 ( .A(n10188), .B(n12177), .ZN(n10576) );
  INV_X1 U12729 ( .A(n10189), .ZN(n10190) );
  NAND2_X1 U12730 ( .A1(n10190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U12731 ( .A1(n10639), .A2(n12190), .ZN(n10198) );
  NAND2_X1 U12732 ( .A1(n10578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12733 ( .A1(n10195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10197) );
  XNOR2_X2 U12734 ( .A(n10197), .B(n10196), .ZN(n14776) );
  NAND2_X1 U12735 ( .A1(n10198), .A2(n12116), .ZN(n10199) );
  INV_X1 U12736 ( .A(n10199), .ZN(n10200) );
  NAND2_X1 U12737 ( .A1(n10201), .A2(n10200), .ZN(n10356) );
  INV_X1 U12738 ( .A(n14776), .ZN(n10597) );
  INV_X1 U12739 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10203) );
  AOI21_X1 U12740 ( .B1(n10597), .B2(n10203), .A(n10202), .ZN(n14287) );
  OAI21_X1 U12741 ( .B1(n10597), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14287), .ZN(
        n10204) );
  XNOR2_X1 U12742 ( .A(n10204), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U12743 ( .A1(n10359), .A2(n10205), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10206) );
  OAI21_X1 U12744 ( .B1(n15064), .B2(n7534), .A(n10206), .ZN(P1_U3243) );
  NAND2_X1 U12745 ( .A1(n12915), .A2(n10665), .ZN(n10207) );
  OAI21_X1 U12746 ( .B1(n10665), .B2(n10208), .A(n10207), .ZN(P3_U3508) );
  NAND2_X1 U12747 ( .A1(n10209), .A2(P1_B_REG_SCAN_IN), .ZN(n10211) );
  MUX2_X1 U12748 ( .A(P1_B_REG_SCAN_IN), .B(n10211), .S(n10210), .Z(n10213) );
  NAND2_X1 U12749 ( .A1(n10214), .A2(n14781), .ZN(n10216) );
  OAI22_X1 U12750 ( .A1(n15143), .A2(P1_D_REG_1__SCAN_IN), .B1(n10065), .B2(
        n10216), .ZN(n10215) );
  INV_X1 U12751 ( .A(n10215), .ZN(P1_U3446) );
  INV_X1 U12752 ( .A(n10210), .ZN(n10217) );
  OAI22_X1 U12753 ( .A1(n15143), .A2(P1_D_REG_0__SCAN_IN), .B1(n10217), .B2(
        n10216), .ZN(n10218) );
  INV_X1 U12754 ( .A(n10218), .ZN(P1_U3445) );
  INV_X1 U12755 ( .A(n11687), .ZN(n11682) );
  INV_X1 U12756 ( .A(n11659), .ZN(n10223) );
  OAI222_X1 U12757 ( .A1(P2_U3088), .A2(n11682), .B1(n14111), .B2(n10223), 
        .C1(n10219), .C2(n14106), .ZN(P2_U3315) );
  NAND2_X1 U12758 ( .A1(n10221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10312) );
  XNOR2_X1 U12759 ( .A(n10312), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11660) );
  INV_X1 U12760 ( .A(n11660), .ZN(n11041) );
  OAI222_X1 U12761 ( .A1(P1_U3086), .A2(n11041), .B1(n14780), .B2(n10223), 
        .C1(n10222), .C2(n14772), .ZN(P1_U3343) );
  INV_X1 U12762 ( .A(n10225), .ZN(n10464) );
  INV_X1 U12763 ( .A(n15401), .ZN(n15417) );
  NOR2_X1 U12764 ( .A1(n10224), .A2(n12400), .ZN(n10455) );
  INV_X1 U12765 ( .A(n15412), .ZN(n15406) );
  NOR2_X1 U12766 ( .A1(n15406), .A2(n14882), .ZN(n10226) );
  NAND2_X1 U12767 ( .A1(n13610), .A2(n13674), .ZN(n12391) );
  OAI21_X1 U12768 ( .B1(n10226), .B2(n10225), .A(n12391), .ZN(n10454) );
  AOI211_X1 U12769 ( .C1(n10464), .C2(n15417), .A(n10455), .B(n10454), .ZN(
        n15364) );
  NAND2_X1 U12770 ( .A1(n15429), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10227) );
  OAI21_X1 U12771 ( .B1(n15364), .B2(n15429), .A(n10227), .ZN(P2_U3499) );
  NAND2_X1 U12772 ( .A1(n11807), .A2(n10665), .ZN(n10228) );
  OAI21_X1 U12773 ( .B1(P3_U3897), .B2(n10229), .A(n10228), .ZN(P3_U3501) );
  NAND2_X1 U12774 ( .A1(n11451), .A2(n10665), .ZN(n10230) );
  OAI21_X1 U12775 ( .B1(P3_U3897), .B2(n10231), .A(n10230), .ZN(P3_U3497) );
  NAND2_X1 U12776 ( .A1(n15528), .A2(n10665), .ZN(n10232) );
  OAI21_X1 U12777 ( .B1(P3_U3897), .B2(n10233), .A(n10232), .ZN(P3_U3500) );
  NAND2_X1 U12778 ( .A1(n13187), .A2(n10665), .ZN(n10234) );
  OAI21_X1 U12779 ( .B1(n10665), .B2(n10235), .A(n10234), .ZN(P3_U3510) );
  NAND2_X1 U12780 ( .A1(n12904), .A2(n10665), .ZN(n10236) );
  OAI21_X1 U12781 ( .B1(n10665), .B2(n10237), .A(n10236), .ZN(P3_U3513) );
  NAND2_X1 U12782 ( .A1(n13204), .A2(n10665), .ZN(n10238) );
  OAI21_X1 U12783 ( .B1(n10665), .B2(n10239), .A(n10238), .ZN(P3_U3511) );
  INV_X1 U12784 ( .A(n13628), .ZN(n13644) );
  OAI21_X1 U12785 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(n10243) );
  NAND2_X1 U12786 ( .A1(n10243), .A2(n13632), .ZN(n10248) );
  OR2_X1 U12787 ( .A1(n10244), .A2(P2_U3088), .ZN(n12393) );
  INV_X1 U12788 ( .A(n13624), .ZN(n13641) );
  NAND2_X1 U12789 ( .A1(n13610), .A2(n7040), .ZN(n10246) );
  NAND2_X1 U12790 ( .A1(n13551), .A2(n9756), .ZN(n10245) );
  NAND2_X1 U12791 ( .A1(n10246), .A2(n10245), .ZN(n11089) );
  AOI22_X1 U12792 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n12393), .B1(n13641), 
        .B2(n11089), .ZN(n10247) );
  OAI211_X1 U12793 ( .C1(n15366), .C2(n13644), .A(n10248), .B(n10247), .ZN(
        P2_U3194) );
  INV_X1 U12794 ( .A(n10258), .ZN(n10344) );
  INV_X1 U12795 ( .A(n10256), .ZN(n15248) );
  XNOR2_X1 U12796 ( .A(n10254), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n15226) );
  AND2_X1 U12797 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10249) );
  XOR2_X1 U12798 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10256), .Z(n15245) );
  NOR2_X1 U12799 ( .A1(n15246), .A2(n15245), .ZN(n15244) );
  XOR2_X1 U12800 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10258), .Z(n10335) );
  XOR2_X1 U12801 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10282), .Z(n10251) );
  OR2_X1 U12802 ( .A1(n10263), .A2(P2_U3088), .ZN(n14099) );
  INV_X1 U12803 ( .A(n14104), .ZN(n10250) );
  AOI211_X1 U12804 ( .C1(n10252), .C2(n10251), .A(n10276), .B(n15298), .ZN(
        n10268) );
  XNOR2_X1 U12805 ( .A(n10254), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n15240) );
  AND3_X1 U12806 ( .A1(n15240), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n15237) );
  AOI21_X1 U12807 ( .B1(n10255), .B2(P2_REG2_REG_1__SCAN_IN), .A(n15237), .ZN(
        n15251) );
  INV_X1 U12808 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10257) );
  MUX2_X1 U12809 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10257), .S(n10256), .Z(
        n15250) );
  NOR2_X1 U12810 ( .A1(n15251), .A2(n15250), .ZN(n15249) );
  AND2_X1 U12811 ( .A1(n15248), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10339) );
  INV_X1 U12812 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10738) );
  MUX2_X1 U12813 ( .A(n10738), .B(P2_REG2_REG_3__SCAN_IN), .S(n10258), .Z(
        n10338) );
  OAI21_X1 U12814 ( .B1(n15249), .B2(n10339), .A(n10338), .ZN(n10337) );
  NAND2_X1 U12815 ( .A1(n10344), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10261) );
  INV_X1 U12816 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10259) );
  MUX2_X1 U12817 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10259), .S(n10282), .Z(
        n10260) );
  AOI21_X1 U12818 ( .B1(n10337), .B2(n10261), .A(n10260), .ZN(n10325) );
  AND3_X1 U12819 ( .A1(n10337), .A2(n10261), .A3(n10260), .ZN(n10262) );
  NOR3_X1 U12820 ( .A1(n15279), .A2(n10325), .A3(n10262), .ZN(n10267) );
  NAND2_X1 U12821 ( .A1(n10263), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10264) );
  NAND2_X1 U12822 ( .A1(n15289), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12823 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10711) );
  OAI211_X1 U12824 ( .C1(n15272), .C2(n10282), .A(n10265), .B(n10711), .ZN(
        n10266) );
  OR3_X1 U12825 ( .A1(n10268), .A2(n10267), .A3(n10266), .ZN(P2_U3218) );
  NAND2_X1 U12826 ( .A1(n12491), .A2(n10665), .ZN(n10269) );
  OAI21_X1 U12827 ( .B1(n10665), .B2(n10270), .A(n10269), .ZN(P3_U3499) );
  NAND2_X1 U12828 ( .A1(n11805), .A2(n10665), .ZN(n10271) );
  OAI21_X1 U12829 ( .B1(n10665), .B2(n10272), .A(n10271), .ZN(P3_U3503) );
  INV_X1 U12830 ( .A(n14826), .ZN(n13043) );
  INV_X1 U12831 ( .A(n10273), .ZN(n10275) );
  INV_X1 U12832 ( .A(SI_18_), .ZN(n10274) );
  OAI222_X1 U12833 ( .A1(n13043), .A2(P3_U3151), .B1(n13439), .B2(n10275), 
        .C1(n10274), .C2(n13430), .ZN(P3_U3277) );
  INV_X1 U12834 ( .A(n10283), .ZN(n10331) );
  INV_X1 U12835 ( .A(n10282), .ZN(n10277) );
  AOI21_X1 U12836 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n10277), .A(n10276), .ZN(
        n10321) );
  XOR2_X1 U12837 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10283), .Z(n10320) );
  NOR2_X1 U12838 ( .A1(n10321), .A2(n10320), .ZN(n10319) );
  INV_X1 U12839 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10278) );
  MUX2_X1 U12840 ( .A(n10278), .B(P2_REG1_REG_6__SCAN_IN), .S(n10284), .Z(
        n10297) );
  NOR2_X1 U12841 ( .A1(n10298), .A2(n10297), .ZN(n10296) );
  INV_X1 U12842 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10279) );
  MUX2_X1 U12843 ( .A(n10279), .B(P2_REG1_REG_7__SCAN_IN), .S(n10397), .Z(
        n10280) );
  AOI211_X1 U12844 ( .C1(n10281), .C2(n10280), .A(n15298), .B(n10393), .ZN(
        n10295) );
  NOR2_X1 U12845 ( .A1(n10282), .A2(n10259), .ZN(n10324) );
  INV_X1 U12846 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10841) );
  MUX2_X1 U12847 ( .A(n10841), .B(P2_REG2_REG_5__SCAN_IN), .S(n10283), .Z(
        n10323) );
  OAI21_X1 U12848 ( .B1(n10325), .B2(n10324), .A(n10323), .ZN(n10322) );
  NAND2_X1 U12849 ( .A1(n10331), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10300) );
  INV_X1 U12850 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10285) );
  MUX2_X1 U12851 ( .A(n10285), .B(P2_REG2_REG_6__SCAN_IN), .S(n10284), .Z(
        n10299) );
  AOI21_X1 U12852 ( .B1(n10322), .B2(n10300), .A(n10299), .ZN(n10302) );
  NOR2_X1 U12853 ( .A1(n10304), .A2(n10285), .ZN(n10288) );
  INV_X1 U12854 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10286) );
  MUX2_X1 U12855 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10286), .S(n10397), .Z(
        n10287) );
  OAI21_X1 U12856 ( .B1(n10302), .B2(n10288), .A(n10287), .ZN(n10401) );
  INV_X1 U12857 ( .A(n10401), .ZN(n10290) );
  NOR3_X1 U12858 ( .A1(n10302), .A2(n10288), .A3(n10287), .ZN(n10289) );
  NOR3_X1 U12859 ( .A1(n15279), .A2(n10290), .A3(n10289), .ZN(n10294) );
  NAND2_X1 U12860 ( .A1(n15289), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U12861 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11410) );
  OAI211_X1 U12862 ( .C1(n15272), .C2(n10292), .A(n10291), .B(n11410), .ZN(
        n10293) );
  OR3_X1 U12863 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(P2_U3221) );
  AND3_X1 U12864 ( .A1(n10322), .A2(n10300), .A3(n10299), .ZN(n10301) );
  NOR3_X1 U12865 ( .A1(n15279), .A2(n10302), .A3(n10301), .ZN(n10306) );
  NAND2_X1 U12866 ( .A1(n15289), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U12867 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11197) );
  OAI211_X1 U12868 ( .C1(n15272), .C2(n10304), .A(n10303), .B(n11197), .ZN(
        n10305) );
  OR3_X1 U12869 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(P2_U3220) );
  OAI222_X1 U12870 ( .A1(n13439), .A2(n10309), .B1(n13441), .B2(n10308), .C1(
        n6665), .C2(n13054), .ZN(P3_U3276) );
  INV_X1 U12871 ( .A(n11849), .ZN(n10311) );
  INV_X1 U12872 ( .A(n11703), .ZN(n10318) );
  OAI222_X1 U12873 ( .A1(P2_U3088), .A2(n10311), .B1(n14111), .B2(n10318), 
        .C1(n10310), .C2(n14106), .ZN(P2_U3314) );
  NAND2_X1 U12874 ( .A1(n10312), .A2(n10046), .ZN(n10313) );
  NAND2_X1 U12875 ( .A1(n10313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U12876 ( .A1(n10315), .A2(n10314), .ZN(n10439) );
  OR2_X1 U12877 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  INV_X1 U12878 ( .A(n11704), .ZN(n14362) );
  OAI222_X1 U12879 ( .A1(P1_U3086), .A2(n14362), .B1(n14780), .B2(n10318), 
        .C1(n10317), .C2(n14772), .ZN(P1_U3342) );
  AOI211_X1 U12880 ( .C1(n10321), .C2(n10320), .A(n10319), .B(n15298), .ZN(
        n10329) );
  INV_X1 U12881 ( .A(n10322), .ZN(n10327) );
  NOR3_X1 U12882 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10326) );
  NOR3_X1 U12883 ( .A1(n15279), .A2(n10327), .A3(n10326), .ZN(n10328) );
  NOR2_X1 U12884 ( .A1(n10329), .A2(n10328), .ZN(n10333) );
  NAND2_X1 U12885 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10868) );
  INV_X1 U12886 ( .A(n10868), .ZN(n10330) );
  AOI21_X1 U12887 ( .B1(n15305), .B2(n10331), .A(n10330), .ZN(n10332) );
  OAI211_X1 U12888 ( .C1(n15313), .C2(n15690), .A(n10333), .B(n10332), .ZN(
        P2_U3219) );
  INV_X1 U12889 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10347) );
  AOI211_X1 U12890 ( .C1(n10336), .C2(n10335), .A(n10334), .B(n15298), .ZN(
        n10343) );
  INV_X1 U12891 ( .A(n10337), .ZN(n10341) );
  NOR3_X1 U12892 ( .A1(n15249), .A2(n10339), .A3(n10338), .ZN(n10340) );
  NOR3_X1 U12893 ( .A1(n15279), .A2(n10341), .A3(n10340), .ZN(n10342) );
  NOR2_X1 U12894 ( .A1(n10343), .A2(n10342), .ZN(n10346) );
  AOI22_X1 U12895 ( .A1(n15305), .A2(n10344), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10345) );
  OAI211_X1 U12896 ( .C1(n15313), .C2(n10347), .A(n10346), .B(n10345), .ZN(
        P2_U3217) );
  INV_X1 U12897 ( .A(n15064), .ZN(n14365) );
  NOR2_X1 U12898 ( .A1(n14365), .A2(n14285), .ZN(P1_U3085) );
  INV_X1 U12899 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15218) );
  MUX2_X1 U12900 ( .A(n15218), .B(P1_REG1_REG_5__SCAN_IN), .S(n10963), .Z(
        n10355) );
  INV_X1 U12901 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10353) );
  AND2_X1 U12902 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14274) );
  INV_X1 U12903 ( .A(n10595), .ZN(n14272) );
  NAND2_X1 U12904 ( .A1(n14272), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12905 ( .A1(n14273), .A2(n10348), .ZN(n14295) );
  XNOR2_X1 U12906 ( .A(n14288), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U12907 ( .A1(n14295), .A2(n14296), .ZN(n14294) );
  INV_X1 U12908 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10349) );
  OR2_X1 U12909 ( .A1(n14288), .A2(n10349), .ZN(n10350) );
  NAND2_X1 U12910 ( .A1(n14294), .A2(n10350), .ZN(n14301) );
  INV_X1 U12911 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10351) );
  XNOR2_X1 U12912 ( .A(n14307), .B(n10351), .ZN(n14302) );
  NAND2_X1 U12913 ( .A1(n14301), .A2(n14302), .ZN(n14300) );
  NAND2_X1 U12914 ( .A1(n14307), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12915 ( .A1(n14300), .A2(n10352), .ZN(n14317) );
  XNOR2_X1 U12916 ( .A(n10923), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U12917 ( .A1(n14317), .A2(n14318), .ZN(n14316) );
  AOI21_X1 U12918 ( .B1(n10355), .B2(n10354), .A(n10467), .ZN(n10372) );
  NAND2_X1 U12919 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U12920 ( .B1(n15064), .B2(n8878), .A(n11552), .ZN(n10357) );
  AOI21_X1 U12921 ( .B1(n10963), .B2(n14398), .A(n10357), .ZN(n10371) );
  NOR2_X1 U12922 ( .A1(n10202), .A2(n14776), .ZN(n10358) );
  INV_X1 U12923 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11423) );
  MUX2_X1 U12924 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11423), .S(n14307), .Z(
        n10362) );
  XNOR2_X1 U12925 ( .A(n10595), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14277) );
  AND2_X1 U12926 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14282) );
  NAND2_X1 U12927 ( .A1(n14277), .A2(n14282), .ZN(n14276) );
  NAND2_X1 U12928 ( .A1(n14272), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U12929 ( .A1(n14276), .A2(n10360), .ZN(n14292) );
  INV_X1 U12930 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11400) );
  MUX2_X1 U12931 ( .A(n11400), .B(P1_REG2_REG_2__SCAN_IN), .S(n14288), .Z(
        n14293) );
  NAND2_X1 U12932 ( .A1(n14292), .A2(n14293), .ZN(n14304) );
  OR2_X1 U12933 ( .A1(n14288), .A2(n11400), .ZN(n14303) );
  NAND2_X1 U12934 ( .A1(n14304), .A2(n14303), .ZN(n10361) );
  NAND2_X1 U12935 ( .A1(n10362), .A2(n10361), .ZN(n14320) );
  NAND2_X1 U12936 ( .A1(n14307), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14319) );
  INV_X1 U12937 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10363) );
  MUX2_X1 U12938 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10363), .S(n10923), .Z(
        n14321) );
  AOI21_X1 U12939 ( .B1(n14320), .B2(n14319), .A(n14321), .ZN(n10365) );
  NOR2_X1 U12940 ( .A1(n10923), .A2(n10363), .ZN(n10366) );
  INV_X1 U12941 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11370) );
  MUX2_X1 U12942 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11370), .S(n10963), .Z(
        n10364) );
  OAI21_X1 U12943 ( .B1(n10365), .B2(n10366), .A(n10364), .ZN(n14338) );
  INV_X1 U12944 ( .A(n10365), .ZN(n14323) );
  INV_X1 U12945 ( .A(n10366), .ZN(n10368) );
  MUX2_X1 U12946 ( .A(n11370), .B(P1_REG2_REG_5__SCAN_IN), .S(n10963), .Z(
        n10367) );
  NAND3_X1 U12947 ( .A1(n14323), .A2(n10368), .A3(n10367), .ZN(n10369) );
  NAND3_X1 U12948 ( .A1(n14400), .A2(n14338), .A3(n10369), .ZN(n10370) );
  OAI211_X1 U12949 ( .C1(n10372), .C2(n14396), .A(n10371), .B(n10370), .ZN(
        P1_U3248) );
  NAND2_X1 U12950 ( .A1(n12873), .A2(n10665), .ZN(n10373) );
  OAI21_X1 U12951 ( .B1(n10665), .B2(n10374), .A(n10373), .ZN(P3_U3514) );
  OAI21_X1 U12952 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n10378) );
  NAND2_X1 U12953 ( .A1(n10378), .A2(n13632), .ZN(n10382) );
  OAI22_X1 U12954 ( .A1(n10380), .A2(n13447), .B1(n13449), .B2(n10379), .ZN(
        n10425) );
  AOI22_X1 U12955 ( .A1(n10425), .A2(n13641), .B1(n12393), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10381) );
  OAI211_X1 U12956 ( .C1(n10422), .C2(n13644), .A(n10382), .B(n10381), .ZN(
        P2_U3209) );
  NAND2_X1 U12957 ( .A1(n15609), .A2(n10665), .ZN(n10383) );
  OAI21_X1 U12958 ( .B1(n10665), .B2(n10384), .A(n10383), .ZN(P3_U3491) );
  NAND2_X1 U12959 ( .A1(n15529), .A2(n10665), .ZN(n10385) );
  OAI21_X1 U12960 ( .B1(n10665), .B2(n10386), .A(n10385), .ZN(P3_U3502) );
  NAND2_X1 U12961 ( .A1(n10557), .A2(n10665), .ZN(n10387) );
  OAI21_X1 U12962 ( .B1(P3_U3897), .B2(n10388), .A(n10387), .ZN(P3_U3494) );
  NAND2_X1 U12963 ( .A1(n15608), .A2(n10665), .ZN(n10389) );
  OAI21_X1 U12964 ( .B1(n10665), .B2(n10390), .A(n10389), .ZN(P3_U3493) );
  NAND2_X1 U12965 ( .A1(n15587), .A2(n10665), .ZN(n10391) );
  OAI21_X1 U12966 ( .B1(n10665), .B2(n10392), .A(n10391), .ZN(P3_U3492) );
  INV_X1 U12967 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10394) );
  MUX2_X1 U12968 ( .A(n10394), .B(P2_REG1_REG_8__SCAN_IN), .S(n11106), .Z(
        n10395) );
  AOI211_X1 U12969 ( .C1(n10396), .C2(n10395), .A(n15298), .B(n11099), .ZN(
        n10406) );
  NAND2_X1 U12970 ( .A1(n10397), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10400) );
  INV_X1 U12971 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10398) );
  MUX2_X1 U12972 ( .A(n10398), .B(P2_REG2_REG_8__SCAN_IN), .S(n11106), .Z(
        n10399) );
  AOI21_X1 U12973 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(n11105) );
  AND3_X1 U12974 ( .A1(n10401), .A2(n10400), .A3(n10399), .ZN(n10402) );
  NOR3_X1 U12975 ( .A1(n15279), .A2(n11105), .A3(n10402), .ZN(n10405) );
  AND2_X1 U12976 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13496) );
  AOI21_X1 U12977 ( .B1(n15305), .B2(n11106), .A(n13496), .ZN(n10403) );
  OAI21_X1 U12978 ( .B1(n15313), .B2(n14797), .A(n10403), .ZN(n10404) );
  OR3_X1 U12979 ( .A1(n10406), .A2(n10405), .A3(n10404), .ZN(P2_U3222) );
  XNOR2_X1 U12980 ( .A(n10408), .B(n10407), .ZN(n10412) );
  OAI22_X1 U12981 ( .A1(n10409), .A2(n13447), .B1(n13449), .B2(n6907), .ZN(
        n10736) );
  AOI22_X1 U12982 ( .A1(n10736), .A2(n13641), .B1(n10742), .B2(n13628), .ZN(
        n10411) );
  MUX2_X1 U12983 ( .A(n13638), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n10410) );
  OAI211_X1 U12984 ( .C1(n10412), .C2(n13630), .A(n10411), .B(n10410), .ZN(
        P2_U3190) );
  NAND2_X1 U12985 ( .A1(n15609), .A2(n10664), .ZN(n12451) );
  INV_X1 U12986 ( .A(n12451), .ZN(n10414) );
  NOR2_X1 U12987 ( .A1(n10413), .A2(n10414), .ZN(n12428) );
  AOI22_X1 U12988 ( .A1(n12936), .A2(n15587), .B1(n12943), .B2(n10447), .ZN(
        n10416) );
  OR2_X1 U12989 ( .A1(n12938), .A2(n6665), .ZN(n12618) );
  NAND2_X1 U12990 ( .A1(n12618), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10415) );
  OAI211_X1 U12991 ( .C1(n12428), .C2(n12945), .A(n10416), .B(n10415), .ZN(
        P3_U3172) );
  NAND2_X1 U12992 ( .A1(n13115), .A2(n10665), .ZN(n10417) );
  OAI21_X1 U12993 ( .B1(n10665), .B2(n10418), .A(n10417), .ZN(P3_U3515) );
  XNOR2_X1 U12994 ( .A(n10419), .B(n10420), .ZN(n15321) );
  INV_X1 U12995 ( .A(n15398), .ZN(n15409) );
  INV_X1 U12996 ( .A(n11093), .ZN(n10421) );
  OAI211_X1 U12997 ( .C1(n10422), .C2(n10421), .A(n9576), .B(n10741), .ZN(
        n15317) );
  OAI21_X1 U12998 ( .B1(n15409), .B2(n10422), .A(n15317), .ZN(n10428) );
  XNOR2_X1 U12999 ( .A(n10423), .B(n10424), .ZN(n10426) );
  AOI21_X1 U13000 ( .B1(n10426), .B2(n14882), .A(n10425), .ZN(n15324) );
  INV_X1 U13001 ( .A(n15324), .ZN(n10427) );
  AOI211_X1 U13002 ( .C1(n15321), .C2(n15370), .A(n10428), .B(n10427), .ZN(
        n15374) );
  NAND2_X1 U13003 ( .A1(n15429), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10429) );
  OAI21_X1 U13004 ( .B1(n15374), .B2(n15429), .A(n10429), .ZN(P2_U3501) );
  INV_X1 U13005 ( .A(n12086), .ZN(n10437) );
  INV_X1 U13006 ( .A(n13703), .ZN(n13695) );
  OAI222_X1 U13007 ( .A1(n14106), .A2(n10430), .B1(n14111), .B2(n10437), .C1(
        n13695), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13008 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U13009 ( .A1(n10432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10434) );
  MUX2_X1 U13010 ( .A(n10434), .B(P1_IR_REG_31__SCAN_IN), .S(n10433), .Z(
        n10435) );
  NAND2_X1 U13011 ( .A1(n10435), .A2(n10055), .ZN(n11756) );
  OAI222_X1 U13012 ( .A1(P1_U3086), .A2(n11756), .B1(n14780), .B2(n10437), 
        .C1(n10436), .C2(n14772), .ZN(P1_U3339) );
  INV_X1 U13013 ( .A(n11915), .ZN(n10442) );
  INV_X1 U13014 ( .A(n13681), .ZN(n11855) );
  OAI222_X1 U13015 ( .A1(n14106), .A2(n10438), .B1(n14111), .B2(n10442), .C1(
        n11855), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U13016 ( .A1(n10439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10440) );
  XNOR2_X1 U13017 ( .A(n10440), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11916) );
  INV_X1 U13018 ( .A(n11916), .ZN(n11742) );
  OAI222_X1 U13019 ( .A1(P1_U3086), .A2(n11742), .B1(n14780), .B2(n10442), 
        .C1(n10441), .C2(n14772), .ZN(P1_U3341) );
  AND2_X1 U13020 ( .A1(n10443), .A2(n15594), .ZN(n10444) );
  OR2_X1 U13021 ( .A1(n12428), .A2(n10444), .ZN(n10446) );
  INV_X1 U13022 ( .A(n15588), .ZN(n15607) );
  NAND2_X1 U13023 ( .A1(n15587), .A2(n15607), .ZN(n10445) );
  NAND2_X1 U13024 ( .A1(n10446), .A2(n10445), .ZN(n10660) );
  AND2_X1 U13025 ( .A1(n10447), .A2(n15583), .ZN(n10448) );
  NOR2_X1 U13026 ( .A1(n10660), .A2(n10448), .ZN(n10553) );
  NAND2_X1 U13027 ( .A1(n15672), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n10449) );
  OAI21_X1 U13028 ( .B1(n10553), .B2(n15672), .A(n10449), .ZN(P3_U3390) );
  NAND2_X1 U13029 ( .A1(n10055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10450) );
  XNOR2_X1 U13030 ( .A(n10450), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14375) );
  INV_X1 U13031 ( .A(n14375), .ZN(n14373) );
  INV_X1 U13032 ( .A(n12090), .ZN(n10452) );
  OAI222_X1 U13033 ( .A1(P1_U3086), .A2(n14373), .B1(n14780), .B2(n10452), 
        .C1(n10451), .C2(n14772), .ZN(P1_U3338) );
  INV_X1 U13034 ( .A(n15304), .ZN(n13697) );
  OAI222_X1 U13035 ( .A1(n14106), .A2(n10453), .B1(n14111), .B2(n10452), .C1(
        n13697), .C2(P2_U3088), .ZN(P2_U3310) );
  AOI21_X1 U13036 ( .B1(n10455), .B2(n9751), .A(n10454), .ZN(n10466) );
  INV_X1 U13037 ( .A(n10456), .ZN(n10458) );
  NAND4_X1 U13038 ( .A1(n10459), .A2(P2_STATE_REG_SCAN_IN), .A3(n10458), .A4(
        n10457), .ZN(n10460) );
  INV_X1 U13039 ( .A(n10461), .ZN(n10731) );
  NOR2_X1 U13040 ( .A1(n6674), .A2(n10731), .ZN(n11298) );
  INV_X1 U13041 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n15235) );
  INV_X1 U13042 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10462) );
  OAI22_X1 U13043 ( .A1(n13963), .A2(n15235), .B1(n10462), .B2(n13957), .ZN(
        n10463) );
  AOI21_X1 U13044 ( .B1(n10464), .B2(n11298), .A(n10463), .ZN(n10465) );
  OAI21_X1 U13045 ( .B1(n10466), .B2(n6674), .A(n10465), .ZN(P2_U3265) );
  INV_X1 U13046 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n15019) );
  MUX2_X1 U13047 ( .A(n15019), .B(P1_REG1_REG_11__SCAN_IN), .S(n11455), .Z(
        n10476) );
  INV_X1 U13048 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10474) );
  INV_X1 U13049 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10473) );
  INV_X1 U13050 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10472) );
  INV_X1 U13051 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10471) );
  INV_X1 U13052 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10469) );
  XOR2_X1 U13053 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10969), .Z(n14334) );
  OAI21_X1 U13054 ( .B1(n14329), .B2(n10469), .A(n14332), .ZN(n14347) );
  MUX2_X1 U13055 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10471), .S(n14350), .Z(
        n14348) );
  NAND2_X1 U13056 ( .A1(n14347), .A2(n14348), .ZN(n14346) );
  OAI21_X1 U13057 ( .B1(n10471), .B2(n10470), .A(n14346), .ZN(n10493) );
  MUX2_X1 U13058 ( .A(n10472), .B(P1_REG1_REG_8__SCAN_IN), .S(n10994), .Z(
        n10494) );
  MUX2_X1 U13059 ( .A(n10473), .B(P1_REG1_REG_9__SCAN_IN), .S(n11265), .Z(
        n10534) );
  MUX2_X1 U13060 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10474), .S(n11471), .Z(
        n10526) );
  NAND2_X1 U13061 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  OAI21_X1 U13062 ( .B1(n10522), .B2(n10474), .A(n10525), .ZN(n10475) );
  AOI21_X1 U13063 ( .B1(n10476), .B2(n10475), .A(n10505), .ZN(n10491) );
  NAND2_X1 U13064 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14982)
         );
  INV_X1 U13065 ( .A(n14982), .ZN(n10478) );
  NOR2_X1 U13066 ( .A1(n15055), .A2(n10512), .ZN(n10477) );
  AOI211_X1 U13067 ( .C1(n14365), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10478), 
        .B(n10477), .ZN(n10490) );
  NAND2_X1 U13068 ( .A1(n10963), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14337) );
  INV_X1 U13069 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10479) );
  MUX2_X1 U13070 ( .A(n10479), .B(P1_REG2_REG_6__SCAN_IN), .S(n10969), .Z(
        n14336) );
  AOI21_X1 U13071 ( .B1(n14338), .B2(n14337), .A(n14336), .ZN(n14335) );
  NOR2_X1 U13072 ( .A1(n14329), .A2(n10479), .ZN(n14349) );
  INV_X1 U13073 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11254) );
  MUX2_X1 U13074 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11254), .S(n14350), .Z(
        n10480) );
  OAI21_X1 U13075 ( .B1(n14335), .B2(n14349), .A(n10480), .ZN(n14355) );
  NAND2_X1 U13076 ( .A1(n14350), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10499) );
  INV_X1 U13077 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10481) );
  MUX2_X1 U13078 ( .A(n10481), .B(P1_REG2_REG_8__SCAN_IN), .S(n10994), .Z(
        n10498) );
  AOI21_X1 U13079 ( .B1(n14355), .B2(n10499), .A(n10498), .ZN(n10543) );
  NOR2_X1 U13080 ( .A1(n10495), .A2(n10481), .ZN(n10538) );
  INV_X1 U13081 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11276) );
  MUX2_X1 U13082 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11276), .S(n11265), .Z(
        n10482) );
  OAI21_X1 U13083 ( .B1(n10543), .B2(n10538), .A(n10482), .ZN(n10541) );
  NAND2_X1 U13084 ( .A1(n11265), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10520) );
  INV_X1 U13085 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10483) );
  MUX2_X1 U13086 ( .A(n10483), .B(P1_REG2_REG_10__SCAN_IN), .S(n11471), .Z(
        n10519) );
  AOI21_X1 U13087 ( .B1(n10541), .B2(n10520), .A(n10519), .ZN(n10531) );
  NOR2_X1 U13088 ( .A1(n10522), .A2(n10483), .ZN(n10487) );
  INV_X1 U13089 ( .A(n10487), .ZN(n10485) );
  INV_X1 U13090 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10511) );
  MUX2_X1 U13091 ( .A(n10511), .B(P1_REG2_REG_11__SCAN_IN), .S(n11455), .Z(
        n10484) );
  NAND2_X1 U13092 ( .A1(n10485), .A2(n10484), .ZN(n10488) );
  MUX2_X1 U13093 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10511), .S(n11455), .Z(
        n10486) );
  OAI21_X1 U13094 ( .B1(n10531), .B2(n10487), .A(n10486), .ZN(n10510) );
  OAI211_X1 U13095 ( .C1(n10531), .C2(n10488), .A(n14400), .B(n10510), .ZN(
        n10489) );
  OAI211_X1 U13096 ( .C1(n10491), .C2(n14396), .A(n10490), .B(n10489), .ZN(
        P1_U3254) );
  AOI21_X1 U13097 ( .B1(n10494), .B2(n10493), .A(n10492), .ZN(n10504) );
  AND2_X1 U13098 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10497) );
  NOR2_X1 U13099 ( .A1(n15055), .A2(n10495), .ZN(n10496) );
  AOI211_X1 U13100 ( .C1(n14365), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10497), .B(
        n10496), .ZN(n10503) );
  INV_X1 U13101 ( .A(n10543), .ZN(n10501) );
  NAND3_X1 U13102 ( .A1(n14355), .A2(n10499), .A3(n10498), .ZN(n10500) );
  NAND3_X1 U13103 ( .A1(n14400), .A2(n10501), .A3(n10500), .ZN(n10502) );
  OAI211_X1 U13104 ( .C1(n10504), .C2(n14396), .A(n10503), .B(n10502), .ZN(
        P1_U3251) );
  INV_X1 U13105 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11702) );
  MUX2_X1 U13106 ( .A(n11702), .B(P1_REG1_REG_12__SCAN_IN), .S(n11660), .Z(
        n10507) );
  AOI21_X1 U13107 ( .B1(n10507), .B2(n10506), .A(n11035), .ZN(n10518) );
  AND2_X1 U13108 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14162) );
  NOR2_X1 U13109 ( .A1(n15055), .A2(n11041), .ZN(n10508) );
  AOI211_X1 U13110 ( .C1(n14365), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n14162), 
        .B(n10508), .ZN(n10517) );
  INV_X1 U13111 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10509) );
  MUX2_X1 U13112 ( .A(n10509), .B(P1_REG2_REG_12__SCAN_IN), .S(n11660), .Z(
        n10514) );
  OAI21_X1 U13113 ( .B1(n10512), .B2(n10511), .A(n10510), .ZN(n10513) );
  NOR2_X1 U13114 ( .A1(n10513), .A2(n10514), .ZN(n11040) );
  AOI21_X1 U13115 ( .B1(n10514), .B2(n10513), .A(n11040), .ZN(n10515) );
  INV_X1 U13116 ( .A(n14400), .ZN(n15057) );
  OR2_X1 U13117 ( .A1(n10515), .A2(n15057), .ZN(n10516) );
  OAI211_X1 U13118 ( .C1(n10518), .C2(n14396), .A(n10517), .B(n10516), .ZN(
        P1_U3255) );
  NAND3_X1 U13119 ( .A1(n10541), .A2(n10520), .A3(n10519), .ZN(n10521) );
  NAND2_X1 U13120 ( .A1(n14400), .A2(n10521), .ZN(n10530) );
  INV_X1 U13121 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n14136) );
  NOR2_X1 U13122 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14136), .ZN(n10524) );
  NOR2_X1 U13123 ( .A1(n15055), .A2(n10522), .ZN(n10523) );
  AOI211_X1 U13124 ( .C1(n14365), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n10524), 
        .B(n10523), .ZN(n10529) );
  OAI211_X1 U13125 ( .C1(n10527), .C2(n10526), .A(n10525), .B(n15060), .ZN(
        n10528) );
  OAI211_X1 U13126 ( .C1(n10531), .C2(n10530), .A(n10529), .B(n10528), .ZN(
        P1_U3253) );
  AOI21_X1 U13127 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n10546) );
  NOR2_X1 U13128 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11007), .ZN(n10537) );
  NOR2_X1 U13129 ( .A1(n15055), .A2(n10535), .ZN(n10536) );
  AOI211_X1 U13130 ( .C1(n14365), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10537), .B(
        n10536), .ZN(n10545) );
  MUX2_X1 U13131 ( .A(n11276), .B(P1_REG2_REG_9__SCAN_IN), .S(n11265), .Z(
        n10540) );
  INV_X1 U13132 ( .A(n10538), .ZN(n10539) );
  NAND2_X1 U13133 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  OAI211_X1 U13134 ( .C1(n10543), .C2(n10542), .A(n14400), .B(n10541), .ZN(
        n10544) );
  OAI211_X1 U13135 ( .C1(n10546), .C2(n14396), .A(n10545), .B(n10544), .ZN(
        P1_U3252) );
  NAND2_X1 U13136 ( .A1(n12874), .A2(n10665), .ZN(n10547) );
  OAI21_X1 U13137 ( .B1(n10665), .B2(n10548), .A(n10547), .ZN(P3_U3516) );
  NAND2_X1 U13138 ( .A1(n6814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10549) );
  XNOR2_X1 U13139 ( .A(n10549), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11921) );
  INV_X1 U13140 ( .A(n11921), .ZN(n15056) );
  INV_X1 U13141 ( .A(n11920), .ZN(n10551) );
  OAI222_X1 U13142 ( .A1(P1_U3086), .A2(n15056), .B1(n14780), .B2(n10551), 
        .C1(n10550), .C2(n14772), .ZN(P1_U3340) );
  OAI222_X1 U13143 ( .A1(n14106), .A2(n10552), .B1(n14111), .B2(n10551), .C1(
        n13684), .C2(P2_U3088), .ZN(P2_U3312) );
  MUX2_X1 U13144 ( .A(n10700), .B(n10553), .S(n15685), .Z(n10554) );
  INV_X1 U13145 ( .A(n10554), .ZN(P3_U3459) );
  OAI21_X1 U13146 ( .B1(n10556), .B2(n10555), .A(n10669), .ZN(n10561) );
  NAND2_X1 U13147 ( .A1(n12618), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13148 ( .A1(n12914), .A2(n15587), .B1(n10557), .B2(n12936), .ZN(
        n10558) );
  OAI211_X1 U13149 ( .C1(n12931), .C2(n15582), .A(n10559), .B(n10558), .ZN(
        n10560) );
  AOI21_X1 U13150 ( .B1(n10561), .B2(n12924), .A(n10560), .ZN(n10562) );
  INV_X1 U13151 ( .A(n10562), .ZN(P3_U3177) );
  INV_X1 U13152 ( .A(n10563), .ZN(n10565) );
  OAI222_X1 U13153 ( .A1(n6665), .A2(n10566), .B1(n13439), .B2(n10565), .C1(
        n10564), .C2(n13430), .ZN(P3_U3275) );
  XNOR2_X2 U13154 ( .A(n10569), .B(n10568), .ZN(n12189) );
  INV_X1 U13155 ( .A(SI_0_), .ZN(n10572) );
  OAI21_X1 U13156 ( .B1(n6673), .B2(n10572), .A(n10571), .ZN(n10573) );
  AND2_X1 U13157 ( .A1(n10574), .A2(n10573), .ZN(n14783) );
  MUX2_X1 U13158 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14783), .S(n10818), .Z(n12213) );
  INV_X1 U13159 ( .A(n10567), .ZN(n10577) );
  NAND2_X1 U13160 ( .A1(n12165), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10586) );
  INV_X1 U13161 ( .A(n12378), .ZN(n10582) );
  AND2_X2 U13162 ( .A1(n10582), .A2(n10581), .ZN(n12124) );
  NAND2_X1 U13163 ( .A1(n12124), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13164 ( .A1(n12125), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10583) );
  INV_X1 U13165 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10587) );
  OAI222_X1 U13166 ( .A1(n10604), .A2(n15148), .B1(n10817), .B2(n15096), .C1(
        n10575), .C2(n10587), .ZN(n10647) );
  AND3_X1 U13167 ( .A1(n10591), .A2(n10590), .A3(n10589), .ZN(n10648) );
  NAND2_X1 U13168 ( .A1(n15149), .A2(n14527), .ZN(n10896) );
  AND2_X1 U13169 ( .A1(n10648), .A2(n11778), .ZN(n10592) );
  AND2_X1 U13170 ( .A1(n6672), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n10596) );
  OAI21_X1 U13171 ( .B1(n14283), .B2(n10597), .A(n10596), .ZN(n10598) );
  NAND2_X1 U13172 ( .A1(n12165), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13173 ( .A1(n6677), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13174 ( .A1(n6679), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13175 ( .A1(n12124), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10599) );
  NOR2_X1 U13176 ( .A1(n10604), .A2(n15107), .ZN(n10605) );
  AOI21_X1 U13177 ( .B1(n11026), .B2(n10887), .A(n10605), .ZN(n10606) );
  NAND2_X1 U13178 ( .A1(n10814), .A2(n10608), .ZN(n10609) );
  NOR2_X1 U13179 ( .A1(n10609), .A2(n10610), .ZN(n10816) );
  AOI21_X1 U13180 ( .B1(n10610), .B2(n10609), .A(n10816), .ZN(n10645) );
  NOR4_X1 U13181 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10614) );
  NOR4_X1 U13182 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10613) );
  NOR4_X1 U13183 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10612) );
  NOR4_X1 U13184 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10611) );
  NAND4_X1 U13185 ( .A1(n10614), .A2(n10613), .A3(n10612), .A4(n10611), .ZN(
        n10620) );
  NOR2_X1 U13186 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10618) );
  NOR4_X1 U13187 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10617) );
  NOR4_X1 U13188 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10616) );
  NOR4_X1 U13189 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10615) );
  NAND4_X1 U13190 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10619) );
  NOR2_X1 U13191 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  OR2_X1 U13192 ( .A1(n10624), .A2(n10621), .ZN(n10636) );
  OR2_X1 U13193 ( .A1(n10624), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10623) );
  NAND2_X1 U13194 ( .A1(n10210), .A2(n14781), .ZN(n10622) );
  OR2_X1 U13195 ( .A1(n10624), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13196 ( .A1(n10209), .A2(n14781), .ZN(n10625) );
  INV_X1 U13197 ( .A(n12189), .ZN(n10628) );
  AND2_X1 U13198 ( .A1(n12194), .A2(n10628), .ZN(n12175) );
  NAND2_X1 U13199 ( .A1(n12175), .A2(n10576), .ZN(n11229) );
  NOR2_X1 U13200 ( .A1(n15156), .A2(n12190), .ZN(n10627) );
  NAND2_X1 U13201 ( .A1(n15149), .A2(n14401), .ZN(n10629) );
  NAND2_X1 U13202 ( .A1(n10570), .A2(n10628), .ZN(n12191) );
  NAND2_X1 U13203 ( .A1(n14645), .A2(n12190), .ZN(n10640) );
  AND2_X1 U13204 ( .A1(n10944), .A2(n11224), .ZN(n10637) );
  NAND2_X1 U13205 ( .A1(n11226), .A2(n10637), .ZN(n14203) );
  INV_X1 U13206 ( .A(n14969), .ZN(n14958) );
  NAND2_X1 U13207 ( .A1(n12124), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13208 ( .A1(n10631), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10634) );
  NAND2_X1 U13209 ( .A1(n12125), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13210 ( .A1(n12165), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10632) );
  NAND4_X1 U13211 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n14269) );
  AOI22_X1 U13212 ( .A1(n14960), .A2(n15091), .B1(n14958), .B2(n14269), .ZN(
        n10644) );
  NAND2_X1 U13213 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  NAND2_X1 U13214 ( .A1(n10638), .A2(n10885), .ZN(n10642) );
  AND2_X1 U13215 ( .A1(n10642), .A2(n11218), .ZN(n14118) );
  AND2_X1 U13216 ( .A1(n10640), .A2(n10639), .ZN(n10641) );
  AND2_X1 U13217 ( .A1(n10575), .A2(n10641), .ZN(n12371) );
  NAND2_X1 U13218 ( .A1(n10642), .A2(n12371), .ZN(n11030) );
  OR2_X1 U13219 ( .A1(n11030), .A2(P1_U3086), .ZN(n10830) );
  AOI22_X1 U13220 ( .A1(n14981), .A2(n10603), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10830), .ZN(n10643) );
  OAI211_X1 U13221 ( .C1(n10645), .C2(n14976), .A(n10644), .B(n10643), .ZN(
        P1_U3222) );
  INV_X1 U13222 ( .A(n14981), .ZN(n14962) );
  AOI21_X1 U13223 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(n14281) );
  NAND2_X1 U13224 ( .A1(n14643), .A2(n10887), .ZN(n15147) );
  OAI22_X1 U13225 ( .A1(n14281), .A2(n14976), .B1(n14203), .B2(n15147), .ZN(
        n10649) );
  AOI21_X1 U13226 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10830), .A(n10649), .ZN(
        n10650) );
  OAI21_X1 U13227 ( .B1(n15148), .B2(n14962), .A(n10650), .ZN(P1_U3232) );
  INV_X1 U13228 ( .A(n10652), .ZN(n13424) );
  INV_X1 U13229 ( .A(n10651), .ZN(n10653) );
  OR2_X1 U13230 ( .A1(n10653), .A2(n10652), .ZN(n10654) );
  OAI21_X1 U13231 ( .B1(n10655), .B2(n13424), .A(n10654), .ZN(n10656) );
  INV_X1 U13232 ( .A(n10656), .ZN(n10657) );
  OR2_X1 U13233 ( .A1(n10661), .A2(n15585), .ZN(n11762) );
  INV_X1 U13234 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10701) );
  AOI21_X1 U13235 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15576), .A(n10660), .ZN(
        n10662) );
  MUX2_X1 U13236 ( .A(n10701), .B(n10662), .S(n15623), .Z(n10663) );
  OAI21_X1 U13237 ( .B1(n13289), .B2(n10664), .A(n10663), .ZN(P3_U3233) );
  NAND2_X1 U13238 ( .A1(n13116), .A2(n10665), .ZN(n10666) );
  OAI21_X1 U13239 ( .B1(n10665), .B2(n10667), .A(n10666), .ZN(P3_U3517) );
  AND2_X1 U13240 ( .A1(n10669), .A2(n10668), .ZN(n10672) );
  OAI211_X1 U13241 ( .C1(n10672), .C2(n10671), .A(n12924), .B(n10670), .ZN(
        n10676) );
  NOR2_X1 U13242 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11309), .ZN(n10797) );
  OAI22_X1 U13243 ( .A1(n10673), .A2(n12941), .B1(n11308), .B2(n12931), .ZN(
        n10674) );
  AOI211_X1 U13244 ( .C1(n12936), .C2(n11301), .A(n10797), .B(n10674), .ZN(
        n10675) );
  OAI211_X1 U13245 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12896), .A(n10676), .B(
        n10675), .ZN(P3_U3158) );
  INV_X1 U13246 ( .A(n12608), .ZN(n10677) );
  OR2_X1 U13247 ( .A1(n10678), .A2(n10677), .ZN(n10690) );
  NAND2_X1 U13248 ( .A1(n12587), .A2(n10679), .ZN(n10680) );
  AND2_X1 U13249 ( .A1(n10681), .A2(n10680), .ZN(n10688) );
  INV_X1 U13250 ( .A(n10695), .ZN(n10682) );
  NAND2_X1 U13251 ( .A1(n10695), .A2(n12990), .ZN(n13051) );
  NAND2_X1 U13252 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10691), .ZN(n10684) );
  INV_X1 U13253 ( .A(n10684), .ZN(n11188) );
  OAI21_X1 U13254 ( .B1(n10747), .B2(n11188), .A(n7758), .ZN(n10686) );
  INV_X1 U13255 ( .A(n10686), .ZN(n10687) );
  INV_X1 U13256 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10685) );
  OR2_X1 U13257 ( .A1(n10686), .A2(n10685), .ZN(n10751) );
  OAI21_X1 U13258 ( .B1(n10687), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10751), .ZN(
        n10699) );
  INV_X1 U13259 ( .A(n10688), .ZN(n10689) );
  INV_X1 U13260 ( .A(n15516), .ZN(n13014) );
  OAI22_X1 U13261 ( .A1(n13014), .A2(n8988), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15619), .ZN(n10698) );
  AND2_X1 U13262 ( .A1(n10691), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U13263 ( .A1(n8230), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10755) );
  OAI21_X1 U13264 ( .B1(n10747), .B2(n11185), .A(n10755), .ZN(n10692) );
  OR2_X1 U13265 ( .A1(n10692), .A2(n8223), .ZN(n10756) );
  NAND2_X1 U13266 ( .A1(n10692), .A2(n8223), .ZN(n10696) );
  INV_X1 U13267 ( .A(n10693), .ZN(n10694) );
  AOI21_X1 U13268 ( .B1(n10756), .B2(n10696), .A(n15523), .ZN(n10697) );
  AOI211_X1 U13269 ( .C1(n15519), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n10704) );
  MUX2_X1 U13270 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12990), .Z(n10748) );
  XNOR2_X1 U13271 ( .A(n10748), .B(n10747), .ZN(n10749) );
  MUX2_X1 U13272 ( .A(n10701), .B(n10700), .S(n12990), .Z(n11189) );
  NAND2_X1 U13273 ( .A1(n11189), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11193) );
  XNOR2_X1 U13274 ( .A(n10749), .B(n11193), .ZN(n10702) );
  NAND2_X1 U13275 ( .A1(n10702), .A2(n15508), .ZN(n10703) );
  OAI211_X1 U13276 ( .C1(n15513), .C2(n10747), .A(n10704), .B(n10703), .ZN(
        P3_U3183) );
  INV_X1 U13277 ( .A(n10705), .ZN(n10706) );
  AOI21_X1 U13278 ( .B1(n10708), .B2(n10707), .A(n10706), .ZN(n10715) );
  NAND2_X1 U13279 ( .A1(n13610), .A2(n13670), .ZN(n10710) );
  NAND2_X1 U13280 ( .A1(n13551), .A2(n13672), .ZN(n10709) );
  AND2_X1 U13281 ( .A1(n10710), .A2(n10709), .ZN(n10721) );
  NAND2_X1 U13282 ( .A1(n13588), .A2(n11056), .ZN(n10712) );
  OAI211_X1 U13283 ( .C1(n10721), .C2(n13624), .A(n10712), .B(n10711), .ZN(
        n10713) );
  AOI21_X1 U13284 ( .B1(n11057), .B2(n13628), .A(n10713), .ZN(n10714) );
  OAI21_X1 U13285 ( .B1(n10715), .B2(n13630), .A(n10714), .ZN(P2_U3202) );
  XNOR2_X1 U13286 ( .A(n10716), .B(n10720), .ZN(n11063) );
  INV_X1 U13287 ( .A(n10740), .ZN(n10718) );
  INV_X1 U13288 ( .A(n10717), .ZN(n10842) );
  AOI211_X1 U13289 ( .C1(n11057), .C2(n10718), .A(n14001), .B(n10842), .ZN(
        n11055) );
  XNOR2_X1 U13290 ( .A(n10719), .B(n10720), .ZN(n10722) );
  OAI21_X1 U13291 ( .B1(n10722), .B2(n13946), .A(n10721), .ZN(n11060) );
  AOI211_X1 U13292 ( .C1(n11063), .C2(n15370), .A(n11055), .B(n11060), .ZN(
        n10730) );
  INV_X1 U13293 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10723) );
  OAI22_X1 U13294 ( .A1(n14046), .A2(n10727), .B1(n15431), .B2(n10723), .ZN(
        n10724) );
  INV_X1 U13295 ( .A(n10724), .ZN(n10725) );
  OAI21_X1 U13296 ( .B1(n10730), .B2(n15429), .A(n10725), .ZN(P2_U3503) );
  INV_X1 U13297 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10726) );
  OAI22_X1 U13298 ( .A1(n14081), .A2(n10727), .B1(n15420), .B2(n10726), .ZN(
        n10728) );
  INV_X1 U13299 ( .A(n10728), .ZN(n10729) );
  OAI21_X1 U13300 ( .B1(n10730), .B2(n15418), .A(n10729), .ZN(P2_U3442) );
  AND2_X1 U13301 ( .A1(n15412), .A2(n10731), .ZN(n10732) );
  XNOR2_X1 U13302 ( .A(n10733), .B(n10735), .ZN(n15375) );
  XNOR2_X1 U13303 ( .A(n10734), .B(n10735), .ZN(n10737) );
  AOI21_X1 U13304 ( .B1(n10737), .B2(n14882), .A(n10736), .ZN(n15378) );
  MUX2_X1 U13305 ( .A(n15378), .B(n10738), .S(n6674), .Z(n10746) );
  AOI211_X1 U13306 ( .C1(n10742), .C2(n10741), .A(n14001), .B(n10740), .ZN(
        n15376) );
  OAI22_X1 U13307 ( .A1(n13918), .A2(n15379), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13957), .ZN(n10744) );
  AOI21_X1 U13308 ( .B1(n15319), .B2(n15376), .A(n10744), .ZN(n10745) );
  OAI211_X1 U13309 ( .C1(n13966), .C2(n15375), .A(n10746), .B(n10745), .ZN(
        P2_U3262) );
  MUX2_X1 U13310 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12990), .Z(n10766) );
  XNOR2_X1 U13311 ( .A(n10766), .B(n10779), .ZN(n10768) );
  OAI22_X1 U13312 ( .A1(n10749), .A2(n11193), .B1(n10748), .B2(n10747), .ZN(
        n10769) );
  XOR2_X1 U13313 ( .A(n10768), .B(n10769), .Z(n10765) );
  INV_X1 U13314 ( .A(n15513), .ZN(n14827) );
  MUX2_X1 U13315 ( .A(n10750), .B(P3_REG1_REG_2__SCAN_IN), .S(n10779), .Z(
        n10753) );
  NAND2_X1 U13316 ( .A1(n10751), .A2(n7758), .ZN(n10752) );
  NAND2_X1 U13317 ( .A1(n10752), .A2(n10753), .ZN(n10778) );
  OAI21_X1 U13318 ( .B1(n10753), .B2(n10752), .A(n10778), .ZN(n10754) );
  INV_X1 U13319 ( .A(n10754), .ZN(n10762) );
  INV_X1 U13320 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15604) );
  MUX2_X1 U13321 ( .A(n15604), .B(P3_REG2_REG_2__SCAN_IN), .S(n10779), .Z(
        n10758) );
  NAND2_X1 U13322 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  NAND2_X1 U13323 ( .A1(n10757), .A2(n10758), .ZN(n10775) );
  OAI21_X1 U13324 ( .B1(n10758), .B2(n10757), .A(n10775), .ZN(n10759) );
  NAND2_X1 U13325 ( .A1(n14837), .A2(n10759), .ZN(n10761) );
  AOI22_X1 U13326 ( .A1(n15516), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(n6665), .ZN(n10760) );
  OAI211_X1 U13327 ( .C1(n10762), .C2(n13051), .A(n10761), .B(n10760), .ZN(
        n10763) );
  AOI21_X1 U13328 ( .B1(n14827), .B2(n10779), .A(n10763), .ZN(n10764) );
  OAI21_X1 U13329 ( .B1(n10765), .B2(n15439), .A(n10764), .ZN(P3_U3184) );
  MUX2_X1 U13330 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12990), .Z(n11139) );
  XNOR2_X1 U13331 ( .A(n11139), .B(n11141), .ZN(n11142) );
  INV_X1 U13332 ( .A(n10766), .ZN(n10767) );
  AOI22_X1 U13333 ( .A1(n10769), .A2(n10768), .B1(n10779), .B2(n10767), .ZN(
        n10794) );
  MUX2_X1 U13334 ( .A(n11306), .B(n10770), .S(n12990), .Z(n10771) );
  XNOR2_X1 U13335 ( .A(n10771), .B(n10805), .ZN(n10795) );
  INV_X1 U13336 ( .A(n10771), .ZN(n10772) );
  XOR2_X1 U13337 ( .A(n11142), .B(n11143), .Z(n10793) );
  NAND2_X1 U13338 ( .A1(n10773), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13339 ( .A1(n11141), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n8268), .B2(
        n11120), .ZN(n11118) );
  XNOR2_X1 U13340 ( .A(n11119), .B(n11118), .ZN(n10791) );
  INV_X1 U13341 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U13342 ( .A1(n11141), .A2(n15676), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n11120), .ZN(n10784) );
  OAI21_X1 U13343 ( .B1(n10779), .B2(n10750), .A(n10778), .ZN(n10781) );
  NAND2_X1 U13344 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  XNOR2_X1 U13345 ( .A(n10781), .B(n10805), .ZN(n10799) );
  NAND2_X1 U13346 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n10799), .ZN(n10798) );
  OAI21_X1 U13347 ( .B1(n10784), .B2(n10783), .A(n11128), .ZN(n10785) );
  NAND2_X1 U13348 ( .A1(n15519), .A2(n10785), .ZN(n10788) );
  INV_X1 U13349 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10786) );
  NOR2_X1 U13350 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10786), .ZN(n10851) );
  INV_X1 U13351 ( .A(n10851), .ZN(n10787) );
  OAI211_X1 U13352 ( .C1(n13014), .C2(n7099), .A(n10788), .B(n10787), .ZN(
        n10790) );
  NOR2_X1 U13353 ( .A1(n15513), .A2(n11120), .ZN(n10789) );
  AOI211_X1 U13354 ( .C1(n14837), .C2(n10791), .A(n10790), .B(n10789), .ZN(
        n10792) );
  OAI21_X1 U13355 ( .B1(n10793), .B2(n15439), .A(n10792), .ZN(P3_U3186) );
  XOR2_X1 U13356 ( .A(n10795), .B(n10794), .Z(n10807) );
  XNOR2_X1 U13357 ( .A(n10796), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10803) );
  AOI21_X1 U13358 ( .B1(n15516), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10797), .ZN(
        n10802) );
  OAI21_X1 U13359 ( .B1(n10799), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10798), .ZN(
        n10800) );
  NAND2_X1 U13360 ( .A1(n15519), .A2(n10800), .ZN(n10801) );
  OAI211_X1 U13361 ( .C1(n15523), .C2(n10803), .A(n10802), .B(n10801), .ZN(
        n10804) );
  AOI21_X1 U13362 ( .B1(n10805), .B2(n14827), .A(n10804), .ZN(n10806) );
  OAI21_X1 U13363 ( .B1(n10807), .B2(n15439), .A(n10806), .ZN(P3_U3185) );
  NAND2_X1 U13364 ( .A1(n12928), .A2(n10665), .ZN(n10808) );
  OAI21_X1 U13365 ( .B1(n10665), .B2(n10809), .A(n10808), .ZN(P3_U3518) );
  INV_X1 U13366 ( .A(n10810), .ZN(n10812) );
  OAI222_X1 U13367 ( .A1(P3_U3151), .A2(n10813), .B1(n13439), .B2(n10812), 
        .C1(n10811), .C2(n13441), .ZN(P3_U3274) );
  INV_X1 U13368 ( .A(n10814), .ZN(n10815) );
  INV_X1 U13369 ( .A(n14269), .ZN(n15101) );
  OR2_X1 U13370 ( .A1(n12162), .A2(n10819), .ZN(n10821) );
  OR2_X1 U13371 ( .A1(n12116), .A2(n14288), .ZN(n10820) );
  INV_X1 U13372 ( .A(n11397), .ZN(n15165) );
  OAI22_X1 U13373 ( .A1(n12726), .A2(n15101), .B1(n15165), .B2(n10604), .ZN(
        n11021) );
  AOI22_X1 U13374 ( .A1(n11546), .A2(n11397), .B1(n11545), .B2(n14269), .ZN(
        n10823) );
  XNOR2_X1 U13375 ( .A(n10823), .B(n11778), .ZN(n11022) );
  AOI21_X1 U13376 ( .B1(n10825), .B2(n10824), .A(n11025), .ZN(n10833) );
  INV_X1 U13377 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13378 ( .A1(n12124), .A2(n10905), .ZN(n10829) );
  NAND2_X1 U13379 ( .A1(n6678), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13380 ( .A1(n10631), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U13381 ( .A1(n12125), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13382 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n14268) );
  OAI22_X1 U13383 ( .A1(n12226), .A2(n15102), .B1(n15097), .B2(n10888), .ZN(
        n11398) );
  AOI22_X1 U13384 ( .A1(n10830), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14214), 
        .B2(n11398), .ZN(n10832) );
  NAND2_X1 U13385 ( .A1(n14981), .A2(n11397), .ZN(n10831) );
  OAI211_X1 U13386 ( .C1(n10833), .C2(n14976), .A(n10832), .B(n10831), .ZN(
        P1_U3237) );
  XNOR2_X1 U13387 ( .A(n10834), .B(n10836), .ZN(n15383) );
  XNOR2_X1 U13388 ( .A(n10835), .B(n10836), .ZN(n10840) );
  NAND2_X1 U13389 ( .A1(n13610), .A2(n13669), .ZN(n10838) );
  NAND2_X1 U13390 ( .A1(n13622), .A2(n13671), .ZN(n10837) );
  AND2_X1 U13391 ( .A1(n10838), .A2(n10837), .ZN(n10870) );
  INV_X1 U13392 ( .A(n10870), .ZN(n10839) );
  AOI21_X1 U13393 ( .B1(n10840), .B2(n14882), .A(n10839), .ZN(n15385) );
  MUX2_X1 U13394 ( .A(n10841), .B(n15385), .S(n13963), .Z(n10847) );
  OAI211_X1 U13395 ( .C1(n10842), .C2(n15386), .A(n9576), .B(n11067), .ZN(
        n15384) );
  INV_X1 U13396 ( .A(n15384), .ZN(n10845) );
  INV_X1 U13397 ( .A(n10867), .ZN(n10843) );
  OAI22_X1 U13398 ( .A1(n13918), .A2(n15386), .B1(n13957), .B2(n10843), .ZN(
        n10844) );
  AOI21_X1 U13399 ( .B1(n15319), .B2(n10845), .A(n10844), .ZN(n10846) );
  OAI211_X1 U13400 ( .C1(n13966), .C2(n15383), .A(n10847), .B(n10846), .ZN(
        P2_U3260) );
  AOI21_X1 U13401 ( .B1(n10849), .B2(n10848), .A(n6836), .ZN(n10855) );
  OAI22_X1 U13402 ( .A1(n15589), .A2(n12941), .B1(n15574), .B2(n12931), .ZN(
        n10850) );
  AOI211_X1 U13403 ( .C1(n12936), .C2(n11505), .A(n10851), .B(n10850), .ZN(
        n10854) );
  INV_X1 U13404 ( .A(n10852), .ZN(n15575) );
  NAND2_X1 U13405 ( .A1(n12938), .A2(n15575), .ZN(n10853) );
  OAI211_X1 U13406 ( .C1(n10855), .C2(n12945), .A(n10854), .B(n10853), .ZN(
        P3_U3170) );
  INV_X1 U13407 ( .A(n13072), .ZN(n10856) );
  NAND2_X1 U13408 ( .A1(n10856), .A2(n10665), .ZN(n10857) );
  OAI21_X1 U13409 ( .B1(P3_U3897), .B2(n10858), .A(n10857), .ZN(P3_U3520) );
  NOR2_X1 U13410 ( .A1(n13441), .A2(SI_22_), .ZN(n10859) );
  AOI21_X1 U13411 ( .B1(n10860), .B2(P3_STATE_REG_SCAN_IN), .A(n10859), .ZN(
        n10861) );
  OAI21_X1 U13412 ( .B1(n10862), .B2(n13439), .A(n10861), .ZN(n10863) );
  INV_X1 U13413 ( .A(n10863), .ZN(P3_U3273) );
  OAI21_X1 U13414 ( .B1(n10866), .B2(n10865), .A(n10864), .ZN(n10873) );
  NOR2_X1 U13415 ( .A1(n13644), .A2(n15386), .ZN(n10872) );
  NAND2_X1 U13416 ( .A1(n13588), .A2(n10867), .ZN(n10869) );
  OAI211_X1 U13417 ( .C1(n10870), .C2(n13624), .A(n10869), .B(n10868), .ZN(
        n10871) );
  AOI211_X1 U13418 ( .C1(n10873), .C2(n13632), .A(n10872), .B(n10871), .ZN(
        n10874) );
  INV_X1 U13419 ( .A(n10874), .ZN(P2_U3199) );
  INV_X1 U13420 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13421 ( .A1(n8224), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10878) );
  INV_X1 U13422 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n10875) );
  OR2_X1 U13423 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  OAI211_X1 U13424 ( .C1(n10879), .C2(n8245), .A(n10878), .B(n10877), .ZN(
        n10880) );
  INV_X1 U13425 ( .A(n10880), .ZN(n10881) );
  AND2_X1 U13426 ( .A1(n10882), .A2(n10881), .ZN(n13058) );
  INV_X1 U13427 ( .A(n13058), .ZN(n12421) );
  NAND2_X1 U13428 ( .A1(n12421), .A2(n10665), .ZN(n10883) );
  OAI21_X1 U13429 ( .B1(P3_U3897), .B2(n10884), .A(n10883), .ZN(P3_U3522) );
  INV_X1 U13430 ( .A(n10885), .ZN(n11217) );
  NOR2_X1 U13431 ( .A1(n11224), .A2(n11217), .ZN(n10886) );
  AND2_X1 U13432 ( .A1(n11226), .A2(n10886), .ZN(n10945) );
  INV_X1 U13433 ( .A(n10944), .ZN(n11225) );
  INV_X1 U13434 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U13435 ( .A1(n10888), .A2(n10603), .ZN(n12215) );
  NAND2_X1 U13436 ( .A1(n15091), .A2(n12213), .ZN(n15085) );
  NAND2_X1 U13437 ( .A1(n10888), .A2(n15107), .ZN(n10889) );
  INV_X1 U13438 ( .A(n12220), .ZN(n11392) );
  NAND2_X1 U13439 ( .A1(n11393), .A2(n11392), .ZN(n11391) );
  NAND2_X1 U13440 ( .A1(n15101), .A2(n15165), .ZN(n10890) );
  NAND2_X1 U13441 ( .A1(n11391), .A2(n10890), .ZN(n10893) );
  INV_X2 U13442 ( .A(n12162), .ZN(n12092) );
  XNOR2_X1 U13443 ( .A(n14268), .B(n12227), .ZN(n12224) );
  INV_X1 U13444 ( .A(n12224), .ZN(n10902) );
  NAND2_X1 U13445 ( .A1(n10893), .A2(n10902), .ZN(n10922) );
  OAI21_X1 U13446 ( .B1(n10893), .B2(n10902), .A(n10922), .ZN(n10913) );
  INV_X1 U13447 ( .A(n10913), .ZN(n11426) );
  NAND2_X1 U13448 ( .A1(n10894), .A2(n14401), .ZN(n15197) );
  OR2_X1 U13449 ( .A1(n10896), .A2(n10895), .ZN(n10897) );
  NAND2_X1 U13450 ( .A1(n14997), .A2(n14527), .ZN(n15198) );
  INV_X1 U13451 ( .A(n15198), .ZN(n15072) );
  NOR2_X1 U13452 ( .A1(n15091), .A2(n15148), .ZN(n10898) );
  NAND2_X1 U13453 ( .A1(n12218), .A2(n10898), .ZN(n10899) );
  NAND2_X1 U13454 ( .A1(n10899), .A2(n12215), .ZN(n12219) );
  NAND2_X1 U13455 ( .A1(n12219), .A2(n12220), .ZN(n10901) );
  NAND2_X1 U13456 ( .A1(n15101), .A2(n11397), .ZN(n10900) );
  NAND2_X1 U13457 ( .A1(n10901), .A2(n10900), .ZN(n10926) );
  XNOR2_X1 U13458 ( .A(n10926), .B(n10902), .ZN(n10903) );
  NOR2_X1 U13459 ( .A1(n10903), .A2(n15145), .ZN(n10912) );
  NAND2_X1 U13460 ( .A1(n12125), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10910) );
  NAND2_X1 U13461 ( .A1(n6678), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10909) );
  INV_X1 U13462 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10904) );
  NAND2_X1 U13463 ( .A1(n10905), .A2(n10904), .ZN(n10906) );
  NAND2_X1 U13464 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10930) );
  AND2_X1 U13465 ( .A1(n10906), .A2(n10930), .ZN(n11355) );
  NAND2_X1 U13466 ( .A1(n12124), .A2(n11355), .ZN(n10908) );
  NAND2_X1 U13467 ( .A1(n10631), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10907) );
  OAI22_X1 U13468 ( .A1(n12235), .A2(n15102), .B1(n15097), .B2(n15101), .ZN(
        n10911) );
  AOI211_X1 U13469 ( .C1(n10913), .C2(n15072), .A(n10912), .B(n10911), .ZN(
        n11422) );
  INV_X1 U13470 ( .A(n12227), .ZN(n10920) );
  OR2_X1 U13471 ( .A1(n15090), .A2(n11397), .ZN(n11394) );
  INV_X1 U13472 ( .A(n11394), .ZN(n10915) );
  NOR2_X1 U13473 ( .A1(n11394), .A2(n12227), .ZN(n10938) );
  INV_X1 U13474 ( .A(n10938), .ZN(n10914) );
  OAI211_X1 U13475 ( .C1(n10920), .C2(n10915), .A(n10914), .B(n15077), .ZN(
        n11420) );
  INV_X1 U13476 ( .A(n11420), .ZN(n10916) );
  AOI21_X1 U13477 ( .B1(n12227), .B2(n15156), .A(n10916), .ZN(n10917) );
  OAI211_X1 U13478 ( .C1(n11426), .C2(n15197), .A(n11422), .B(n10917), .ZN(
        n10946) );
  NAND2_X1 U13479 ( .A1(n10946), .A2(n15212), .ZN(n10918) );
  OAI21_X1 U13480 ( .B1(n15212), .B2(n10919), .A(n10918), .ZN(P1_U3468) );
  INV_X1 U13481 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U13482 ( .A1(n12226), .A2(n10920), .ZN(n10921) );
  OR2_X1 U13483 ( .A1(n10109), .A2(n11914), .ZN(n10925) );
  INV_X1 U13484 ( .A(n10923), .ZN(n14315) );
  AOI22_X1 U13485 ( .A1(n12092), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12091), 
        .B2(n14315), .ZN(n10924) );
  XNOR2_X1 U13486 ( .A(n10960), .B(n12231), .ZN(n11361) );
  NAND2_X1 U13487 ( .A1(n10926), .A2(n12224), .ZN(n10928) );
  NAND2_X1 U13488 ( .A1(n12226), .A2(n12227), .ZN(n10927) );
  NAND2_X1 U13489 ( .A1(n10928), .A2(n10927), .ZN(n11005) );
  XNOR2_X1 U13490 ( .A(n11005), .B(n12231), .ZN(n10937) );
  NAND2_X1 U13491 ( .A1(n12125), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13492 ( .A1(n6678), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10934) );
  NOR2_X1 U13493 ( .A1(n10930), .A2(n10929), .ZN(n10972) );
  AND2_X1 U13494 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  NOR2_X1 U13495 ( .A1(n10972), .A2(n10931), .ZN(n11555) );
  NAND2_X1 U13496 ( .A1(n12124), .A2(n11555), .ZN(n10933) );
  NAND2_X1 U13497 ( .A1(n10631), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10932) );
  OR2_X1 U13498 ( .A1(n15102), .A2(n12241), .ZN(n10936) );
  OAI21_X1 U13499 ( .B1(n15097), .B2(n12226), .A(n10936), .ZN(n11492) );
  AOI21_X1 U13500 ( .B1(n10937), .B2(n14645), .A(n11492), .ZN(n11358) );
  INV_X1 U13501 ( .A(n12234), .ZN(n12233) );
  OAI21_X1 U13502 ( .B1(n10938), .B2(n12234), .A(n15077), .ZN(n10939) );
  OR2_X1 U13503 ( .A1(n11363), .A2(n10939), .ZN(n11356) );
  INV_X1 U13504 ( .A(n11356), .ZN(n10940) );
  AOI21_X1 U13505 ( .B1(n12233), .B2(n15156), .A(n10940), .ZN(n10941) );
  OAI211_X1 U13506 ( .C1(n11361), .C2(n15146), .A(n11358), .B(n10941), .ZN(
        n10948) );
  NAND2_X1 U13507 ( .A1(n10948), .A2(n15212), .ZN(n10942) );
  OAI21_X1 U13508 ( .B1(n15212), .B2(n10943), .A(n10942), .ZN(P1_U3471) );
  NAND2_X1 U13509 ( .A1(n10946), .A2(n15225), .ZN(n10947) );
  OAI21_X1 U13510 ( .B1(n15225), .B2(n10351), .A(n10947), .ZN(P1_U3531) );
  NAND2_X1 U13511 ( .A1(n10948), .A2(n15225), .ZN(n10949) );
  OAI21_X1 U13512 ( .B1(n15225), .B2(n10353), .A(n10949), .ZN(P1_U3532) );
  INV_X1 U13513 ( .A(n12115), .ZN(n10955) );
  INV_X1 U13514 ( .A(n13718), .ZN(n13711) );
  OAI222_X1 U13515 ( .A1(n14106), .A2(n10950), .B1(n14111), .B2(n10955), .C1(
        P2_U3088), .C2(n13711), .ZN(P2_U3309) );
  NAND2_X1 U13516 ( .A1(n6818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10951) );
  MUX2_X1 U13517 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10951), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n10954) );
  INV_X1 U13518 ( .A(n10952), .ZN(n10953) );
  NAND2_X1 U13519 ( .A1(n10954), .A2(n10953), .ZN(n14379) );
  OAI222_X1 U13520 ( .A1(n14379), .A2(P1_U3086), .B1(n14780), .B2(n10955), 
        .C1(n12117), .C2(n14772), .ZN(P1_U3337) );
  NAND2_X1 U13521 ( .A1(n10956), .A2(n10665), .ZN(n10957) );
  OAI21_X1 U13522 ( .B1(P3_U3897), .B2(n10958), .A(n10957), .ZN(P3_U3519) );
  INV_X1 U13523 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11018) );
  INV_X1 U13524 ( .A(n12235), .ZN(n14267) );
  NAND2_X1 U13525 ( .A1(n12233), .A2(n14267), .ZN(n10959) );
  NAND2_X1 U13526 ( .A1(n12234), .A2(n12235), .ZN(n10961) );
  INV_X2 U13527 ( .A(n11914), .ZN(n12161) );
  NAND2_X1 U13528 ( .A1(n10962), .A2(n12161), .ZN(n10965) );
  AOI22_X1 U13529 ( .A1(n12092), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12091), 
        .B2(n10963), .ZN(n10964) );
  INV_X1 U13530 ( .A(n12241), .ZN(n14266) );
  XNOR2_X1 U13531 ( .A(n15174), .B(n14266), .ZN(n12101) );
  NAND2_X1 U13532 ( .A1(n15174), .A2(n12241), .ZN(n10966) );
  NAND2_X1 U13533 ( .A1(n10967), .A2(n10966), .ZN(n15066) );
  NAND2_X1 U13534 ( .A1(n10968), .A2(n12161), .ZN(n10971) );
  AOI22_X1 U13535 ( .A1(n12092), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12091), 
        .B2(n10969), .ZN(n10970) );
  NAND2_X1 U13536 ( .A1(n6678), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U13537 ( .A1(n12125), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13538 ( .A1(n10972), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10985) );
  OR2_X1 U13539 ( .A1(n10972), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10973) );
  AND2_X1 U13540 ( .A1(n10985), .A2(n10973), .ZN(n15073) );
  NAND2_X1 U13541 ( .A1(n12124), .A2(n15073), .ZN(n10975) );
  NAND2_X1 U13542 ( .A1(n10631), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10974) );
  XNOR2_X1 U13543 ( .A(n15180), .B(n14265), .ZN(n15068) );
  NAND2_X1 U13544 ( .A1(n15066), .A2(n15068), .ZN(n10979) );
  NAND2_X1 U13545 ( .A1(n15180), .A2(n11634), .ZN(n10978) );
  NAND2_X1 U13546 ( .A1(n10980), .A2(n12161), .ZN(n10982) );
  AOI22_X1 U13547 ( .A1(n12092), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12091), 
        .B2(n14350), .ZN(n10981) );
  NAND2_X1 U13548 ( .A1(n12125), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U13549 ( .A1(n6678), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10989) );
  INV_X1 U13550 ( .A(n12124), .ZN(n10983) );
  NAND2_X1 U13551 ( .A1(n10985), .A2(n10984), .ZN(n10986) );
  AND2_X1 U13552 ( .A1(n10997), .A2(n10986), .ZN(n11256) );
  NAND2_X1 U13553 ( .A1(n12056), .A2(n11256), .ZN(n10988) );
  NAND2_X1 U13554 ( .A1(n10631), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10987) );
  XNOR2_X1 U13555 ( .A(n11782), .B(n11777), .ZN(n12104) );
  INV_X1 U13556 ( .A(n12104), .ZN(n10991) );
  NAND2_X1 U13557 ( .A1(n11782), .A2(n11777), .ZN(n10992) );
  AOI22_X1 U13558 ( .A1(n12092), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12091), 
        .B2(n10994), .ZN(n10995) );
  NAND2_X1 U13559 ( .A1(n12156), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11002) );
  NAND2_X1 U13560 ( .A1(n6678), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U13561 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NAND2_X1 U13562 ( .A1(n11008), .A2(n10998), .ZN(n11969) );
  INV_X1 U13563 ( .A(n11969), .ZN(n11219) );
  NAND2_X1 U13564 ( .A1(n12124), .A2(n11219), .ZN(n11000) );
  NAND2_X1 U13565 ( .A1(n10631), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U13566 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n14263) );
  XNOR2_X1 U13567 ( .A(n11261), .B(n12105), .ZN(n11230) );
  INV_X1 U13568 ( .A(n11777), .ZN(n14264) );
  INV_X1 U13569 ( .A(n15180), .ZN(n15075) );
  INV_X1 U13570 ( .A(n15174), .ZN(n12242) );
  NAND2_X1 U13571 ( .A1(n14267), .A2(n12234), .ZN(n11004) );
  NOR2_X1 U13572 ( .A1(n14267), .A2(n12234), .ZN(n11003) );
  OAI21_X1 U13573 ( .B1(n11782), .B2(n14264), .A(n11249), .ZN(n11006) );
  INV_X1 U13574 ( .A(n12105), .ZN(n11260) );
  XNOR2_X1 U13575 ( .A(n11268), .B(n11260), .ZN(n11015) );
  NAND2_X1 U13576 ( .A1(n12156), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11013) );
  NAND2_X1 U13577 ( .A1(n6678), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11012) );
  AND2_X1 U13578 ( .A1(n11008), .A2(n11007), .ZN(n11009) );
  NOR2_X1 U13579 ( .A1(n11461), .A2(n11009), .ZN(n14193) );
  NAND2_X1 U13580 ( .A1(n12056), .A2(n14193), .ZN(n11011) );
  NAND2_X1 U13581 ( .A1(n10631), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11010) );
  NAND4_X1 U13582 ( .A1(n11013), .A2(n11012), .A3(n11011), .A4(n11010), .ZN(
        n14262) );
  INV_X1 U13583 ( .A(n14262), .ZN(n14138) );
  OR2_X1 U13584 ( .A1(n15102), .A2(n14138), .ZN(n11014) );
  OAI21_X1 U13585 ( .B1(n15097), .B2(n11777), .A(n11014), .ZN(n11967) );
  AOI21_X1 U13586 ( .B1(n11015), .B2(n14645), .A(n11967), .ZN(n11223) );
  AND2_X2 U13587 ( .A1(n11363), .A2(n15174), .ZN(n15078) );
  AOI21_X1 U13588 ( .B1(n12255), .B2(n11255), .A(n11278), .ZN(n11221) );
  AOI22_X1 U13589 ( .A1(n11221), .A2(n15077), .B1(n12255), .B2(n15156), .ZN(
        n11016) );
  OAI211_X1 U13590 ( .C1(n15146), .C2(n11230), .A(n11223), .B(n11016), .ZN(
        n11019) );
  NAND2_X1 U13591 ( .A1(n11019), .A2(n15212), .ZN(n11017) );
  OAI21_X1 U13592 ( .B1(n15212), .B2(n11018), .A(n11017), .ZN(P1_U3483) );
  NAND2_X1 U13593 ( .A1(n11019), .A2(n15225), .ZN(n11020) );
  OAI21_X1 U13594 ( .B1(n15225), .B2(n10472), .A(n11020), .ZN(P1_U3536) );
  AOI22_X1 U13595 ( .A1(n12767), .A2(n14268), .B1(n11545), .B2(n12227), .ZN(
        n11490) );
  AOI22_X1 U13596 ( .A1(n11545), .A2(n14268), .B1(n12770), .B2(n12227), .ZN(
        n11027) );
  OAI211_X1 U13597 ( .C1(n11029), .C2(n11028), .A(n11491), .B(n14965), .ZN(
        n11034) );
  INV_X1 U13598 ( .A(n14960), .ZN(n14972) );
  OAI22_X1 U13599 ( .A1(n14972), .A2(n15101), .B1(n12235), .B2(n14969), .ZN(
        n11032) );
  MUX2_X1 U13600 ( .A(n14244), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n11031) );
  AOI211_X1 U13601 ( .C1(n14981), .C2(n12227), .A(n11032), .B(n11031), .ZN(
        n11033) );
  NAND2_X1 U13602 ( .A1(n11034), .A2(n11033), .ZN(P1_U3218) );
  INV_X1 U13603 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15012) );
  MUX2_X1 U13604 ( .A(n15012), .B(P1_REG1_REG_14__SCAN_IN), .S(n11916), .Z(
        n11037) );
  INV_X1 U13605 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11834) );
  MUX2_X1 U13606 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11834), .S(n11704), .Z(
        n14360) );
  NAND2_X1 U13607 ( .A1(n14361), .A2(n14360), .ZN(n14359) );
  OAI21_X1 U13608 ( .B1(n14362), .B2(n11834), .A(n14359), .ZN(n11036) );
  AOI21_X1 U13609 ( .B1(n11037), .B2(n11036), .A(n11741), .ZN(n11050) );
  NAND2_X1 U13610 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14939)
         );
  INV_X1 U13611 ( .A(n14939), .ZN(n11039) );
  NOR2_X1 U13612 ( .A1(n15055), .A2(n11742), .ZN(n11038) );
  AOI211_X1 U13613 ( .C1(n14365), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11039), 
        .B(n11038), .ZN(n11049) );
  AOI21_X1 U13614 ( .B1(n10509), .B2(n11041), .A(n11040), .ZN(n14368) );
  INV_X1 U13615 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11042) );
  MUX2_X1 U13616 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11042), .S(n11704), .Z(
        n14367) );
  NAND2_X1 U13617 ( .A1(n14368), .A2(n14367), .ZN(n14366) );
  NAND2_X1 U13618 ( .A1(n11704), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11045) );
  INV_X1 U13619 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U13620 ( .A(n11043), .B(P1_REG2_REG_14__SCAN_IN), .S(n11916), .Z(
        n11044) );
  AOI21_X1 U13621 ( .B1(n14366), .B2(n11045), .A(n11044), .ZN(n11746) );
  INV_X1 U13622 ( .A(n11746), .ZN(n11047) );
  NAND3_X1 U13623 ( .A1(n14366), .A2(n11045), .A3(n11044), .ZN(n11046) );
  NAND3_X1 U13624 ( .A1(n11047), .A2(n14400), .A3(n11046), .ZN(n11048) );
  OAI211_X1 U13625 ( .C1(n11050), .C2(n14396), .A(n11049), .B(n11048), .ZN(
        P1_U3257) );
  NAND2_X1 U13626 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  OAI211_X1 U13627 ( .C1(n11054), .C2(n13441), .A(n11053), .B(n12608), .ZN(
        P3_U3272) );
  INV_X1 U13628 ( .A(n11055), .ZN(n11059) );
  AOI22_X1 U13629 ( .A1(n15314), .A2(n11057), .B1(n15316), .B2(n11056), .ZN(
        n11058) );
  OAI21_X1 U13630 ( .B1(n11059), .B2(n13961), .A(n11058), .ZN(n11062) );
  MUX2_X1 U13631 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11060), .S(n13963), .Z(
        n11061) );
  AOI211_X1 U13632 ( .C1(n15320), .C2(n11063), .A(n11062), .B(n11061), .ZN(
        n11064) );
  INV_X1 U13633 ( .A(n11064), .ZN(P2_U3261) );
  XNOR2_X1 U13634 ( .A(n11066), .B(n11065), .ZN(n11214) );
  AOI211_X1 U13635 ( .C1(n11208), .C2(n11067), .A(n14001), .B(n11234), .ZN(
        n11206) );
  XNOR2_X1 U13636 ( .A(n11068), .B(n11069), .ZN(n11072) );
  NAND2_X1 U13637 ( .A1(n13610), .A2(n13668), .ZN(n11071) );
  NAND2_X1 U13638 ( .A1(n13551), .A2(n13670), .ZN(n11070) );
  AND2_X1 U13639 ( .A1(n11071), .A2(n11070), .ZN(n11199) );
  OAI21_X1 U13640 ( .B1(n11072), .B2(n13946), .A(n11199), .ZN(n11211) );
  AOI211_X1 U13641 ( .C1(n15370), .C2(n11214), .A(n11206), .B(n11211), .ZN(
        n11079) );
  OAI22_X1 U13642 ( .A1(n14046), .A2(n11076), .B1(n15431), .B2(n10278), .ZN(
        n11073) );
  INV_X1 U13643 ( .A(n11073), .ZN(n11074) );
  OAI21_X1 U13644 ( .B1(n11079), .B2(n15429), .A(n11074), .ZN(P2_U3505) );
  INV_X1 U13645 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11075) );
  OAI22_X1 U13646 ( .A1(n14081), .A2(n11076), .B1(n15420), .B2(n11075), .ZN(
        n11077) );
  INV_X1 U13647 ( .A(n11077), .ZN(n11078) );
  OAI21_X1 U13648 ( .B1(n11079), .B2(n15418), .A(n11078), .ZN(P2_U3448) );
  AOI21_X1 U13649 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n11087) );
  NOR2_X1 U13650 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8277), .ZN(n15442) );
  INV_X1 U13651 ( .A(n12936), .ZN(n12917) );
  OAI22_X1 U13652 ( .A1(n15555), .A2(n12917), .B1(n12931), .B2(n15561), .ZN(
        n11083) );
  AOI211_X1 U13653 ( .C1(n12914), .C2(n11301), .A(n15442), .B(n11083), .ZN(
        n11086) );
  INV_X1 U13654 ( .A(n11084), .ZN(n15562) );
  NAND2_X1 U13655 ( .A1(n12938), .A2(n15562), .ZN(n11085) );
  OAI211_X1 U13656 ( .C1(n11087), .C2(n12945), .A(n11086), .B(n11085), .ZN(
        P3_U3167) );
  XNOR2_X1 U13657 ( .A(n11088), .B(n11092), .ZN(n11090) );
  AOI21_X1 U13658 ( .B1(n11090), .B2(n14882), .A(n11089), .ZN(n15367) );
  XNOR2_X1 U13659 ( .A(n11092), .B(n11091), .ZN(n15371) );
  OAI211_X1 U13660 ( .C1(n15366), .C2(n12400), .A(n9576), .B(n11093), .ZN(
        n15365) );
  NAND2_X1 U13661 ( .A1(n15314), .A2(n11094), .ZN(n11096) );
  AOI22_X1 U13662 ( .A1(n6674), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n15316), .ZN(n11095) );
  OAI211_X1 U13663 ( .C1(n15365), .C2(n13961), .A(n11096), .B(n11095), .ZN(
        n11097) );
  AOI21_X1 U13664 ( .B1(n15320), .B2(n15371), .A(n11097), .ZN(n11098) );
  OAI21_X1 U13665 ( .B1(n6674), .B2(n15367), .A(n11098), .ZN(P2_U3264) );
  INV_X1 U13666 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11100) );
  MUX2_X1 U13667 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11100), .S(n15267), .Z(
        n15261) );
  OAI21_X1 U13668 ( .B1(n15267), .B2(P2_REG1_REG_9__SCAN_IN), .A(n15260), .ZN(
        n15274) );
  INV_X1 U13669 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11101) );
  MUX2_X1 U13670 ( .A(n11101), .B(P2_REG1_REG_10__SCAN_IN), .S(n11108), .Z(
        n15275) );
  NOR2_X1 U13671 ( .A1(n15274), .A2(n15275), .ZN(n15273) );
  INV_X1 U13672 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11102) );
  MUX2_X1 U13673 ( .A(n11102), .B(P2_REG1_REG_11__SCAN_IN), .S(n11332), .Z(
        n11103) );
  AOI211_X1 U13674 ( .C1(n11104), .C2(n11103), .A(n15298), .B(n11331), .ZN(
        n11117) );
  INV_X1 U13675 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11115) );
  AOI21_X1 U13676 ( .B1(n11106), .B2(P2_REG2_REG_8__SCAN_IN), .A(n11105), .ZN(
        n15258) );
  INV_X1 U13677 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11437) );
  MUX2_X1 U13678 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11437), .S(n15267), .Z(
        n15257) );
  NAND2_X1 U13679 ( .A1(n15258), .A2(n15257), .ZN(n15256) );
  OAI21_X1 U13680 ( .B1(n15267), .B2(P2_REG2_REG_9__SCAN_IN), .A(n15256), .ZN(
        n15280) );
  INV_X1 U13681 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11107) );
  MUX2_X1 U13682 ( .A(n11107), .B(P2_REG2_REG_10__SCAN_IN), .S(n11108), .Z(
        n15281) );
  NOR2_X1 U13683 ( .A1(n15280), .A2(n15281), .ZN(n15278) );
  AOI21_X1 U13684 ( .B1(n11108), .B2(P2_REG2_REG_10__SCAN_IN), .A(n15278), 
        .ZN(n11110) );
  INV_X1 U13685 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11339) );
  MUX2_X1 U13686 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11339), .S(n11332), .Z(
        n11109) );
  NOR2_X1 U13687 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  AND2_X1 U13688 ( .A1(n11110), .A2(n11109), .ZN(n11337) );
  OAI21_X1 U13689 ( .B1(n11111), .B2(n11337), .A(n15307), .ZN(n11114) );
  NOR2_X1 U13690 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13600), .ZN(n11112) );
  AOI21_X1 U13691 ( .B1(n15305), .B2(n11332), .A(n11112), .ZN(n11113) );
  OAI211_X1 U13692 ( .C1(n15313), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        n11116) );
  OR2_X1 U13693 ( .A1(n11117), .A2(n11116), .ZN(P2_U3225) );
  NOR2_X1 U13694 ( .A1(n7476), .A2(n11121), .ZN(n11122) );
  NOR2_X1 U13695 ( .A1(n15564), .A2(n15433), .ZN(n15432) );
  AOI22_X1 U13696 ( .A1(n11147), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11146), 
        .B2(n15458), .ZN(n15450) );
  NOR2_X1 U13697 ( .A1(n11153), .A2(n11123), .ZN(n11124) );
  NOR2_X1 U13698 ( .A1(n11152), .A2(n15469), .ZN(n15468) );
  NOR2_X1 U13699 ( .A1(n11124), .A2(n15468), .ZN(n15486) );
  AOI22_X1 U13700 ( .A1(n11160), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11159), 
        .B2(n15493), .ZN(n15485) );
  NOR2_X1 U13701 ( .A1(n15486), .A2(n15485), .ZN(n15484) );
  NOR2_X1 U13702 ( .A1(n11166), .A2(n11125), .ZN(n11126) );
  AOI22_X1 U13703 ( .A1(n11381), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n11172), 
        .B2(n11374), .ZN(n11127) );
  AOI21_X1 U13704 ( .B1(n6827), .B2(n11127), .A(n11373), .ZN(n11183) );
  AOI22_X1 U13705 ( .A1(n11381), .A2(n11171), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11374), .ZN(n11136) );
  AOI22_X1 U13706 ( .A1(n11160), .A2(n11158), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15493), .ZN(n15497) );
  AOI22_X1 U13707 ( .A1(n11147), .A2(n11145), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15458), .ZN(n15462) );
  NAND2_X1 U13708 ( .A1(n15438), .A2(n11129), .ZN(n11130) );
  NAND2_X1 U13709 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15444), .ZN(n15443) );
  NAND2_X1 U13710 ( .A1(n15475), .A2(n11131), .ZN(n11132) );
  NAND2_X1 U13711 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15479), .ZN(n15478) );
  NAND2_X1 U13712 ( .A1(n15512), .A2(n11133), .ZN(n11134) );
  NAND2_X1 U13713 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15518), .ZN(n15517) );
  OAI21_X1 U13714 ( .B1(n11136), .B2(n11135), .A(n11380), .ZN(n11181) );
  NOR2_X1 U13715 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11137), .ZN(n11585) );
  AOI21_X1 U13716 ( .B1(n15516), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11585), 
        .ZN(n11138) );
  OAI21_X1 U13717 ( .B1(n15513), .B2(n11374), .A(n11138), .ZN(n11180) );
  INV_X1 U13718 ( .A(n11139), .ZN(n11140) );
  AOI22_X1 U13719 ( .A1(n11143), .A2(n11142), .B1(n11141), .B2(n11140), .ZN(
        n15436) );
  MUX2_X1 U13720 ( .A(n15564), .B(n15678), .S(n12990), .Z(n11144) );
  NOR2_X1 U13721 ( .A1(n11144), .A2(n7476), .ZN(n15434) );
  NOR2_X1 U13722 ( .A1(n15436), .A2(n15434), .ZN(n15454) );
  AND2_X1 U13723 ( .A1(n11144), .A2(n7476), .ZN(n15453) );
  MUX2_X1 U13724 ( .A(n11146), .B(n11145), .S(n12990), .Z(n11148) );
  NAND2_X1 U13725 ( .A1(n11148), .A2(n11147), .ZN(n15471) );
  INV_X1 U13726 ( .A(n11148), .ZN(n11149) );
  NAND2_X1 U13727 ( .A1(n11149), .A2(n15458), .ZN(n11150) );
  AND2_X1 U13728 ( .A1(n15471), .A2(n11150), .ZN(n15452) );
  OAI21_X1 U13729 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15472) );
  MUX2_X1 U13730 ( .A(n11152), .B(n11151), .S(n12990), .Z(n11154) );
  NAND2_X1 U13731 ( .A1(n11154), .A2(n11153), .ZN(n11157) );
  INV_X1 U13732 ( .A(n11154), .ZN(n11155) );
  NAND2_X1 U13733 ( .A1(n11155), .A2(n15475), .ZN(n11156) );
  NAND2_X1 U13734 ( .A1(n11157), .A2(n11156), .ZN(n15470) );
  AOI21_X1 U13735 ( .B1(n15472), .B2(n15471), .A(n15470), .ZN(n15489) );
  INV_X1 U13736 ( .A(n11157), .ZN(n15488) );
  MUX2_X1 U13737 ( .A(n11159), .B(n11158), .S(n12990), .Z(n11161) );
  NAND2_X1 U13738 ( .A1(n11161), .A2(n11160), .ZN(n15506) );
  INV_X1 U13739 ( .A(n11161), .ZN(n11162) );
  NAND2_X1 U13740 ( .A1(n11162), .A2(n15493), .ZN(n11163) );
  AND2_X1 U13741 ( .A1(n15506), .A2(n11163), .ZN(n15487) );
  OAI21_X1 U13742 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15507) );
  MUX2_X1 U13743 ( .A(n11165), .B(n11164), .S(n12990), .Z(n11167) );
  NAND2_X1 U13744 ( .A1(n11167), .A2(n11166), .ZN(n11170) );
  INV_X1 U13745 ( .A(n11167), .ZN(n11168) );
  NAND2_X1 U13746 ( .A1(n11168), .A2(n15512), .ZN(n11169) );
  NAND2_X1 U13747 ( .A1(n11170), .A2(n11169), .ZN(n15505) );
  AOI21_X1 U13748 ( .B1(n15507), .B2(n15506), .A(n15505), .ZN(n15510) );
  INV_X1 U13749 ( .A(n11170), .ZN(n11177) );
  MUX2_X1 U13750 ( .A(n11172), .B(n11171), .S(n12990), .Z(n11173) );
  NAND2_X1 U13751 ( .A1(n11173), .A2(n11381), .ZN(n11376) );
  INV_X1 U13752 ( .A(n11173), .ZN(n11174) );
  NAND2_X1 U13753 ( .A1(n11174), .A2(n11374), .ZN(n11175) );
  AND2_X1 U13754 ( .A1(n11376), .A2(n11175), .ZN(n11176) );
  OAI21_X1 U13755 ( .B1(n15510), .B2(n11177), .A(n11176), .ZN(n11377) );
  OR3_X1 U13756 ( .A1(n15510), .A2(n11177), .A3(n11176), .ZN(n11178) );
  AOI21_X1 U13757 ( .B1(n11377), .B2(n11178), .A(n15439), .ZN(n11179) );
  AOI211_X1 U13758 ( .C1(n15519), .C2(n11181), .A(n11180), .B(n11179), .ZN(
        n11182) );
  OAI21_X1 U13759 ( .B1(n11183), .B2(n15523), .A(n11182), .ZN(P3_U3192) );
  NOR3_X1 U13760 ( .A1(n15519), .A2(n14837), .A3(n15508), .ZN(n11194) );
  OAI22_X1 U13761 ( .A1(n13014), .A2(n9033), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11184), .ZN(n11187) );
  AND2_X1 U13762 ( .A1(n14837), .A2(n11185), .ZN(n11186) );
  AOI211_X1 U13763 ( .C1(n15519), .C2(n11188), .A(n11187), .B(n11186), .ZN(
        n11192) );
  OR2_X1 U13764 ( .A1(n15439), .A2(n11189), .ZN(n11190) );
  MUX2_X1 U13765 ( .A(n11190), .B(n15513), .S(P3_IR_REG_0__SCAN_IN), .Z(n11191) );
  OAI211_X1 U13766 ( .C1(n11194), .C2(n11193), .A(n11192), .B(n11191), .ZN(
        P3_U3182) );
  INV_X1 U13767 ( .A(n12073), .ZN(n11195) );
  OAI222_X1 U13768 ( .A1(P1_U3086), .A2(n14527), .B1(n14780), .B2(n11195), 
        .C1(n12074), .C2(n14772), .ZN(P1_U3336) );
  OAI222_X1 U13769 ( .A1(n14106), .A2(n11196), .B1(n14111), .B2(n11195), .C1(
        n13726), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13770 ( .A1(n13588), .A2(n11207), .ZN(n11198) );
  OAI211_X1 U13771 ( .C1(n11199), .C2(n13624), .A(n11198), .B(n11197), .ZN(
        n11204) );
  XNOR2_X1 U13772 ( .A(n11201), .B(n11200), .ZN(n11202) );
  NOR2_X1 U13773 ( .A1(n11202), .A2(n13630), .ZN(n11203) );
  AOI211_X1 U13774 ( .C1(n11208), .C2(n13628), .A(n11204), .B(n11203), .ZN(
        n11205) );
  INV_X1 U13775 ( .A(n11205), .ZN(P2_U3211) );
  INV_X1 U13776 ( .A(n11206), .ZN(n11210) );
  AOI22_X1 U13777 ( .A1(n15314), .A2(n11208), .B1(n15316), .B2(n11207), .ZN(
        n11209) );
  OAI21_X1 U13778 ( .B1(n11210), .B2(n13961), .A(n11209), .ZN(n11213) );
  MUX2_X1 U13779 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11211), .S(n13963), .Z(
        n11212) );
  AOI211_X1 U13780 ( .C1(n15320), .C2(n11214), .A(n11213), .B(n11212), .ZN(
        n11215) );
  INV_X1 U13781 ( .A(n11215), .ZN(P2_U3259) );
  INV_X1 U13782 ( .A(n11216), .ZN(n11220) );
  AOI22_X1 U13783 ( .A1(n11221), .A2(n11220), .B1(n11219), .B2(n15099), .ZN(
        n11222) );
  NAND2_X1 U13784 ( .A1(n11223), .A2(n11222), .ZN(n11228) );
  AND2_X1 U13785 ( .A1(n11225), .A2(n11224), .ZN(n11227) );
  MUX2_X1 U13786 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11228), .S(n15103), .Z(
        n11232) );
  INV_X1 U13787 ( .A(n11229), .ZN(n14990) );
  OAI22_X1 U13788 ( .A1(n11230), .A2(n14623), .B1(n7013), .B2(n15106), .ZN(
        n11231) );
  OR2_X1 U13789 ( .A1(n11232), .A2(n11231), .ZN(P1_U3285) );
  XOR2_X1 U13790 ( .A(n11233), .B(n11237), .Z(n11353) );
  OAI21_X1 U13791 ( .B1(n11234), .B2(n11244), .A(n9576), .ZN(n11235) );
  NOR2_X1 U13792 ( .A1(n11235), .A2(n11294), .ZN(n11347) );
  XNOR2_X1 U13793 ( .A(n11236), .B(n11237), .ZN(n11240) );
  NAND2_X1 U13794 ( .A1(n13610), .A2(n13667), .ZN(n11239) );
  NAND2_X1 U13795 ( .A1(n13622), .A2(n13669), .ZN(n11238) );
  AND2_X1 U13796 ( .A1(n11239), .A2(n11238), .ZN(n11412) );
  OAI21_X1 U13797 ( .B1(n11240), .B2(n13946), .A(n11412), .ZN(n11350) );
  AOI211_X1 U13798 ( .C1(n15370), .C2(n11353), .A(n11347), .B(n11350), .ZN(
        n11247) );
  INV_X1 U13799 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11241) );
  OAI22_X1 U13800 ( .A1(n14081), .A2(n11244), .B1(n15420), .B2(n11241), .ZN(
        n11242) );
  INV_X1 U13801 ( .A(n11242), .ZN(n11243) );
  OAI21_X1 U13802 ( .B1(n11247), .B2(n15418), .A(n11243), .ZN(P2_U3451) );
  OAI22_X1 U13803 ( .A1(n14046), .A2(n11244), .B1(n15431), .B2(n10279), .ZN(
        n11245) );
  INV_X1 U13804 ( .A(n11245), .ZN(n11246) );
  OAI21_X1 U13805 ( .B1(n11247), .B2(n15429), .A(n11246), .ZN(P2_U3506) );
  XNOR2_X1 U13806 ( .A(n11248), .B(n12104), .ZN(n15187) );
  XNOR2_X1 U13807 ( .A(n11249), .B(n12104), .ZN(n11252) );
  OR2_X1 U13808 ( .A1(n15097), .A2(n11634), .ZN(n11251) );
  INV_X1 U13809 ( .A(n14263), .ZN(n11274) );
  OR2_X1 U13810 ( .A1(n15102), .A2(n11274), .ZN(n11250) );
  AND2_X1 U13811 ( .A1(n11251), .A2(n11250), .ZN(n11783) );
  OAI21_X1 U13812 ( .B1(n11252), .B2(n15145), .A(n11783), .ZN(n15191) );
  INV_X1 U13813 ( .A(n15191), .ZN(n11253) );
  MUX2_X1 U13814 ( .A(n11254), .B(n11253), .S(n15103), .Z(n11259) );
  INV_X1 U13815 ( .A(n15077), .ZN(n15159) );
  AOI211_X1 U13816 ( .C1(n12251), .C2(n15076), .A(n15159), .B(n7014), .ZN(
        n15188) );
  INV_X1 U13817 ( .A(n11256), .ZN(n11787) );
  OAI22_X1 U13818 ( .A1(n15106), .A2(n11782), .B1(n14648), .B2(n11787), .ZN(
        n11257) );
  AOI21_X1 U13819 ( .B1(n15080), .B2(n15188), .A(n11257), .ZN(n11258) );
  OAI211_X1 U13820 ( .C1(n14623), .C2(n15187), .A(n11259), .B(n11258), .ZN(
        P1_U3286) );
  OR2_X1 U13821 ( .A1(n12255), .A2(n14263), .ZN(n11262) );
  NAND2_X1 U13822 ( .A1(n11264), .A2(n12161), .ZN(n11267) );
  AOI22_X1 U13823 ( .A1(n12091), .A2(n11265), .B1(n12092), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n11266) );
  XNOR2_X1 U13824 ( .A(n11468), .B(n12106), .ZN(n15196) );
  XNOR2_X1 U13825 ( .A(n11475), .B(n12106), .ZN(n11275) );
  NAND2_X1 U13826 ( .A1(n12156), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U13827 ( .A1(n6678), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11271) );
  XNOR2_X1 U13828 ( .A(n11461), .B(n14136), .ZN(n14141) );
  NAND2_X1 U13829 ( .A1(n12056), .A2(n14141), .ZN(n11270) );
  NAND2_X1 U13830 ( .A1(n10631), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U13831 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n14261) );
  OR2_X1 U13832 ( .A1(n15102), .A2(n14971), .ZN(n11273) );
  OAI21_X1 U13833 ( .B1(n15097), .B2(n11274), .A(n11273), .ZN(n14191) );
  AOI21_X1 U13834 ( .B1(n11275), .B2(n14645), .A(n14191), .ZN(n15194) );
  MUX2_X1 U13835 ( .A(n11276), .B(n15194), .S(n15103), .Z(n11283) );
  INV_X1 U13836 ( .A(n14192), .ZN(n15195) );
  INV_X1 U13837 ( .A(n11532), .ZN(n11277) );
  OAI211_X1 U13838 ( .C1(n15195), .C2(n11278), .A(n11277), .B(n15077), .ZN(
        n15193) );
  INV_X1 U13839 ( .A(n15193), .ZN(n11281) );
  INV_X1 U13840 ( .A(n14193), .ZN(n11279) );
  OAI22_X1 U13841 ( .A1(n15106), .A2(n15195), .B1(n14648), .B2(n11279), .ZN(
        n11280) );
  AOI21_X1 U13842 ( .B1(n15080), .B2(n11281), .A(n11280), .ZN(n11282) );
  OAI211_X1 U13843 ( .C1(n14623), .C2(n15196), .A(n11283), .B(n11282), .ZN(
        P1_U3284) );
  XNOR2_X1 U13844 ( .A(n11285), .B(n11284), .ZN(n15393) );
  NAND2_X1 U13845 ( .A1(n15393), .A2(n15406), .ZN(n11293) );
  NAND2_X1 U13846 ( .A1(n6830), .A2(n11286), .ZN(n11287) );
  NAND2_X1 U13847 ( .A1(n11288), .A2(n11287), .ZN(n11291) );
  NAND2_X1 U13848 ( .A1(n13610), .A2(n13666), .ZN(n11290) );
  NAND2_X1 U13849 ( .A1(n13622), .A2(n13668), .ZN(n11289) );
  NAND2_X1 U13850 ( .A1(n11290), .A2(n11289), .ZN(n13499) );
  AOI21_X1 U13851 ( .B1(n11291), .B2(n14882), .A(n13499), .ZN(n11292) );
  OAI211_X1 U13852 ( .C1(n11294), .C2(n15391), .A(n9576), .B(n11435), .ZN(
        n15390) );
  AOI22_X1 U13853 ( .A1(n6674), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n13497), .B2(
        n15316), .ZN(n11296) );
  NAND2_X1 U13854 ( .A1(n15314), .A2(n13498), .ZN(n11295) );
  OAI211_X1 U13855 ( .C1(n15390), .C2(n13961), .A(n11296), .B(n11295), .ZN(
        n11297) );
  AOI21_X1 U13856 ( .B1(n15393), .B2(n11298), .A(n11297), .ZN(n11299) );
  OAI21_X1 U13857 ( .B1(n15395), .B2(n6674), .A(n11299), .ZN(P2_U3257) );
  XNOR2_X1 U13858 ( .A(n11303), .B(n11300), .ZN(n15634) );
  AND2_X1 U13859 ( .A1(n12449), .A2(n15585), .ZN(n15602) );
  INV_X1 U13860 ( .A(n13156), .ZN(n15620) );
  INV_X1 U13861 ( .A(n15599), .ZN(n15616) );
  AOI22_X1 U13862 ( .A1(n15610), .A2(n15608), .B1(n11301), .B2(n15607), .ZN(
        n11305) );
  OAI211_X1 U13863 ( .C1(n6831), .C2(n11303), .A(n11302), .B(n15612), .ZN(
        n11304) );
  OAI211_X1 U13864 ( .C1(n15634), .C2(n15616), .A(n11305), .B(n11304), .ZN(
        n15635) );
  INV_X1 U13865 ( .A(n15635), .ZN(n11307) );
  MUX2_X1 U13866 ( .A(n11307), .B(n11306), .S(n15625), .Z(n11311) );
  NOR2_X1 U13867 ( .A1(n11308), .A2(n15605), .ZN(n15636) );
  AOI22_X1 U13868 ( .A1(n15577), .A2(n15636), .B1(n15576), .B2(n11309), .ZN(
        n11310) );
  OAI211_X1 U13869 ( .C1(n15634), .C2(n15620), .A(n11311), .B(n11310), .ZN(
        P3_U3230) );
  INV_X1 U13870 ( .A(n11312), .ZN(n11313) );
  NOR2_X1 U13871 ( .A1(n11080), .A2(n11313), .ZN(n11316) );
  XNOR2_X1 U13872 ( .A(n15555), .B(n11314), .ZN(n11315) );
  NAND2_X1 U13873 ( .A1(n11316), .A2(n11315), .ZN(n11447) );
  OAI211_X1 U13874 ( .C1(n11316), .C2(n11315), .A(n11447), .B(n12924), .ZN(
        n11322) );
  NOR2_X1 U13875 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11317), .ZN(n15460) );
  OAI22_X1 U13876 ( .A1(n11319), .A2(n12917), .B1(n11318), .B2(n12931), .ZN(
        n11320) );
  AOI211_X1 U13877 ( .C1(n12914), .C2(n11505), .A(n15460), .B(n11320), .ZN(
        n11321) );
  OAI211_X1 U13878 ( .C1(n11502), .C2(n12896), .A(n11322), .B(n11321), .ZN(
        P3_U3179) );
  AOI21_X1 U13879 ( .B1(n11325), .B2(n11324), .A(n11323), .ZN(n11330) );
  AND2_X1 U13880 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15515) );
  INV_X1 U13881 ( .A(n11807), .ZN(n14862) );
  OAI22_X1 U13882 ( .A1(n14862), .A2(n12917), .B1(n12931), .B2(n11651), .ZN(
        n11326) );
  AOI211_X1 U13883 ( .C1(n12914), .C2(n12491), .A(n15515), .B(n11326), .ZN(
        n11329) );
  INV_X1 U13884 ( .A(n11327), .ZN(n11652) );
  NAND2_X1 U13885 ( .A1(n12938), .A2(n11652), .ZN(n11328) );
  OAI211_X1 U13886 ( .C1(n11330), .C2(n12945), .A(n11329), .B(n11328), .ZN(
        P3_U3171) );
  INV_X1 U13887 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11333) );
  MUX2_X1 U13888 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11333), .S(n11687), .Z(
        n11334) );
  OAI21_X1 U13889 ( .B1(n11335), .B2(n11334), .A(n11686), .ZN(n11336) );
  NAND2_X1 U13890 ( .A1(n11336), .A2(n15265), .ZN(n11346) );
  AOI21_X1 U13891 ( .B1(n11339), .B2(n11338), .A(n11337), .ZN(n11342) );
  INV_X1 U13892 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11340) );
  MUX2_X1 U13893 ( .A(n11340), .B(P2_REG2_REG_12__SCAN_IN), .S(n11687), .Z(
        n11341) );
  NOR2_X1 U13894 ( .A1(n11342), .A2(n11341), .ZN(n11681) );
  AOI21_X1 U13895 ( .B1(n11342), .B2(n11341), .A(n11681), .ZN(n11343) );
  OAI22_X1 U13896 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9361), .B1(n11343), .B2(
        n15279), .ZN(n11344) );
  AOI21_X1 U13897 ( .B1(n15305), .B2(n11687), .A(n11344), .ZN(n11345) );
  OAI211_X1 U13898 ( .C1(n15313), .C2(n7517), .A(n11346), .B(n11345), .ZN(
        P2_U3226) );
  INV_X1 U13899 ( .A(n11347), .ZN(n11349) );
  AOI22_X1 U13900 ( .A1(n15314), .A2(n11418), .B1(n15316), .B2(n11409), .ZN(
        n11348) );
  OAI21_X1 U13901 ( .B1(n11349), .B2(n13961), .A(n11348), .ZN(n11352) );
  MUX2_X1 U13902 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11350), .S(n13963), .Z(
        n11351) );
  AOI211_X1 U13903 ( .C1(n15320), .C2(n11353), .A(n11352), .B(n11351), .ZN(
        n11354) );
  INV_X1 U13904 ( .A(n11354), .ZN(P2_U3258) );
  INV_X1 U13905 ( .A(n11355), .ZN(n11495) );
  OAI22_X1 U13906 ( .A1(n14577), .A2(n11356), .B1(n11495), .B2(n14648), .ZN(
        n11357) );
  AOI21_X1 U13907 ( .B1(n15074), .B2(n12233), .A(n11357), .ZN(n11360) );
  MUX2_X1 U13908 ( .A(n10363), .B(n11358), .S(n15103), .Z(n11359) );
  OAI211_X1 U13909 ( .C1(n14623), .C2(n11361), .A(n11360), .B(n11359), .ZN(
        P1_U3289) );
  XOR2_X1 U13910 ( .A(n11362), .B(n12101), .Z(n15171) );
  OAI21_X1 U13911 ( .B1(n11363), .B2(n15174), .A(n15077), .ZN(n11364) );
  OR2_X1 U13912 ( .A1(n15078), .A2(n11364), .ZN(n15173) );
  INV_X1 U13913 ( .A(n11555), .ZN(n11365) );
  OAI22_X1 U13914 ( .A1(n14577), .A2(n15173), .B1(n11365), .B2(n14648), .ZN(
        n11366) );
  AOI21_X1 U13915 ( .B1(n15074), .B2(n12242), .A(n11366), .ZN(n11372) );
  XNOR2_X1 U13916 ( .A(n11367), .B(n12101), .ZN(n11369) );
  OR2_X1 U13917 ( .A1(n15102), .A2(n11634), .ZN(n11368) );
  OAI21_X1 U13918 ( .B1(n15097), .B2(n12235), .A(n11368), .ZN(n11551) );
  AOI21_X1 U13919 ( .B1(n11369), .B2(n14645), .A(n11551), .ZN(n15172) );
  MUX2_X1 U13920 ( .A(n11370), .B(n15172), .S(n15103), .Z(n11371) );
  OAI211_X1 U13921 ( .C1(n14623), .C2(n15171), .A(n11372), .B(n11371), .ZN(
        P1_U3288) );
  AOI21_X1 U13922 ( .B1(n8374), .B2(n11375), .A(n11559), .ZN(n11390) );
  NAND2_X1 U13923 ( .A1(n11377), .A2(n11376), .ZN(n11379) );
  MUX2_X1 U13924 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12990), .Z(n11571) );
  XNOR2_X1 U13925 ( .A(n11571), .B(n11572), .ZN(n11378) );
  NAND2_X1 U13926 ( .A1(n11379), .A2(n11378), .ZN(n11577) );
  OAI21_X1 U13927 ( .B1(n11379), .B2(n11378), .A(n11577), .ZN(n11388) );
  NAND2_X1 U13928 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11382), .ZN(n11565) );
  OAI21_X1 U13929 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11382), .A(n11565), 
        .ZN(n11383) );
  NAND2_X1 U13930 ( .A1(n11383), .A2(n15519), .ZN(n11386) );
  NOR2_X1 U13931 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11384), .ZN(n11804) );
  AOI21_X1 U13932 ( .B1(n15516), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11804), 
        .ZN(n11385) );
  OAI211_X1 U13933 ( .C1(n15513), .C2(n11564), .A(n11386), .B(n11385), .ZN(
        n11387) );
  AOI21_X1 U13934 ( .B1(n11388), .B2(n15508), .A(n11387), .ZN(n11389) );
  OAI21_X1 U13935 ( .B1(n11390), .B2(n15523), .A(n11389), .ZN(P3_U3193) );
  OAI21_X1 U13936 ( .B1(n11393), .B2(n11392), .A(n11391), .ZN(n15169) );
  INV_X1 U13937 ( .A(n15169), .ZN(n11403) );
  INV_X1 U13938 ( .A(n15090), .ZN(n11395) );
  OAI211_X1 U13939 ( .C1(n15165), .C2(n11395), .A(n15077), .B(n11394), .ZN(
        n15164) );
  INV_X1 U13940 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14289) );
  OAI22_X1 U13941 ( .A1(n14577), .A2(n15164), .B1(n14289), .B2(n14648), .ZN(
        n11396) );
  AOI21_X1 U13942 ( .B1(n15074), .B2(n11397), .A(n11396), .ZN(n11402) );
  XNOR2_X1 U13943 ( .A(n12220), .B(n12219), .ZN(n11399) );
  AOI21_X1 U13944 ( .B1(n14645), .B2(n11399), .A(n11398), .ZN(n15166) );
  MUX2_X1 U13945 ( .A(n11400), .B(n15166), .S(n15103), .Z(n11401) );
  OAI211_X1 U13946 ( .C1(n14623), .C2(n11403), .A(n11402), .B(n11401), .ZN(
        P1_U3291) );
  AOI21_X1 U13947 ( .B1(n14645), .B2(n15103), .A(n14654), .ZN(n11408) );
  OAI21_X1 U13948 ( .B1(n15091), .B2(n12213), .A(n15085), .ZN(n15144) );
  INV_X1 U13949 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11404) );
  OAI22_X1 U13950 ( .A1(n15112), .A2(n15147), .B1(n11404), .B2(n14648), .ZN(
        n11405) );
  AOI21_X1 U13951 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15112), .A(n11405), .ZN(
        n11407) );
  NOR2_X1 U13952 ( .A1(n14577), .A2(n15159), .ZN(n15100) );
  OAI21_X1 U13953 ( .B1(n15100), .B2(n15074), .A(n12213), .ZN(n11406) );
  OAI211_X1 U13954 ( .C1(n11408), .C2(n15144), .A(n11407), .B(n11406), .ZN(
        P1_U3293) );
  NAND2_X1 U13955 ( .A1(n13588), .A2(n11409), .ZN(n11411) );
  OAI211_X1 U13956 ( .C1(n11412), .C2(n13624), .A(n11411), .B(n11410), .ZN(
        n11417) );
  XNOR2_X1 U13957 ( .A(n11414), .B(n11413), .ZN(n11415) );
  NOR2_X1 U13958 ( .A1(n11415), .A2(n13630), .ZN(n11416) );
  AOI211_X1 U13959 ( .C1(n11418), .C2(n13628), .A(n11417), .B(n11416), .ZN(
        n11419) );
  INV_X1 U13960 ( .A(n11419), .ZN(P2_U3185) );
  NAND2_X1 U13961 ( .A1(n12214), .A2(n14401), .ZN(n15084) );
  NOR2_X1 U13962 ( .A1(n15112), .A2(n15084), .ZN(n15081) );
  INV_X1 U13963 ( .A(n15081), .ZN(n11427) );
  OAI22_X1 U13964 ( .A1(n14577), .A2(n11420), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14648), .ZN(n11421) );
  AOI21_X1 U13965 ( .B1(n15074), .B2(n12227), .A(n11421), .ZN(n11425) );
  MUX2_X1 U13966 ( .A(n11423), .B(n11422), .S(n15103), .Z(n11424) );
  OAI211_X1 U13967 ( .C1(n11427), .C2(n11426), .A(n11425), .B(n11424), .ZN(
        P1_U3290) );
  XNOR2_X1 U13968 ( .A(n11428), .B(n11429), .ZN(n15402) );
  XNOR2_X1 U13969 ( .A(n11430), .B(n11429), .ZN(n11433) );
  NAND2_X1 U13970 ( .A1(n13610), .A2(n13665), .ZN(n11432) );
  NAND2_X1 U13971 ( .A1(n13622), .A2(n13667), .ZN(n11431) );
  AND2_X1 U13972 ( .A1(n11432), .A2(n11431), .ZN(n11614) );
  OAI21_X1 U13973 ( .B1(n11433), .B2(n13946), .A(n11614), .ZN(n15403) );
  NAND2_X1 U13974 ( .A1(n15403), .A2(n13963), .ZN(n11441) );
  INV_X1 U13975 ( .A(n11519), .ZN(n11434) );
  AOI211_X1 U13976 ( .C1(n15399), .C2(n11435), .A(n14001), .B(n11434), .ZN(
        n15397) );
  NOR2_X1 U13977 ( .A1(n13918), .A2(n7344), .ZN(n11439) );
  INV_X1 U13978 ( .A(n11612), .ZN(n11436) );
  OAI22_X1 U13979 ( .A1(n13963), .A2(n11437), .B1(n11436), .B2(n13957), .ZN(
        n11438) );
  AOI211_X1 U13980 ( .C1(n15397), .C2(n15319), .A(n11439), .B(n11438), .ZN(
        n11440) );
  OAI211_X1 U13981 ( .C1(n15402), .C2(n13966), .A(n11441), .B(n11440), .ZN(
        P2_U3256) );
  INV_X1 U13982 ( .A(n11442), .ZN(n11444) );
  OAI222_X1 U13983 ( .A1(n11445), .A2(n6665), .B1(n13439), .B2(n11444), .C1(
        n11443), .C2(n13441), .ZN(P3_U3271) );
  NAND2_X1 U13984 ( .A1(n11447), .A2(n11446), .ZN(n12819) );
  XNOR2_X1 U13985 ( .A(n12819), .B(n11448), .ZN(n11449) );
  NAND2_X1 U13986 ( .A1(n11449), .A2(n12924), .ZN(n11453) );
  AND2_X1 U13987 ( .A1(n6665), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15477) );
  OAI22_X1 U13988 ( .A1(n15542), .A2(n12917), .B1(n15546), .B2(n12931), .ZN(
        n11450) );
  AOI211_X1 U13989 ( .C1(n12914), .C2(n11451), .A(n15477), .B(n11450), .ZN(
        n11452) );
  OAI211_X1 U13990 ( .C1(n15547), .C2(n12896), .A(n11453), .B(n11452), .ZN(
        P3_U3153) );
  NAND2_X1 U13991 ( .A1(n11454), .A2(n12161), .ZN(n11457) );
  AOI22_X1 U13992 ( .A1(n11455), .A2(n12091), .B1(n12092), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U13993 ( .A1(n6678), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U13994 ( .A1(n11461), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11459) );
  INV_X1 U13995 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11458) );
  NAND2_X1 U13996 ( .A1(n11459), .A2(n11458), .ZN(n11462) );
  AND2_X1 U13997 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n11460) );
  NAND2_X1 U13998 ( .A1(n11461), .A2(n11460), .ZN(n11477) );
  NAND2_X1 U13999 ( .A1(n11462), .A2(n11477), .ZN(n14984) );
  INV_X1 U14000 ( .A(n14984), .ZN(n11463) );
  NAND2_X1 U14001 ( .A1(n12056), .A2(n11463), .ZN(n11466) );
  NAND2_X1 U14002 ( .A1(n10631), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11465) );
  NAND2_X1 U14003 ( .A1(n12156), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11464) );
  NAND4_X1 U14004 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n14260) );
  XNOR2_X1 U14005 ( .A(n15013), .B(n14137), .ZN(n12110) );
  OR2_X1 U14006 ( .A1(n14192), .A2(n14262), .ZN(n11469) );
  NAND2_X1 U14007 ( .A1(n11470), .A2(n12161), .ZN(n11473) );
  AOI22_X1 U14008 ( .A1(n11471), .A2(n12091), .B1(n12092), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14009 ( .A1(n11473), .A2(n11472), .ZN(n12638) );
  XNOR2_X1 U14010 ( .A(n12638), .B(n14971), .ZN(n12109) );
  OR2_X1 U14011 ( .A1(n12638), .A2(n14261), .ZN(n11474) );
  XOR2_X1 U14012 ( .A(n11674), .B(n12110), .Z(n15016) );
  INV_X1 U14013 ( .A(n12109), .ZN(n11529) );
  XOR2_X1 U14014 ( .A(n12110), .B(n11657), .Z(n11483) );
  NAND2_X1 U14015 ( .A1(n12156), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14016 ( .A1(n6678), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14017 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  AND2_X1 U14018 ( .A1(n11664), .A2(n11478), .ZN(n14161) );
  NAND2_X1 U14019 ( .A1(n12056), .A2(n14161), .ZN(n11480) );
  NAND2_X1 U14020 ( .A1(n10631), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14021 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n14259) );
  OAI222_X1 U14022 ( .A1(n15097), .A2(n14971), .B1(n11483), .B2(n15145), .C1(
        n15102), .C2(n14970), .ZN(n15018) );
  NAND2_X1 U14023 ( .A1(n15018), .A2(n15103), .ZN(n11487) );
  OAI22_X1 U14024 ( .A1(n15103), .A2(n10511), .B1(n14984), .B2(n14648), .ZN(
        n11485) );
  INV_X1 U14025 ( .A(n12638), .ZN(n15205) );
  INV_X1 U14026 ( .A(n15013), .ZN(n11658) );
  OAI211_X1 U14027 ( .C1(n11534), .C2(n11658), .A(n15077), .B(n11672), .ZN(
        n15014) );
  NOR2_X1 U14028 ( .A1(n15014), .A2(n14577), .ZN(n11484) );
  AOI211_X1 U14029 ( .C1(n15074), .C2(n15013), .A(n11485), .B(n11484), .ZN(
        n11486) );
  OAI211_X1 U14030 ( .C1(n14623), .C2(n15016), .A(n11487), .B(n11486), .ZN(
        P1_U3282) );
  AOI22_X1 U14031 ( .A1(n12770), .A2(n12233), .B1(n12768), .B2(n14267), .ZN(
        n11488) );
  XOR2_X1 U14032 ( .A(n11778), .B(n11488), .Z(n11543) );
  OAI22_X1 U14033 ( .A1(n12726), .A2(n12235), .B1(n12234), .B2(n10604), .ZN(
        n11540) );
  XOR2_X1 U14034 ( .A(n11544), .B(n11543), .Z(n11497) );
  NAND2_X1 U14035 ( .A1(n14981), .A2(n12233), .ZN(n11494) );
  AND2_X1 U14036 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14312) );
  AOI21_X1 U14037 ( .B1(n14214), .B2(n11492), .A(n14312), .ZN(n11493) );
  OAI211_X1 U14038 ( .C1(n14985), .C2(n11495), .A(n11494), .B(n11493), .ZN(
        n11496) );
  AOI21_X1 U14039 ( .B1(n11497), .B2(n14965), .A(n11496), .ZN(n11498) );
  INV_X1 U14040 ( .A(n11498), .ZN(P1_U3230) );
  XNOR2_X1 U14041 ( .A(n11500), .B(n11499), .ZN(n15649) );
  NAND2_X1 U14042 ( .A1(n11501), .A2(n15583), .ZN(n15646) );
  OAI22_X1 U14043 ( .A1(n11762), .A2(n15646), .B1(n15618), .B2(n11502), .ZN(
        n11510) );
  OAI211_X1 U14044 ( .C1(n11504), .C2(n12429), .A(n11503), .B(n15612), .ZN(
        n11508) );
  AOI22_X1 U14045 ( .A1(n15610), .A2(n11505), .B1(n12951), .B2(n15607), .ZN(
        n11507) );
  NAND2_X1 U14046 ( .A1(n15649), .A2(n15599), .ZN(n11506) );
  NAND3_X1 U14047 ( .A1(n11508), .A2(n11507), .A3(n11506), .ZN(n15647) );
  MUX2_X1 U14048 ( .A(n15647), .B(P3_REG2_REG_6__SCAN_IN), .S(n15625), .Z(
        n11509) );
  AOI211_X1 U14049 ( .C1(n15649), .C2(n13156), .A(n11510), .B(n11509), .ZN(
        n11511) );
  INV_X1 U14050 ( .A(n11511), .ZN(P3_U3227) );
  INV_X1 U14051 ( .A(n12061), .ZN(n11525) );
  XNOR2_X1 U14052 ( .A(n11512), .B(n7258), .ZN(n11516) );
  OAI22_X1 U14053 ( .A1(n11514), .A2(n13447), .B1(n13449), .B2(n11513), .ZN(
        n11629) );
  INV_X1 U14054 ( .A(n11629), .ZN(n11515) );
  OAI21_X1 U14055 ( .B1(n11516), .B2(n13946), .A(n11515), .ZN(n11730) );
  INV_X1 U14056 ( .A(n11730), .ZN(n11524) );
  XNOR2_X1 U14057 ( .A(n11517), .B(n11518), .ZN(n11732) );
  INV_X1 U14058 ( .A(n11737), .ZN(n11734) );
  AOI211_X1 U14059 ( .C1(n11737), .C2(n11519), .A(n14001), .B(n11606), .ZN(
        n11731) );
  NAND2_X1 U14060 ( .A1(n11731), .A2(n15319), .ZN(n11521) );
  AOI22_X1 U14061 ( .A1(n6674), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11626), 
        .B2(n15316), .ZN(n11520) );
  OAI211_X1 U14062 ( .C1(n11734), .C2(n13918), .A(n11521), .B(n11520), .ZN(
        n11522) );
  AOI21_X1 U14063 ( .B1(n11732), .B2(n15320), .A(n11522), .ZN(n11523) );
  OAI21_X1 U14064 ( .B1(n11524), .B2(n6674), .A(n11523), .ZN(P2_U3255) );
  OAI222_X1 U14065 ( .A1(n14106), .A2(n11526), .B1(P2_U3088), .B2(n8122), .C1(
        n14111), .C2(n11525), .ZN(P2_U3307) );
  XNOR2_X1 U14066 ( .A(n11527), .B(n12109), .ZN(n15209) );
  INV_X1 U14067 ( .A(n15209), .ZN(n11539) );
  OAI211_X1 U14068 ( .C1(n11530), .C2(n11529), .A(n11528), .B(n14645), .ZN(
        n11531) );
  OAI21_X1 U14069 ( .B1(n14138), .B2(n15097), .A(n11531), .ZN(n15206) );
  OAI21_X1 U14070 ( .B1(n11532), .B2(n15205), .A(n15077), .ZN(n11533) );
  OR2_X1 U14071 ( .A1(n11534), .A2(n11533), .ZN(n15203) );
  NAND2_X1 U14072 ( .A1(n14643), .A2(n14260), .ZN(n15202) );
  AOI21_X1 U14073 ( .B1(n15203), .B2(n15202), .A(n14577), .ZN(n11537) );
  AOI22_X1 U14074 ( .A1(n15112), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n14141), 
        .B2(n15099), .ZN(n11535) );
  OAI21_X1 U14075 ( .B1(n15205), .B2(n15106), .A(n11535), .ZN(n11536) );
  AOI211_X1 U14076 ( .C1(n15206), .C2(n15103), .A(n11537), .B(n11536), .ZN(
        n11538) );
  OAI21_X1 U14077 ( .B1(n14623), .B2(n11539), .A(n11538), .ZN(P1_U3283) );
  OAI22_X1 U14078 ( .A1(n12241), .A2(n10604), .B1(n12727), .B2(n15174), .ZN(
        n11547) );
  XNOR2_X1 U14079 ( .A(n11547), .B(n12756), .ZN(n11549) );
  OAI22_X1 U14080 ( .A1(n12726), .A2(n12241), .B1(n15174), .B2(n10604), .ZN(
        n11548) );
  NAND2_X1 U14081 ( .A1(n11549), .A2(n11548), .ZN(n11632) );
  NAND2_X1 U14082 ( .A1(n6834), .A2(n11632), .ZN(n11550) );
  XNOR2_X1 U14083 ( .A(n11633), .B(n11550), .ZN(n11557) );
  NAND2_X1 U14084 ( .A1(n14214), .A2(n11551), .ZN(n11553) );
  OAI211_X1 U14085 ( .C1(n14962), .C2(n15174), .A(n11553), .B(n11552), .ZN(
        n11554) );
  AOI21_X1 U14086 ( .B1(n11555), .B2(n14244), .A(n11554), .ZN(n11556) );
  OAI21_X1 U14087 ( .B1(n11557), .B2(n14976), .A(n11556), .ZN(P1_U3227) );
  NOR2_X1 U14088 ( .A1(n11572), .A2(n11558), .ZN(n11560) );
  NAND2_X1 U14089 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11899), .ZN(n11561) );
  OAI21_X1 U14090 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11899), .A(n11561), 
        .ZN(n11562) );
  AOI21_X1 U14091 ( .B1(n6815), .B2(n11562), .A(n11894), .ZN(n11584) );
  AOI22_X1 U14092 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11899), .B1(n11574), 
        .B2(n8389), .ZN(n11568) );
  NAND2_X1 U14093 ( .A1(n11564), .A2(n11563), .ZN(n11566) );
  OAI21_X1 U14094 ( .B1(n11568), .B2(n11567), .A(n11896), .ZN(n11582) );
  NOR2_X1 U14095 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11569), .ZN(n11862) );
  AOI21_X1 U14096 ( .B1(n15516), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11862), 
        .ZN(n11570) );
  OAI21_X1 U14097 ( .B1(n15513), .B2(n11899), .A(n11570), .ZN(n11581) );
  INV_X1 U14098 ( .A(n11571), .ZN(n11573) );
  NAND2_X1 U14099 ( .A1(n11573), .A2(n11572), .ZN(n11576) );
  MUX2_X1 U14100 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12990), .Z(n11900) );
  XNOR2_X1 U14101 ( .A(n11900), .B(n11574), .ZN(n11575) );
  NAND3_X1 U14102 ( .A1(n11577), .A2(n11576), .A3(n11575), .ZN(n11903) );
  INV_X1 U14103 ( .A(n11903), .ZN(n11579) );
  AOI21_X1 U14104 ( .B1(n11577), .B2(n11576), .A(n11575), .ZN(n11578) );
  NOR3_X1 U14105 ( .A1(n11579), .A2(n11578), .A3(n15439), .ZN(n11580) );
  AOI211_X1 U14106 ( .C1(n15519), .C2(n11582), .A(n11581), .B(n11580), .ZN(
        n11583) );
  OAI21_X1 U14107 ( .B1(n11584), .B2(n15523), .A(n11583), .ZN(P3_U3194) );
  AOI21_X1 U14108 ( .B1(n15529), .B2(n12936), .A(n11585), .ZN(n11587) );
  NAND2_X1 U14109 ( .A1(n12914), .A2(n15528), .ZN(n11586) );
  OAI211_X1 U14110 ( .C1(n12931), .C2(n15534), .A(n11587), .B(n11586), .ZN(
        n11593) );
  OR2_X1 U14111 ( .A1(n11323), .A2(n11588), .ZN(n11590) );
  AOI211_X1 U14112 ( .C1(n11591), .C2(n11590), .A(n12945), .B(n11589), .ZN(
        n11592) );
  AOI211_X1 U14113 ( .C1(n15531), .C2(n12938), .A(n11593), .B(n11592), .ZN(
        n11594) );
  INV_X1 U14114 ( .A(n11594), .ZN(P3_U3157) );
  INV_X1 U14115 ( .A(n11595), .ZN(n11596) );
  OAI222_X1 U14116 ( .A1(n6665), .A2(n11598), .B1(n13441), .B2(n11597), .C1(
        n13439), .C2(n11596), .ZN(P3_U3270) );
  XNOR2_X1 U14117 ( .A(n11599), .B(n11603), .ZN(n11602) );
  NAND2_X1 U14118 ( .A1(n13610), .A2(n13663), .ZN(n11601) );
  NAND2_X1 U14119 ( .A1(n13622), .A2(n13665), .ZN(n11600) );
  NAND2_X1 U14120 ( .A1(n11601), .A2(n11600), .ZN(n13603) );
  AOI21_X1 U14121 ( .B1(n11602), .B2(n14882), .A(n13603), .ZN(n15411) );
  XOR2_X1 U14122 ( .A(n11604), .B(n11603), .Z(n15413) );
  INV_X1 U14123 ( .A(n15413), .ZN(n15416) );
  INV_X1 U14124 ( .A(n11794), .ZN(n11605) );
  OAI211_X1 U14125 ( .C1(n15410), .C2(n11606), .A(n11605), .B(n9576), .ZN(
        n15408) );
  AOI22_X1 U14126 ( .A1(n6674), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n13599), 
        .B2(n15316), .ZN(n11609) );
  NAND2_X1 U14127 ( .A1(n11607), .A2(n15314), .ZN(n11608) );
  OAI211_X1 U14128 ( .C1(n15408), .C2(n13961), .A(n11609), .B(n11608), .ZN(
        n11610) );
  AOI21_X1 U14129 ( .B1(n15416), .B2(n15320), .A(n11610), .ZN(n11611) );
  OAI21_X1 U14130 ( .B1(n6674), .B2(n15411), .A(n11611), .ZN(P2_U3254) );
  NAND2_X1 U14131 ( .A1(n13588), .A2(n11612), .ZN(n11613) );
  NAND2_X1 U14132 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n15263) );
  OAI211_X1 U14133 ( .C1(n11614), .C2(n13624), .A(n11613), .B(n15263), .ZN(
        n11620) );
  NAND2_X1 U14134 ( .A1(n11615), .A2(n11616), .ZN(n11617) );
  AOI21_X1 U14135 ( .B1(n11618), .B2(n11617), .A(n13630), .ZN(n11619) );
  AOI211_X1 U14136 ( .C1(n15399), .C2(n13628), .A(n11620), .B(n11619), .ZN(
        n11621) );
  INV_X1 U14137 ( .A(n11621), .ZN(P2_U3203) );
  INV_X1 U14138 ( .A(n12041), .ZN(n12609) );
  OAI222_X1 U14139 ( .A1(P1_U3086), .A2(n12194), .B1(n14775), .B2(n12609), 
        .C1(n12042), .C2(n14772), .ZN(P1_U3334) );
  AOI21_X1 U14140 ( .B1(n11623), .B2(n11622), .A(n13630), .ZN(n11625) );
  NAND2_X1 U14141 ( .A1(n11625), .A2(n11624), .ZN(n11631) );
  INV_X1 U14142 ( .A(n11626), .ZN(n11627) );
  OAI22_X1 U14143 ( .A1(n13638), .A2(n11627), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9343), .ZN(n11628) );
  AOI21_X1 U14144 ( .B1(n13641), .B2(n11629), .A(n11628), .ZN(n11630) );
  OAI211_X1 U14145 ( .C1(n11734), .C2(n13644), .A(n11631), .B(n11630), .ZN(
        P2_U3189) );
  INV_X1 U14146 ( .A(n15073), .ZN(n11643) );
  OAI22_X1 U14147 ( .A1(n15180), .A2(n12727), .B1(n10604), .B2(n11634), .ZN(
        n11635) );
  XNOR2_X1 U14148 ( .A(n11635), .B(n11778), .ZN(n11773) );
  AOI22_X1 U14149 ( .A1(n12767), .A2(n14265), .B1(n12769), .B2(n15075), .ZN(
        n11775) );
  XNOR2_X1 U14150 ( .A(n11773), .B(n11775), .ZN(n11636) );
  OAI211_X1 U14151 ( .C1(n11637), .C2(n11636), .A(n11776), .B(n14965), .ZN(
        n11642) );
  INV_X1 U14152 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n14328) );
  OR2_X1 U14153 ( .A1(n15102), .A2(n11777), .ZN(n11638) );
  OAI21_X1 U14154 ( .B1(n15097), .B2(n12241), .A(n11638), .ZN(n15071) );
  NAND2_X1 U14155 ( .A1(n14214), .A2(n15071), .ZN(n11639) );
  OAI21_X1 U14156 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n14328), .A(n11639), .ZN(
        n11640) );
  AOI21_X1 U14157 ( .B1(n14981), .B2(n15075), .A(n11640), .ZN(n11641) );
  OAI211_X1 U14158 ( .C1(n14985), .C2(n11643), .A(n11642), .B(n11641), .ZN(
        P1_U3239) );
  XNOR2_X1 U14159 ( .A(n11644), .B(n12430), .ZN(n11650) );
  AND2_X1 U14160 ( .A1(n11765), .A2(n11645), .ZN(n11647) );
  NAND2_X1 U14161 ( .A1(n11765), .A2(n11646), .ZN(n15526) );
  OAI211_X1 U14162 ( .C1(n11647), .C2(n12430), .A(n15612), .B(n15526), .ZN(
        n11649) );
  AOI22_X1 U14163 ( .A1(n15610), .A2(n12491), .B1(n11807), .B2(n15607), .ZN(
        n11648) );
  OAI211_X1 U14164 ( .C1(n15616), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n15660) );
  INV_X1 U14165 ( .A(n15660), .ZN(n11656) );
  INV_X1 U14166 ( .A(n11650), .ZN(n15663) );
  NOR2_X1 U14167 ( .A1(n11651), .A2(n15605), .ZN(n15661) );
  AOI22_X1 U14168 ( .A1(n15577), .A2(n15661), .B1(n15576), .B2(n11652), .ZN(
        n11653) );
  OAI21_X1 U14169 ( .B1(n11165), .B2(n15623), .A(n11653), .ZN(n11654) );
  AOI21_X1 U14170 ( .B1(n15663), .B2(n13156), .A(n11654), .ZN(n11655) );
  OAI21_X1 U14171 ( .B1(n11656), .B2(n15625), .A(n11655), .ZN(P3_U3224) );
  NAND2_X1 U14172 ( .A1(n11659), .A2(n12161), .ZN(n11662) );
  AOI22_X1 U14173 ( .A1(n11660), .A2(n12091), .B1(n12092), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11661) );
  XNOR2_X1 U14174 ( .A(n14172), .B(n14970), .ZN(n12111) );
  XNOR2_X1 U14175 ( .A(n11709), .B(n12111), .ZN(n11671) );
  NAND2_X1 U14176 ( .A1(n6678), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11669) );
  AND2_X1 U14177 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  NOR2_X1 U14178 ( .A1(n11711), .A2(n11665), .ZN(n14212) );
  NAND2_X1 U14179 ( .A1(n12056), .A2(n14212), .ZN(n11668) );
  NAND2_X1 U14180 ( .A1(n10631), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14181 ( .A1(n12156), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14182 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n14258) );
  INV_X1 U14183 ( .A(n14258), .ZN(n14930) );
  OR2_X1 U14184 ( .A1(n15102), .A2(n14930), .ZN(n11670) );
  OAI21_X1 U14185 ( .B1(n15097), .B2(n14137), .A(n11670), .ZN(n14163) );
  AOI21_X1 U14186 ( .B1(n11671), .B2(n14645), .A(n14163), .ZN(n11696) );
  AOI211_X1 U14187 ( .C1(n14172), .C2(n11672), .A(n15159), .B(n7015), .ZN(
        n11694) );
  INV_X1 U14188 ( .A(n14172), .ZN(n11707) );
  AOI22_X1 U14189 ( .A1(n15112), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14161), 
        .B2(n15099), .ZN(n11673) );
  OAI21_X1 U14190 ( .B1(n11707), .B2(n15106), .A(n11673), .ZN(n11678) );
  INV_X1 U14191 ( .A(n12111), .ZN(n11708) );
  NAND2_X1 U14192 ( .A1(n15013), .A2(n14260), .ZN(n11675) );
  AOI21_X1 U14193 ( .B1(n11708), .B2(n11676), .A(n6817), .ZN(n11697) );
  NOR2_X1 U14194 ( .A1(n11697), .A2(n14623), .ZN(n11677) );
  AOI211_X1 U14195 ( .C1(n11694), .C2(n15080), .A(n11678), .B(n11677), .ZN(
        n11679) );
  OAI21_X1 U14196 ( .B1(n11696), .B2(n15112), .A(n11679), .ZN(P1_U3281) );
  INV_X1 U14197 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11680) );
  MUX2_X1 U14198 ( .A(n11680), .B(P2_REG2_REG_13__SCAN_IN), .S(n11849), .Z(
        n11850) );
  AOI21_X1 U14199 ( .B1(n11340), .B2(n11682), .A(n11681), .ZN(n11852) );
  XOR2_X1 U14200 ( .A(n11850), .B(n11852), .Z(n11693) );
  NAND2_X1 U14201 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n13581)
         );
  INV_X1 U14202 ( .A(n13581), .ZN(n11683) );
  AOI21_X1 U14203 ( .B1(n15305), .B2(n11849), .A(n11683), .ZN(n11684) );
  INV_X1 U14204 ( .A(n11684), .ZN(n11691) );
  INV_X1 U14205 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11685) );
  MUX2_X1 U14206 ( .A(n11685), .B(P2_REG1_REG_13__SCAN_IN), .S(n11849), .Z(
        n11689) );
  OAI21_X1 U14207 ( .B1(n11687), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11686), 
        .ZN(n11688) );
  NOR2_X1 U14208 ( .A1(n11688), .A2(n11689), .ZN(n11843) );
  AOI211_X1 U14209 ( .C1(n11689), .C2(n11688), .A(n15298), .B(n11843), .ZN(
        n11690) );
  AOI211_X1 U14210 ( .C1(n15289), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n11691), 
        .B(n11690), .ZN(n11692) );
  OAI21_X1 U14211 ( .B1(n11693), .B2(n15279), .A(n11692), .ZN(P2_U3227) );
  INV_X1 U14212 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11699) );
  AOI21_X1 U14213 ( .B1(n14172), .B2(n15156), .A(n11694), .ZN(n11695) );
  OAI211_X1 U14214 ( .C1(n15146), .C2(n11697), .A(n11696), .B(n11695), .ZN(
        n11700) );
  NAND2_X1 U14215 ( .A1(n11700), .A2(n15212), .ZN(n11698) );
  OAI21_X1 U14216 ( .B1(n15212), .B2(n11699), .A(n11698), .ZN(P1_U3495) );
  NAND2_X1 U14217 ( .A1(n11700), .A2(n15225), .ZN(n11701) );
  OAI21_X1 U14218 ( .B1(n15225), .B2(n11702), .A(n11701), .ZN(P1_U3540) );
  NAND2_X1 U14219 ( .A1(n11703), .A2(n12161), .ZN(n11706) );
  AOI22_X1 U14220 ( .A1(n11704), .A2(n12091), .B1(n12092), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11705) );
  XNOR2_X1 U14221 ( .A(n12662), .B(n14258), .ZN(n12112) );
  AOI211_X1 U14222 ( .C1(n11719), .C2(n11710), .A(n15145), .B(n11931), .ZN(
        n11718) );
  NOR2_X1 U14223 ( .A1(n11711), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11712) );
  OR2_X1 U14224 ( .A1(n11924), .A2(n11712), .ZN(n14941) );
  INV_X1 U14225 ( .A(n14941), .ZN(n11947) );
  NAND2_X1 U14226 ( .A1(n11947), .A2(n12056), .ZN(n11716) );
  NAND2_X1 U14227 ( .A1(n6678), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14228 ( .A1(n10631), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U14229 ( .A1(n12156), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14230 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n14257) );
  INV_X1 U14231 ( .A(n14257), .ZN(n12667) );
  OR2_X1 U14232 ( .A1(n15102), .A2(n12667), .ZN(n11717) );
  OAI21_X1 U14233 ( .B1(n15097), .B2(n14970), .A(n11717), .ZN(n14213) );
  NOR2_X1 U14234 ( .A1(n11718), .A2(n14213), .ZN(n11831) );
  OAI21_X1 U14235 ( .B1(n11720), .B2(n11719), .A(n11913), .ZN(n11828) );
  AOI211_X1 U14236 ( .C1(n12662), .C2(n11721), .A(n15159), .B(n6824), .ZN(
        n11829) );
  NAND2_X1 U14237 ( .A1(n11829), .A2(n15080), .ZN(n11723) );
  AOI22_X1 U14238 ( .A1(n15112), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n14212), 
        .B2(n15099), .ZN(n11722) );
  OAI211_X1 U14239 ( .C1(n7313), .C2(n15106), .A(n11723), .B(n11722), .ZN(
        n11724) );
  AOI21_X1 U14240 ( .B1(n11828), .B2(n14654), .A(n11724), .ZN(n11725) );
  OAI21_X1 U14241 ( .B1(n11831), .B2(n15112), .A(n11725), .ZN(P1_U3280) );
  INV_X1 U14242 ( .A(n11726), .ZN(n11727) );
  OAI222_X1 U14243 ( .A1(P3_U3151), .A2(n11729), .B1(n13441), .B2(n11728), 
        .C1(n12381), .C2(n11727), .ZN(P3_U3269) );
  AOI211_X1 U14244 ( .C1(n15370), .C2(n11732), .A(n11731), .B(n11730), .ZN(
        n11739) );
  INV_X1 U14245 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11733) );
  OAI22_X1 U14246 ( .A1(n11734), .A2(n14081), .B1(n15420), .B2(n11733), .ZN(
        n11735) );
  INV_X1 U14247 ( .A(n11735), .ZN(n11736) );
  OAI21_X1 U14248 ( .B1(n11739), .B2(n15418), .A(n11736), .ZN(P2_U3460) );
  AOI22_X1 U14249 ( .A1(n9569), .A2(n11737), .B1(n15429), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11738) );
  OAI21_X1 U14250 ( .B1(n11739), .B2(n15429), .A(n11738), .ZN(P2_U3509) );
  INV_X1 U14251 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15007) );
  NOR2_X1 U14252 ( .A1(n12087), .A2(n15007), .ZN(n11740) );
  AOI21_X1 U14253 ( .B1(n12087), .B2(n15007), .A(n11740), .ZN(n11745) );
  INV_X1 U14254 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15051) );
  OAI21_X1 U14255 ( .B1(n11743), .B2(n11921), .A(n15050), .ZN(n11744) );
  NOR2_X1 U14256 ( .A1(n11744), .A2(n11745), .ZN(n11872) );
  AOI211_X1 U14257 ( .C1(n11745), .C2(n11744), .A(n14396), .B(n11872), .ZN(
        n11759) );
  INV_X1 U14258 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11749) );
  MUX2_X1 U14259 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11749), .S(n11756), .Z(
        n11753) );
  AOI21_X1 U14260 ( .B1(n11916), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11746), 
        .ZN(n11747) );
  NAND2_X1 U14261 ( .A1(n11747), .A2(n15056), .ZN(n11751) );
  XNOR2_X1 U14262 ( .A(n11747), .B(n15056), .ZN(n15054) );
  NOR2_X1 U14263 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15054), .ZN(n15053) );
  INV_X1 U14264 ( .A(n15053), .ZN(n11748) );
  NAND2_X1 U14265 ( .A1(n11751), .A2(n11748), .ZN(n11752) );
  AOI21_X1 U14266 ( .B1(n11756), .B2(n11749), .A(n15053), .ZN(n11750) );
  OAI211_X1 U14267 ( .C1(n11749), .C2(n11756), .A(n11751), .B(n11750), .ZN(
        n11877) );
  INV_X1 U14268 ( .A(n11877), .ZN(n11881) );
  AOI211_X1 U14269 ( .C1(n11753), .C2(n11752), .A(n15057), .B(n11881), .ZN(
        n11758) );
  NAND2_X1 U14270 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14952)
         );
  INV_X1 U14271 ( .A(n14952), .ZN(n11754) );
  AOI21_X1 U14272 ( .B1(n14365), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11754), 
        .ZN(n11755) );
  OAI21_X1 U14273 ( .B1(n15055), .B2(n11756), .A(n11755), .ZN(n11757) );
  OR3_X1 U14274 ( .A1(n11759), .A2(n11758), .A3(n11757), .ZN(P1_U3259) );
  XNOR2_X1 U14275 ( .A(n11760), .B(n8334), .ZN(n11769) );
  INV_X1 U14276 ( .A(n11769), .ZN(n15658) );
  NAND2_X1 U14277 ( .A1(n12824), .A2(n15583), .ZN(n15655) );
  OAI22_X1 U14278 ( .A1(n11762), .A2(n15655), .B1(n15618), .B2(n11761), .ZN(
        n11771) );
  NAND2_X1 U14279 ( .A1(n11763), .A2(n12488), .ZN(n11764) );
  NAND2_X1 U14280 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  NAND2_X1 U14281 ( .A1(n11766), .A2(n15612), .ZN(n11768) );
  AOI22_X1 U14282 ( .A1(n15610), .A2(n12951), .B1(n15528), .B2(n15607), .ZN(
        n11767) );
  OAI211_X1 U14283 ( .C1(n15616), .C2(n11769), .A(n11768), .B(n11767), .ZN(
        n15656) );
  MUX2_X1 U14284 ( .A(n15656), .B(P3_REG2_REG_8__SCAN_IN), .S(n15625), .Z(
        n11770) );
  AOI211_X1 U14285 ( .C1(n13156), .C2(n15658), .A(n11771), .B(n11770), .ZN(
        n11772) );
  INV_X1 U14286 ( .A(n11772), .ZN(P3_U3225) );
  INV_X1 U14287 ( .A(n11773), .ZN(n11774) );
  OAI22_X1 U14288 ( .A1(n11782), .A2(n12727), .B1(n10604), .B2(n11777), .ZN(
        n11779) );
  XNOR2_X1 U14289 ( .A(n11779), .B(n11778), .ZN(n11959) );
  AOI22_X1 U14290 ( .A1(n12767), .A2(n14264), .B1(n12768), .B2(n12251), .ZN(
        n11961) );
  XNOR2_X1 U14291 ( .A(n11959), .B(n11961), .ZN(n11780) );
  OAI211_X1 U14292 ( .C1(n11781), .C2(n11780), .A(n11962), .B(n14965), .ZN(
        n11786) );
  NOR2_X1 U14293 ( .A1(n15204), .A2(n11782), .ZN(n15189) );
  NAND2_X1 U14294 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14343) );
  OAI21_X1 U14295 ( .B1(n14203), .B2(n11783), .A(n14343), .ZN(n11784) );
  AOI21_X1 U14296 ( .B1(n14118), .B2(n15189), .A(n11784), .ZN(n11785) );
  OAI211_X1 U14297 ( .C1(n14985), .C2(n11787), .A(n11786), .B(n11785), .ZN(
        P1_U3213) );
  XOR2_X1 U14298 ( .A(n11793), .B(n11788), .Z(n11791) );
  NAND2_X1 U14299 ( .A1(n13610), .A2(n13662), .ZN(n11790) );
  NAND2_X1 U14300 ( .A1(n13551), .A2(n13664), .ZN(n11789) );
  NAND2_X1 U14301 ( .A1(n11790), .A2(n11789), .ZN(n13521) );
  AOI21_X1 U14302 ( .B1(n11791), .B2(n14882), .A(n13521), .ZN(n14917) );
  XOR2_X1 U14303 ( .A(n11793), .B(n11792), .Z(n14918) );
  INV_X1 U14304 ( .A(n14918), .ZN(n14921) );
  OAI211_X1 U14305 ( .C1(n11794), .C2(n14916), .A(n9576), .B(n11822), .ZN(
        n14915) );
  AOI22_X1 U14306 ( .A1(n6674), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n13518), 
        .B2(n15316), .ZN(n11797) );
  NAND2_X1 U14307 ( .A1(n11795), .A2(n15314), .ZN(n11796) );
  OAI211_X1 U14308 ( .C1(n14915), .C2(n13961), .A(n11797), .B(n11796), .ZN(
        n11798) );
  AOI21_X1 U14309 ( .B1(n14921), .B2(n15320), .A(n11798), .ZN(n11799) );
  OAI21_X1 U14310 ( .B1(n6674), .B2(n14917), .A(n11799), .ZN(P2_U3253) );
  INV_X1 U14311 ( .A(n11800), .ZN(n11802) );
  OAI222_X1 U14312 ( .A1(n6665), .A2(n12990), .B1(n13439), .B2(n11802), .C1(
        n11801), .C2(n13441), .ZN(P3_U3268) );
  XNOR2_X1 U14313 ( .A(n11803), .B(n15529), .ZN(n11813) );
  AOI21_X1 U14314 ( .B1(n11805), .B2(n12936), .A(n11804), .ZN(n11811) );
  NAND2_X1 U14315 ( .A1(n12943), .A2(n12507), .ZN(n11810) );
  INV_X1 U14316 ( .A(n11806), .ZN(n14866) );
  NAND2_X1 U14317 ( .A1(n12938), .A2(n14866), .ZN(n11809) );
  NAND2_X1 U14318 ( .A1(n12914), .A2(n11807), .ZN(n11808) );
  NAND4_X1 U14319 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  AOI21_X1 U14320 ( .B1(n11813), .B2(n12924), .A(n11812), .ZN(n11814) );
  INV_X1 U14321 ( .A(n11814), .ZN(P3_U3176) );
  XNOR2_X1 U14322 ( .A(n11815), .B(n11820), .ZN(n11818) );
  NAND2_X1 U14323 ( .A1(n13610), .A2(n13661), .ZN(n11817) );
  NAND2_X1 U14324 ( .A1(n13551), .A2(n13663), .ZN(n11816) );
  NAND2_X1 U14325 ( .A1(n11817), .A2(n11816), .ZN(n13584) );
  AOI21_X1 U14326 ( .B1(n11818), .B2(n14882), .A(n13584), .ZN(n14911) );
  XOR2_X1 U14327 ( .A(n11820), .B(n11819), .Z(n14914) );
  INV_X1 U14328 ( .A(n11823), .ZN(n14910) );
  INV_X1 U14329 ( .A(n11821), .ZN(n14892) );
  AOI211_X1 U14330 ( .C1(n11823), .C2(n11822), .A(n14001), .B(n14892), .ZN(
        n14908) );
  NAND2_X1 U14331 ( .A1(n14908), .A2(n15319), .ZN(n11825) );
  AOI22_X1 U14332 ( .A1(n6674), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13580), 
        .B2(n15316), .ZN(n11824) );
  OAI211_X1 U14333 ( .C1(n14910), .C2(n13918), .A(n11825), .B(n11824), .ZN(
        n11826) );
  AOI21_X1 U14334 ( .B1(n14914), .B2(n15320), .A(n11826), .ZN(n11827) );
  OAI21_X1 U14335 ( .B1(n6674), .B2(n14911), .A(n11827), .ZN(P2_U3252) );
  INV_X1 U14336 ( .A(n11828), .ZN(n11832) );
  AOI21_X1 U14337 ( .B1(n12662), .B2(n15156), .A(n11829), .ZN(n11830) );
  OAI211_X1 U14338 ( .C1(n15146), .C2(n11832), .A(n11831), .B(n11830), .ZN(
        n11835) );
  NAND2_X1 U14339 ( .A1(n11835), .A2(n15225), .ZN(n11833) );
  OAI21_X1 U14340 ( .B1(n15225), .B2(n11834), .A(n11833), .ZN(P1_U3541) );
  INV_X1 U14341 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U14342 ( .A1(n11835), .A2(n15212), .ZN(n11836) );
  OAI21_X1 U14343 ( .B1(n15212), .B2(n11837), .A(n11836), .ZN(P1_U3498) );
  INV_X1 U14344 ( .A(n11838), .ZN(n11839) );
  OAI222_X1 U14345 ( .A1(n14106), .A2(n11840), .B1(n14111), .B2(n11839), .C1(
        n6685), .C2(P2_U3088), .ZN(P2_U3305) );
  AND2_X1 U14346 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n11841) );
  AOI21_X1 U14347 ( .B1(n15305), .B2(n13681), .A(n11841), .ZN(n11842) );
  INV_X1 U14348 ( .A(n11842), .ZN(n11848) );
  INV_X1 U14349 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11844) );
  MUX2_X1 U14350 ( .A(n11844), .B(P2_REG1_REG_14__SCAN_IN), .S(n13681), .Z(
        n11845) );
  AOI211_X1 U14351 ( .C1(n11846), .C2(n11845), .A(n13675), .B(n15298), .ZN(
        n11847) );
  AOI211_X1 U14352 ( .C1(n15289), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11848), 
        .B(n11847), .ZN(n11858) );
  NAND2_X1 U14353 ( .A1(n11849), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11854) );
  INV_X1 U14354 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U14355 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U14356 ( .A1(n11854), .A2(n11853), .ZN(n13680) );
  XNOR2_X1 U14357 ( .A(n13680), .B(n11855), .ZN(n11856) );
  NAND2_X1 U14358 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n11856), .ZN(n13682) );
  OAI211_X1 U14359 ( .C1(n11856), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15307), 
        .B(n13682), .ZN(n11857) );
  NAND2_X1 U14360 ( .A1(n11858), .A2(n11857), .ZN(P2_U3228) );
  NAND2_X1 U14361 ( .A1(n7223), .A2(n11860), .ZN(n11861) );
  XNOR2_X1 U14362 ( .A(n11859), .B(n11861), .ZN(n11869) );
  AOI21_X1 U14363 ( .B1(n14851), .B2(n12936), .A(n11862), .ZN(n11867) );
  NAND2_X1 U14364 ( .A1(n14854), .A2(n12943), .ZN(n11866) );
  INV_X1 U14365 ( .A(n11863), .ZN(n14855) );
  NAND2_X1 U14366 ( .A1(n12938), .A2(n14855), .ZN(n11865) );
  NAND2_X1 U14367 ( .A1(n12914), .A2(n15529), .ZN(n11864) );
  NAND4_X1 U14368 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  AOI21_X1 U14369 ( .B1(n11869), .B2(n12924), .A(n11868), .ZN(n11870) );
  INV_X1 U14370 ( .A(n11870), .ZN(P3_U3164) );
  NOR2_X1 U14371 ( .A1(n14373), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11871) );
  AOI21_X1 U14372 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14373), .A(n11871), 
        .ZN(n11874) );
  AOI21_X1 U14373 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n12087), .A(n11872), 
        .ZN(n11873) );
  NOR2_X1 U14374 ( .A1(n11873), .A2(n11874), .ZN(n14374) );
  AOI211_X1 U14375 ( .C1(n11874), .C2(n11873), .A(n14396), .B(n14374), .ZN(
        n11886) );
  INV_X1 U14376 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14999) );
  OR2_X1 U14377 ( .A1(n14375), .A2(n14999), .ZN(n11875) );
  NAND2_X1 U14378 ( .A1(n12087), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11876) );
  OAI211_X1 U14379 ( .C1(n14373), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11875), 
        .B(n11876), .ZN(n11880) );
  NAND2_X1 U14380 ( .A1(n11877), .A2(n11876), .ZN(n11879) );
  NAND2_X1 U14381 ( .A1(n14375), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11878) );
  OAI211_X1 U14382 ( .C1(n14375), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11879), 
        .B(n11878), .ZN(n14372) );
  OAI211_X1 U14383 ( .C1(n11881), .C2(n11880), .A(n14372), .B(n14400), .ZN(
        n11884) );
  NAND2_X1 U14384 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14967)
         );
  INV_X1 U14385 ( .A(n14967), .ZN(n11882) );
  AOI21_X1 U14386 ( .B1(n14365), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11882), 
        .ZN(n11883) );
  OAI211_X1 U14387 ( .C1(n15055), .C2(n14373), .A(n11884), .B(n11883), .ZN(
        n11885) );
  OR2_X1 U14388 ( .A1(n11886), .A2(n11885), .ZN(P1_U3260) );
  NAND2_X1 U14389 ( .A1(n12144), .A2(n14098), .ZN(n11888) );
  OAI211_X1 U14390 ( .C1(n11889), .C2(n14106), .A(n11888), .B(n11887), .ZN(
        P2_U3304) );
  INV_X1 U14391 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U14392 ( .A1(n12144), .A2(n11890), .ZN(n11891) );
  OAI211_X1 U14393 ( .C1(n12145), .C2(n14777), .A(n11891), .B(n12374), .ZN(
        P1_U3332) );
  INV_X1 U14394 ( .A(n12134), .ZN(n12376) );
  OAI222_X1 U14395 ( .A1(n14106), .A2(n11893), .B1(n14111), .B2(n12376), .C1(
        n11892), .C2(P2_U3088), .ZN(P2_U3303) );
  XOR2_X1 U14396 ( .A(n12958), .B(n12952), .Z(n11895) );
  NOR2_X1 U14397 ( .A1(n13291), .A2(n11895), .ZN(n12953) );
  AOI21_X1 U14398 ( .B1(n13291), .B2(n11895), .A(n12953), .ZN(n11911) );
  INV_X1 U14399 ( .A(n12958), .ZN(n12964) );
  NAND2_X1 U14400 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11899), .ZN(n11897) );
  NAND2_X1 U14401 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11898), .ZN(n12959) );
  OAI21_X1 U14402 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11898), .A(n12959), 
        .ZN(n11909) );
  NAND2_X1 U14403 ( .A1(n11900), .A2(n11899), .ZN(n11902) );
  MUX2_X1 U14404 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12990), .Z(n12963) );
  XNOR2_X1 U14405 ( .A(n12963), .B(n12964), .ZN(n11901) );
  NAND3_X1 U14406 ( .A1(n11903), .A2(n11902), .A3(n11901), .ZN(n12970) );
  INV_X1 U14407 ( .A(n12970), .ZN(n11905) );
  AOI21_X1 U14408 ( .B1(n11903), .B2(n11902), .A(n11901), .ZN(n11904) );
  OAI21_X1 U14409 ( .B1(n11905), .B2(n11904), .A(n15508), .ZN(n11907) );
  NOR2_X1 U14410 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8417), .ZN(n12893) );
  AOI21_X1 U14411 ( .B1(n15516), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12893), 
        .ZN(n11906) );
  OAI211_X1 U14412 ( .C1(n15513), .C2(n12958), .A(n11907), .B(n11906), .ZN(
        n11908) );
  AOI21_X1 U14413 ( .B1(n15519), .B2(n11909), .A(n11908), .ZN(n11910) );
  OAI21_X1 U14414 ( .B1(n11911), .B2(n15523), .A(n11910), .ZN(P3_U3195) );
  OR2_X1 U14415 ( .A1(n12662), .A2(n14258), .ZN(n11912) );
  NAND2_X1 U14416 ( .A1(n11913), .A2(n11912), .ZN(n11950) );
  NAND2_X1 U14417 ( .A1(n11915), .A2(n12161), .ZN(n11918) );
  AOI22_X1 U14418 ( .A1(n11916), .A2(n12091), .B1(n12092), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11917) );
  OR2_X1 U14419 ( .A1(n14938), .A2(n12667), .ZN(n12279) );
  NAND2_X1 U14420 ( .A1(n14938), .A2(n12667), .ZN(n12283) );
  NAND2_X1 U14421 ( .A1(n12279), .A2(n12283), .ZN(n12278) );
  INV_X1 U14422 ( .A(n12278), .ZN(n12290) );
  NAND2_X1 U14423 ( .A1(n14938), .A2(n14257), .ZN(n11919) );
  NAND2_X1 U14424 ( .A1(n11920), .A2(n12161), .ZN(n11923) );
  AOI22_X1 U14425 ( .A1(n12092), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12091), 
        .B2(n11921), .ZN(n11922) );
  OR2_X1 U14426 ( .A1(n11924), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U14427 ( .A1(n11935), .A2(n11925), .ZN(n14250) );
  NAND2_X1 U14428 ( .A1(n12156), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U14429 ( .A1(n6678), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11926) );
  AND2_X1 U14430 ( .A1(n11927), .A2(n11926), .ZN(n11929) );
  NAND2_X1 U14431 ( .A1(n10631), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11928) );
  OAI211_X1 U14432 ( .C1(n14250), .C2(n10983), .A(n11929), .B(n11928), .ZN(
        n14642) );
  INV_X1 U14433 ( .A(n14642), .ZN(n14943) );
  NAND2_X1 U14434 ( .A1(n14416), .A2(n14943), .ZN(n12287) );
  NAND2_X1 U14435 ( .A1(n14431), .A2(n12287), .ZN(n14415) );
  XNOR2_X1 U14436 ( .A(n14414), .B(n7582), .ZN(n11978) );
  INV_X1 U14437 ( .A(n11978), .ZN(n11945) );
  NAND2_X1 U14438 ( .A1(n14416), .A2(n11951), .ZN(n11930) );
  NAND2_X1 U14439 ( .A1(n14647), .A2(n11930), .ZN(n11976) );
  INV_X1 U14440 ( .A(n12283), .ZN(n11932) );
  XNOR2_X1 U14441 ( .A(n14433), .B(n14415), .ZN(n11933) );
  NAND2_X1 U14442 ( .A1(n11933), .A2(n14645), .ZN(n11975) );
  INV_X1 U14443 ( .A(n14250), .ZN(n11940) );
  INV_X1 U14444 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14445 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  NAND2_X1 U14446 ( .A1(n12096), .A2(n11936), .ZN(n14954) );
  AOI22_X1 U14447 ( .A1(n10631), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n12156), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U14448 ( .A1(n6678), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11937) );
  OAI211_X1 U14449 ( .C1(n14954), .C2(n10983), .A(n11938), .B(n11937), .ZN(
        n14959) );
  INV_X1 U14450 ( .A(n14959), .ZN(n14738) );
  OR2_X1 U14451 ( .A1(n15102), .A2(n14738), .ZN(n11939) );
  OAI21_X1 U14452 ( .B1(n15097), .B2(n12667), .A(n11939), .ZN(n11973) );
  AOI21_X1 U14453 ( .B1(n15099), .B2(n11940), .A(n11973), .ZN(n11941) );
  OAI211_X1 U14454 ( .C1(n11216), .C2(n11976), .A(n11975), .B(n11941), .ZN(
        n11942) );
  NAND2_X1 U14455 ( .A1(n11942), .A2(n15103), .ZN(n11944) );
  AOI22_X1 U14456 ( .A1(n14416), .A2(n15074), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n15112), .ZN(n11943) );
  OAI211_X1 U14457 ( .C1(n11945), .C2(n14623), .A(n11944), .B(n11943), .ZN(
        P1_U3278) );
  XNOR2_X1 U14458 ( .A(n6709), .B(n12278), .ZN(n11946) );
  OAI222_X1 U14459 ( .A1(n15102), .A2(n14943), .B1(n15097), .B2(n14930), .C1(
        n11946), .C2(n15145), .ZN(n15009) );
  AOI21_X1 U14460 ( .B1(n11947), .B2(n15099), .A(n15009), .ZN(n11955) );
  INV_X1 U14461 ( .A(n11948), .ZN(n11949) );
  AOI21_X1 U14462 ( .B1(n12290), .B2(n11950), .A(n11949), .ZN(n15011) );
  OAI211_X1 U14463 ( .C1(n7312), .C2(n6824), .A(n15077), .B(n11951), .ZN(
        n15008) );
  AOI22_X1 U14464 ( .A1(n14938), .A2(n15074), .B1(n15112), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n11952) );
  OAI21_X1 U14465 ( .B1(n15008), .B2(n14577), .A(n11952), .ZN(n11953) );
  AOI21_X1 U14466 ( .B1(n15011), .B2(n14654), .A(n11953), .ZN(n11954) );
  OAI21_X1 U14467 ( .B1(n11955), .B2(n15112), .A(n11954), .ZN(P1_U3279) );
  AOI22_X1 U14468 ( .A1(n12767), .A2(n14263), .B1(n12769), .B2(n12255), .ZN(
        n12627) );
  NAND2_X1 U14469 ( .A1(n12255), .A2(n12770), .ZN(n11957) );
  NAND2_X1 U14470 ( .A1(n12769), .A2(n14263), .ZN(n11956) );
  NAND2_X1 U14471 ( .A1(n11957), .A2(n11956), .ZN(n11958) );
  XNOR2_X1 U14472 ( .A(n11958), .B(n12756), .ZN(n12626) );
  XOR2_X1 U14473 ( .A(n12627), .B(n12626), .Z(n11966) );
  INV_X1 U14474 ( .A(n11959), .ZN(n11960) );
  INV_X1 U14475 ( .A(n12630), .ZN(n11964) );
  AOI21_X1 U14476 ( .B1(n11966), .B2(n11965), .A(n11964), .ZN(n11972) );
  AOI22_X1 U14477 ( .A1(n14214), .A2(n11967), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11968) );
  OAI21_X1 U14478 ( .B1(n14985), .B2(n11969), .A(n11968), .ZN(n11970) );
  AOI21_X1 U14479 ( .B1(n14981), .B2(n12255), .A(n11970), .ZN(n11971) );
  OAI21_X1 U14480 ( .B1(n11972), .B2(n14976), .A(n11971), .ZN(P1_U3221) );
  AOI21_X1 U14481 ( .B1(n14416), .B2(n15156), .A(n11973), .ZN(n11974) );
  OAI211_X1 U14482 ( .C1(n15159), .C2(n11976), .A(n11975), .B(n11974), .ZN(
        n11977) );
  AOI21_X1 U14483 ( .B1(n11978), .B2(n15208), .A(n11977), .ZN(n11982) );
  NAND2_X1 U14484 ( .A1(n15223), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11979) );
  OAI21_X1 U14485 ( .B1(n11982), .B2(n15223), .A(n11979), .ZN(P1_U3543) );
  INV_X1 U14486 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11980) );
  OR2_X1 U14487 ( .A1(n15212), .A2(n11980), .ZN(n11981) );
  OAI21_X1 U14488 ( .B1(n11982), .B2(n15210), .A(n11981), .ZN(P1_U3504) );
  XNOR2_X1 U14489 ( .A(n11983), .B(n6913), .ZN(n11984) );
  NAND2_X1 U14490 ( .A1(n11984), .A2(n14882), .ZN(n11988) );
  NAND2_X1 U14491 ( .A1(n13610), .A2(n13659), .ZN(n11986) );
  NAND2_X1 U14492 ( .A1(n13551), .A2(n13661), .ZN(n11985) );
  NAND2_X1 U14493 ( .A1(n11986), .A2(n11985), .ZN(n13640) );
  INV_X1 U14494 ( .A(n13640), .ZN(n11987) );
  NAND2_X1 U14495 ( .A1(n11988), .A2(n11987), .ZN(n14900) );
  AOI21_X1 U14496 ( .B1(n13636), .B2(n15316), .A(n14900), .ZN(n11997) );
  NAND2_X1 U14497 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  NAND2_X1 U14498 ( .A1(n11992), .A2(n11991), .ZN(n14896) );
  OAI211_X1 U14499 ( .C1(n14890), .C2(n14899), .A(n9576), .B(n13952), .ZN(
        n14897) );
  AOI22_X1 U14500 ( .A1(n11993), .A2(n15314), .B1(n6674), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n11994) );
  OAI21_X1 U14501 ( .B1(n14897), .B2(n13961), .A(n11994), .ZN(n11995) );
  AOI21_X1 U14502 ( .B1(n14896), .B2(n15320), .A(n11995), .ZN(n11996) );
  OAI21_X1 U14503 ( .B1(n11997), .B2(n6674), .A(n11996), .ZN(P2_U3250) );
  INV_X1 U14504 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11998) );
  OR2_X1 U14505 ( .A1(n12162), .A2(n11998), .ZN(n11999) );
  NAND2_X1 U14506 ( .A1(n6678), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U14507 ( .A1(n6680), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U14508 ( .A1(n12156), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12000) );
  AND3_X1 U14509 ( .A1(n12002), .A2(n12001), .A3(n12000), .ZN(n12176) );
  INV_X1 U14510 ( .A(n12176), .ZN(n14406) );
  XNOR2_X1 U14511 ( .A(n14407), .B(n14406), .ZN(n12203) );
  NAND2_X1 U14512 ( .A1(n14769), .A2(n12161), .ZN(n12004) );
  OR2_X1 U14513 ( .A1(n12162), .A2(n14770), .ZN(n12003) );
  NAND2_X1 U14514 ( .A1(n12156), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U14515 ( .A1(n6678), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12010) );
  INV_X1 U14516 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U14517 ( .A1(n12121), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12123) );
  INV_X1 U14518 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12078) );
  INV_X1 U14519 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U14520 ( .A1(n12066), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12055) );
  INV_X1 U14521 ( .A(n12055), .ZN(n12005) );
  NAND2_X1 U14522 ( .A1(n12005), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12149) );
  NAND2_X1 U14523 ( .A1(n12054), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U14524 ( .A1(n12148), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12032) );
  INV_X1 U14525 ( .A(n12032), .ZN(n12137) );
  NAND2_X1 U14526 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n12137), .ZN(n12034) );
  INV_X1 U14527 ( .A(n12034), .ZN(n12006) );
  NAND2_X1 U14528 ( .A1(n12006), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12024) );
  INV_X1 U14529 ( .A(n12024), .ZN(n12007) );
  NAND2_X1 U14530 ( .A1(n12007), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12167) );
  XNOR2_X1 U14531 ( .A(n12167), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U14532 ( .A1(n12056), .A2(n14473), .ZN(n12009) );
  NAND2_X1 U14533 ( .A1(n10631), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12008) );
  NAND4_X1 U14534 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n14447) );
  XNOR2_X1 U14535 ( .A(n14477), .B(n14488), .ZN(n14466) );
  NAND2_X1 U14536 ( .A1(n14102), .A2(n12161), .ZN(n12013) );
  OR2_X1 U14537 ( .A1(n12162), .A2(n14773), .ZN(n12012) );
  NAND2_X1 U14538 ( .A1(n12156), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U14539 ( .A1(n6678), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12018) );
  INV_X1 U14540 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U14541 ( .A1(n12024), .A2(n12014), .ZN(n12015) );
  NAND2_X1 U14542 ( .A1(n12056), .A2(n14496), .ZN(n12017) );
  NAND2_X1 U14543 ( .A1(n10631), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U14544 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n14505) );
  INV_X1 U14545 ( .A(n14505), .ZN(n14468) );
  XNOR2_X1 U14546 ( .A(n14497), .B(n14468), .ZN(n14486) );
  NAND2_X1 U14547 ( .A1(n14105), .A2(n12161), .ZN(n12021) );
  INV_X1 U14548 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14778) );
  OR2_X1 U14549 ( .A1(n12162), .A2(n14778), .ZN(n12020) );
  NAND2_X1 U14550 ( .A1(n12156), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U14551 ( .A1(n6678), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12027) );
  INV_X1 U14552 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n12022) );
  NAND2_X1 U14553 ( .A1(n12034), .A2(n12022), .ZN(n12023) );
  AND2_X1 U14554 ( .A1(n12024), .A2(n12023), .ZN(n14510) );
  NAND2_X1 U14555 ( .A1(n12056), .A2(n14510), .ZN(n12026) );
  NAND2_X1 U14556 ( .A1(n6680), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U14557 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n14524) );
  INV_X1 U14558 ( .A(n14524), .ZN(n14489) );
  NAND2_X1 U14559 ( .A1(n14507), .A2(n14489), .ZN(n14446) );
  OR2_X1 U14560 ( .A1(n14507), .A2(n14489), .ZN(n12029) );
  NAND2_X1 U14561 ( .A1(n14446), .A2(n12029), .ZN(n14445) );
  NAND2_X1 U14562 ( .A1(n12624), .A2(n12161), .ZN(n12031) );
  OR2_X1 U14563 ( .A1(n12162), .A2(n12625), .ZN(n12030) );
  NAND2_X1 U14564 ( .A1(n12156), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12039) );
  NAND2_X1 U14565 ( .A1(n6678), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12038) );
  INV_X1 U14566 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U14567 ( .A1(n12033), .A2(n12032), .ZN(n12035) );
  AND2_X1 U14568 ( .A1(n12035), .A2(n12034), .ZN(n14531) );
  NAND2_X1 U14569 ( .A1(n12056), .A2(n14531), .ZN(n12037) );
  NAND2_X1 U14570 ( .A1(n10631), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U14571 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n14504) );
  INV_X1 U14572 ( .A(n14504), .ZN(n14538) );
  NAND2_X1 U14573 ( .A1(n14518), .A2(n14538), .ZN(n14444) );
  OR2_X1 U14574 ( .A1(n14518), .A2(n14538), .ZN(n12040) );
  NAND2_X1 U14575 ( .A1(n14444), .A2(n12040), .ZN(n14529) );
  NAND2_X1 U14576 ( .A1(n12041), .A2(n12161), .ZN(n12044) );
  OR2_X1 U14577 ( .A1(n12162), .A2(n12042), .ZN(n12043) );
  OR2_X1 U14578 ( .A1(n12066), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U14579 ( .A1(n12045), .A2(n12055), .ZN(n14587) );
  OR2_X1 U14580 ( .A1(n14587), .A2(n10983), .ZN(n12051) );
  INV_X1 U14581 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U14582 ( .A1(n12156), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U14583 ( .A1(n10631), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12046) );
  OAI211_X1 U14584 ( .C1(n6669), .C2(n12048), .A(n12047), .B(n12046), .ZN(
        n12049) );
  INV_X1 U14585 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U14586 ( .A1(n12051), .A2(n12050), .ZN(n14565) );
  INV_X1 U14587 ( .A(n14565), .ZN(n14225) );
  XNOR2_X1 U14588 ( .A(n14709), .B(n14225), .ZN(n14581) );
  NAND2_X1 U14589 ( .A1(n6678), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U14590 ( .A1(n10631), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12059) );
  INV_X1 U14591 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14224) );
  AOI21_X1 U14592 ( .B1(n14224), .B2(n12055), .A(n12054), .ZN(n14573) );
  NAND2_X1 U14593 ( .A1(n12056), .A2(n14573), .ZN(n12058) );
  NAND2_X1 U14594 ( .A1(n12156), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n12057) );
  XNOR2_X1 U14595 ( .A(n14572), .B(n14585), .ZN(n14569) );
  NAND2_X1 U14596 ( .A1(n12061), .A2(n12161), .ZN(n12064) );
  OR2_X1 U14597 ( .A1(n12162), .A2(n12062), .ZN(n12063) );
  AND2_X1 U14598 ( .A1(n12080), .A2(n14202), .ZN(n12065) );
  OR2_X1 U14599 ( .A1(n12066), .A2(n12065), .ZN(n14602) );
  INV_X1 U14600 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n12069) );
  NAND2_X1 U14601 ( .A1(n12156), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U14602 ( .A1(n10631), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12067) );
  OAI211_X1 U14603 ( .C1(n6669), .C2(n12069), .A(n12068), .B(n12067), .ZN(
        n12070) );
  INV_X1 U14604 ( .A(n12070), .ZN(n12071) );
  OAI21_X1 U14605 ( .B1(n14602), .B2(n10983), .A(n12071), .ZN(n14584) );
  INV_X1 U14606 ( .A(n14584), .ZN(n14612) );
  OR2_X1 U14607 ( .A1(n14714), .A2(n14612), .ZN(n14437) );
  NAND2_X1 U14608 ( .A1(n14714), .A2(n14612), .ZN(n12072) );
  NAND2_X1 U14609 ( .A1(n12073), .A2(n12161), .ZN(n12077) );
  OAI22_X1 U14610 ( .A1(n14527), .A2(n12116), .B1(n12162), .B2(n12074), .ZN(
        n12075) );
  INV_X1 U14611 ( .A(n12075), .ZN(n12076) );
  NAND2_X1 U14612 ( .A1(n12123), .A2(n12078), .ZN(n12079) );
  NAND2_X1 U14613 ( .A1(n12080), .A2(n12079), .ZN(n14616) );
  OR2_X1 U14614 ( .A1(n14616), .A2(n10983), .ZN(n12085) );
  INV_X1 U14615 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U14616 ( .A1(n12156), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U14617 ( .A1(n10631), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12081) );
  OAI211_X1 U14618 ( .C1(n6669), .C2(n14387), .A(n12082), .B(n12081), .ZN(
        n12083) );
  INV_X1 U14619 ( .A(n12083), .ZN(n12084) );
  NAND2_X1 U14620 ( .A1(n12085), .A2(n12084), .ZN(n14627) );
  INV_X1 U14621 ( .A(n14627), .ZN(n14233) );
  OR2_X1 U14622 ( .A1(n14721), .A2(n14233), .ZN(n12304) );
  NAND2_X1 U14623 ( .A1(n14721), .A2(n14233), .ZN(n14436) );
  NAND2_X1 U14624 ( .A1(n12304), .A2(n14436), .ZN(n14422) );
  NAND2_X1 U14625 ( .A1(n12086), .A2(n12161), .ZN(n12089) );
  AOI22_X1 U14626 ( .A1(n12092), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12091), 
        .B2(n12087), .ZN(n12088) );
  XNOR2_X1 U14627 ( .A(n14951), .B(n14738), .ZN(n14652) );
  NAND2_X1 U14628 ( .A1(n12090), .A2(n12161), .ZN(n12094) );
  AOI22_X1 U14629 ( .A1(n12092), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12091), 
        .B2(n14375), .ZN(n12093) );
  AND2_X1 U14630 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  OR2_X1 U14631 ( .A1(n12097), .A2(n12121), .ZN(n14988) );
  AOI22_X1 U14632 ( .A1(n6678), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n10631), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n12099) );
  NAND2_X1 U14633 ( .A1(n12156), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12098) );
  OAI211_X1 U14634 ( .C1(n14988), .C2(n10983), .A(n12099), .B(n12098), .ZN(
        n14644) );
  NOR2_X1 U14635 ( .A1(n14991), .A2(n14644), .ZN(n14419) );
  NAND2_X1 U14636 ( .A1(n14991), .A2(n14644), .ZN(n14420) );
  NAND2_X1 U14637 ( .A1(n7566), .A2(n14420), .ZN(n14733) );
  INV_X1 U14638 ( .A(n12231), .ZN(n12103) );
  NAND4_X1 U14639 ( .A1(n15092), .A2(n12224), .A3(n12220), .A4(n15144), .ZN(
        n12102) );
  NOR4_X1 U14640 ( .A1(n12103), .A2(n15068), .A3(n12102), .A4(n12101), .ZN(
        n12107) );
  NAND4_X1 U14641 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12108) );
  NOR4_X1 U14642 ( .A1(n12111), .A2(n12110), .A3(n12109), .A4(n12108), .ZN(
        n12113) );
  NAND3_X1 U14643 ( .A1(n14733), .A2(n12113), .A3(n12112), .ZN(n12114) );
  NOR4_X1 U14644 ( .A1(n14652), .A2(n14415), .A3(n12114), .A4(n12278), .ZN(
        n12132) );
  NAND2_X1 U14645 ( .A1(n12115), .A2(n12161), .ZN(n12120) );
  OAI22_X1 U14646 ( .A1(n12162), .A2(n12117), .B1(n14379), .B2(n12116), .ZN(
        n12118) );
  INV_X1 U14647 ( .A(n12118), .ZN(n12119) );
  OR2_X1 U14648 ( .A1(n12121), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12122) );
  AND2_X1 U14649 ( .A1(n12123), .A2(n12122), .ZN(n14633) );
  NAND2_X1 U14650 ( .A1(n14633), .A2(n12124), .ZN(n12131) );
  INV_X1 U14651 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U14652 ( .A1(n12156), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U14653 ( .A1(n10631), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n12126) );
  OAI211_X1 U14654 ( .C1(n6669), .C2(n12128), .A(n12127), .B(n12126), .ZN(
        n12129) );
  INV_X1 U14655 ( .A(n12129), .ZN(n12130) );
  NAND2_X1 U14656 ( .A1(n12131), .A2(n12130), .ZN(n14957) );
  INV_X1 U14657 ( .A(n14957), .ZN(n14739) );
  XNOR2_X1 U14658 ( .A(n14727), .B(n14739), .ZN(n12299) );
  NAND4_X1 U14659 ( .A1(n14596), .A2(n14609), .A3(n12132), .A4(n14625), .ZN(
        n12133) );
  NOR4_X1 U14660 ( .A1(n14529), .A2(n14581), .A3(n14569), .A4(n12133), .ZN(
        n12154) );
  NAND2_X1 U14661 ( .A1(n12134), .A2(n12161), .ZN(n12136) );
  OR2_X1 U14662 ( .A1(n12162), .A2(n12375), .ZN(n12135) );
  NAND2_X1 U14663 ( .A1(n12156), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U14664 ( .A1(n6678), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12142) );
  INV_X1 U14665 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n12139) );
  AOI21_X1 U14666 ( .B1(n12139), .B2(n12138), .A(n12137), .ZN(n14548) );
  NAND2_X1 U14667 ( .A1(n12124), .A2(n14548), .ZN(n12141) );
  NAND2_X1 U14668 ( .A1(n10631), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U14669 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n14523) );
  XNOR2_X1 U14670 ( .A(n14549), .B(n14523), .ZN(n14442) );
  NAND2_X1 U14671 ( .A1(n12144), .A2(n12161), .ZN(n12147) );
  OR2_X1 U14672 ( .A1(n12162), .A2(n12145), .ZN(n12146) );
  NAND2_X1 U14673 ( .A1(n12156), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U14674 ( .A1(n6678), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12152) );
  INV_X1 U14675 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14127) );
  AOI21_X1 U14676 ( .B1(n14127), .B2(n12149), .A(n12148), .ZN(n14558) );
  NAND2_X1 U14677 ( .A1(n12124), .A2(n14558), .ZN(n12151) );
  NAND2_X1 U14678 ( .A1(n10631), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U14679 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n14566) );
  XNOR2_X1 U14680 ( .A(n14562), .B(n14566), .ZN(n14441) );
  NAND3_X1 U14681 ( .A1(n12154), .A2(n14442), .A3(n14441), .ZN(n12155) );
  NOR4_X1 U14682 ( .A1(n14466), .A2(n14486), .A3(n14445), .A4(n12155), .ZN(
        n12173) );
  NAND2_X1 U14683 ( .A1(n6678), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12159) );
  NAND2_X1 U14684 ( .A1(n10631), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U14685 ( .A1(n12156), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12157) );
  NAND3_X1 U14686 ( .A1(n12159), .A2(n12158), .A3(n12157), .ZN(n14454) );
  INV_X1 U14687 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12403) );
  NOR2_X1 U14688 ( .A1(n12162), .A2(n12403), .ZN(n12160) );
  XOR2_X1 U14689 ( .A(n14454), .B(n14660), .Z(n12172) );
  NAND2_X1 U14690 ( .A1(n14095), .A2(n12161), .ZN(n12164) );
  INV_X1 U14691 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14766) );
  OR2_X1 U14692 ( .A1(n12162), .A2(n14766), .ZN(n12163) );
  INV_X1 U14693 ( .A(n14661), .ZN(n14462) );
  NAND2_X1 U14694 ( .A1(n12156), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U14695 ( .A1(n6678), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12170) );
  INV_X1 U14696 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12166) );
  NOR2_X1 U14697 ( .A1(n12167), .A2(n12166), .ZN(n14456) );
  NAND2_X1 U14698 ( .A1(n12056), .A2(n14456), .ZN(n12169) );
  NAND2_X1 U14699 ( .A1(n10631), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12168) );
  XNOR2_X1 U14700 ( .A(n14462), .B(n14469), .ZN(n14448) );
  NAND4_X1 U14701 ( .A1(n12203), .A2(n12173), .A3(n12172), .A4(n14448), .ZN(
        n12174) );
  XNOR2_X1 U14702 ( .A(n12174), .B(n14527), .ZN(n12212) );
  INV_X1 U14703 ( .A(n12175), .ZN(n12211) );
  NAND2_X1 U14704 ( .A1(n12177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U14705 ( .A1(n14760), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n12178) );
  AND2_X1 U14706 ( .A1(n12179), .A2(n12178), .ZN(n12184) );
  INV_X1 U14707 ( .A(n12184), .ZN(n12183) );
  NAND2_X1 U14708 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n12180) );
  OAI211_X1 U14709 ( .C1(P1_IR_REG_22__SCAN_IN), .C2(P1_IR_REG_20__SCAN_IN), 
        .A(P1_IR_REG_31__SCAN_IN), .B(n12180), .ZN(n12181) );
  NOR2_X1 U14710 ( .A1(n10567), .A2(n12181), .ZN(n12182) );
  AOI21_X1 U14711 ( .B1(n12186), .B2(n12183), .A(n12182), .ZN(n12188) );
  NAND2_X1 U14712 ( .A1(n10567), .A2(n12184), .ZN(n12185) );
  NAND2_X1 U14713 ( .A1(n12188), .A2(n12187), .ZN(n12193) );
  OAI21_X1 U14714 ( .B1(n12190), .B2(n10894), .A(n15084), .ZN(n12208) );
  AND2_X1 U14715 ( .A1(n12208), .A2(n12211), .ZN(n12204) );
  NAND2_X1 U14716 ( .A1(n12206), .A2(n12204), .ZN(n12361) );
  INV_X1 U14717 ( .A(n12361), .ZN(n12202) );
  OAI21_X1 U14718 ( .B1(n12191), .B2(n14406), .A(n14454), .ZN(n12192) );
  MUX2_X1 U14719 ( .A(n12192), .B(n14660), .S(n12350), .Z(n12201) );
  INV_X1 U14720 ( .A(n14454), .ZN(n12198) );
  AOI22_X1 U14721 ( .A1(n12350), .A2(n14406), .B1(n12194), .B2(n12193), .ZN(
        n12197) );
  INV_X1 U14722 ( .A(n14660), .ZN(n12195) );
  NAND2_X1 U14723 ( .A1(n12195), .A2(n6682), .ZN(n12196) );
  OAI21_X1 U14724 ( .B1(n12198), .B2(n12197), .A(n12196), .ZN(n12200) );
  NOR2_X1 U14725 ( .A1(n12201), .A2(n12200), .ZN(n12364) );
  INV_X1 U14726 ( .A(n12208), .ZN(n12199) );
  AND2_X1 U14727 ( .A1(n12203), .A2(n12199), .ZN(n12363) );
  AND2_X1 U14728 ( .A1(n12201), .A2(n12200), .ZN(n12362) );
  AOI22_X1 U14729 ( .A1(n12202), .A2(n12364), .B1(n12363), .B2(n12362), .ZN(
        n12210) );
  INV_X1 U14730 ( .A(n12203), .ZN(n12205) );
  NAND2_X1 U14731 ( .A1(n12205), .A2(n12204), .ZN(n12207) );
  MUX2_X1 U14732 ( .A(n12208), .B(n12207), .S(n12206), .Z(n12209) );
  AOI21_X1 U14733 ( .B1(n15096), .B2(n12214), .A(n12213), .ZN(n12217) );
  NOR2_X1 U14734 ( .A1(n15096), .A2(n12214), .ZN(n12216) );
  NAND2_X1 U14735 ( .A1(n12350), .A2(n15101), .ZN(n12222) );
  NAND2_X1 U14736 ( .A1(n6682), .A2(n14269), .ZN(n12221) );
  MUX2_X1 U14737 ( .A(n12222), .B(n12221), .S(n15165), .Z(n12223) );
  NAND2_X1 U14738 ( .A1(n12350), .A2(n14268), .ZN(n12229) );
  NAND2_X1 U14739 ( .A1(n6682), .A2(n12226), .ZN(n12228) );
  MUX2_X1 U14740 ( .A(n12229), .B(n12228), .S(n12227), .Z(n12230) );
  NAND3_X1 U14741 ( .A1(n12232), .A2(n12231), .A3(n12230), .ZN(n12239) );
  OAI21_X1 U14742 ( .B1(n6682), .B2(n14267), .A(n12233), .ZN(n12237) );
  OAI21_X1 U14743 ( .B1(n12350), .B2(n12235), .A(n12234), .ZN(n12236) );
  NAND2_X1 U14744 ( .A1(n12237), .A2(n12236), .ZN(n12238) );
  NAND2_X1 U14745 ( .A1(n12239), .A2(n12238), .ZN(n12245) );
  MUX2_X1 U14746 ( .A(n15174), .B(n12241), .S(n12350), .Z(n12244) );
  MUX2_X1 U14747 ( .A(n14266), .B(n12242), .S(n12350), .Z(n12243) );
  NAND2_X1 U14748 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  NAND2_X1 U14749 ( .A1(n12247), .A2(n12246), .ZN(n12249) );
  MUX2_X1 U14750 ( .A(n14265), .B(n15075), .S(n12350), .Z(n12250) );
  MUX2_X1 U14751 ( .A(n14264), .B(n12251), .S(n6682), .Z(n12253) );
  MUX2_X1 U14752 ( .A(n14264), .B(n12251), .S(n12350), .Z(n12252) );
  INV_X1 U14753 ( .A(n12253), .ZN(n12254) );
  MUX2_X1 U14754 ( .A(n14263), .B(n12255), .S(n12350), .Z(n12259) );
  NAND2_X1 U14755 ( .A1(n12258), .A2(n12259), .ZN(n12257) );
  INV_X1 U14756 ( .A(n12258), .ZN(n12261) );
  INV_X1 U14757 ( .A(n12259), .ZN(n12260) );
  NAND2_X1 U14758 ( .A1(n12261), .A2(n12260), .ZN(n12262) );
  MUX2_X1 U14759 ( .A(n14262), .B(n14192), .S(n6682), .Z(n12264) );
  MUX2_X1 U14760 ( .A(n14262), .B(n14192), .S(n12350), .Z(n12263) );
  MUX2_X1 U14761 ( .A(n14261), .B(n12638), .S(n12350), .Z(n12266) );
  INV_X1 U14762 ( .A(n12266), .ZN(n12267) );
  MUX2_X1 U14763 ( .A(n14260), .B(n15013), .S(n6682), .Z(n12271) );
  NAND2_X1 U14764 ( .A1(n12270), .A2(n12271), .ZN(n12269) );
  MUX2_X1 U14765 ( .A(n14260), .B(n15013), .S(n12350), .Z(n12268) );
  NAND2_X1 U14766 ( .A1(n12269), .A2(n12268), .ZN(n12275) );
  INV_X1 U14767 ( .A(n12271), .ZN(n12272) );
  NAND2_X1 U14768 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  MUX2_X1 U14769 ( .A(n14259), .B(n14172), .S(n12350), .Z(n12277) );
  MUX2_X1 U14770 ( .A(n14258), .B(n12662), .S(n6682), .Z(n12285) );
  OR2_X1 U14771 ( .A1(n12278), .A2(n12285), .ZN(n12281) );
  AND2_X1 U14772 ( .A1(n14431), .A2(n12279), .ZN(n12280) );
  OAI22_X1 U14773 ( .A1(n12286), .A2(n12281), .B1(n12350), .B2(n12280), .ZN(
        n12282) );
  NAND2_X1 U14774 ( .A1(n12282), .A2(n12287), .ZN(n12294) );
  NAND2_X1 U14775 ( .A1(n12287), .A2(n12283), .ZN(n12284) );
  NAND2_X1 U14776 ( .A1(n12284), .A2(n12350), .ZN(n12293) );
  NAND2_X1 U14777 ( .A1(n12286), .A2(n12285), .ZN(n12291) );
  AND2_X1 U14778 ( .A1(n12287), .A2(n14258), .ZN(n12288) );
  MUX2_X1 U14779 ( .A(n12662), .B(n12288), .S(n6682), .Z(n12289) );
  NAND3_X1 U14780 ( .A1(n12291), .A2(n12290), .A3(n12289), .ZN(n12292) );
  OR2_X1 U14781 ( .A1(n14431), .A2(n6682), .ZN(n12295) );
  MUX2_X1 U14782 ( .A(n14959), .B(n14951), .S(n6682), .Z(n12297) );
  MUX2_X1 U14783 ( .A(n14959), .B(n14951), .S(n12350), .Z(n12296) );
  NOR2_X1 U14784 ( .A1(n14422), .A2(n12299), .ZN(n12300) );
  MUX2_X1 U14785 ( .A(n14644), .B(n14991), .S(n12350), .Z(n12301) );
  OR2_X1 U14786 ( .A1(n14727), .A2(n14739), .ZN(n14435) );
  NAND3_X1 U14787 ( .A1(n14727), .A2(n14739), .A3(n12350), .ZN(n12302) );
  OAI21_X1 U14788 ( .B1(n14435), .B2(n12350), .A(n12302), .ZN(n12303) );
  INV_X1 U14789 ( .A(n12303), .ZN(n12306) );
  MUX2_X1 U14790 ( .A(n14436), .B(n12304), .S(n6682), .Z(n12305) );
  OAI21_X1 U14791 ( .B1(n14422), .B2(n12306), .A(n12305), .ZN(n12307) );
  INV_X1 U14792 ( .A(n12307), .ZN(n12308) );
  INV_X1 U14793 ( .A(n14714), .ZN(n14208) );
  MUX2_X1 U14794 ( .A(n14612), .B(n14208), .S(n6682), .Z(n12310) );
  MUX2_X1 U14795 ( .A(n14584), .B(n14714), .S(n12350), .Z(n12309) );
  NAND2_X1 U14796 ( .A1(n12311), .A2(n12310), .ZN(n12312) );
  MUX2_X1 U14797 ( .A(n14565), .B(n14709), .S(n12350), .Z(n12316) );
  NAND2_X1 U14798 ( .A1(n12315), .A2(n12316), .ZN(n12314) );
  NAND2_X1 U14799 ( .A1(n12314), .A2(n12313), .ZN(n12320) );
  INV_X1 U14800 ( .A(n12315), .ZN(n12318) );
  INV_X1 U14801 ( .A(n12316), .ZN(n12317) );
  NAND2_X1 U14802 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  NAND2_X1 U14803 ( .A1(n12320), .A2(n12319), .ZN(n12323) );
  INV_X1 U14804 ( .A(n14572), .ZN(n14574) );
  MUX2_X1 U14805 ( .A(n14440), .B(n14572), .S(n12350), .Z(n12321) );
  AOI21_X1 U14806 ( .B1(n12323), .B2(n12322), .A(n12321), .ZN(n12325) );
  NOR2_X1 U14807 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  MUX2_X1 U14808 ( .A(n14566), .B(n14562), .S(n12350), .Z(n12327) );
  MUX2_X1 U14809 ( .A(n14566), .B(n14562), .S(n6682), .Z(n12326) );
  MUX2_X1 U14810 ( .A(n14523), .B(n14549), .S(n6682), .Z(n12331) );
  NAND2_X1 U14811 ( .A1(n12330), .A2(n12331), .ZN(n12329) );
  MUX2_X1 U14812 ( .A(n14523), .B(n14549), .S(n12350), .Z(n12328) );
  NAND2_X1 U14813 ( .A1(n12329), .A2(n12328), .ZN(n12335) );
  INV_X1 U14814 ( .A(n12330), .ZN(n12333) );
  INV_X1 U14815 ( .A(n12331), .ZN(n12332) );
  NAND2_X1 U14816 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  NAND2_X1 U14817 ( .A1(n12335), .A2(n12334), .ZN(n12337) );
  MUX2_X1 U14818 ( .A(n14504), .B(n14518), .S(n12350), .Z(n12338) );
  MUX2_X1 U14819 ( .A(n14524), .B(n14507), .S(n6682), .Z(n12340) );
  MUX2_X1 U14820 ( .A(n14524), .B(n14507), .S(n12350), .Z(n12339) );
  INV_X1 U14821 ( .A(n12340), .ZN(n12341) );
  MUX2_X1 U14822 ( .A(n14505), .B(n14497), .S(n12350), .Z(n12345) );
  NAND2_X1 U14823 ( .A1(n12344), .A2(n12345), .ZN(n12343) );
  NAND2_X1 U14824 ( .A1(n12343), .A2(n12342), .ZN(n12349) );
  INV_X1 U14825 ( .A(n12344), .ZN(n12347) );
  INV_X1 U14826 ( .A(n12345), .ZN(n12346) );
  NAND2_X1 U14827 ( .A1(n12347), .A2(n12346), .ZN(n12348) );
  NAND2_X1 U14828 ( .A1(n12349), .A2(n12348), .ZN(n12353) );
  MUX2_X1 U14829 ( .A(n14477), .B(n14447), .S(n12350), .Z(n12354) );
  NAND2_X1 U14830 ( .A1(n12353), .A2(n12354), .ZN(n12352) );
  MUX2_X1 U14831 ( .A(n14447), .B(n14477), .S(n12350), .Z(n12351) );
  NAND2_X1 U14832 ( .A1(n12352), .A2(n12351), .ZN(n12358) );
  INV_X1 U14833 ( .A(n12353), .ZN(n12356) );
  INV_X1 U14834 ( .A(n12354), .ZN(n12355) );
  NAND2_X1 U14835 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  INV_X1 U14836 ( .A(n14469), .ZN(n14256) );
  MUX2_X1 U14837 ( .A(n14256), .B(n14661), .S(n12350), .Z(n12360) );
  MUX2_X1 U14838 ( .A(n14256), .B(n14661), .S(n6682), .Z(n12359) );
  INV_X1 U14839 ( .A(n12363), .ZN(n12365) );
  NOR2_X1 U14840 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  NOR2_X1 U14841 ( .A1(n14776), .A2(P1_U3086), .ZN(n12370) );
  NAND3_X1 U14842 ( .A1(n12371), .A2(n14641), .A3(n12370), .ZN(n12372) );
  OAI211_X1 U14843 ( .C1(n15149), .C2(n12374), .A(n12372), .B(P1_B_REG_SCAN_IN), .ZN(n12373) );
  OAI222_X1 U14844 ( .A1(P1_U3086), .A2(n10210), .B1(n14775), .B2(n12376), 
        .C1(n12375), .C2(n14772), .ZN(P1_U3331) );
  INV_X1 U14845 ( .A(n12377), .ZN(n14094) );
  OAI222_X1 U14846 ( .A1(n14775), .A2(n14094), .B1(n12378), .B2(P1_U3086), 
        .C1(n12403), .C2(n14777), .ZN(P1_U3325) );
  INV_X1 U14847 ( .A(n12379), .ZN(n12380) );
  OAI222_X1 U14848 ( .A1(n13441), .A2(n12383), .B1(P3_U3151), .B2(n12382), 
        .C1(n12381), .C2(n12380), .ZN(P3_U3267) );
  NAND2_X1 U14849 ( .A1(n15307), .A2(n15235), .ZN(n12386) );
  INV_X1 U14850 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U14851 ( .A1(n15265), .A2(n12384), .ZN(n12385) );
  AND3_X1 U14852 ( .A1(n12386), .A2(n15272), .A3(n12385), .ZN(n12388) );
  AOI22_X1 U14853 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15307), .B1(n15265), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n12387) );
  MUX2_X1 U14854 ( .A(n12388), .B(n12387), .S(n15236), .Z(n12390) );
  AOI22_X1 U14855 ( .A1(n15289), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n12389) );
  NAND2_X1 U14856 ( .A1(n12390), .A2(n12389), .ZN(P2_U3214) );
  INV_X1 U14857 ( .A(n12391), .ZN(n12392) );
  AOI22_X1 U14858 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n12393), .B1(n13641), 
        .B2(n12392), .ZN(n12399) );
  NOR2_X1 U14859 ( .A1(n12395), .A2(n12394), .ZN(n12397) );
  OAI21_X1 U14860 ( .B1(n12397), .B2(n12396), .A(n13632), .ZN(n12398) );
  OAI211_X1 U14861 ( .C1(n13644), .C2(n12400), .A(n12399), .B(n12398), .ZN(
        P2_U3204) );
  NAND2_X1 U14862 ( .A1(n14091), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12405) );
  NAND2_X1 U14863 ( .A1(n12403), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12404) );
  AND2_X1 U14864 ( .A1(n12405), .A2(n12404), .ZN(n12409) );
  NAND2_X1 U14865 ( .A1(n12408), .A2(n12409), .ZN(n12413) );
  NAND2_X1 U14866 ( .A1(n12413), .A2(n12405), .ZN(n12407) );
  XOR2_X1 U14867 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .Z(n12406) );
  XNOR2_X1 U14868 ( .A(n12407), .B(n12406), .ZN(n13435) );
  INV_X1 U14869 ( .A(SI_31_), .ZN(n13431) );
  INV_X1 U14870 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14871 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14872 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  NOR2_X1 U14873 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  INV_X1 U14874 ( .A(n12418), .ZN(n12947) );
  OAI22_X1 U14875 ( .A1(n13365), .A2(n13058), .B1(n13369), .B2(n12947), .ZN(
        n12443) );
  OAI21_X1 U14876 ( .B1(n13369), .B2(n12421), .A(n12588), .ZN(n12419) );
  INV_X1 U14877 ( .A(n13365), .ZN(n13297) );
  INV_X1 U14878 ( .A(n12424), .ZN(n12601) );
  INV_X1 U14879 ( .A(n13158), .ZN(n13163) );
  INV_X1 U14880 ( .A(n12425), .ZN(n12516) );
  OR2_X1 U14881 ( .A1(n12517), .A2(n12516), .ZN(n13283) );
  NOR2_X1 U14882 ( .A1(n15568), .A2(n15553), .ZN(n12426) );
  AND4_X1 U14883 ( .A1(n12428), .A2(n12427), .A3(n8370), .A4(n12426), .ZN(
        n12434) );
  NOR2_X1 U14884 ( .A1(n15611), .A2(n12429), .ZN(n12432) );
  NOR2_X1 U14885 ( .A1(n15540), .A2(n12463), .ZN(n12431) );
  INV_X1 U14886 ( .A(n12430), .ZN(n12495) );
  AND4_X1 U14887 ( .A1(n12432), .A2(n12431), .A3(n12495), .A4(n12488), .ZN(
        n12433) );
  NAND4_X1 U14888 ( .A1(n12434), .A2(n14859), .A3(n12433), .A4(n14845), .ZN(
        n12435) );
  NOR4_X1 U14889 ( .A1(n13258), .A2(n13276), .A3(n13283), .A4(n12435), .ZN(
        n12436) );
  AND4_X1 U14890 ( .A1(n13208), .A2(n13250), .A3(n13238), .A4(n12436), .ZN(
        n12437) );
  INV_X1 U14891 ( .A(n13190), .ZN(n13186) );
  NAND4_X1 U14892 ( .A1(n13177), .A2(n13220), .A3(n12437), .A4(n13186), .ZN(
        n12438) );
  OR4_X1 U14893 ( .A1(n13132), .A2(n8569), .A3(n13163), .A4(n12438), .ZN(
        n12439) );
  NOR2_X1 U14894 ( .A1(n13113), .A2(n12439), .ZN(n12440) );
  INV_X1 U14895 ( .A(n12443), .ZN(n12596) );
  INV_X1 U14896 ( .A(n12444), .ZN(n12445) );
  NAND2_X1 U14897 ( .A1(n12483), .A2(n12447), .ZN(n12448) );
  NAND2_X1 U14898 ( .A1(n12448), .A2(n12587), .ZN(n12477) );
  INV_X1 U14899 ( .A(n12477), .ZN(n12484) );
  OAI22_X1 U14900 ( .A1(n10413), .A2(n12449), .B1(n12587), .B2(n12450), .ZN(
        n12454) );
  NAND2_X1 U14901 ( .A1(n12450), .A2(n12451), .ZN(n12452) );
  AOI22_X1 U14902 ( .A1(n12452), .A2(n12606), .B1(n12451), .B2(n12578), .ZN(
        n12453) );
  OR2_X1 U14903 ( .A1(n12454), .A2(n12453), .ZN(n12456) );
  MUX2_X1 U14904 ( .A(n12587), .B(n12456), .S(n12455), .Z(n12464) );
  NAND2_X1 U14905 ( .A1(n12466), .A2(n12457), .ZN(n12460) );
  NAND2_X1 U14906 ( .A1(n12465), .A2(n12458), .ZN(n12459) );
  MUX2_X1 U14907 ( .A(n12460), .B(n12459), .S(n12587), .Z(n12461) );
  INV_X1 U14908 ( .A(n12461), .ZN(n12462) );
  OAI21_X1 U14909 ( .B1(n12464), .B2(n12463), .A(n12462), .ZN(n12468) );
  MUX2_X1 U14910 ( .A(n12466), .B(n12465), .S(n12578), .Z(n12467) );
  NAND3_X1 U14911 ( .A1(n12468), .A2(n15566), .A3(n12467), .ZN(n12473) );
  MUX2_X1 U14912 ( .A(n12470), .B(n12469), .S(n12587), .Z(n12471) );
  NAND3_X1 U14913 ( .A1(n12473), .A2(n12472), .A3(n12471), .ZN(n12478) );
  NAND2_X1 U14914 ( .A1(n12479), .A2(n12474), .ZN(n12475) );
  NAND2_X1 U14915 ( .A1(n12475), .A2(n12578), .ZN(n12476) );
  NAND3_X1 U14916 ( .A1(n12478), .A2(n12477), .A3(n12476), .ZN(n12482) );
  NOR2_X1 U14917 ( .A1(n12479), .A2(n12578), .ZN(n12480) );
  NOR2_X1 U14918 ( .A1(n12480), .A2(n15540), .ZN(n12481) );
  OAI211_X1 U14919 ( .C1(n12484), .C2(n12483), .A(n12482), .B(n12481), .ZN(
        n12489) );
  MUX2_X1 U14920 ( .A(n12486), .B(n12485), .S(n12587), .Z(n12487) );
  NAND3_X1 U14921 ( .A1(n12489), .A2(n12488), .A3(n12487), .ZN(n12496) );
  INV_X1 U14922 ( .A(n12824), .ZN(n12490) );
  NAND2_X1 U14923 ( .A1(n12491), .A2(n12490), .ZN(n12493) );
  MUX2_X1 U14924 ( .A(n12493), .B(n12492), .S(n12578), .Z(n12494) );
  NAND3_X1 U14925 ( .A1(n12496), .A2(n12495), .A3(n12494), .ZN(n12500) );
  MUX2_X1 U14926 ( .A(n12498), .B(n12497), .S(n12587), .Z(n12499) );
  NAND2_X1 U14927 ( .A1(n12500), .A2(n12499), .ZN(n12505) );
  MUX2_X1 U14928 ( .A(n12502), .B(n12501), .S(n12578), .Z(n12503) );
  NAND2_X1 U14929 ( .A1(n12503), .A2(n14859), .ZN(n12504) );
  AOI21_X1 U14930 ( .B1(n12505), .B2(n8370), .A(n12504), .ZN(n12515) );
  NAND2_X1 U14931 ( .A1(n12511), .A2(n12506), .ZN(n12510) );
  OAI21_X1 U14932 ( .B1(n12508), .B2(n12507), .A(n12512), .ZN(n12509) );
  MUX2_X1 U14933 ( .A(n12510), .B(n12509), .S(n12587), .Z(n12514) );
  INV_X1 U14934 ( .A(n13283), .ZN(n13288) );
  MUX2_X1 U14935 ( .A(n12512), .B(n12511), .S(n12587), .Z(n12513) );
  OAI211_X1 U14936 ( .C1(n12515), .C2(n12514), .A(n13288), .B(n12513), .ZN(
        n12520) );
  MUX2_X1 U14937 ( .A(n12517), .B(n12516), .S(n12587), .Z(n12518) );
  INV_X1 U14938 ( .A(n12518), .ZN(n12519) );
  NAND3_X1 U14939 ( .A1(n12520), .A2(n8654), .A3(n12519), .ZN(n12521) );
  OAI21_X1 U14940 ( .B1(n12578), .B2(n12522), .A(n12521), .ZN(n12523) );
  NAND2_X1 U14941 ( .A1(n12523), .A2(n13262), .ZN(n12529) );
  OAI211_X1 U14942 ( .C1(n13258), .C2(n12525), .A(n12532), .B(n12524), .ZN(
        n12526) );
  NAND2_X1 U14943 ( .A1(n12526), .A2(n12578), .ZN(n12528) );
  INV_X1 U14944 ( .A(n12531), .ZN(n12527) );
  AOI21_X1 U14945 ( .B1(n12529), .B2(n12528), .A(n12527), .ZN(n12534) );
  AOI21_X1 U14946 ( .B1(n12531), .B2(n12530), .A(n12578), .ZN(n12533) );
  OAI22_X1 U14947 ( .A1(n12534), .A2(n12533), .B1(n12532), .B2(n12578), .ZN(
        n12537) );
  NOR2_X1 U14948 ( .A1(n12535), .A2(n12587), .ZN(n12536) );
  AOI21_X1 U14949 ( .B1(n12537), .B2(n13238), .A(n12536), .ZN(n12546) );
  NAND2_X1 U14950 ( .A1(n12548), .A2(n12538), .ZN(n12543) );
  INV_X1 U14951 ( .A(n12538), .ZN(n12541) );
  OAI211_X1 U14952 ( .C1(n12541), .C2(n12540), .A(n12547), .B(n12539), .ZN(
        n12542) );
  MUX2_X1 U14953 ( .A(n12543), .B(n12542), .S(n12587), .Z(n12544) );
  INV_X1 U14954 ( .A(n12544), .ZN(n12545) );
  OAI21_X1 U14955 ( .B1(n12546), .B2(n8502), .A(n12545), .ZN(n12550) );
  MUX2_X1 U14956 ( .A(n12548), .B(n12547), .S(n12578), .Z(n12549) );
  NAND3_X1 U14957 ( .A1(n12550), .A2(n13186), .A3(n12549), .ZN(n12554) );
  NAND2_X1 U14958 ( .A1(n13332), .A2(n13175), .ZN(n12552) );
  MUX2_X1 U14959 ( .A(n12552), .B(n12551), .S(n12587), .Z(n12553) );
  NAND3_X1 U14960 ( .A1(n12554), .A2(n13177), .A3(n12553), .ZN(n12558) );
  MUX2_X1 U14961 ( .A(n12556), .B(n12555), .S(n12578), .Z(n12557) );
  NAND3_X1 U14962 ( .A1(n12558), .A2(n13158), .A3(n12557), .ZN(n12561) );
  NAND3_X1 U14963 ( .A1(n12561), .A2(n13149), .A3(n12559), .ZN(n12565) );
  NAND3_X1 U14964 ( .A1(n12561), .A2(n13149), .A3(n12560), .ZN(n12563) );
  AND2_X1 U14965 ( .A1(n12563), .A2(n12562), .ZN(n12564) );
  MUX2_X1 U14966 ( .A(n12565), .B(n12564), .S(n12587), .Z(n12573) );
  NAND2_X1 U14967 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  NAND2_X1 U14968 ( .A1(n12568), .A2(n12578), .ZN(n12570) );
  MUX2_X1 U14969 ( .A(n12578), .B(n12570), .S(n12569), .Z(n12571) );
  OAI211_X1 U14970 ( .C1(n12573), .C2(n13132), .A(n12572), .B(n12571), .ZN(
        n12577) );
  MUX2_X1 U14971 ( .A(n12575), .B(n12574), .S(n12587), .Z(n12576) );
  NAND3_X1 U14972 ( .A1(n13102), .A2(n12577), .A3(n12576), .ZN(n12582) );
  MUX2_X1 U14973 ( .A(n12580), .B(n12579), .S(n12578), .Z(n12581) );
  NAND2_X1 U14974 ( .A1(n12582), .A2(n12581), .ZN(n12583) );
  NAND2_X1 U14975 ( .A1(n13088), .A2(n12583), .ZN(n12589) );
  NAND2_X1 U14976 ( .A1(n13378), .A2(n12928), .ZN(n12584) );
  NAND2_X1 U14977 ( .A1(n13076), .A2(n12587), .ZN(n12590) );
  OAI21_X1 U14978 ( .B1(n12590), .B2(n12589), .A(n12588), .ZN(n12593) );
  OAI211_X1 U14979 ( .C1(n12594), .C2(n12593), .A(n12592), .B(n12591), .ZN(
        n12597) );
  AOI21_X1 U14980 ( .B1(n12597), .B2(n12596), .A(n12595), .ZN(n12598) );
  MUX2_X1 U14981 ( .A(n15585), .B(n12599), .S(n12598), .Z(n12600) );
  NAND2_X1 U14982 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  OAI211_X1 U14983 ( .C1(n12606), .C2(n12608), .A(n12605), .B(P3_B_REG_SCAN_IN), .ZN(n12607) );
  OAI222_X1 U14984 ( .A1(n14106), .A2(n12610), .B1(n14111), .B2(n12609), .C1(
        n9752), .C2(P2_U3088), .ZN(P2_U3306) );
  NOR3_X1 U14985 ( .A1(n6939), .A2(n10413), .A3(n7688), .ZN(n12613) );
  AOI211_X1 U14986 ( .C1(n12615), .C2(n12611), .A(n12614), .B(n12613), .ZN(
        n12620) );
  AOI22_X1 U14987 ( .A1(n12914), .A2(n15609), .B1(n15608), .B2(n12936), .ZN(
        n12616) );
  OAI21_X1 U14988 ( .B1(n15606), .B2(n12931), .A(n12616), .ZN(n12617) );
  AOI21_X1 U14989 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n12618), .A(n12617), .ZN(
        n12619) );
  OAI21_X1 U14990 ( .B1(n12620), .B2(n12945), .A(n12619), .ZN(P3_U3162) );
  INV_X1 U14991 ( .A(n12621), .ZN(n12622) );
  OAI222_X1 U14992 ( .A1(P3_U3151), .A2(n12623), .B1(n13439), .B2(n12622), 
        .C1(n13430), .C2(n12414), .ZN(P3_U3265) );
  INV_X1 U14993 ( .A(n12624), .ZN(n14110) );
  OAI222_X1 U14994 ( .A1(P1_U3086), .A2(n10209), .B1(n14775), .B2(n14110), 
        .C1(n12625), .C2(n14777), .ZN(P1_U3330) );
  INV_X1 U14995 ( .A(n12626), .ZN(n12628) );
  NAND2_X1 U14996 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  AOI22_X1 U14997 ( .A1(n14192), .A2(n12769), .B1(n12767), .B2(n14262), .ZN(
        n12632) );
  AOI22_X1 U14998 ( .A1(n14192), .A2(n12770), .B1(n12769), .B2(n14262), .ZN(
        n12631) );
  XNOR2_X1 U14999 ( .A(n12631), .B(n12756), .ZN(n12633) );
  XOR2_X1 U15000 ( .A(n12632), .B(n12633), .Z(n14189) );
  INV_X1 U15001 ( .A(n12632), .ZN(n12635) );
  NOR2_X1 U15002 ( .A1(n12726), .A2(n14971), .ZN(n12637) );
  AOI21_X1 U15003 ( .B1(n12638), .B2(n12769), .A(n12637), .ZN(n12645) );
  AOI22_X1 U15004 ( .A1(n12638), .A2(n12770), .B1(n12769), .B2(n14261), .ZN(
        n12639) );
  XNOR2_X1 U15005 ( .A(n12639), .B(n12756), .ZN(n12644) );
  XOR2_X1 U15006 ( .A(n12645), .B(n12644), .Z(n14134) );
  NAND2_X1 U15007 ( .A1(n14135), .A2(n14134), .ZN(n14133) );
  NAND2_X1 U15008 ( .A1(n15013), .A2(n12770), .ZN(n12641) );
  NAND2_X1 U15009 ( .A1(n12769), .A2(n14260), .ZN(n12640) );
  NAND2_X1 U15010 ( .A1(n12641), .A2(n12640), .ZN(n12642) );
  INV_X2 U15011 ( .A(n6708), .ZN(n12756) );
  XNOR2_X1 U15012 ( .A(n12642), .B(n12756), .ZN(n12651) );
  NOR2_X1 U15013 ( .A1(n12726), .A2(n14137), .ZN(n12643) );
  AOI21_X1 U15014 ( .B1(n15013), .B2(n12769), .A(n12643), .ZN(n12649) );
  XNOR2_X1 U15015 ( .A(n12651), .B(n12649), .ZN(n14973) );
  INV_X1 U15016 ( .A(n12644), .ZN(n12647) );
  INV_X1 U15017 ( .A(n12645), .ZN(n12646) );
  NAND2_X1 U15018 ( .A1(n12647), .A2(n12646), .ZN(n14974) );
  INV_X1 U15019 ( .A(n12649), .ZN(n12650) );
  OR2_X1 U15020 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  NOR2_X1 U15021 ( .A1(n12726), .A2(n14970), .ZN(n12653) );
  AOI21_X1 U15022 ( .B1(n14172), .B2(n12769), .A(n12653), .ZN(n12657) );
  NAND2_X1 U15023 ( .A1(n14172), .A2(n12770), .ZN(n12655) );
  NAND2_X1 U15024 ( .A1(n12769), .A2(n14259), .ZN(n12654) );
  NAND2_X1 U15025 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  XNOR2_X1 U15026 ( .A(n12656), .B(n12756), .ZN(n12659) );
  XOR2_X1 U15027 ( .A(n12657), .B(n12659), .Z(n14169) );
  INV_X1 U15028 ( .A(n12657), .ZN(n12658) );
  NAND2_X1 U15029 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  NAND2_X1 U15030 ( .A1(n14166), .A2(n12660), .ZN(n14210) );
  NOR2_X1 U15031 ( .A1(n12726), .A2(n14930), .ZN(n12661) );
  AOI21_X1 U15032 ( .B1(n12662), .B2(n12769), .A(n12661), .ZN(n12669) );
  AOI22_X1 U15033 ( .A1(n12662), .A2(n12770), .B1(n12769), .B2(n14258), .ZN(
        n12663) );
  XNOR2_X1 U15034 ( .A(n12663), .B(n12756), .ZN(n12670) );
  XOR2_X1 U15035 ( .A(n12669), .B(n12670), .Z(n14211) );
  NAND2_X1 U15036 ( .A1(n14210), .A2(n14211), .ZN(n14209) );
  NAND2_X1 U15037 ( .A1(n14938), .A2(n12770), .ZN(n12665) );
  NAND2_X1 U15038 ( .A1(n12769), .A2(n14257), .ZN(n12664) );
  NAND2_X1 U15039 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  XNOR2_X1 U15040 ( .A(n12666), .B(n6708), .ZN(n12672) );
  NOR2_X1 U15041 ( .A1(n12726), .A2(n12667), .ZN(n12668) );
  AOI21_X1 U15042 ( .B1(n14938), .B2(n12769), .A(n12668), .ZN(n12673) );
  XNOR2_X1 U15043 ( .A(n12672), .B(n12673), .ZN(n14931) );
  NOR2_X1 U15044 ( .A1(n12670), .A2(n12669), .ZN(n14932) );
  NOR2_X1 U15045 ( .A1(n14931), .A2(n14932), .ZN(n12671) );
  NAND2_X1 U15046 ( .A1(n14209), .A2(n12671), .ZN(n14934) );
  INV_X1 U15047 ( .A(n12672), .ZN(n12675) );
  INV_X1 U15048 ( .A(n12673), .ZN(n12674) );
  NAND2_X1 U15049 ( .A1(n14416), .A2(n12770), .ZN(n12677) );
  NAND2_X1 U15050 ( .A1(n12769), .A2(n14642), .ZN(n12676) );
  NAND2_X1 U15051 ( .A1(n12677), .A2(n12676), .ZN(n12678) );
  XNOR2_X1 U15052 ( .A(n12678), .B(n12756), .ZN(n12680) );
  INV_X1 U15053 ( .A(n14416), .ZN(n14255) );
  OAI22_X1 U15054 ( .A1(n14255), .A2(n10604), .B1(n14943), .B2(n12726), .ZN(
        n14248) );
  INV_X1 U15055 ( .A(n12679), .ZN(n12681) );
  NAND2_X1 U15056 ( .A1(n14951), .A2(n12770), .ZN(n12683) );
  NAND2_X1 U15057 ( .A1(n12769), .A2(n14959), .ZN(n12682) );
  NAND2_X1 U15058 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  XNOR2_X1 U15059 ( .A(n12684), .B(n6708), .ZN(n12688) );
  NOR2_X1 U15060 ( .A1(n12726), .A2(n14738), .ZN(n12685) );
  AOI21_X1 U15061 ( .B1(n14951), .B2(n12769), .A(n12685), .ZN(n12687) );
  XNOR2_X1 U15062 ( .A(n12688), .B(n12687), .ZN(n14944) );
  NAND2_X1 U15063 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U15064 ( .A1(n14947), .A2(n12689), .ZN(n14956) );
  NAND2_X1 U15065 ( .A1(n14991), .A2(n12770), .ZN(n12691) );
  NAND2_X1 U15066 ( .A1(n12768), .A2(n14644), .ZN(n12690) );
  NAND2_X1 U15067 ( .A1(n12691), .A2(n12690), .ZN(n12692) );
  XNOR2_X1 U15068 ( .A(n12692), .B(n12756), .ZN(n12693) );
  AOI22_X1 U15069 ( .A1(n14991), .A2(n12769), .B1(n12767), .B2(n14644), .ZN(
        n12694) );
  XNOR2_X1 U15070 ( .A(n12693), .B(n12694), .ZN(n14955) );
  NAND2_X1 U15071 ( .A1(n14956), .A2(n14955), .ZN(n12697) );
  INV_X1 U15072 ( .A(n12693), .ZN(n12695) );
  NAND2_X1 U15073 ( .A1(n12695), .A2(n12694), .ZN(n12696) );
  NAND2_X1 U15074 ( .A1(n12697), .A2(n12696), .ZN(n14231) );
  NAND2_X1 U15075 ( .A1(n14727), .A2(n12770), .ZN(n12699) );
  NAND2_X1 U15076 ( .A1(n12769), .A2(n14957), .ZN(n12698) );
  NAND2_X1 U15077 ( .A1(n12699), .A2(n12698), .ZN(n12700) );
  XNOR2_X1 U15078 ( .A(n12700), .B(n12756), .ZN(n12701) );
  AOI22_X1 U15079 ( .A1(n14727), .A2(n12769), .B1(n12767), .B2(n14957), .ZN(
        n12702) );
  XNOR2_X1 U15080 ( .A(n12701), .B(n12702), .ZN(n14230) );
  INV_X1 U15081 ( .A(n12701), .ZN(n12703) );
  NAND2_X1 U15082 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  NOR2_X1 U15083 ( .A1(n12726), .A2(n14233), .ZN(n12705) );
  AOI21_X1 U15084 ( .B1(n14721), .B2(n12768), .A(n12705), .ZN(n12710) );
  NAND2_X1 U15085 ( .A1(n14721), .A2(n12770), .ZN(n12707) );
  NAND2_X1 U15086 ( .A1(n12768), .A2(n14627), .ZN(n12706) );
  NAND2_X1 U15087 ( .A1(n12707), .A2(n12706), .ZN(n12708) );
  XNOR2_X1 U15088 ( .A(n12708), .B(n12756), .ZN(n12712) );
  XOR2_X1 U15089 ( .A(n12710), .B(n12712), .Z(n14144) );
  INV_X1 U15090 ( .A(n14144), .ZN(n12709) );
  INV_X1 U15091 ( .A(n12710), .ZN(n12711) );
  NAND2_X1 U15092 ( .A1(n12712), .A2(n12711), .ZN(n12713) );
  NAND2_X1 U15093 ( .A1(n14714), .A2(n12770), .ZN(n12715) );
  NAND2_X1 U15094 ( .A1(n14584), .A2(n12769), .ZN(n12714) );
  NAND2_X1 U15095 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  XNOR2_X1 U15096 ( .A(n12716), .B(n12756), .ZN(n12719) );
  AOI22_X1 U15097 ( .A1(n14714), .A2(n12769), .B1(n12767), .B2(n14584), .ZN(
        n12717) );
  XNOR2_X1 U15098 ( .A(n12719), .B(n12717), .ZN(n14199) );
  INV_X1 U15099 ( .A(n12717), .ZN(n12718) );
  NAND2_X1 U15100 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  AOI22_X1 U15101 ( .A1(n14709), .A2(n12770), .B1(n12768), .B2(n14565), .ZN(
        n12721) );
  XNOR2_X1 U15102 ( .A(n12721), .B(n12756), .ZN(n12724) );
  AOI22_X1 U15103 ( .A1(n14709), .A2(n12769), .B1(n12767), .B2(n14565), .ZN(
        n12723) );
  XNOR2_X1 U15104 ( .A(n12724), .B(n12723), .ZN(n14155) );
  NAND2_X1 U15105 ( .A1(n12724), .A2(n12723), .ZN(n12725) );
  OAI22_X1 U15106 ( .A1(n14572), .A2(n10604), .B1(n14440), .B2(n12726), .ZN(
        n12730) );
  OAI22_X1 U15107 ( .A1(n14572), .A2(n12727), .B1(n14440), .B2(n10604), .ZN(
        n12728) );
  XNOR2_X1 U15108 ( .A(n12728), .B(n12756), .ZN(n12729) );
  XOR2_X1 U15109 ( .A(n12730), .B(n12729), .Z(n14222) );
  INV_X1 U15110 ( .A(n12729), .ZN(n12732) );
  INV_X1 U15111 ( .A(n12730), .ZN(n12731) );
  NAND2_X1 U15112 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  NAND2_X1 U15113 ( .A1(n14562), .A2(n12770), .ZN(n12735) );
  NAND2_X1 U15114 ( .A1(n12768), .A2(n14566), .ZN(n12734) );
  NAND2_X1 U15115 ( .A1(n12735), .A2(n12734), .ZN(n12736) );
  XNOR2_X1 U15116 ( .A(n12736), .B(n12756), .ZN(n12737) );
  AOI22_X1 U15117 ( .A1(n14562), .A2(n12769), .B1(n12767), .B2(n14566), .ZN(
        n12738) );
  XNOR2_X1 U15118 ( .A(n12737), .B(n12738), .ZN(n14124) );
  INV_X1 U15119 ( .A(n12737), .ZN(n12739) );
  NAND2_X1 U15120 ( .A1(n12739), .A2(n12738), .ZN(n12740) );
  NAND2_X1 U15121 ( .A1(n14549), .A2(n12770), .ZN(n12742) );
  NAND2_X1 U15122 ( .A1(n12768), .A2(n14523), .ZN(n12741) );
  NAND2_X1 U15123 ( .A1(n12742), .A2(n12741), .ZN(n12743) );
  XNOR2_X1 U15124 ( .A(n12743), .B(n12756), .ZN(n12744) );
  AOI22_X1 U15125 ( .A1(n14549), .A2(n12769), .B1(n12767), .B2(n14523), .ZN(
        n12745) );
  XNOR2_X1 U15126 ( .A(n12744), .B(n12745), .ZN(n14182) );
  INV_X1 U15127 ( .A(n12744), .ZN(n12746) );
  NAND2_X1 U15128 ( .A1(n14518), .A2(n12770), .ZN(n12748) );
  NAND2_X1 U15129 ( .A1(n12768), .A2(n14504), .ZN(n12747) );
  NAND2_X1 U15130 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  XNOR2_X1 U15131 ( .A(n12749), .B(n12756), .ZN(n12750) );
  AOI22_X1 U15132 ( .A1(n14518), .A2(n12769), .B1(n12767), .B2(n14504), .ZN(
        n12751) );
  XNOR2_X1 U15133 ( .A(n12750), .B(n12751), .ZN(n14175) );
  INV_X1 U15134 ( .A(n12750), .ZN(n12752) );
  NAND2_X1 U15135 ( .A1(n12752), .A2(n12751), .ZN(n12753) );
  NAND2_X1 U15136 ( .A1(n14507), .A2(n12770), .ZN(n12755) );
  NAND2_X1 U15137 ( .A1(n12768), .A2(n14524), .ZN(n12754) );
  NAND2_X1 U15138 ( .A1(n12755), .A2(n12754), .ZN(n12757) );
  XNOR2_X1 U15139 ( .A(n12757), .B(n12756), .ZN(n12758) );
  AOI22_X1 U15140 ( .A1(n14507), .A2(n12768), .B1(n12767), .B2(n14524), .ZN(
        n12759) );
  XNOR2_X1 U15141 ( .A(n12758), .B(n12759), .ZN(n14239) );
  INV_X1 U15142 ( .A(n12758), .ZN(n12760) );
  NAND2_X1 U15143 ( .A1(n14497), .A2(n12770), .ZN(n12762) );
  NAND2_X1 U15144 ( .A1(n12768), .A2(n14505), .ZN(n12761) );
  NAND2_X1 U15145 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  XNOR2_X1 U15146 ( .A(n12763), .B(n12756), .ZN(n12764) );
  AOI22_X1 U15147 ( .A1(n14497), .A2(n12769), .B1(n12767), .B2(n14505), .ZN(
        n12765) );
  XNOR2_X1 U15148 ( .A(n12764), .B(n12765), .ZN(n14116) );
  INV_X1 U15149 ( .A(n12764), .ZN(n12766) );
  AOI22_X1 U15150 ( .A1(n14477), .A2(n12768), .B1(n12767), .B2(n14447), .ZN(
        n12773) );
  AOI22_X1 U15151 ( .A1(n14477), .A2(n12770), .B1(n12769), .B2(n14447), .ZN(
        n12771) );
  XNOR2_X1 U15152 ( .A(n12771), .B(n12756), .ZN(n12772) );
  XOR2_X1 U15153 ( .A(n12773), .B(n12772), .Z(n12774) );
  XNOR2_X1 U15154 ( .A(n12775), .B(n12774), .ZN(n12780) );
  NAND2_X1 U15155 ( .A1(n14244), .A2(n14473), .ZN(n12777) );
  AOI22_X1 U15156 ( .A1(n14960), .A2(n14505), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12776) );
  OAI211_X1 U15157 ( .C1(n14469), .C2(n14969), .A(n12777), .B(n12776), .ZN(
        n12778) );
  AOI21_X1 U15158 ( .B1(n14477), .B2(n14981), .A(n12778), .ZN(n12779) );
  OAI21_X1 U15159 ( .B1(n12780), .B2(n14976), .A(n12779), .ZN(P1_U3220) );
  AOI21_X1 U15160 ( .B1(n12782), .B2(n12781), .A(n6816), .ZN(n12790) );
  INV_X1 U15161 ( .A(n13418), .ZN(n12788) );
  NOR2_X1 U15162 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12783), .ZN(n12973) );
  AOI21_X1 U15163 ( .B1(n14851), .B2(n12914), .A(n12973), .ZN(n12786) );
  INV_X1 U15164 ( .A(n12784), .ZN(n13278) );
  NAND2_X1 U15165 ( .A1(n12938), .A2(n13278), .ZN(n12785) );
  OAI211_X1 U15166 ( .C1(n13275), .C2(n12917), .A(n12786), .B(n12785), .ZN(
        n12787) );
  AOI21_X1 U15167 ( .B1(n12788), .B2(n12943), .A(n12787), .ZN(n12789) );
  OAI21_X1 U15168 ( .B1(n12790), .B2(n12945), .A(n12789), .ZN(P3_U3155) );
  AOI21_X1 U15169 ( .B1(n12873), .B2(n12792), .A(n12870), .ZN(n12797) );
  AOI22_X1 U15170 ( .A1(n12904), .A2(n12914), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12794) );
  NAND2_X1 U15171 ( .A1(n13152), .A2(n12938), .ZN(n12793) );
  OAI211_X1 U15172 ( .C1(n13145), .C2(n12917), .A(n12794), .B(n12793), .ZN(
        n12795) );
  AOI21_X1 U15173 ( .B1(n13319), .B2(n12943), .A(n12795), .ZN(n12796) );
  OAI21_X1 U15174 ( .B1(n12797), .B2(n12945), .A(n12796), .ZN(P3_U3156) );
  INV_X1 U15175 ( .A(n12798), .ZN(n13398) );
  NAND2_X1 U15176 ( .A1(n12799), .A2(n12800), .ZN(n12880) );
  OAI211_X1 U15177 ( .C1(n12799), .C2(n12800), .A(n12880), .B(n12924), .ZN(
        n12804) );
  NAND2_X1 U15178 ( .A1(n13203), .A2(n12914), .ZN(n12801) );
  NAND2_X1 U15179 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13053)
         );
  OAI211_X1 U15180 ( .C1(n13175), .C2(n12917), .A(n12801), .B(n13053), .ZN(
        n12802) );
  AOI21_X1 U15181 ( .B1(n13209), .B2(n12938), .A(n12802), .ZN(n12803) );
  OAI211_X1 U15182 ( .C1(n13398), .C2(n12931), .A(n12804), .B(n12803), .ZN(
        P3_U3159) );
  XNOR2_X1 U15183 ( .A(n13076), .B(n7688), .ZN(n12811) );
  INV_X1 U15184 ( .A(n12811), .ZN(n12805) );
  NAND2_X1 U15185 ( .A1(n12805), .A2(n12924), .ZN(n12817) );
  INV_X1 U15186 ( .A(n12806), .ZN(n12807) );
  NAND4_X1 U15187 ( .A1(n12816), .A2(n12924), .A3(n12807), .A4(n12811), .ZN(
        n12815) );
  AOI22_X1 U15188 ( .A1(n13079), .A2(n12938), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12809) );
  NAND2_X1 U15189 ( .A1(n12928), .A2(n12914), .ZN(n12808) );
  OAI211_X1 U15190 ( .C1(n13072), .C2(n12917), .A(n12809), .B(n12808), .ZN(
        n12813) );
  NOR4_X1 U15191 ( .A1(n12811), .A2(n12810), .A3(n12945), .A4(n12928), .ZN(
        n12812) );
  AOI211_X1 U15192 ( .C1(n12943), .C2(n7039), .A(n12813), .B(n12812), .ZN(
        n12814) );
  OAI211_X1 U15193 ( .C1(n12817), .C2(n12816), .A(n12815), .B(n12814), .ZN(
        P3_U3160) );
  MUX2_X1 U15194 ( .A(n12951), .B(n12819), .S(n12818), .Z(n12821) );
  XNOR2_X1 U15195 ( .A(n12821), .B(n12820), .ZN(n12822) );
  NAND2_X1 U15196 ( .A1(n12822), .A2(n12924), .ZN(n12829) );
  NOR2_X1 U15197 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12823), .ZN(n15495) );
  AOI21_X1 U15198 ( .B1(n12914), .B2(n12951), .A(n15495), .ZN(n12828) );
  AOI22_X1 U15199 ( .A1(n12936), .A2(n15528), .B1(n12943), .B2(n12824), .ZN(
        n12827) );
  NAND2_X1 U15200 ( .A1(n12938), .A2(n12825), .ZN(n12826) );
  NAND4_X1 U15201 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        P3_U3161) );
  INV_X1 U15202 ( .A(n12830), .ZN(n12831) );
  AOI21_X1 U15203 ( .B1(n12833), .B2(n12832), .A(n12831), .ZN(n12839) );
  OAI22_X1 U15204 ( .A1(n13175), .A2(n12941), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12834), .ZN(n12836) );
  NOR2_X1 U15205 ( .A1(n13176), .A2(n12917), .ZN(n12835) );
  AOI211_X1 U15206 ( .C1(n13180), .C2(n12938), .A(n12836), .B(n12835), .ZN(
        n12838) );
  NAND2_X1 U15207 ( .A1(n13179), .A2(n12943), .ZN(n12837) );
  OAI211_X1 U15208 ( .C1(n12839), .C2(n12945), .A(n12838), .B(n12837), .ZN(
        P3_U3163) );
  AOI22_X1 U15209 ( .A1(n13115), .A2(n12914), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12841) );
  NAND2_X1 U15210 ( .A1(n13121), .A2(n12938), .ZN(n12840) );
  OAI211_X1 U15211 ( .C1(n13090), .C2(n12917), .A(n12841), .B(n12840), .ZN(
        n12847) );
  NAND3_X1 U15212 ( .A1(n12842), .A2(n12844), .A3(n6921), .ZN(n12845) );
  INV_X1 U15213 ( .A(n12848), .ZN(P3_U3165) );
  INV_X1 U15214 ( .A(n12849), .ZN(n13410) );
  OAI211_X1 U15215 ( .C1(n12852), .C2(n12851), .A(n12850), .B(n12924), .ZN(
        n12856) );
  NAND2_X1 U15216 ( .A1(n12949), .A2(n12914), .ZN(n12853) );
  NAND2_X1 U15217 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13012)
         );
  OAI211_X1 U15218 ( .C1(n13249), .C2(n12917), .A(n12853), .B(n13012), .ZN(
        n12854) );
  AOI21_X1 U15219 ( .B1(n13252), .B2(n12938), .A(n12854), .ZN(n12855) );
  OAI211_X1 U15220 ( .C1(n13410), .C2(n12931), .A(n12856), .B(n12855), .ZN(
        P3_U3166) );
  INV_X1 U15221 ( .A(n12857), .ZN(n12858) );
  AOI21_X1 U15222 ( .B1(n12860), .B2(n12859), .A(n12858), .ZN(n12866) );
  NOR2_X1 U15223 ( .A1(n13260), .A2(n12941), .ZN(n12863) );
  OAI22_X1 U15224 ( .A1(n13236), .A2(n12917), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12861), .ZN(n12862) );
  AOI211_X1 U15225 ( .C1(n13241), .C2(n12938), .A(n12863), .B(n12862), .ZN(
        n12865) );
  NAND2_X1 U15226 ( .A1(n13240), .A2(n12943), .ZN(n12864) );
  OAI211_X1 U15227 ( .C1(n12866), .C2(n12945), .A(n12865), .B(n12864), .ZN(
        P3_U3168) );
  INV_X1 U15228 ( .A(n12867), .ZN(n12869) );
  NOR3_X1 U15229 ( .A1(n12870), .A2(n12869), .A3(n12868), .ZN(n12872) );
  INV_X1 U15230 ( .A(n12842), .ZN(n12871) );
  OAI21_X1 U15231 ( .B1(n12872), .B2(n12871), .A(n12924), .ZN(n12878) );
  AOI22_X1 U15232 ( .A1(n13137), .A2(n12938), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12877) );
  AOI22_X1 U15233 ( .A1(n12874), .A2(n12936), .B1(n12914), .B2(n12873), .ZN(
        n12876) );
  NAND2_X1 U15234 ( .A1(n13314), .A2(n12943), .ZN(n12875) );
  NAND4_X1 U15235 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        P3_U3169) );
  NAND2_X1 U15236 ( .A1(n12880), .A2(n12879), .ZN(n12883) );
  XNOR2_X1 U15237 ( .A(n12881), .B(n13204), .ZN(n12882) );
  XNOR2_X1 U15238 ( .A(n12883), .B(n12882), .ZN(n12888) );
  AOI22_X1 U15239 ( .A1(n13188), .A2(n12936), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(n6665), .ZN(n12885) );
  NAND2_X1 U15240 ( .A1(n12938), .A2(n13194), .ZN(n12884) );
  OAI211_X1 U15241 ( .C1(n13222), .C2(n12941), .A(n12885), .B(n12884), .ZN(
        n12886) );
  AOI21_X1 U15242 ( .B1(n13332), .B2(n12943), .A(n12886), .ZN(n12887) );
  OAI21_X1 U15243 ( .B1(n12888), .B2(n12945), .A(n12887), .ZN(P3_U3173) );
  XNOR2_X1 U15244 ( .A(n12889), .B(n14851), .ZN(n12890) );
  XNOR2_X1 U15245 ( .A(n12891), .B(n12890), .ZN(n12900) );
  INV_X1 U15246 ( .A(n13422), .ZN(n12898) );
  NOR2_X1 U15247 ( .A1(n14863), .A2(n12941), .ZN(n12892) );
  AOI211_X1 U15248 ( .C1(n12936), .C2(n12894), .A(n12893), .B(n12892), .ZN(
        n12895) );
  OAI21_X1 U15249 ( .B1(n13290), .B2(n12896), .A(n12895), .ZN(n12897) );
  AOI21_X1 U15250 ( .B1(n12898), .B2(n12943), .A(n12897), .ZN(n12899) );
  OAI21_X1 U15251 ( .B1(n12900), .B2(n12945), .A(n12899), .ZN(P3_U3174) );
  INV_X1 U15252 ( .A(n12901), .ZN(n12902) );
  AOI21_X1 U15253 ( .B1(n12904), .B2(n12903), .A(n12902), .ZN(n12909) );
  AOI22_X1 U15254 ( .A1(n13188), .A2(n12914), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(n6665), .ZN(n12906) );
  NAND2_X1 U15255 ( .A1(n13166), .A2(n12938), .ZN(n12905) );
  OAI211_X1 U15256 ( .C1(n13161), .C2(n12917), .A(n12906), .B(n12905), .ZN(
        n12907) );
  AOI21_X1 U15257 ( .B1(n13165), .B2(n12943), .A(n12907), .ZN(n12908) );
  OAI21_X1 U15258 ( .B1(n12909), .B2(n12945), .A(n12908), .ZN(P3_U3175) );
  INV_X1 U15259 ( .A(n13228), .ZN(n13402) );
  AOI21_X1 U15260 ( .B1(n12911), .B2(n12910), .A(n12945), .ZN(n12913) );
  NAND2_X1 U15261 ( .A1(n12913), .A2(n12912), .ZN(n12920) );
  NAND2_X1 U15262 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U15263 ( .A1(n6665), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14841) );
  OAI211_X1 U15264 ( .C1(n13222), .C2(n12917), .A(n12916), .B(n14841), .ZN(
        n12918) );
  AOI21_X1 U15265 ( .B1(n13223), .B2(n12938), .A(n12918), .ZN(n12919) );
  OAI211_X1 U15266 ( .C1(n13402), .C2(n12931), .A(n12920), .B(n12919), .ZN(
        P3_U3178) );
  INV_X1 U15267 ( .A(n13306), .ZN(n13108) );
  OAI21_X1 U15268 ( .B1(n12923), .B2(n12922), .A(n12921), .ZN(n12925) );
  NAND2_X1 U15269 ( .A1(n12925), .A2(n12924), .ZN(n12930) );
  AOI22_X1 U15270 ( .A1(n13106), .A2(n12938), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12926) );
  OAI21_X1 U15271 ( .B1(n13130), .B2(n12941), .A(n12926), .ZN(n12927) );
  AOI21_X1 U15272 ( .B1(n12928), .B2(n12936), .A(n12927), .ZN(n12929) );
  OAI211_X1 U15273 ( .C1(n13108), .C2(n12931), .A(n12930), .B(n12929), .ZN(
        P3_U3180) );
  XNOR2_X1 U15274 ( .A(n12933), .B(n12949), .ZN(n12934) );
  XNOR2_X1 U15275 ( .A(n12932), .B(n12934), .ZN(n12946) );
  NOR2_X1 U15276 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12935), .ZN(n12995) );
  AOI21_X1 U15277 ( .B1(n12948), .B2(n12936), .A(n12995), .ZN(n12940) );
  INV_X1 U15278 ( .A(n12937), .ZN(n13265) );
  NAND2_X1 U15279 ( .A1(n12938), .A2(n13265), .ZN(n12939) );
  OAI211_X1 U15280 ( .C1(n13286), .C2(n12941), .A(n12940), .B(n12939), .ZN(
        n12942) );
  AOI21_X1 U15281 ( .B1(n13264), .B2(n12943), .A(n12942), .ZN(n12944) );
  OAI21_X1 U15282 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(P3_U3181) );
  MUX2_X1 U15283 ( .A(n12947), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12950), .Z(
        P3_U3521) );
  MUX2_X1 U15284 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13188), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15285 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13203), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15286 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12948), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15287 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12949), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15288 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14851), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15289 ( .A(n12951), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12950), .Z(
        P3_U3498) );
  NOR2_X1 U15290 ( .A1(n12964), .A2(n12952), .ZN(n12954) );
  NAND2_X1 U15291 ( .A1(n12976), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12987) );
  OR2_X1 U15292 ( .A1(n12976), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12955) );
  NAND2_X1 U15293 ( .A1(n12987), .A2(n12955), .ZN(n12966) );
  AOI21_X1 U15294 ( .B1(n12956), .B2(n12966), .A(n12981), .ZN(n12980) );
  NAND2_X1 U15295 ( .A1(n12958), .A2(n12957), .ZN(n12960) );
  NAND2_X1 U15296 ( .A1(n12976), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12986) );
  OR2_X1 U15297 ( .A1(n12976), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12961) );
  AND2_X1 U15298 ( .A1(n12986), .A2(n12961), .ZN(n12967) );
  OAI21_X1 U15299 ( .B1(n12962), .B2(n12967), .A(n12984), .ZN(n12978) );
  INV_X1 U15300 ( .A(n12963), .ZN(n12965) );
  NAND2_X1 U15301 ( .A1(n12965), .A2(n12964), .ZN(n12969) );
  AND2_X1 U15302 ( .A1(n12970), .A2(n12969), .ZN(n12972) );
  INV_X1 U15303 ( .A(n12966), .ZN(n12968) );
  MUX2_X1 U15304 ( .A(n12968), .B(n12967), .S(n12990), .Z(n12971) );
  NAND3_X1 U15305 ( .A1(n12970), .A2(n12969), .A3(n12971), .ZN(n12989) );
  OAI211_X1 U15306 ( .C1(n12972), .C2(n12971), .A(n15508), .B(n12989), .ZN(
        n12975) );
  AOI21_X1 U15307 ( .B1(n15516), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12973), 
        .ZN(n12974) );
  OAI211_X1 U15308 ( .C1(n15513), .C2(n12976), .A(n12975), .B(n12974), .ZN(
        n12977) );
  AOI21_X1 U15309 ( .B1(n15519), .B2(n12978), .A(n12977), .ZN(n12979) );
  OAI21_X1 U15310 ( .B1(n12980), .B2(n15523), .A(n12979), .ZN(P3_U3196) );
  AOI21_X1 U15311 ( .B1(n12983), .B2(n12982), .A(n13003), .ZN(n13001) );
  NAND2_X1 U15312 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12985), .ZN(n13008) );
  OAI21_X1 U15313 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12985), .A(n13008), 
        .ZN(n12999) );
  MUX2_X1 U15314 ( .A(n12987), .B(n12986), .S(n12990), .Z(n12988) );
  NAND2_X1 U15315 ( .A1(n12989), .A2(n12988), .ZN(n13018) );
  XNOR2_X1 U15316 ( .A(n13018), .B(n13007), .ZN(n12992) );
  MUX2_X1 U15317 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12990), .Z(n12991) );
  NOR2_X1 U15318 ( .A1(n12992), .A2(n12991), .ZN(n13019) );
  AOI21_X1 U15319 ( .B1(n12992), .B2(n12991), .A(n13019), .ZN(n12997) );
  NOR2_X1 U15320 ( .A1(n13014), .A2(n12993), .ZN(n12994) );
  AOI211_X1 U15321 ( .C1(n14827), .C2(n13020), .A(n12995), .B(n12994), .ZN(
        n12996) );
  OAI21_X1 U15322 ( .B1(n12997), .B2(n15439), .A(n12996), .ZN(n12998) );
  AOI21_X1 U15323 ( .B1(n15519), .B2(n12999), .A(n12998), .ZN(n13000) );
  OAI21_X1 U15324 ( .B1(n13001), .B2(n15523), .A(n13000), .ZN(P3_U3197) );
  AND2_X1 U15325 ( .A1(n13007), .A2(n13002), .ZN(n13004) );
  AOI22_X1 U15326 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13045), .B1(n13031), 
        .B2(n13022), .ZN(n13005) );
  AOI21_X1 U15327 ( .B1(n6744), .B2(n13005), .A(n13030), .ZN(n13029) );
  AOI22_X1 U15328 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13031), .B1(n13045), 
        .B2(n13351), .ZN(n13011) );
  NAND2_X1 U15329 ( .A1(n13007), .A2(n13006), .ZN(n13009) );
  NAND2_X1 U15330 ( .A1(n13009), .A2(n13008), .ZN(n13010) );
  NAND2_X1 U15331 ( .A1(n13011), .A2(n13010), .ZN(n13044) );
  OAI21_X1 U15332 ( .B1(n13011), .B2(n13010), .A(n13044), .ZN(n13017) );
  NOR2_X1 U15333 ( .A1(n15513), .A2(n13031), .ZN(n13016) );
  OAI21_X1 U15334 ( .B1(n13014), .B2(n13013), .A(n13012), .ZN(n13015) );
  AOI211_X1 U15335 ( .C1(n13017), .C2(n15519), .A(n13016), .B(n13015), .ZN(
        n13028) );
  INV_X1 U15336 ( .A(n13018), .ZN(n13021) );
  AOI21_X1 U15337 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(n13035) );
  MUX2_X1 U15338 ( .A(n13022), .B(n13351), .S(n12990), .Z(n13023) );
  NOR2_X1 U15339 ( .A1(n13023), .A2(n13045), .ZN(n13034) );
  INV_X1 U15340 ( .A(n13034), .ZN(n13024) );
  NAND2_X1 U15341 ( .A1(n13023), .A2(n13045), .ZN(n13033) );
  NAND2_X1 U15342 ( .A1(n13024), .A2(n13033), .ZN(n13025) );
  XNOR2_X1 U15343 ( .A(n13035), .B(n13025), .ZN(n13026) );
  NAND2_X1 U15344 ( .A1(n13026), .A2(n15508), .ZN(n13027) );
  OAI211_X1 U15345 ( .C1(n13029), .C2(n15523), .A(n13028), .B(n13027), .ZN(
        P3_U3198) );
  AOI21_X1 U15346 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13031), .A(n13030), 
        .ZN(n13032) );
  XOR2_X1 U15347 ( .A(n13046), .B(n13032), .Z(n14819) );
  AOI22_X1 U15348 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14826), .B1(n13043), 
        .B2(n13225), .ZN(n14838) );
  XNOR2_X1 U15349 ( .A(n13039), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13038) );
  MUX2_X1 U15350 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12990), .Z(n13036) );
  OAI21_X1 U15351 ( .B1(n13035), .B2(n13034), .A(n13033), .ZN(n14815) );
  XNOR2_X1 U15352 ( .A(n13036), .B(n13046), .ZN(n14816) );
  NOR2_X1 U15353 ( .A1(n14815), .A2(n14816), .ZN(n14814) );
  AOI21_X1 U15354 ( .B1(n13036), .B2(n13046), .A(n14814), .ZN(n13037) );
  XNOR2_X1 U15355 ( .A(n13037), .B(n14826), .ZN(n14832) );
  MUX2_X1 U15356 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12990), .Z(n14833) );
  NOR2_X1 U15357 ( .A1(n14832), .A2(n14833), .ZN(n14831) );
  AOI21_X1 U15358 ( .B1(n13037), .B2(n14826), .A(n14831), .ZN(n13042) );
  INV_X1 U15359 ( .A(n13038), .ZN(n13040) );
  XNOR2_X1 U15360 ( .A(n13039), .B(n13339), .ZN(n13049) );
  MUX2_X1 U15361 ( .A(n13040), .B(n13049), .S(n12990), .Z(n13041) );
  XNOR2_X1 U15362 ( .A(n13042), .B(n13041), .ZN(n13056) );
  AOI22_X1 U15363 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n13043), .B1(n14826), 
        .B2(n13343), .ZN(n14830) );
  OAI21_X1 U15364 ( .B1(n13045), .B2(n13351), .A(n13044), .ZN(n13047) );
  NAND2_X1 U15365 ( .A1(n13046), .A2(n13047), .ZN(n13048) );
  XNOR2_X1 U15366 ( .A(n14811), .B(n13047), .ZN(n14813) );
  NAND2_X1 U15367 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14813), .ZN(n14812) );
  NAND2_X1 U15368 ( .A1(n13048), .A2(n14812), .ZN(n14829) );
  NAND2_X1 U15369 ( .A1(n14830), .A2(n14829), .ZN(n14828) );
  OAI21_X1 U15370 ( .B1(n14826), .B2(n13343), .A(n14828), .ZN(n13050) );
  NAND2_X1 U15371 ( .A1(n15516), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13052) );
  OAI211_X1 U15372 ( .C1(n15513), .C2(n13054), .A(n13053), .B(n13052), .ZN(
        n13055) );
  NAND2_X1 U15373 ( .A1(n13064), .A2(n15576), .ZN(n13059) );
  OR2_X1 U15374 ( .A1(n13058), .A2(n13057), .ZN(n13366) );
  AOI21_X1 U15375 ( .B1(n13059), .B2(n13366), .A(n15625), .ZN(n13061) );
  AOI21_X1 U15376 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15625), .A(n13061), 
        .ZN(n13060) );
  OAI21_X1 U15377 ( .B1(n13297), .B2(n13289), .A(n13060), .ZN(P3_U3202) );
  AOI21_X1 U15378 ( .B1(n15625), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13061), 
        .ZN(n13062) );
  OAI21_X1 U15379 ( .B1(n13369), .B2(n13289), .A(n13062), .ZN(P3_U3203) );
  INV_X1 U15380 ( .A(n13063), .ZN(n13070) );
  OR2_X1 U15381 ( .A1(n15599), .A2(n15602), .ZN(n14864) );
  AOI22_X1 U15382 ( .A1(n13064), .A2(n15576), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15625), .ZN(n13065) );
  OAI21_X1 U15383 ( .B1(n13066), .B2(n13289), .A(n13065), .ZN(n13067) );
  AOI21_X1 U15384 ( .B1(n13068), .B2(n15535), .A(n13067), .ZN(n13069) );
  OAI21_X1 U15385 ( .B1(n13070), .B2(n15625), .A(n13069), .ZN(P3_U3204) );
  OAI22_X1 U15386 ( .A1(n13072), .A2(n15588), .B1(n13101), .B2(n15590), .ZN(
        n13073) );
  INV_X1 U15387 ( .A(n13073), .ZN(n13074) );
  INV_X1 U15388 ( .A(n13301), .ZN(n13083) );
  NAND2_X1 U15389 ( .A1(n13087), .A2(n13075), .ZN(n13077) );
  XNOR2_X1 U15390 ( .A(n13077), .B(n13076), .ZN(n13300) );
  AOI22_X1 U15391 ( .A1(n13079), .A2(n15576), .B1(n15625), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13080) );
  OAI21_X1 U15392 ( .B1(n13375), .B2(n13289), .A(n13080), .ZN(n13081) );
  AOI21_X1 U15393 ( .B1(n13300), .B2(n15535), .A(n13081), .ZN(n13082) );
  OAI21_X1 U15394 ( .B1(n13083), .B2(n15625), .A(n13082), .ZN(P3_U3205) );
  INV_X1 U15395 ( .A(n13084), .ZN(n13085) );
  AOI21_X1 U15396 ( .B1(n13088), .B2(n13086), .A(n13085), .ZN(n13094) );
  OAI21_X1 U15397 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13304) );
  OAI22_X1 U15398 ( .A1(n13091), .A2(n15588), .B1(n13090), .B2(n15590), .ZN(
        n13092) );
  AOI21_X1 U15399 ( .B1(n13304), .B2(n15599), .A(n13092), .ZN(n13093) );
  INV_X1 U15400 ( .A(n13303), .ZN(n13099) );
  AOI22_X1 U15401 ( .A1(n13095), .A2(n15576), .B1(n15625), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13096) );
  OAI21_X1 U15402 ( .B1(n13378), .B2(n13289), .A(n13096), .ZN(n13097) );
  AOI21_X1 U15403 ( .B1(n13304), .B2(n13156), .A(n13097), .ZN(n13098) );
  OAI21_X1 U15404 ( .B1(n13099), .B2(n15625), .A(n13098), .ZN(P3_U3206) );
  XNOR2_X1 U15405 ( .A(n13100), .B(n13102), .ZN(n13307) );
  OAI22_X1 U15406 ( .A1(n13101), .A2(n15588), .B1(n13130), .B2(n15590), .ZN(
        n13105) );
  AOI211_X1 U15407 ( .C1(n13307), .C2(n15599), .A(n13105), .B(n13104), .ZN(
        n13309) );
  AOI22_X1 U15408 ( .A1(n13106), .A2(n15576), .B1(n15625), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13107) );
  OAI21_X1 U15409 ( .B1(n13108), .B2(n13289), .A(n13107), .ZN(n13109) );
  AOI21_X1 U15410 ( .B1(n13307), .B2(n13156), .A(n13109), .ZN(n13110) );
  OAI21_X1 U15411 ( .B1(n13309), .B2(n15625), .A(n13110), .ZN(P3_U3207) );
  XNOR2_X1 U15412 ( .A(n13111), .B(n13113), .ZN(n13119) );
  OAI211_X1 U15413 ( .C1(n13114), .C2(n13113), .A(n13112), .B(n15612), .ZN(
        n13118) );
  AOI22_X1 U15414 ( .A1(n13116), .A2(n15607), .B1(n13115), .B2(n15610), .ZN(
        n13117) );
  OAI211_X1 U15415 ( .C1(n15616), .C2(n13119), .A(n13118), .B(n13117), .ZN(
        n13310) );
  INV_X1 U15416 ( .A(n13310), .ZN(n13125) );
  INV_X1 U15417 ( .A(n13119), .ZN(n13311) );
  INV_X1 U15418 ( .A(n13120), .ZN(n13383) );
  AOI22_X1 U15419 ( .A1(n13121), .A2(n15576), .B1(n15625), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13122) );
  OAI21_X1 U15420 ( .B1(n13383), .B2(n13289), .A(n13122), .ZN(n13123) );
  AOI21_X1 U15421 ( .B1(n13311), .B2(n13156), .A(n13123), .ZN(n13124) );
  OAI21_X1 U15422 ( .B1(n13125), .B2(n15625), .A(n13124), .ZN(P3_U3208) );
  INV_X1 U15423 ( .A(n13126), .ZN(n13143) );
  OAI21_X1 U15424 ( .B1(n13143), .B2(n13127), .A(n13132), .ZN(n13129) );
  NAND2_X1 U15425 ( .A1(n13129), .A2(n13128), .ZN(n13315) );
  OAI22_X1 U15426 ( .A1(n13130), .A2(n15588), .B1(n13161), .B2(n15590), .ZN(
        n13136) );
  OAI211_X1 U15427 ( .C1(n13133), .C2(n13132), .A(n13131), .B(n15612), .ZN(
        n13134) );
  INV_X1 U15428 ( .A(n13134), .ZN(n13135) );
  AOI211_X1 U15429 ( .C1(n15599), .C2(n13315), .A(n13136), .B(n13135), .ZN(
        n13317) );
  INV_X1 U15430 ( .A(n13314), .ZN(n13139) );
  AOI22_X1 U15431 ( .A1(n13137), .A2(n15576), .B1(n15625), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13138) );
  OAI21_X1 U15432 ( .B1(n13139), .B2(n13289), .A(n13138), .ZN(n13140) );
  AOI21_X1 U15433 ( .B1(n13315), .B2(n13156), .A(n13140), .ZN(n13141) );
  OAI21_X1 U15434 ( .B1(n13317), .B2(n15625), .A(n13141), .ZN(P3_U3209) );
  INV_X1 U15435 ( .A(n13142), .ZN(n13144) );
  AOI21_X1 U15436 ( .B1(n13144), .B2(n8569), .A(n13143), .ZN(n13318) );
  OAI22_X1 U15437 ( .A1(n13145), .A2(n15588), .B1(n13176), .B2(n15590), .ZN(
        n13151) );
  INV_X1 U15438 ( .A(n13146), .ZN(n13147) );
  AOI211_X1 U15439 ( .C1(n13149), .C2(n13148), .A(n15594), .B(n13147), .ZN(
        n13150) );
  AOI211_X1 U15440 ( .C1(n13318), .C2(n15599), .A(n13151), .B(n13150), .ZN(
        n13321) );
  INV_X1 U15441 ( .A(n13319), .ZN(n13154) );
  AOI22_X1 U15442 ( .A1(n13152), .A2(n15576), .B1(P3_REG2_REG_23__SCAN_IN), 
        .B2(n15625), .ZN(n13153) );
  OAI21_X1 U15443 ( .B1(n13154), .B2(n13289), .A(n13153), .ZN(n13155) );
  AOI21_X1 U15444 ( .B1(n13318), .B2(n13156), .A(n13155), .ZN(n13157) );
  OAI21_X1 U15445 ( .B1(n13321), .B2(n15625), .A(n13157), .ZN(P3_U3210) );
  XNOR2_X1 U15446 ( .A(n13159), .B(n13158), .ZN(n13160) );
  OAI222_X1 U15447 ( .A1(n15590), .A2(n13162), .B1(n15588), .B2(n13161), .C1(
        n15594), .C2(n13160), .ZN(n13324) );
  INV_X1 U15448 ( .A(n13324), .ZN(n13170) );
  XNOR2_X1 U15449 ( .A(n13164), .B(n13163), .ZN(n13325) );
  INV_X1 U15450 ( .A(n13165), .ZN(n13389) );
  AOI22_X1 U15451 ( .A1(n15576), .A2(n13166), .B1(n15625), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13167) );
  OAI21_X1 U15452 ( .B1(n13389), .B2(n13289), .A(n13167), .ZN(n13168) );
  AOI21_X1 U15453 ( .B1(n13325), .B2(n15535), .A(n13168), .ZN(n13169) );
  OAI21_X1 U15454 ( .B1(n13170), .B2(n15625), .A(n13169), .ZN(P3_U3211) );
  INV_X1 U15455 ( .A(n13171), .ZN(n13172) );
  AOI21_X1 U15456 ( .B1(n13177), .B2(n13173), .A(n13172), .ZN(n13174) );
  OAI222_X1 U15457 ( .A1(n15588), .A2(n13176), .B1(n15590), .B2(n13175), .C1(
        n15594), .C2(n13174), .ZN(n13328) );
  INV_X1 U15458 ( .A(n13328), .ZN(n13184) );
  XOR2_X1 U15459 ( .A(n13178), .B(n13177), .Z(n13329) );
  INV_X1 U15460 ( .A(n13179), .ZN(n13393) );
  AOI22_X1 U15461 ( .A1(n15625), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15576), 
        .B2(n13180), .ZN(n13181) );
  OAI21_X1 U15462 ( .B1(n13393), .B2(n13289), .A(n13181), .ZN(n13182) );
  AOI21_X1 U15463 ( .B1(n13329), .B2(n15535), .A(n13182), .ZN(n13183) );
  OAI21_X1 U15464 ( .B1(n13184), .B2(n15625), .A(n13183), .ZN(P3_U3212) );
  XNOR2_X1 U15465 ( .A(n13185), .B(n13186), .ZN(n13189) );
  AOI222_X1 U15466 ( .A1(n15612), .A2(n13189), .B1(n13188), .B2(n15607), .C1(
        n13187), .C2(n15610), .ZN(n13334) );
  NAND2_X1 U15467 ( .A1(n13191), .A2(n13190), .ZN(n13192) );
  NAND2_X1 U15468 ( .A1(n13193), .A2(n13192), .ZN(n13335) );
  INV_X1 U15469 ( .A(n15535), .ZN(n13231) );
  AOI22_X1 U15470 ( .A1(n15625), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15576), 
        .B2(n13194), .ZN(n13196) );
  INV_X1 U15471 ( .A(n13289), .ZN(n13227) );
  NAND2_X1 U15472 ( .A1(n13332), .A2(n13227), .ZN(n13195) );
  OAI211_X1 U15473 ( .C1(n13335), .C2(n13231), .A(n13196), .B(n13195), .ZN(
        n13197) );
  INV_X1 U15474 ( .A(n13197), .ZN(n13198) );
  OAI21_X1 U15475 ( .B1(n13334), .B2(n15625), .A(n13198), .ZN(P3_U3213) );
  INV_X1 U15476 ( .A(n13199), .ZN(n13202) );
  INV_X1 U15477 ( .A(n13208), .ZN(n13201) );
  OAI211_X1 U15478 ( .C1(n13202), .C2(n13201), .A(n15612), .B(n13200), .ZN(
        n13206) );
  AOI22_X1 U15479 ( .A1(n13204), .A2(n15607), .B1(n15610), .B2(n13203), .ZN(
        n13205) );
  NAND2_X1 U15480 ( .A1(n13206), .A2(n13205), .ZN(n13337) );
  INV_X1 U15481 ( .A(n13337), .ZN(n13213) );
  XOR2_X1 U15482 ( .A(n13207), .B(n13208), .Z(n13338) );
  AOI22_X1 U15483 ( .A1(n15625), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15576), 
        .B2(n13209), .ZN(n13210) );
  OAI21_X1 U15484 ( .B1(n13398), .B2(n13289), .A(n13210), .ZN(n13211) );
  AOI21_X1 U15485 ( .B1(n13338), .B2(n15535), .A(n13211), .ZN(n13212) );
  OAI21_X1 U15486 ( .B1(n13213), .B2(n15625), .A(n13212), .ZN(P3_U3214) );
  NAND2_X1 U15487 ( .A1(n13214), .A2(n8502), .ZN(n13215) );
  INV_X1 U15488 ( .A(n13342), .ZN(n13232) );
  INV_X1 U15489 ( .A(n13217), .ZN(n13218) );
  AOI21_X1 U15490 ( .B1(n13220), .B2(n13219), .A(n13218), .ZN(n13221) );
  OAI222_X1 U15491 ( .A1(n15588), .A2(n13222), .B1(n15590), .B2(n13249), .C1(
        n15594), .C2(n13221), .ZN(n13341) );
  NAND2_X1 U15492 ( .A1(n13341), .A2(n15623), .ZN(n13230) );
  INV_X1 U15493 ( .A(n13223), .ZN(n13224) );
  OAI22_X1 U15494 ( .A1(n15623), .A2(n13225), .B1(n13224), .B2(n15618), .ZN(
        n13226) );
  AOI21_X1 U15495 ( .B1(n13228), .B2(n13227), .A(n13226), .ZN(n13229) );
  OAI211_X1 U15496 ( .C1(n13232), .C2(n13231), .A(n13230), .B(n13229), .ZN(
        P3_U3215) );
  XNOR2_X1 U15497 ( .A(n13233), .B(n13234), .ZN(n13235) );
  OAI222_X1 U15498 ( .A1(n15588), .A2(n13236), .B1(n15590), .B2(n13260), .C1(
        n13235), .C2(n15594), .ZN(n13345) );
  INV_X1 U15499 ( .A(n13345), .ZN(n13245) );
  OAI21_X1 U15500 ( .B1(n13239), .B2(n13238), .A(n13237), .ZN(n13346) );
  INV_X1 U15501 ( .A(n13240), .ZN(n13406) );
  AOI22_X1 U15502 ( .A1(n15625), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15576), 
        .B2(n13241), .ZN(n13242) );
  OAI21_X1 U15503 ( .B1(n13406), .B2(n13289), .A(n13242), .ZN(n13243) );
  AOI21_X1 U15504 ( .B1(n13346), .B2(n15535), .A(n13243), .ZN(n13244) );
  OAI21_X1 U15505 ( .B1(n13245), .B2(n15625), .A(n13244), .ZN(P3_U3216) );
  XNOR2_X1 U15506 ( .A(n13246), .B(n13247), .ZN(n13248) );
  OAI222_X1 U15507 ( .A1(n15588), .A2(n13249), .B1(n15590), .B2(n13275), .C1(
        n13248), .C2(n15594), .ZN(n13349) );
  INV_X1 U15508 ( .A(n13349), .ZN(n13256) );
  XNOR2_X1 U15509 ( .A(n13251), .B(n13250), .ZN(n13350) );
  AOI22_X1 U15510 ( .A1(n15625), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15576), 
        .B2(n13252), .ZN(n13253) );
  OAI21_X1 U15511 ( .B1(n13410), .B2(n13289), .A(n13253), .ZN(n13254) );
  AOI21_X1 U15512 ( .B1(n13350), .B2(n15535), .A(n13254), .ZN(n13255) );
  OAI21_X1 U15513 ( .B1(n13256), .B2(n15625), .A(n13255), .ZN(P3_U3217) );
  XNOR2_X1 U15514 ( .A(n13257), .B(n13258), .ZN(n13259) );
  OAI222_X1 U15515 ( .A1(n15588), .A2(n13260), .B1(n15590), .B2(n13286), .C1(
        n13259), .C2(n15594), .ZN(n13353) );
  INV_X1 U15516 ( .A(n13353), .ZN(n13269) );
  OAI21_X1 U15517 ( .B1(n13263), .B2(n13262), .A(n13261), .ZN(n13354) );
  INV_X1 U15518 ( .A(n13264), .ZN(n13414) );
  AOI22_X1 U15519 ( .A1(n15625), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15576), 
        .B2(n13265), .ZN(n13266) );
  OAI21_X1 U15520 ( .B1(n13414), .B2(n13289), .A(n13266), .ZN(n13267) );
  AOI21_X1 U15521 ( .B1(n13354), .B2(n15535), .A(n13267), .ZN(n13268) );
  OAI21_X1 U15522 ( .B1(n13269), .B2(n15625), .A(n13268), .ZN(P3_U3218) );
  NAND2_X1 U15523 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  XNOR2_X1 U15524 ( .A(n13272), .B(n13276), .ZN(n13273) );
  OAI222_X1 U15525 ( .A1(n15588), .A2(n13275), .B1(n15590), .B2(n13274), .C1(
        n13273), .C2(n15594), .ZN(n13357) );
  INV_X1 U15526 ( .A(n13357), .ZN(n13282) );
  XNOR2_X1 U15527 ( .A(n13277), .B(n13276), .ZN(n13358) );
  AOI22_X1 U15528 ( .A1(n15625), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15576), 
        .B2(n13278), .ZN(n13279) );
  OAI21_X1 U15529 ( .B1(n13418), .B2(n13289), .A(n13279), .ZN(n13280) );
  AOI21_X1 U15530 ( .B1(n13358), .B2(n15535), .A(n13280), .ZN(n13281) );
  OAI21_X1 U15531 ( .B1(n13282), .B2(n15625), .A(n13281), .ZN(P3_U3219) );
  XNOR2_X1 U15532 ( .A(n13284), .B(n13283), .ZN(n13285) );
  OAI222_X1 U15533 ( .A1(n15588), .A2(n13286), .B1(n15590), .B2(n14863), .C1(
        n13285), .C2(n15594), .ZN(n13361) );
  INV_X1 U15534 ( .A(n13361), .ZN(n13295) );
  XNOR2_X1 U15535 ( .A(n13287), .B(n13288), .ZN(n13362) );
  NOR2_X1 U15536 ( .A1(n13422), .A2(n13289), .ZN(n13293) );
  OAI22_X1 U15537 ( .A1(n15623), .A2(n13291), .B1(n13290), .B2(n15618), .ZN(
        n13292) );
  AOI211_X1 U15538 ( .C1(n13362), .C2(n15535), .A(n13293), .B(n13292), .ZN(
        n13294) );
  OAI21_X1 U15539 ( .B1(n13295), .B2(n15625), .A(n13294), .ZN(P3_U3220) );
  NOR2_X1 U15540 ( .A1(n13366), .A2(n8704), .ZN(n13298) );
  AOI21_X1 U15541 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n8704), .A(n13298), .ZN(
        n13296) );
  OAI21_X1 U15542 ( .B1(n13297), .B2(n13364), .A(n13296), .ZN(P3_U3490) );
  AOI21_X1 U15543 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n8704), .A(n13298), .ZN(
        n13299) );
  OAI21_X1 U15544 ( .B1(n13369), .B2(n13364), .A(n13299), .ZN(P3_U3489) );
  INV_X1 U15545 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13302) );
  INV_X1 U15546 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U15547 ( .A1(n13307), .A2(n15662), .B1(n15583), .B2(n13306), .ZN(
        n13308) );
  NAND2_X1 U15548 ( .A1(n13309), .A2(n13308), .ZN(n13379) );
  MUX2_X1 U15549 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13379), .S(n15685), .Z(
        P3_U3485) );
  INV_X1 U15550 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13312) );
  AOI21_X1 U15551 ( .B1(n15662), .B2(n13311), .A(n13310), .ZN(n13380) );
  MUX2_X1 U15552 ( .A(n13312), .B(n13380), .S(n15685), .Z(n13313) );
  OAI21_X1 U15553 ( .B1(n13383), .B2(n13364), .A(n13313), .ZN(P3_U3484) );
  AOI22_X1 U15554 ( .A1(n13315), .A2(n15662), .B1(n15583), .B2(n13314), .ZN(
        n13316) );
  NAND2_X1 U15555 ( .A1(n13317), .A2(n13316), .ZN(n13384) );
  MUX2_X1 U15556 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13384), .S(n15685), .Z(
        P3_U3483) );
  INV_X1 U15557 ( .A(n13318), .ZN(n13323) );
  INV_X1 U15558 ( .A(n15662), .ZN(n13322) );
  NAND2_X1 U15559 ( .A1(n13319), .A2(n15583), .ZN(n13320) );
  OAI211_X1 U15560 ( .C1(n13323), .C2(n13322), .A(n13321), .B(n13320), .ZN(
        n13385) );
  MUX2_X1 U15561 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13385), .S(n15685), .Z(
        P3_U3482) );
  INV_X1 U15562 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13326) );
  AOI21_X1 U15563 ( .B1(n15669), .B2(n13325), .A(n13324), .ZN(n13386) );
  MUX2_X1 U15564 ( .A(n13326), .B(n13386), .S(n15685), .Z(n13327) );
  OAI21_X1 U15565 ( .B1(n13389), .B2(n13364), .A(n13327), .ZN(P3_U3481) );
  INV_X1 U15566 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13330) );
  AOI21_X1 U15567 ( .B1(n15669), .B2(n13329), .A(n13328), .ZN(n13390) );
  MUX2_X1 U15568 ( .A(n13330), .B(n13390), .S(n15685), .Z(n13331) );
  OAI21_X1 U15569 ( .B1(n13393), .B2(n13364), .A(n13331), .ZN(P3_U3480) );
  INV_X1 U15570 ( .A(n15669), .ZN(n13336) );
  NAND2_X1 U15571 ( .A1(n13332), .A2(n15583), .ZN(n13333) );
  OAI211_X1 U15572 ( .C1(n13336), .C2(n13335), .A(n13334), .B(n13333), .ZN(
        n13394) );
  MUX2_X1 U15573 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13394), .S(n15685), .Z(
        P3_U3479) );
  AOI21_X1 U15574 ( .B1(n15669), .B2(n13338), .A(n13337), .ZN(n13395) );
  MUX2_X1 U15575 ( .A(n13339), .B(n13395), .S(n15685), .Z(n13340) );
  OAI21_X1 U15576 ( .B1(n13398), .B2(n13364), .A(n13340), .ZN(P3_U3478) );
  AOI21_X1 U15577 ( .B1(n13342), .B2(n15669), .A(n13341), .ZN(n13399) );
  MUX2_X1 U15578 ( .A(n13343), .B(n13399), .S(n15685), .Z(n13344) );
  OAI21_X1 U15579 ( .B1(n13402), .B2(n13364), .A(n13344), .ZN(P3_U3477) );
  AOI21_X1 U15580 ( .B1(n15669), .B2(n13346), .A(n13345), .ZN(n13403) );
  MUX2_X1 U15581 ( .A(n13347), .B(n13403), .S(n15685), .Z(n13348) );
  OAI21_X1 U15582 ( .B1(n13406), .B2(n13364), .A(n13348), .ZN(P3_U3476) );
  AOI21_X1 U15583 ( .B1(n13350), .B2(n15669), .A(n13349), .ZN(n13407) );
  MUX2_X1 U15584 ( .A(n13351), .B(n13407), .S(n15685), .Z(n13352) );
  OAI21_X1 U15585 ( .B1(n13410), .B2(n13364), .A(n13352), .ZN(P3_U3475) );
  INV_X1 U15586 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13355) );
  AOI21_X1 U15587 ( .B1(n15669), .B2(n13354), .A(n13353), .ZN(n13411) );
  MUX2_X1 U15588 ( .A(n13355), .B(n13411), .S(n15685), .Z(n13356) );
  OAI21_X1 U15589 ( .B1(n13414), .B2(n13364), .A(n13356), .ZN(P3_U3474) );
  INV_X1 U15590 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13359) );
  AOI21_X1 U15591 ( .B1(n15669), .B2(n13358), .A(n13357), .ZN(n13415) );
  MUX2_X1 U15592 ( .A(n13359), .B(n13415), .S(n15685), .Z(n13360) );
  OAI21_X1 U15593 ( .B1(n13364), .B2(n13418), .A(n13360), .ZN(P3_U3473) );
  AOI21_X1 U15594 ( .B1(n13362), .B2(n15669), .A(n13361), .ZN(n13419) );
  MUX2_X1 U15595 ( .A(n8416), .B(n13419), .S(n15685), .Z(n13363) );
  OAI21_X1 U15596 ( .B1(n13364), .B2(n13422), .A(n13363), .ZN(P3_U3472) );
  NAND2_X1 U15597 ( .A1(n13365), .A2(n8719), .ZN(n13368) );
  INV_X1 U15598 ( .A(n13366), .ZN(n13367) );
  NAND2_X1 U15599 ( .A1(n13367), .A2(n15670), .ZN(n13371) );
  OAI211_X1 U15600 ( .C1(n10879), .C2(n15670), .A(n13368), .B(n13371), .ZN(
        P3_U3458) );
  INV_X1 U15601 ( .A(n13369), .ZN(n13370) );
  NAND2_X1 U15602 ( .A1(n13370), .A2(n8719), .ZN(n13372) );
  OAI211_X1 U15603 ( .C1(n8642), .C2(n15670), .A(n13372), .B(n13371), .ZN(
        P3_U3457) );
  MUX2_X1 U15604 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13379), .S(n15670), .Z(
        P3_U3453) );
  MUX2_X1 U15605 ( .A(n13381), .B(n13380), .S(n15670), .Z(n13382) );
  OAI21_X1 U15606 ( .B1(n13383), .B2(n13423), .A(n13382), .ZN(P3_U3452) );
  MUX2_X1 U15607 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13384), .S(n15670), .Z(
        P3_U3451) );
  MUX2_X1 U15608 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13385), .S(n15670), .Z(
        P3_U3450) );
  MUX2_X1 U15609 ( .A(n13387), .B(n13386), .S(n15670), .Z(n13388) );
  OAI21_X1 U15610 ( .B1(n13389), .B2(n13423), .A(n13388), .ZN(P3_U3449) );
  INV_X1 U15611 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13391) );
  MUX2_X1 U15612 ( .A(n13391), .B(n13390), .S(n15670), .Z(n13392) );
  OAI21_X1 U15613 ( .B1(n13393), .B2(n13423), .A(n13392), .ZN(P3_U3448) );
  MUX2_X1 U15614 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13394), .S(n15670), .Z(
        P3_U3447) );
  INV_X1 U15615 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13396) );
  MUX2_X1 U15616 ( .A(n13396), .B(n13395), .S(n15670), .Z(n13397) );
  OAI21_X1 U15617 ( .B1(n13398), .B2(n13423), .A(n13397), .ZN(P3_U3446) );
  MUX2_X1 U15618 ( .A(n13400), .B(n13399), .S(n15670), .Z(n13401) );
  OAI21_X1 U15619 ( .B1(n13402), .B2(n13423), .A(n13401), .ZN(P3_U3444) );
  MUX2_X1 U15620 ( .A(n13404), .B(n13403), .S(n15670), .Z(n13405) );
  OAI21_X1 U15621 ( .B1(n13406), .B2(n13423), .A(n13405), .ZN(P3_U3441) );
  INV_X1 U15622 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13408) );
  MUX2_X1 U15623 ( .A(n13408), .B(n13407), .S(n15670), .Z(n13409) );
  OAI21_X1 U15624 ( .B1(n13410), .B2(n13423), .A(n13409), .ZN(P3_U3438) );
  MUX2_X1 U15625 ( .A(n13412), .B(n13411), .S(n15670), .Z(n13413) );
  OAI21_X1 U15626 ( .B1(n13414), .B2(n13423), .A(n13413), .ZN(P3_U3435) );
  MUX2_X1 U15627 ( .A(n13416), .B(n13415), .S(n15670), .Z(n13417) );
  OAI21_X1 U15628 ( .B1(n13423), .B2(n13418), .A(n13417), .ZN(P3_U3432) );
  INV_X1 U15629 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13420) );
  MUX2_X1 U15630 ( .A(n13420), .B(n13419), .S(n15670), .Z(n13421) );
  OAI21_X1 U15631 ( .B1(n13423), .B2(n13422), .A(n13421), .ZN(P3_U3429) );
  MUX2_X1 U15632 ( .A(P3_D_REG_1__SCAN_IN), .B(n13424), .S(n13426), .Z(
        P3_U3377) );
  INV_X1 U15633 ( .A(n13425), .ZN(n13427) );
  MUX2_X1 U15634 ( .A(P3_D_REG_0__SCAN_IN), .B(n13427), .S(n13426), .Z(
        P3_U3376) );
  NAND3_X1 U15635 ( .A1(n13429), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13432) );
  OAI22_X1 U15636 ( .A1(n13428), .A2(n13432), .B1(n13431), .B2(n13430), .ZN(
        n13433) );
  INV_X1 U15637 ( .A(n13433), .ZN(n13434) );
  OAI21_X1 U15638 ( .B1(n13435), .B2(n13439), .A(n13434), .ZN(P3_U3264) );
  INV_X1 U15639 ( .A(n13436), .ZN(n13438) );
  OAI222_X1 U15640 ( .A1(n13441), .A2(n13440), .B1(n13439), .B2(n13438), .C1(
        n13437), .C2(n6665), .ZN(P3_U3266) );
  MUX2_X1 U15641 ( .A(n13442), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15642 ( .B1(n13443), .B2(n13444), .A(n13630), .ZN(n13446) );
  NAND2_X1 U15643 ( .A1(n13446), .A2(n13445), .ZN(n13455) );
  OAI22_X1 U15644 ( .A1(n13450), .A2(n13449), .B1(n13448), .B2(n13447), .ZN(
        n13772) );
  INV_X1 U15645 ( .A(n13779), .ZN(n13452) );
  OAI22_X1 U15646 ( .A1(n13452), .A2(n13638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13451), .ZN(n13453) );
  AOI21_X1 U15647 ( .B1(n13772), .B2(n13641), .A(n13453), .ZN(n13454) );
  OAI211_X1 U15648 ( .C1(n13456), .C2(n13644), .A(n13455), .B(n13454), .ZN(
        P2_U3186) );
  INV_X1 U15649 ( .A(n13457), .ZN(n13458) );
  AOI21_X1 U15650 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(n13466) );
  NAND2_X1 U15651 ( .A1(n13610), .A2(n13660), .ZN(n13462) );
  NAND2_X1 U15652 ( .A1(n13551), .A2(n13662), .ZN(n13461) );
  AND2_X1 U15653 ( .A1(n13462), .A2(n13461), .ZN(n14880) );
  AOI22_X1 U15654 ( .A1(n13588), .A2(n14884), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13463) );
  OAI21_X1 U15655 ( .B1(n14880), .B2(n13624), .A(n13463), .ZN(n13464) );
  AOI21_X1 U15656 ( .B1(n14889), .B2(n13628), .A(n13464), .ZN(n13465) );
  OAI21_X1 U15657 ( .B1(n13466), .B2(n13630), .A(n13465), .ZN(P2_U3187) );
  INV_X1 U15658 ( .A(n13467), .ZN(n13592) );
  NOR2_X1 U15659 ( .A1(n13592), .A2(n13591), .ZN(n13590) );
  NOR2_X1 U15660 ( .A1(n13590), .A2(n13468), .ZN(n13470) );
  XNOR2_X1 U15661 ( .A(n13470), .B(n13469), .ZN(n13472) );
  AOI21_X1 U15662 ( .B1(n13472), .B2(n13473), .A(n13630), .ZN(n13471) );
  OAI21_X1 U15663 ( .B1(n13473), .B2(n13472), .A(n13471), .ZN(n13480) );
  NAND2_X1 U15664 ( .A1(n13651), .A2(n13610), .ZN(n13475) );
  NAND2_X1 U15665 ( .A1(n13653), .A2(n13622), .ZN(n13474) );
  NAND2_X1 U15666 ( .A1(n13475), .A2(n13474), .ZN(n13839) );
  INV_X1 U15667 ( .A(n13476), .ZN(n13845) );
  OAI22_X1 U15668 ( .A1(n13638), .A2(n13845), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13477), .ZN(n13478) );
  AOI21_X1 U15669 ( .B1(n13839), .B2(n13641), .A(n13478), .ZN(n13479) );
  OAI211_X1 U15670 ( .C1(n7361), .C2(n13644), .A(n13480), .B(n13479), .ZN(
        P2_U3188) );
  OAI21_X1 U15671 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(n13484) );
  NAND2_X1 U15672 ( .A1(n13484), .A2(n13632), .ZN(n13490) );
  NAND2_X1 U15673 ( .A1(n13655), .A2(n13610), .ZN(n13486) );
  NAND2_X1 U15674 ( .A1(n13551), .A2(n13657), .ZN(n13485) );
  NAND2_X1 U15675 ( .A1(n13486), .A2(n13485), .ZN(n13901) );
  INV_X1 U15676 ( .A(n13487), .ZN(n13905) );
  NAND2_X1 U15677 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13729)
         );
  OAI21_X1 U15678 ( .B1(n13638), .B2(n13905), .A(n13729), .ZN(n13488) );
  AOI21_X1 U15679 ( .B1(n13641), .B2(n13901), .A(n13488), .ZN(n13489) );
  OAI211_X1 U15680 ( .C1(n14072), .C2(n13644), .A(n13490), .B(n13489), .ZN(
        P2_U3191) );
  NAND2_X1 U15681 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  XNOR2_X1 U15682 ( .A(n13491), .B(n13494), .ZN(n13495) );
  NAND2_X1 U15683 ( .A1(n13495), .A2(n13632), .ZN(n13503) );
  AOI21_X1 U15684 ( .B1(n13588), .B2(n13497), .A(n13496), .ZN(n13502) );
  NAND2_X1 U15685 ( .A1(n13628), .A2(n13498), .ZN(n13501) );
  NAND2_X1 U15686 ( .A1(n13641), .A2(n13499), .ZN(n13500) );
  NAND4_X1 U15687 ( .A1(n13503), .A2(n13502), .A3(n13501), .A4(n13500), .ZN(
        P2_U3193) );
  AOI21_X1 U15688 ( .B1(n13504), .B2(n13505), .A(n13630), .ZN(n13507) );
  NAND2_X1 U15689 ( .A1(n13507), .A2(n13506), .ZN(n13513) );
  NAND2_X1 U15690 ( .A1(n13653), .A2(n13610), .ZN(n13509) );
  NAND2_X1 U15691 ( .A1(n13655), .A2(n13622), .ZN(n13508) );
  NAND2_X1 U15692 ( .A1(n13509), .A2(n13508), .ZN(n13869) );
  OAI22_X1 U15693 ( .A1(n13638), .A2(n13875), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13510), .ZN(n13511) );
  AOI21_X1 U15694 ( .B1(n13641), .B2(n13869), .A(n13511), .ZN(n13512) );
  OAI211_X1 U15695 ( .C1(n7358), .C2(n13644), .A(n13513), .B(n13512), .ZN(
        P2_U3195) );
  OAI21_X1 U15696 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13517) );
  NAND2_X1 U15697 ( .A1(n13517), .A2(n13632), .ZN(n13523) );
  INV_X1 U15698 ( .A(n13518), .ZN(n13519) );
  OAI22_X1 U15699 ( .A1(n13638), .A2(n13519), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9361), .ZN(n13520) );
  AOI21_X1 U15700 ( .B1(n13641), .B2(n13521), .A(n13520), .ZN(n13522) );
  OAI211_X1 U15701 ( .C1(n14916), .C2(n13644), .A(n13523), .B(n13522), .ZN(
        P2_U3196) );
  OAI211_X1 U15702 ( .C1(n13524), .C2(n13526), .A(n13525), .B(n13632), .ZN(
        n13532) );
  NAND2_X1 U15703 ( .A1(n13649), .A2(n13610), .ZN(n13528) );
  NAND2_X1 U15704 ( .A1(n13651), .A2(n13622), .ZN(n13527) );
  NAND2_X1 U15705 ( .A1(n13528), .A2(n13527), .ZN(n13802) );
  OAI22_X1 U15706 ( .A1(n13809), .A2(n13638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13529), .ZN(n13530) );
  AOI21_X1 U15707 ( .B1(n13802), .B2(n13641), .A(n13530), .ZN(n13531) );
  OAI211_X1 U15708 ( .C1(n14059), .C2(n13644), .A(n13532), .B(n13531), .ZN(
        P2_U3197) );
  INV_X1 U15709 ( .A(n13959), .ZN(n14082) );
  OAI21_X1 U15710 ( .B1(n13535), .B2(n13534), .A(n13533), .ZN(n13536) );
  NAND2_X1 U15711 ( .A1(n13536), .A2(n13632), .ZN(n13543) );
  NAND2_X1 U15712 ( .A1(n13610), .A2(n13658), .ZN(n13538) );
  NAND2_X1 U15713 ( .A1(n13551), .A2(n13660), .ZN(n13537) );
  NAND2_X1 U15714 ( .A1(n13538), .A2(n13537), .ZN(n13949) );
  INV_X1 U15715 ( .A(n13539), .ZN(n13956) );
  OAI22_X1 U15716 ( .A1(n13638), .A2(n13956), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13540), .ZN(n13541) );
  AOI21_X1 U15717 ( .B1(n13641), .B2(n13949), .A(n13541), .ZN(n13542) );
  OAI211_X1 U15718 ( .C1(n14082), .C2(n13644), .A(n13543), .B(n13542), .ZN(
        P2_U3198) );
  INV_X1 U15719 ( .A(n13533), .ZN(n13547) );
  INV_X1 U15720 ( .A(n13544), .ZN(n13546) );
  NOR3_X1 U15721 ( .A1(n13547), .A2(n13546), .A3(n13545), .ZN(n13550) );
  INV_X1 U15722 ( .A(n13548), .ZN(n13549) );
  OAI21_X1 U15723 ( .B1(n13550), .B2(n13549), .A(n13632), .ZN(n13557) );
  NAND2_X1 U15724 ( .A1(n13610), .A2(n13657), .ZN(n13553) );
  NAND2_X1 U15725 ( .A1(n13551), .A2(n13659), .ZN(n13552) );
  NAND2_X1 U15726 ( .A1(n13553), .A2(n13552), .ZN(n13928) );
  INV_X1 U15727 ( .A(n13935), .ZN(n13554) );
  OAI22_X1 U15728 ( .A1(n13638), .A2(n13554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15297), .ZN(n13555) );
  AOI21_X1 U15729 ( .B1(n13641), .B2(n13928), .A(n13555), .ZN(n13556) );
  OAI211_X1 U15730 ( .C1(n14077), .C2(n13644), .A(n13557), .B(n13556), .ZN(
        P2_U3200) );
  INV_X1 U15731 ( .A(n13524), .ZN(n13564) );
  INV_X1 U15732 ( .A(n13558), .ZN(n13560) );
  NAND2_X1 U15733 ( .A1(n13560), .A2(n13559), .ZN(n13562) );
  AOI22_X1 U15734 ( .A1(n13564), .A2(n13563), .B1(n13562), .B2(n13561), .ZN(
        n13569) );
  AOI22_X1 U15735 ( .A1(n13650), .A2(n13610), .B1(n13622), .B2(n13652), .ZN(
        n13819) );
  INV_X1 U15736 ( .A(n13565), .ZN(n13828) );
  AOI22_X1 U15737 ( .A1(n13828), .A2(n13588), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13566) );
  OAI21_X1 U15738 ( .B1(n13819), .B2(n13624), .A(n13566), .ZN(n13567) );
  AOI21_X1 U15739 ( .B1(n13996), .B2(n13628), .A(n13567), .ZN(n13568) );
  OAI21_X1 U15740 ( .B1(n13569), .B2(n13630), .A(n13568), .ZN(P2_U3201) );
  XOR2_X1 U15741 ( .A(n13571), .B(n13570), .Z(n13576) );
  AOI22_X1 U15742 ( .A1(n13654), .A2(n13610), .B1(n13622), .B2(n13656), .ZN(
        n13886) );
  INV_X1 U15743 ( .A(n13891), .ZN(n13572) );
  AOI22_X1 U15744 ( .A1(n13588), .A2(n13572), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13573) );
  OAI21_X1 U15745 ( .B1(n13886), .B2(n13624), .A(n13573), .ZN(n13574) );
  AOI21_X1 U15746 ( .B1(n14022), .B2(n13628), .A(n13574), .ZN(n13575) );
  OAI21_X1 U15747 ( .B1(n13576), .B2(n13630), .A(n13575), .ZN(P2_U3205) );
  OAI211_X1 U15748 ( .C1(n13579), .C2(n13578), .A(n13577), .B(n13632), .ZN(
        n13586) );
  INV_X1 U15749 ( .A(n13580), .ZN(n13582) );
  OAI21_X1 U15750 ( .B1(n13638), .B2(n13582), .A(n13581), .ZN(n13583) );
  AOI21_X1 U15751 ( .B1(n13641), .B2(n13584), .A(n13583), .ZN(n13585) );
  OAI211_X1 U15752 ( .C1(n14910), .C2(n13644), .A(n13586), .B(n13585), .ZN(
        P2_U3206) );
  AOI22_X1 U15753 ( .A1(n13652), .A2(n13610), .B1(n13622), .B2(n13654), .ZN(
        n13851) );
  INV_X1 U15754 ( .A(n13858), .ZN(n13587) );
  AOI22_X1 U15755 ( .A1(n13588), .A2(n13587), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13589) );
  OAI21_X1 U15756 ( .B1(n13851), .B2(n13624), .A(n13589), .ZN(n13594) );
  AOI211_X1 U15757 ( .C1(n13592), .C2(n13591), .A(n13630), .B(n13590), .ZN(
        n13593) );
  AOI211_X1 U15758 ( .C1(n14010), .C2(n13628), .A(n13594), .B(n13593), .ZN(
        n13595) );
  INV_X1 U15759 ( .A(n13595), .ZN(P2_U3207) );
  OAI211_X1 U15760 ( .C1(n13598), .C2(n13597), .A(n13596), .B(n13632), .ZN(
        n13605) );
  INV_X1 U15761 ( .A(n13599), .ZN(n13601) );
  OAI22_X1 U15762 ( .A1(n13638), .A2(n13601), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13600), .ZN(n13602) );
  AOI21_X1 U15763 ( .B1(n13641), .B2(n13603), .A(n13602), .ZN(n13604) );
  OAI211_X1 U15764 ( .C1(n15410), .C2(n13644), .A(n13605), .B(n13604), .ZN(
        P2_U3208) );
  INV_X1 U15765 ( .A(n14031), .ZN(n13919) );
  AOI21_X1 U15766 ( .B1(n13607), .B2(n13606), .A(n13630), .ZN(n13609) );
  NAND2_X1 U15767 ( .A1(n13609), .A2(n13608), .ZN(n13617) );
  NAND2_X1 U15768 ( .A1(n13622), .A2(n13658), .ZN(n13612) );
  NAND2_X1 U15769 ( .A1(n13610), .A2(n13656), .ZN(n13611) );
  NAND2_X1 U15770 ( .A1(n13612), .A2(n13611), .ZN(n13913) );
  INV_X1 U15771 ( .A(n13916), .ZN(n13614) );
  OAI22_X1 U15772 ( .A1(n13638), .A2(n13614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13613), .ZN(n13615) );
  AOI21_X1 U15773 ( .B1(n13641), .B2(n13913), .A(n13615), .ZN(n13616) );
  OAI211_X1 U15774 ( .C1(n13919), .C2(n13644), .A(n13617), .B(n13616), .ZN(
        P2_U3210) );
  INV_X1 U15775 ( .A(n13618), .ZN(n13619) );
  AOI21_X1 U15776 ( .B1(n13621), .B2(n13620), .A(n13619), .ZN(n13631) );
  AND2_X1 U15777 ( .A1(n13650), .A2(n13622), .ZN(n13623) );
  AOI21_X1 U15778 ( .B1(n13648), .B2(n13610), .A(n13623), .ZN(n13793) );
  NOR2_X1 U15779 ( .A1(n13793), .A2(n13624), .ZN(n13627) );
  OAI22_X1 U15780 ( .A1(n13789), .A2(n13638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13625), .ZN(n13626) );
  AOI211_X1 U15781 ( .C1(n13986), .C2(n13628), .A(n13627), .B(n13626), .ZN(
        n13629) );
  OAI21_X1 U15782 ( .B1(n13631), .B2(n13630), .A(n13629), .ZN(P2_U3212) );
  OAI211_X1 U15783 ( .C1(n13635), .C2(n13634), .A(n13633), .B(n13632), .ZN(
        n13643) );
  INV_X1 U15784 ( .A(n13636), .ZN(n13637) );
  NAND2_X1 U15785 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15295)
         );
  OAI21_X1 U15786 ( .B1(n13638), .B2(n13637), .A(n15295), .ZN(n13639) );
  AOI21_X1 U15787 ( .B1(n13641), .B2(n13640), .A(n13639), .ZN(n13642) );
  OAI211_X1 U15788 ( .C1(n14899), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        P2_U3213) );
  MUX2_X1 U15789 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13645), .S(n6675), .Z(
        P2_U3562) );
  MUX2_X1 U15790 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13646), .S(n6675), .Z(
        P2_U3561) );
  MUX2_X1 U15791 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13647), .S(n6675), .Z(
        P2_U3560) );
  MUX2_X1 U15792 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9494), .S(n6675), .Z(
        P2_U3559) );
  MUX2_X1 U15793 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13648), .S(n6675), .Z(
        P2_U3558) );
  MUX2_X1 U15794 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13649), .S(n6675), .Z(
        P2_U3557) );
  MUX2_X1 U15795 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13650), .S(n6675), .Z(
        P2_U3556) );
  MUX2_X1 U15796 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13651), .S(n6675), .Z(
        P2_U3555) );
  MUX2_X1 U15797 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13652), .S(n6675), .Z(
        P2_U3554) );
  MUX2_X1 U15798 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13653), .S(n6675), .Z(
        P2_U3553) );
  MUX2_X1 U15799 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13654), .S(n6675), .Z(
        P2_U3552) );
  MUX2_X1 U15800 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13655), .S(n6675), .Z(
        P2_U3551) );
  MUX2_X1 U15801 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13656), .S(n6675), .Z(
        P2_U3550) );
  MUX2_X1 U15802 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13657), .S(n6675), .Z(
        P2_U3549) );
  MUX2_X1 U15803 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13658), .S(n6675), .Z(
        P2_U3548) );
  MUX2_X1 U15804 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13659), .S(n6675), .Z(
        P2_U3547) );
  MUX2_X1 U15805 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13660), .S(n6675), .Z(
        P2_U3546) );
  MUX2_X1 U15806 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13661), .S(n6675), .Z(
        P2_U3545) );
  MUX2_X1 U15807 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13662), .S(n6675), .Z(
        P2_U3544) );
  MUX2_X1 U15808 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13663), .S(n6675), .Z(
        P2_U3543) );
  MUX2_X1 U15809 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13664), .S(n6675), .Z(
        P2_U3542) );
  MUX2_X1 U15810 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13665), .S(n6675), .Z(
        P2_U3541) );
  MUX2_X1 U15811 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13666), .S(n6675), .Z(
        P2_U3540) );
  MUX2_X1 U15812 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13667), .S(n6675), .Z(
        P2_U3539) );
  MUX2_X1 U15813 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13668), .S(n6675), .Z(
        P2_U3538) );
  MUX2_X1 U15814 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13669), .S(n6675), .Z(
        P2_U3537) );
  MUX2_X1 U15815 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13670), .S(n6675), .Z(
        P2_U3536) );
  MUX2_X1 U15816 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13671), .S(n6675), .Z(
        P2_U3535) );
  MUX2_X1 U15817 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13672), .S(n6675), .Z(
        P2_U3534) );
  MUX2_X1 U15818 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7040), .S(n6675), .Z(
        P2_U3533) );
  MUX2_X1 U15819 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13674), .S(n6675), .Z(
        P2_U3532) );
  MUX2_X1 U15820 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9756), .S(n6675), .Z(
        P2_U3531) );
  NOR2_X1 U15821 ( .A1(n13676), .A2(n13684), .ZN(n13677) );
  INV_X1 U15822 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15286) );
  NOR2_X1 U15823 ( .A1(n15286), .A2(n15287), .ZN(n15285) );
  NOR2_X1 U15824 ( .A1(n13677), .A2(n15285), .ZN(n13679) );
  XNOR2_X1 U15825 ( .A(n13703), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13678) );
  NOR2_X1 U15826 ( .A1(n13679), .A2(n13678), .ZN(n13702) );
  AOI211_X1 U15827 ( .C1(n13679), .C2(n13678), .A(n13702), .B(n15298), .ZN(
        n13693) );
  NAND2_X1 U15828 ( .A1(n13681), .A2(n13680), .ZN(n13683) );
  NAND2_X1 U15829 ( .A1(n13683), .A2(n13682), .ZN(n13685) );
  NAND2_X1 U15830 ( .A1(n15292), .A2(n13685), .ZN(n13686) );
  XNOR2_X1 U15831 ( .A(n13685), .B(n13684), .ZN(n15291) );
  NAND2_X1 U15832 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15291), .ZN(n15290) );
  NAND2_X1 U15833 ( .A1(n13686), .A2(n15290), .ZN(n13688) );
  INV_X1 U15834 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U15835 ( .A1(n13703), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13696), 
        .B2(n13695), .ZN(n13687) );
  NAND2_X1 U15836 ( .A1(n13687), .A2(n13688), .ZN(n13694) );
  OAI211_X1 U15837 ( .C1(n13688), .C2(n13687), .A(n15307), .B(n13694), .ZN(
        n13691) );
  AND2_X1 U15838 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13689) );
  AOI21_X1 U15839 ( .B1(n15305), .B2(n13703), .A(n13689), .ZN(n13690) );
  OAI211_X1 U15840 ( .C1(n15313), .C2(n7529), .A(n13691), .B(n13690), .ZN(
        n13692) );
  OR2_X1 U15841 ( .A1(n13693), .A2(n13692), .ZN(P2_U3230) );
  INV_X1 U15842 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U15843 ( .A1(n15304), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13698), 
        .B2(n13697), .ZN(n15309) );
  OAI21_X1 U15844 ( .B1(n13696), .B2(n13695), .A(n13694), .ZN(n15308) );
  NAND2_X1 U15845 ( .A1(n15309), .A2(n15308), .ZN(n15306) );
  OAI21_X1 U15846 ( .B1(n13698), .B2(n13697), .A(n15306), .ZN(n13717) );
  XOR2_X1 U15847 ( .A(n13717), .B(n13711), .Z(n13699) );
  NOR2_X1 U15848 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13699), .ZN(n13719) );
  AOI21_X1 U15849 ( .B1(n13699), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13719), 
        .ZN(n13710) );
  AND2_X1 U15850 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13701) );
  NOR2_X1 U15851 ( .A1(n15272), .A2(n13711), .ZN(n13700) );
  AOI211_X1 U15852 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15289), .A(n13701), 
        .B(n13700), .ZN(n13709) );
  XNOR2_X1 U15853 ( .A(n15304), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15300) );
  INV_X1 U15854 ( .A(n13704), .ZN(n13707) );
  INV_X1 U15855 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13705) );
  INV_X1 U15856 ( .A(n13714), .ZN(n13706) );
  OAI211_X1 U15857 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13707), .A(n15265), 
        .B(n13706), .ZN(n13708) );
  OAI211_X1 U15858 ( .C1(n13710), .C2(n15279), .A(n13709), .B(n13708), .ZN(
        P2_U3232) );
  NOR2_X1 U15859 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  NOR2_X1 U15860 ( .A1(n13714), .A2(n13713), .ZN(n13716) );
  INV_X1 U15861 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13715) );
  XOR2_X1 U15862 ( .A(n13716), .B(n13715), .Z(n13725) );
  INV_X1 U15863 ( .A(n13725), .ZN(n13723) );
  NOR2_X1 U15864 ( .A1(n13718), .A2(n13717), .ZN(n13720) );
  NOR2_X1 U15865 ( .A1(n13720), .A2(n13719), .ZN(n13721) );
  XOR2_X1 U15866 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13721), .Z(n13724) );
  OAI21_X1 U15867 ( .B1(n13724), .B2(n15279), .A(n15272), .ZN(n13722) );
  AOI21_X1 U15868 ( .B1(n13723), .B2(n15265), .A(n13722), .ZN(n13728) );
  AOI22_X1 U15869 ( .A1(n13725), .A2(n15265), .B1(n15307), .B2(n13724), .ZN(
        n13727) );
  MUX2_X1 U15870 ( .A(n13728), .B(n13727), .S(n13726), .Z(n13730) );
  OAI211_X1 U15871 ( .C1(n15313), .C2(n13731), .A(n13730), .B(n13729), .ZN(
        P2_U3233) );
  NAND2_X1 U15872 ( .A1(n13732), .A2(n15319), .ZN(n13735) );
  INV_X1 U15873 ( .A(n13733), .ZN(n13967) );
  NOR2_X1 U15874 ( .A1(n13967), .A2(n6674), .ZN(n13740) );
  AOI21_X1 U15875 ( .B1(n6674), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13740), .ZN(
        n13734) );
  OAI211_X1 U15876 ( .C1(n13736), .C2(n13918), .A(n13735), .B(n13734), .ZN(
        P2_U3234) );
  OAI211_X1 U15877 ( .C1(n14050), .C2(n13738), .A(n9576), .B(n13737), .ZN(
        n13968) );
  NOR2_X1 U15878 ( .A1(n13963), .A2(n13739), .ZN(n13741) );
  AOI211_X1 U15879 ( .C1(n13742), .C2(n15314), .A(n13741), .B(n13740), .ZN(
        n13743) );
  OAI21_X1 U15880 ( .B1(n13968), .B2(n13961), .A(n13743), .ZN(P2_U3235) );
  INV_X1 U15881 ( .A(n13744), .ZN(n13754) );
  NAND3_X1 U15882 ( .A1(n13745), .A2(n15316), .A3(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n13747) );
  NAND2_X1 U15883 ( .A1(n6674), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13746) );
  OAI211_X1 U15884 ( .C1(n13748), .C2(n13918), .A(n13747), .B(n13746), .ZN(
        n13749) );
  AOI21_X1 U15885 ( .B1(n13750), .B2(n15319), .A(n13749), .ZN(n13753) );
  NAND2_X1 U15886 ( .A1(n13751), .A2(n13963), .ZN(n13752) );
  OAI211_X1 U15887 ( .C1(n13754), .C2(n13966), .A(n13753), .B(n13752), .ZN(
        P2_U3236) );
  NOR2_X1 U15888 ( .A1(n14053), .A2(n13778), .ZN(n13758) );
  NOR3_X1 U15889 ( .A1(n13759), .A2(n13758), .A3(n14001), .ZN(n13973) );
  AOI22_X1 U15890 ( .A1(n13760), .A2(n15316), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n6674), .ZN(n13761) );
  OAI21_X1 U15891 ( .B1(n14053), .B2(n13918), .A(n13761), .ZN(n13762) );
  AOI21_X1 U15892 ( .B1(n13973), .B2(n15319), .A(n13762), .ZN(n13769) );
  OAI211_X1 U15893 ( .C1(n13765), .C2(n13764), .A(n13763), .B(n14882), .ZN(
        n13767) );
  NAND2_X1 U15894 ( .A1(n13767), .A2(n13766), .ZN(n13972) );
  NAND2_X1 U15895 ( .A1(n13972), .A2(n13963), .ZN(n13768) );
  OAI211_X1 U15896 ( .C1(n13971), .C2(n13966), .A(n13769), .B(n13768), .ZN(
        P2_U3237) );
  XNOR2_X1 U15897 ( .A(n13771), .B(n13770), .ZN(n13773) );
  AOI21_X1 U15898 ( .B1(n13773), .B2(n14882), .A(n13772), .ZN(n13982) );
  OR2_X1 U15899 ( .A1(n13775), .A2(n13774), .ZN(n13978) );
  NAND3_X1 U15900 ( .A1(n13978), .A2(n13977), .A3(n15320), .ZN(n13784) );
  NAND2_X1 U15901 ( .A1(n13980), .A2(n13785), .ZN(n13776) );
  NAND2_X1 U15902 ( .A1(n13776), .A2(n9576), .ZN(n13777) );
  NOR2_X1 U15903 ( .A1(n13778), .A2(n13777), .ZN(n13979) );
  NAND2_X1 U15904 ( .A1(n13980), .A2(n15314), .ZN(n13781) );
  AOI22_X1 U15905 ( .A1(n13779), .A2(n15316), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n6674), .ZN(n13780) );
  NAND2_X1 U15906 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  AOI21_X1 U15907 ( .B1(n13979), .B2(n15319), .A(n13782), .ZN(n13783) );
  OAI211_X1 U15908 ( .C1(n6674), .C2(n13982), .A(n13784), .B(n13783), .ZN(
        P2_U3238) );
  XNOR2_X1 U15909 ( .A(n6792), .B(n13792), .ZN(n13988) );
  INV_X1 U15910 ( .A(n13785), .ZN(n13786) );
  AOI211_X1 U15911 ( .C1(n13986), .C2(n13807), .A(n14001), .B(n13786), .ZN(
        n13985) );
  NOR2_X1 U15912 ( .A1(n13787), .A2(n13918), .ZN(n13791) );
  OAI22_X1 U15913 ( .A1(n13789), .A2(n13957), .B1(n13788), .B2(n13963), .ZN(
        n13790) );
  AOI211_X1 U15914 ( .C1(n13985), .C2(n15319), .A(n13791), .B(n13790), .ZN(
        n13796) );
  XOR2_X1 U15915 ( .A(n13792), .B(n6788), .Z(n13794) );
  OAI21_X1 U15916 ( .B1(n13794), .B2(n13946), .A(n13793), .ZN(n13984) );
  NAND2_X1 U15917 ( .A1(n13984), .A2(n13963), .ZN(n13795) );
  OAI211_X1 U15918 ( .C1(n13988), .C2(n13966), .A(n13796), .B(n13795), .ZN(
        P2_U3239) );
  AND3_X1 U15919 ( .A1(n13797), .A2(n13799), .A3(n13798), .ZN(n13800) );
  OR2_X1 U15920 ( .A1(n13801), .A2(n13800), .ZN(n13803) );
  AOI21_X1 U15921 ( .B1(n13803), .B2(n14882), .A(n13802), .ZN(n13990) );
  AND2_X1 U15922 ( .A1(n13804), .A2(n7556), .ZN(n13805) );
  OR2_X1 U15923 ( .A1(n13806), .A2(n13805), .ZN(n13992) );
  OAI211_X1 U15924 ( .C1(n13827), .C2(n14059), .A(n9576), .B(n13807), .ZN(
        n13989) );
  OAI22_X1 U15925 ( .A1(n13809), .A2(n13957), .B1(n13963), .B2(n13808), .ZN(
        n13810) );
  AOI21_X1 U15926 ( .B1(n13811), .B2(n15314), .A(n13810), .ZN(n13812) );
  OAI21_X1 U15927 ( .B1(n13989), .B2(n13961), .A(n13812), .ZN(n13813) );
  AOI21_X1 U15928 ( .B1(n13992), .B2(n15320), .A(n13813), .ZN(n13814) );
  OAI21_X1 U15929 ( .B1(n6674), .B2(n13990), .A(n13814), .ZN(P2_U3240) );
  INV_X1 U15930 ( .A(n13815), .ZN(n13817) );
  OAI21_X1 U15931 ( .B1(n13817), .B2(n13816), .A(n13823), .ZN(n13818) );
  AOI21_X1 U15932 ( .B1(n13818), .B2(n13797), .A(n13946), .ZN(n13821) );
  INV_X1 U15933 ( .A(n13819), .ZN(n13820) );
  NOR2_X1 U15934 ( .A1(n13821), .A2(n13820), .ZN(n13998) );
  OAI21_X1 U15935 ( .B1(n13824), .B2(n13823), .A(n13822), .ZN(n13999) );
  INV_X1 U15936 ( .A(n13999), .ZN(n13833) );
  INV_X1 U15937 ( .A(n13996), .ZN(n13831) );
  NAND2_X1 U15938 ( .A1(n13844), .A2(n13996), .ZN(n13825) );
  NAND2_X1 U15939 ( .A1(n13825), .A2(n9576), .ZN(n13826) );
  NOR2_X1 U15940 ( .A1(n13827), .A2(n13826), .ZN(n13995) );
  NAND2_X1 U15941 ( .A1(n13995), .A2(n15319), .ZN(n13830) );
  AOI22_X1 U15942 ( .A1(n13828), .A2(n15316), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n6674), .ZN(n13829) );
  OAI211_X1 U15943 ( .C1(n13831), .C2(n13918), .A(n13830), .B(n13829), .ZN(
        n13832) );
  AOI21_X1 U15944 ( .B1(n13833), .B2(n15320), .A(n13832), .ZN(n13834) );
  OAI21_X1 U15945 ( .B1(n6674), .B2(n13998), .A(n13834), .ZN(P2_U3241) );
  XNOR2_X1 U15946 ( .A(n13836), .B(n13835), .ZN(n14000) );
  INV_X1 U15947 ( .A(n14000), .ZN(n13849) );
  AOI22_X1 U15948 ( .A1(n13842), .A2(n15314), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n6674), .ZN(n13848) );
  OAI211_X1 U15949 ( .C1(n13838), .C2(n13837), .A(n13815), .B(n14882), .ZN(
        n13841) );
  INV_X1 U15950 ( .A(n13839), .ZN(n13840) );
  NAND2_X1 U15951 ( .A1(n13841), .A2(n13840), .ZN(n14004) );
  NAND2_X1 U15952 ( .A1(n13842), .A2(n13860), .ZN(n13843) );
  NAND2_X1 U15953 ( .A1(n13844), .A2(n13843), .ZN(n14002) );
  OAI22_X1 U15954 ( .A1(n14002), .A2(n6681), .B1(n13845), .B2(n13957), .ZN(
        n13846) );
  OAI21_X1 U15955 ( .B1(n14004), .B2(n13846), .A(n13963), .ZN(n13847) );
  OAI211_X1 U15956 ( .C1(n13849), .C2(n13966), .A(n13848), .B(n13847), .ZN(
        P2_U3242) );
  INV_X1 U15957 ( .A(n13855), .ZN(n13850) );
  OAI21_X1 U15958 ( .B1(n6700), .B2(n13850), .A(n7275), .ZN(n13853) );
  INV_X1 U15959 ( .A(n13851), .ZN(n13852) );
  AOI21_X1 U15960 ( .B1(n13853), .B2(n14882), .A(n13852), .ZN(n14012) );
  OAI21_X1 U15961 ( .B1(n13856), .B2(n13855), .A(n13854), .ZN(n14013) );
  NAND2_X1 U15962 ( .A1(n6674), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13857) );
  OAI21_X1 U15963 ( .B1(n13957), .B2(n13858), .A(n13857), .ZN(n13859) );
  AOI21_X1 U15964 ( .B1(n14010), .B2(n15314), .A(n13859), .ZN(n13863) );
  AOI21_X1 U15965 ( .B1(n14010), .B2(n13873), .A(n14001), .ZN(n13861) );
  AND2_X1 U15966 ( .A1(n13861), .A2(n13860), .ZN(n14009) );
  NAND2_X1 U15967 ( .A1(n14009), .A2(n15319), .ZN(n13862) );
  OAI211_X1 U15968 ( .C1(n14013), .C2(n13966), .A(n13863), .B(n13862), .ZN(
        n13864) );
  INV_X1 U15969 ( .A(n13864), .ZN(n13865) );
  OAI21_X1 U15970 ( .B1(n6674), .B2(n14012), .A(n13865), .ZN(P2_U3243) );
  OR2_X1 U15971 ( .A1(n13866), .A2(n13885), .ZN(n13883) );
  NAND2_X1 U15972 ( .A1(n13883), .A2(n13867), .ZN(n13868) );
  XNOR2_X1 U15973 ( .A(n13868), .B(n13871), .ZN(n13870) );
  AOI21_X1 U15974 ( .B1(n13870), .B2(n14882), .A(n13869), .ZN(n14017) );
  XNOR2_X1 U15975 ( .A(n13872), .B(n13871), .ZN(n14014) );
  AOI21_X1 U15976 ( .B1(n13877), .B2(n13888), .A(n14001), .ZN(n13874) );
  NAND2_X1 U15977 ( .A1(n13874), .A2(n13873), .ZN(n14015) );
  INV_X1 U15978 ( .A(n13875), .ZN(n13876) );
  AOI22_X1 U15979 ( .A1(n6674), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13876), 
        .B2(n15316), .ZN(n13879) );
  NAND2_X1 U15980 ( .A1(n13877), .A2(n15314), .ZN(n13878) );
  OAI211_X1 U15981 ( .C1(n14015), .C2(n13961), .A(n13879), .B(n13878), .ZN(
        n13880) );
  AOI21_X1 U15982 ( .B1(n14014), .B2(n15320), .A(n13880), .ZN(n13881) );
  OAI21_X1 U15983 ( .B1(n14017), .B2(n6674), .A(n13881), .ZN(P2_U3244) );
  XNOR2_X1 U15984 ( .A(n13882), .B(n13885), .ZN(n14024) );
  INV_X1 U15985 ( .A(n13883), .ZN(n13884) );
  AOI21_X1 U15986 ( .B1(n13866), .B2(n13885), .A(n13884), .ZN(n13887) );
  OAI21_X1 U15987 ( .B1(n13887), .B2(n13946), .A(n13886), .ZN(n14020) );
  AOI21_X1 U15988 ( .B1(n14022), .B2(n13903), .A(n14001), .ZN(n13889) );
  AND2_X1 U15989 ( .A1(n13889), .A2(n13888), .ZN(n14021) );
  NAND2_X1 U15990 ( .A1(n14021), .A2(n15319), .ZN(n13894) );
  NAND2_X1 U15991 ( .A1(n6674), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13890) );
  OAI21_X1 U15992 ( .B1(n13957), .B2(n13891), .A(n13890), .ZN(n13892) );
  AOI21_X1 U15993 ( .B1(n14022), .B2(n15314), .A(n13892), .ZN(n13893) );
  NAND2_X1 U15994 ( .A1(n13894), .A2(n13893), .ZN(n13895) );
  AOI21_X1 U15995 ( .B1(n14020), .B2(n13963), .A(n13895), .ZN(n13896) );
  OAI21_X1 U15996 ( .B1(n13966), .B2(n14024), .A(n13896), .ZN(P2_U3245) );
  INV_X1 U15997 ( .A(n13899), .ZN(n13897) );
  XNOR2_X1 U15998 ( .A(n13898), .B(n13897), .ZN(n14027) );
  XNOR2_X1 U15999 ( .A(n13900), .B(n13899), .ZN(n13902) );
  AOI21_X1 U16000 ( .B1(n13902), .B2(n14882), .A(n13901), .ZN(n14026) );
  INV_X1 U16001 ( .A(n14026), .ZN(n13910) );
  OAI211_X1 U16002 ( .C1(n13915), .C2(n14072), .A(n9576), .B(n13903), .ZN(
        n14025) );
  NAND2_X1 U16003 ( .A1(n6674), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U16004 ( .B1(n13957), .B2(n13905), .A(n13904), .ZN(n13906) );
  AOI21_X1 U16005 ( .B1(n13907), .B2(n15314), .A(n13906), .ZN(n13908) );
  OAI21_X1 U16006 ( .B1(n14025), .B2(n13961), .A(n13908), .ZN(n13909) );
  AOI21_X1 U16007 ( .B1(n13910), .B2(n13963), .A(n13909), .ZN(n13911) );
  OAI21_X1 U16008 ( .B1(n13966), .B2(n14027), .A(n13911), .ZN(P2_U3246) );
  XNOR2_X1 U16009 ( .A(n13912), .B(n13923), .ZN(n13914) );
  AOI21_X1 U16010 ( .B1(n13914), .B2(n14882), .A(n13913), .ZN(n14033) );
  AOI211_X1 U16011 ( .C1(n14031), .C2(n13933), .A(n14001), .B(n13915), .ZN(
        n14030) );
  AOI22_X1 U16012 ( .A1(n6674), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13916), 
        .B2(n15316), .ZN(n13917) );
  OAI21_X1 U16013 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n13925) );
  INV_X1 U16014 ( .A(n13920), .ZN(n13921) );
  AOI21_X1 U16015 ( .B1(n13923), .B2(n13922), .A(n13921), .ZN(n14034) );
  NOR2_X1 U16016 ( .A1(n14034), .A2(n13966), .ZN(n13924) );
  AOI211_X1 U16017 ( .C1(n14030), .C2(n15319), .A(n13925), .B(n13924), .ZN(
        n13926) );
  OAI21_X1 U16018 ( .B1(n6674), .B2(n14033), .A(n13926), .ZN(P2_U3247) );
  XNOR2_X1 U16019 ( .A(n13927), .B(n13931), .ZN(n13929) );
  AOI21_X1 U16020 ( .B1(n13929), .B2(n14882), .A(n13928), .ZN(n14036) );
  OAI21_X1 U16021 ( .B1(n13932), .B2(n13931), .A(n13930), .ZN(n14037) );
  INV_X1 U16022 ( .A(n14037), .ZN(n13940) );
  AOI21_X1 U16023 ( .B1(n13953), .B2(n13936), .A(n14001), .ZN(n13934) );
  NAND2_X1 U16024 ( .A1(n13934), .A2(n13933), .ZN(n14035) );
  AOI22_X1 U16025 ( .A1(n6674), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13935), 
        .B2(n15316), .ZN(n13938) );
  NAND2_X1 U16026 ( .A1(n13936), .A2(n15314), .ZN(n13937) );
  OAI211_X1 U16027 ( .C1(n14035), .C2(n13961), .A(n13938), .B(n13937), .ZN(
        n13939) );
  AOI21_X1 U16028 ( .B1(n13940), .B2(n15320), .A(n13939), .ZN(n13941) );
  OAI21_X1 U16029 ( .B1(n14036), .B2(n6674), .A(n13941), .ZN(P2_U3248) );
  NAND2_X1 U16030 ( .A1(n13943), .A2(n13942), .ZN(n13944) );
  NAND2_X1 U16031 ( .A1(n13945), .A2(n13944), .ZN(n14042) );
  AOI21_X1 U16032 ( .B1(n13948), .B2(n13947), .A(n13946), .ZN(n13951) );
  AOI21_X1 U16033 ( .B1(n13951), .B2(n13950), .A(n13949), .ZN(n14041) );
  INV_X1 U16034 ( .A(n14041), .ZN(n13964) );
  AOI21_X1 U16035 ( .B1(n13952), .B2(n13959), .A(n14001), .ZN(n13954) );
  NAND2_X1 U16036 ( .A1(n13954), .A2(n13953), .ZN(n14040) );
  NAND2_X1 U16037 ( .A1(n6674), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13955) );
  OAI21_X1 U16038 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(n13958) );
  AOI21_X1 U16039 ( .B1(n13959), .B2(n15314), .A(n13958), .ZN(n13960) );
  OAI21_X1 U16040 ( .B1(n14040), .B2(n13961), .A(n13960), .ZN(n13962) );
  AOI21_X1 U16041 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n13965) );
  OAI21_X1 U16042 ( .B1(n13966), .B2(n14042), .A(n13965), .ZN(P2_U3249) );
  INV_X1 U16043 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13969) );
  AND2_X1 U16044 ( .A1(n13968), .A2(n13967), .ZN(n14047) );
  MUX2_X1 U16045 ( .A(n13969), .B(n14047), .S(n15431), .Z(n13970) );
  OAI21_X1 U16046 ( .B1(n14050), .B2(n14046), .A(n13970), .ZN(P2_U3529) );
  INV_X1 U16047 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13975) );
  INV_X1 U16048 ( .A(n13971), .ZN(n13974) );
  OAI21_X1 U16049 ( .B1(n14053), .B2(n14046), .A(n13976), .ZN(P2_U3527) );
  NAND3_X1 U16050 ( .A1(n13978), .A2(n13977), .A3(n15370), .ZN(n13983) );
  AOI21_X1 U16051 ( .B1(n13980), .B2(n15398), .A(n13979), .ZN(n13981) );
  NAND3_X1 U16052 ( .A1(n13983), .A2(n13982), .A3(n13981), .ZN(n14054) );
  MUX2_X1 U16053 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14054), .S(n15431), .Z(
        P2_U3526) );
  AOI211_X1 U16054 ( .C1(n13986), .C2(n15398), .A(n13985), .B(n13984), .ZN(
        n13987) );
  OAI21_X1 U16055 ( .B1(n14043), .B2(n13988), .A(n13987), .ZN(n14055) );
  MUX2_X1 U16056 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14055), .S(n15431), .Z(
        P2_U3525) );
  INV_X1 U16057 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U16058 ( .A1(n13990), .A2(n13989), .ZN(n13991) );
  AOI21_X1 U16059 ( .B1(n13992), .B2(n15370), .A(n13991), .ZN(n14056) );
  MUX2_X1 U16060 ( .A(n13993), .B(n14056), .S(n15431), .Z(n13994) );
  OAI21_X1 U16061 ( .B1(n14059), .B2(n14046), .A(n13994), .ZN(P2_U3524) );
  AOI21_X1 U16062 ( .B1(n13996), .B2(n15398), .A(n13995), .ZN(n13997) );
  OAI211_X1 U16063 ( .C1(n13999), .C2(n14043), .A(n13998), .B(n13997), .ZN(
        n14060) );
  MUX2_X1 U16064 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14060), .S(n15431), .Z(
        P2_U3523) );
  NAND2_X1 U16065 ( .A1(n14000), .A2(n15370), .ZN(n14006) );
  NOR2_X1 U16066 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  NOR2_X1 U16067 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  NAND2_X1 U16068 ( .A1(n14006), .A2(n14005), .ZN(n14061) );
  MUX2_X1 U16069 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14061), .S(n15431), .Z(
        n14007) );
  INV_X1 U16070 ( .A(n14007), .ZN(n14008) );
  OAI21_X1 U16071 ( .B1(n7361), .B2(n14046), .A(n14008), .ZN(P2_U3522) );
  AOI21_X1 U16072 ( .B1(n14010), .B2(n15398), .A(n14009), .ZN(n14011) );
  OAI211_X1 U16073 ( .C1(n14013), .C2(n14043), .A(n14012), .B(n14011), .ZN(
        n14064) );
  MUX2_X1 U16074 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14064), .S(n15431), .Z(
        P2_U3521) );
  NAND2_X1 U16075 ( .A1(n14014), .A2(n15370), .ZN(n14016) );
  NAND3_X1 U16076 ( .A1(n14017), .A2(n14016), .A3(n14015), .ZN(n14065) );
  MUX2_X1 U16077 ( .A(n14065), .B(P2_REG1_REG_21__SCAN_IN), .S(n15429), .Z(
        n14018) );
  INV_X1 U16078 ( .A(n14018), .ZN(n14019) );
  OAI21_X1 U16079 ( .B1(n7358), .B2(n14046), .A(n14019), .ZN(P2_U3520) );
  AOI211_X1 U16080 ( .C1(n14022), .C2(n15398), .A(n14021), .B(n14020), .ZN(
        n14023) );
  OAI21_X1 U16081 ( .B1(n14043), .B2(n14024), .A(n14023), .ZN(n14068) );
  MUX2_X1 U16082 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14068), .S(n15431), .Z(
        P2_U3519) );
  OAI211_X1 U16083 ( .C1(n14043), .C2(n14027), .A(n14026), .B(n14025), .ZN(
        n14069) );
  MUX2_X1 U16084 ( .A(n14069), .B(P2_REG1_REG_19__SCAN_IN), .S(n15429), .Z(
        n14028) );
  INV_X1 U16085 ( .A(n14028), .ZN(n14029) );
  OAI21_X1 U16086 ( .B1(n14072), .B2(n14046), .A(n14029), .ZN(P2_U3518) );
  AOI21_X1 U16087 ( .B1(n14031), .B2(n15398), .A(n14030), .ZN(n14032) );
  OAI211_X1 U16088 ( .C1(n14034), .C2(n14043), .A(n14033), .B(n14032), .ZN(
        n14073) );
  MUX2_X1 U16089 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14073), .S(n15431), .Z(
        P2_U3517) );
  OAI211_X1 U16090 ( .C1(n14043), .C2(n14037), .A(n14036), .B(n14035), .ZN(
        n14074) );
  MUX2_X1 U16091 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14074), .S(n15431), .Z(
        n14038) );
  INV_X1 U16092 ( .A(n14038), .ZN(n14039) );
  OAI21_X1 U16093 ( .B1(n14077), .B2(n14046), .A(n14039), .ZN(P2_U3516) );
  OAI211_X1 U16094 ( .C1(n14043), .C2(n14042), .A(n14041), .B(n14040), .ZN(
        n14078) );
  MUX2_X1 U16095 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14078), .S(n15431), .Z(
        n14044) );
  INV_X1 U16096 ( .A(n14044), .ZN(n14045) );
  OAI21_X1 U16097 ( .B1(n14082), .B2(n14046), .A(n14045), .ZN(P2_U3515) );
  INV_X1 U16098 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14048) );
  MUX2_X1 U16099 ( .A(n14048), .B(n14047), .S(n15420), .Z(n14049) );
  OAI21_X1 U16100 ( .B1(n14050), .B2(n14081), .A(n14049), .ZN(P2_U3497) );
  INV_X1 U16101 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14051) );
  MUX2_X1 U16102 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14054), .S(n15420), .Z(
        P2_U3494) );
  MUX2_X1 U16103 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14055), .S(n15420), .Z(
        P2_U3493) );
  INV_X1 U16104 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14057) );
  MUX2_X1 U16105 ( .A(n14057), .B(n14056), .S(n15420), .Z(n14058) );
  OAI21_X1 U16106 ( .B1(n14059), .B2(n14081), .A(n14058), .ZN(P2_U3492) );
  MUX2_X1 U16107 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14060), .S(n15420), .Z(
        P2_U3491) );
  MUX2_X1 U16108 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14061), .S(n15420), .Z(
        n14062) );
  INV_X1 U16109 ( .A(n14062), .ZN(n14063) );
  OAI21_X1 U16110 ( .B1(n7361), .B2(n14081), .A(n14063), .ZN(P2_U3490) );
  MUX2_X1 U16111 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14064), .S(n15420), .Z(
        P2_U3489) );
  MUX2_X1 U16112 ( .A(n14065), .B(P2_REG0_REG_21__SCAN_IN), .S(n15418), .Z(
        n14066) );
  INV_X1 U16113 ( .A(n14066), .ZN(n14067) );
  OAI21_X1 U16114 ( .B1(n7358), .B2(n14081), .A(n14067), .ZN(P2_U3488) );
  MUX2_X1 U16115 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14068), .S(n15420), .Z(
        P2_U3487) );
  MUX2_X1 U16116 ( .A(n14069), .B(P2_REG0_REG_19__SCAN_IN), .S(n15418), .Z(
        n14070) );
  INV_X1 U16117 ( .A(n14070), .ZN(n14071) );
  OAI21_X1 U16118 ( .B1(n14072), .B2(n14081), .A(n14071), .ZN(P2_U3486) );
  MUX2_X1 U16119 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14073), .S(n15420), .Z(
        P2_U3484) );
  MUX2_X1 U16120 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14074), .S(n15420), .Z(
        n14075) );
  INV_X1 U16121 ( .A(n14075), .ZN(n14076) );
  OAI21_X1 U16122 ( .B1(n14077), .B2(n14081), .A(n14076), .ZN(P2_U3481) );
  MUX2_X1 U16123 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14078), .S(n15420), .Z(
        n14079) );
  INV_X1 U16124 ( .A(n14079), .ZN(n14080) );
  OAI21_X1 U16125 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(P2_U3478) );
  INV_X1 U16126 ( .A(n14083), .ZN(n14765) );
  INV_X1 U16127 ( .A(n14084), .ZN(n14086) );
  NOR4_X1 U16128 ( .A1(n14086), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14085), .A4(
        P2_U3088), .ZN(n14087) );
  AOI21_X1 U16129 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n14088), .A(n14087), 
        .ZN(n14089) );
  OAI21_X1 U16130 ( .B1(n14765), .B2(n14111), .A(n14089), .ZN(P2_U3296) );
  INV_X1 U16131 ( .A(n14090), .ZN(n14092) );
  OAI222_X1 U16132 ( .A1(n14111), .A2(n14094), .B1(P2_U3088), .B2(n14092), 
        .C1(n14091), .C2(n14106), .ZN(P2_U3297) );
  INV_X1 U16133 ( .A(n14095), .ZN(n14768) );
  OAI222_X1 U16134 ( .A1(n14111), .A2(n14768), .B1(P2_U3088), .B2(n14097), 
        .C1(n14096), .C2(n14106), .ZN(P2_U3298) );
  NAND2_X1 U16135 ( .A1(n14769), .A2(n14098), .ZN(n14100) );
  OAI211_X1 U16136 ( .C1(n14106), .C2(n14101), .A(n14100), .B(n14099), .ZN(
        P2_U3299) );
  INV_X1 U16137 ( .A(n14102), .ZN(n14774) );
  OAI222_X1 U16138 ( .A1(n14104), .A2(P2_U3088), .B1(n14111), .B2(n14774), 
        .C1(n14103), .C2(n14106), .ZN(P2_U3300) );
  INV_X1 U16139 ( .A(n14105), .ZN(n14779) );
  OAI222_X1 U16140 ( .A1(n14108), .A2(P2_U3088), .B1(n14111), .B2(n14779), 
        .C1(n14107), .C2(n14106), .ZN(P2_U3301) );
  OAI222_X1 U16141 ( .A1(n14106), .A2(n14112), .B1(n14111), .B2(n14110), .C1(
        n14109), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U16142 ( .A(n14113), .ZN(n14114) );
  MUX2_X1 U16143 ( .A(n14114), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16144 ( .A(n14116), .B(n14115), .Z(n14122) );
  AOI22_X1 U16145 ( .A1(n14960), .A2(n14524), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14117) );
  OAI21_X1 U16146 ( .B1(n14488), .B2(n14969), .A(n14117), .ZN(n14120) );
  NAND2_X1 U16147 ( .A1(n14497), .A2(n15156), .ZN(n14679) );
  NOR2_X1 U16148 ( .A1(n14679), .A2(n14241), .ZN(n14119) );
  AOI211_X1 U16149 ( .C1(n14244), .C2(n14496), .A(n14120), .B(n14119), .ZN(
        n14121) );
  OAI21_X1 U16150 ( .B1(n14122), .B2(n14976), .A(n14121), .ZN(P1_U3214) );
  XOR2_X1 U16151 ( .A(n14124), .B(n14123), .Z(n14132) );
  OR2_X1 U16152 ( .A1(n15097), .A2(n14440), .ZN(n14126) );
  INV_X1 U16153 ( .A(n14523), .ZN(n14443) );
  OR2_X1 U16154 ( .A1(n15102), .A2(n14443), .ZN(n14125) );
  NAND2_X1 U16155 ( .A1(n14126), .A2(n14125), .ZN(n14698) );
  INV_X1 U16156 ( .A(n14698), .ZN(n14128) );
  OAI22_X1 U16157 ( .A1(n14203), .A2(n14128), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14127), .ZN(n14130) );
  NAND2_X1 U16158 ( .A1(n14562), .A2(n15156), .ZN(n14697) );
  NOR2_X1 U16159 ( .A1(n14697), .A2(n14241), .ZN(n14129) );
  AOI211_X1 U16160 ( .C1(n14244), .C2(n14558), .A(n14130), .B(n14129), .ZN(
        n14131) );
  OAI21_X1 U16161 ( .B1(n14132), .B2(n14976), .A(n14131), .ZN(P1_U3216) );
  OAI211_X1 U16162 ( .C1(n14135), .C2(n14134), .A(n14133), .B(n14965), .ZN(
        n14143) );
  OAI22_X1 U16163 ( .A1(n14969), .A2(n14137), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14136), .ZN(n14140) );
  NOR2_X1 U16164 ( .A1(n14972), .A2(n14138), .ZN(n14139) );
  AOI211_X1 U16165 ( .C1(n14244), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14142) );
  OAI211_X1 U16166 ( .C1(n15205), .C2(n14962), .A(n14143), .B(n14142), .ZN(
        P1_U3217) );
  INV_X1 U16167 ( .A(n14721), .ZN(n14619) );
  AOI21_X1 U16168 ( .B1(n14145), .B2(n14144), .A(n14976), .ZN(n14147) );
  NAND2_X1 U16169 ( .A1(n14147), .A2(n14146), .ZN(n14151) );
  NAND2_X1 U16170 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14403)
         );
  OAI21_X1 U16171 ( .B1(n14969), .B2(n14612), .A(n14403), .ZN(n14149) );
  NOR2_X1 U16172 ( .A1(n14985), .A2(n14616), .ZN(n14148) );
  AOI211_X1 U16173 ( .C1(n14960), .C2(n14957), .A(n14149), .B(n14148), .ZN(
        n14150) );
  OAI211_X1 U16174 ( .C1(n14619), .C2(n14962), .A(n14151), .B(n14150), .ZN(
        P1_U3219) );
  INV_X1 U16175 ( .A(n14152), .ZN(n14153) );
  AOI21_X1 U16176 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14160) );
  AOI22_X1 U16177 ( .A1(n14958), .A2(n14585), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14157) );
  NAND2_X1 U16178 ( .A1(n14960), .A2(n14584), .ZN(n14156) );
  OAI211_X1 U16179 ( .C1(n14985), .C2(n14587), .A(n14157), .B(n14156), .ZN(
        n14158) );
  AOI21_X1 U16180 ( .B1(n14709), .B2(n14981), .A(n14158), .ZN(n14159) );
  OAI21_X1 U16181 ( .B1(n14160), .B2(n14976), .A(n14159), .ZN(P1_U3223) );
  INV_X1 U16182 ( .A(n14161), .ZN(n14165) );
  AOI21_X1 U16183 ( .B1(n14214), .B2(n14163), .A(n14162), .ZN(n14164) );
  OAI21_X1 U16184 ( .B1(n14985), .B2(n14165), .A(n14164), .ZN(n14171) );
  INV_X1 U16185 ( .A(n14166), .ZN(n14167) );
  AOI211_X1 U16186 ( .C1(n14169), .C2(n14168), .A(n14976), .B(n14167), .ZN(
        n14170) );
  AOI211_X1 U16187 ( .C1(n14981), .C2(n14172), .A(n14171), .B(n14170), .ZN(
        n14173) );
  INV_X1 U16188 ( .A(n14173), .ZN(P1_U3224) );
  XOR2_X1 U16189 ( .A(n14175), .B(n14174), .Z(n14180) );
  AOI22_X1 U16190 ( .A1(n14960), .A2(n14523), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14176) );
  OAI21_X1 U16191 ( .B1(n14489), .B2(n14969), .A(n14176), .ZN(n14178) );
  NAND2_X1 U16192 ( .A1(n14518), .A2(n15156), .ZN(n14686) );
  NOR2_X1 U16193 ( .A1(n14686), .A2(n14241), .ZN(n14177) );
  AOI211_X1 U16194 ( .C1(n14244), .C2(n14531), .A(n14178), .B(n14177), .ZN(
        n14179) );
  OAI21_X1 U16195 ( .B1(n14180), .B2(n14976), .A(n14179), .ZN(P1_U3225) );
  XOR2_X1 U16196 ( .A(n14182), .B(n14181), .Z(n14187) );
  AOI22_X1 U16197 ( .A1(n14960), .A2(n14566), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14183) );
  OAI21_X1 U16198 ( .B1(n14538), .B2(n14969), .A(n14183), .ZN(n14185) );
  NAND2_X1 U16199 ( .A1(n14549), .A2(n15156), .ZN(n14695) );
  NOR2_X1 U16200 ( .A1(n14695), .A2(n14241), .ZN(n14184) );
  AOI211_X1 U16201 ( .C1(n14244), .C2(n14548), .A(n14185), .B(n14184), .ZN(
        n14186) );
  OAI21_X1 U16202 ( .B1(n14187), .B2(n14976), .A(n14186), .ZN(P1_U3229) );
  OAI211_X1 U16203 ( .C1(n14190), .C2(n14189), .A(n14188), .B(n14965), .ZN(
        n14197) );
  AOI22_X1 U16204 ( .A1(n14214), .A2(n14191), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14196) );
  NAND2_X1 U16205 ( .A1(n14981), .A2(n14192), .ZN(n14195) );
  NAND2_X1 U16206 ( .A1(n14244), .A2(n14193), .ZN(n14194) );
  NAND4_X1 U16207 ( .A1(n14197), .A2(n14196), .A3(n14195), .A4(n14194), .ZN(
        P1_U3231) );
  OAI211_X1 U16208 ( .C1(n14200), .C2(n14199), .A(n14198), .B(n14965), .ZN(
        n14207) );
  INV_X1 U16209 ( .A(n14602), .ZN(n14205) );
  AND2_X1 U16210 ( .A1(n14627), .A2(n14641), .ZN(n14201) );
  AOI21_X1 U16211 ( .B1(n14565), .B2(n14643), .A(n14201), .ZN(n14598) );
  OAI22_X1 U16212 ( .A1(n14203), .A2(n14598), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14202), .ZN(n14204) );
  AOI21_X1 U16213 ( .B1(n14244), .B2(n14205), .A(n14204), .ZN(n14206) );
  OAI211_X1 U16214 ( .C1(n14208), .C2(n14962), .A(n14207), .B(n14206), .ZN(
        P1_U3233) );
  OAI211_X1 U16215 ( .C1(n14211), .C2(n14210), .A(n14209), .B(n14965), .ZN(
        n14219) );
  INV_X1 U16216 ( .A(n14212), .ZN(n14216) );
  AND2_X1 U16217 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14364) );
  AOI21_X1 U16218 ( .B1(n14214), .B2(n14213), .A(n14364), .ZN(n14215) );
  OAI21_X1 U16219 ( .B1(n14985), .B2(n14216), .A(n14215), .ZN(n14217) );
  INV_X1 U16220 ( .A(n14217), .ZN(n14218) );
  OAI211_X1 U16221 ( .C1(n7313), .C2(n14962), .A(n14219), .B(n14218), .ZN(
        P1_U3234) );
  OAI21_X1 U16222 ( .B1(n14222), .B2(n14221), .A(n14220), .ZN(n14223) );
  NAND2_X1 U16223 ( .A1(n14223), .A2(n14965), .ZN(n14229) );
  INV_X1 U16224 ( .A(n14566), .ZN(n14539) );
  OAI22_X1 U16225 ( .A1(n14969), .A2(n14539), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14224), .ZN(n14227) );
  NOR2_X1 U16226 ( .A1(n14972), .A2(n14225), .ZN(n14226) );
  AOI211_X1 U16227 ( .C1(n14244), .C2(n14573), .A(n14227), .B(n14226), .ZN(
        n14228) );
  OAI211_X1 U16228 ( .C1(n14707), .C2(n14241), .A(n14229), .B(n14228), .ZN(
        P1_U3235) );
  XOR2_X1 U16229 ( .A(n14231), .B(n14230), .Z(n14237) );
  NAND2_X1 U16230 ( .A1(n14960), .A2(n14644), .ZN(n14232) );
  NAND2_X1 U16231 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14380)
         );
  OAI211_X1 U16232 ( .C1(n14233), .C2(n14969), .A(n14232), .B(n14380), .ZN(
        n14235) );
  INV_X1 U16233 ( .A(n14727), .ZN(n14636) );
  NOR2_X1 U16234 ( .A1(n14636), .A2(n14962), .ZN(n14234) );
  AOI211_X1 U16235 ( .C1(n14244), .C2(n14633), .A(n14235), .B(n14234), .ZN(
        n14236) );
  OAI21_X1 U16236 ( .B1(n14237), .B2(n14976), .A(n14236), .ZN(P1_U3238) );
  XOR2_X1 U16237 ( .A(n14239), .B(n14238), .Z(n14246) );
  AOI22_X1 U16238 ( .A1(n14960), .A2(n14504), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14240) );
  OAI21_X1 U16239 ( .B1(n14468), .B2(n14969), .A(n14240), .ZN(n14243) );
  NAND2_X1 U16240 ( .A1(n14507), .A2(n15156), .ZN(n14684) );
  NOR2_X1 U16241 ( .A1(n14684), .A2(n14241), .ZN(n14242) );
  AOI211_X1 U16242 ( .C1(n14244), .C2(n14510), .A(n14243), .B(n14242), .ZN(
        n14245) );
  OAI21_X1 U16243 ( .B1(n14246), .B2(n14976), .A(n14245), .ZN(P1_U3240) );
  OAI211_X1 U16244 ( .C1(n14249), .C2(n14248), .A(n14247), .B(n14965), .ZN(
        n14254) );
  NAND2_X1 U16245 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15062)
         );
  OAI21_X1 U16246 ( .B1(n14969), .B2(n14738), .A(n15062), .ZN(n14252) );
  NOR2_X1 U16247 ( .A1(n14985), .A2(n14250), .ZN(n14251) );
  AOI211_X1 U16248 ( .C1(n14960), .C2(n14257), .A(n14252), .B(n14251), .ZN(
        n14253) );
  OAI211_X1 U16249 ( .C1(n14255), .C2(n14962), .A(n14254), .B(n14253), .ZN(
        P1_U3241) );
  MUX2_X1 U16250 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14406), .S(n14285), .Z(
        P1_U3591) );
  MUX2_X1 U16251 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14454), .S(n14285), .Z(
        P1_U3590) );
  MUX2_X1 U16252 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14256), .S(n14285), .Z(
        P1_U3589) );
  MUX2_X1 U16253 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14447), .S(n14285), .Z(
        P1_U3588) );
  MUX2_X1 U16254 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14505), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16255 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14524), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16256 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14504), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16257 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14523), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16258 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14566), .S(n14285), .Z(
        P1_U3583) );
  MUX2_X1 U16259 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14585), .S(n14285), .Z(
        P1_U3582) );
  MUX2_X1 U16260 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14565), .S(n14285), .Z(
        P1_U3581) );
  MUX2_X1 U16261 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14584), .S(n14285), .Z(
        P1_U3580) );
  MUX2_X1 U16262 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14627), .S(n14285), .Z(
        P1_U3579) );
  MUX2_X1 U16263 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14957), .S(n14285), .Z(
        P1_U3578) );
  MUX2_X1 U16264 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14644), .S(n14285), .Z(
        P1_U3577) );
  MUX2_X1 U16265 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14959), .S(n14285), .Z(
        P1_U3576) );
  MUX2_X1 U16266 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14642), .S(n14285), .Z(
        P1_U3575) );
  MUX2_X1 U16267 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14257), .S(n14285), .Z(
        P1_U3574) );
  MUX2_X1 U16268 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14258), .S(n14285), .Z(
        P1_U3573) );
  MUX2_X1 U16269 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14259), .S(n14285), .Z(
        P1_U3572) );
  MUX2_X1 U16270 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14260), .S(n14285), .Z(
        P1_U3571) );
  MUX2_X1 U16271 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14261), .S(n14285), .Z(
        P1_U3570) );
  MUX2_X1 U16272 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14262), .S(n14285), .Z(
        P1_U3569) );
  MUX2_X1 U16273 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14263), .S(n14285), .Z(
        P1_U3568) );
  MUX2_X1 U16274 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14264), .S(n14285), .Z(
        P1_U3567) );
  MUX2_X1 U16275 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14265), .S(n14285), .Z(
        P1_U3566) );
  MUX2_X1 U16276 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14266), .S(n14285), .Z(
        P1_U3565) );
  MUX2_X1 U16277 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14267), .S(n14285), .Z(
        P1_U3564) );
  MUX2_X1 U16278 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14268), .S(n14285), .Z(
        P1_U3563) );
  MUX2_X1 U16279 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14269), .S(n14285), .Z(
        P1_U3562) );
  MUX2_X1 U16280 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10887), .S(n14285), .Z(
        P1_U3561) );
  MUX2_X1 U16281 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15091), .S(n14285), .Z(
        P1_U3560) );
  INV_X1 U16282 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14270) );
  OAI22_X1 U16283 ( .A1(n15064), .A2(n7087), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14270), .ZN(n14271) );
  AOI21_X1 U16284 ( .B1(n14272), .B2(n14398), .A(n14271), .ZN(n14280) );
  OAI211_X1 U16285 ( .C1(n14275), .C2(n14274), .A(n15060), .B(n14273), .ZN(
        n14279) );
  OAI211_X1 U16286 ( .C1(n14277), .C2(n14282), .A(n14400), .B(n14276), .ZN(
        n14278) );
  NAND3_X1 U16287 ( .A1(n14280), .A2(n14279), .A3(n14278), .ZN(P1_U3244) );
  MUX2_X1 U16288 ( .A(n14282), .B(n14281), .S(n14776), .Z(n14284) );
  NAND2_X1 U16289 ( .A1(n14284), .A2(n14283), .ZN(n14286) );
  OAI211_X1 U16290 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14287), .A(n14286), .B(
        n14285), .ZN(n14327) );
  INV_X1 U16291 ( .A(n14288), .ZN(n14291) );
  OAI22_X1 U16292 ( .A1(n15064), .A2(n7085), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14289), .ZN(n14290) );
  AOI21_X1 U16293 ( .B1(n14291), .B2(n14398), .A(n14290), .ZN(n14299) );
  OAI211_X1 U16294 ( .C1(n14293), .C2(n14292), .A(n14400), .B(n14304), .ZN(
        n14298) );
  OAI211_X1 U16295 ( .C1(n14296), .C2(n14295), .A(n15060), .B(n14294), .ZN(
        n14297) );
  NAND4_X1 U16296 ( .A1(n14327), .A2(n14299), .A3(n14298), .A4(n14297), .ZN(
        P1_U3245) );
  OAI211_X1 U16297 ( .C1(n14302), .C2(n14301), .A(n15060), .B(n14300), .ZN(
        n14311) );
  MUX2_X1 U16298 ( .A(n11423), .B(P1_REG2_REG_3__SCAN_IN), .S(n14307), .Z(
        n14305) );
  NAND3_X1 U16299 ( .A1(n14305), .A2(n14304), .A3(n14303), .ZN(n14306) );
  NAND3_X1 U16300 ( .A1(n14400), .A2(n14320), .A3(n14306), .ZN(n14310) );
  AOI22_X1 U16301 ( .A1(n14365), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14309) );
  NAND2_X1 U16302 ( .A1(n14398), .A2(n14307), .ZN(n14308) );
  NAND4_X1 U16303 ( .A1(n14311), .A2(n14310), .A3(n14309), .A4(n14308), .ZN(
        P1_U3246) );
  INV_X1 U16304 ( .A(n14312), .ZN(n14313) );
  OAI21_X1 U16305 ( .B1(n15064), .B2(n8862), .A(n14313), .ZN(n14314) );
  AOI21_X1 U16306 ( .B1(n14315), .B2(n14398), .A(n14314), .ZN(n14326) );
  OAI211_X1 U16307 ( .C1(n14318), .C2(n14317), .A(n15060), .B(n14316), .ZN(
        n14325) );
  NAND3_X1 U16308 ( .A1(n14321), .A2(n14320), .A3(n14319), .ZN(n14322) );
  NAND3_X1 U16309 ( .A1(n14400), .A2(n14323), .A3(n14322), .ZN(n14324) );
  NAND4_X1 U16310 ( .A1(n14327), .A2(n14326), .A3(n14325), .A4(n14324), .ZN(
        P1_U3247) );
  NOR2_X1 U16311 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14328), .ZN(n14331) );
  NOR2_X1 U16312 ( .A1(n15055), .A2(n14329), .ZN(n14330) );
  AOI211_X1 U16313 ( .C1(n14365), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n14331), .B(
        n14330), .ZN(n14342) );
  OAI211_X1 U16314 ( .C1(n14334), .C2(n14333), .A(n15060), .B(n14332), .ZN(
        n14341) );
  INV_X1 U16315 ( .A(n14335), .ZN(n14353) );
  NAND3_X1 U16316 ( .A1(n14338), .A2(n14337), .A3(n14336), .ZN(n14339) );
  NAND3_X1 U16317 ( .A1(n14400), .A2(n14353), .A3(n14339), .ZN(n14340) );
  NAND3_X1 U16318 ( .A1(n14342), .A2(n14341), .A3(n14340), .ZN(P1_U3249) );
  INV_X1 U16319 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14344) );
  OAI21_X1 U16320 ( .B1(n15064), .B2(n14344), .A(n14343), .ZN(n14345) );
  AOI21_X1 U16321 ( .B1(n14350), .B2(n14398), .A(n14345), .ZN(n14358) );
  OAI211_X1 U16322 ( .C1(n14348), .C2(n14347), .A(n15060), .B(n14346), .ZN(
        n14357) );
  INV_X1 U16323 ( .A(n14349), .ZN(n14352) );
  MUX2_X1 U16324 ( .A(n11254), .B(P1_REG2_REG_7__SCAN_IN), .S(n14350), .Z(
        n14351) );
  NAND3_X1 U16325 ( .A1(n14353), .A2(n14352), .A3(n14351), .ZN(n14354) );
  NAND3_X1 U16326 ( .A1(n14400), .A2(n14355), .A3(n14354), .ZN(n14356) );
  NAND3_X1 U16327 ( .A1(n14358), .A2(n14357), .A3(n14356), .ZN(P1_U3250) );
  OAI211_X1 U16328 ( .C1(n14361), .C2(n14360), .A(n14359), .B(n15060), .ZN(
        n14371) );
  NOR2_X1 U16329 ( .A1(n15055), .A2(n14362), .ZN(n14363) );
  AOI211_X1 U16330 ( .C1(n14365), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n14364), 
        .B(n14363), .ZN(n14370) );
  OAI211_X1 U16331 ( .C1(n14368), .C2(n14367), .A(n14366), .B(n14400), .ZN(
        n14369) );
  NAND3_X1 U16332 ( .A1(n14371), .A2(n14370), .A3(n14369), .ZN(P1_U3256) );
  OAI21_X1 U16333 ( .B1(n14999), .B2(n14373), .A(n14372), .ZN(n14390) );
  XNOR2_X1 U16334 ( .A(n14390), .B(n14379), .ZN(n14391) );
  XNOR2_X1 U16335 ( .A(n14391), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14384) );
  AOI21_X1 U16336 ( .B1(n14375), .B2(P1_REG1_REG_17__SCAN_IN), .A(n14374), 
        .ZN(n14376) );
  NOR2_X1 U16337 ( .A1(n14376), .A2(n14379), .ZN(n14386) );
  AOI21_X1 U16338 ( .B1(n14376), .B2(n14379), .A(n14386), .ZN(n14378) );
  AND2_X1 U16339 ( .A1(n14378), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14385) );
  INV_X1 U16340 ( .A(n14385), .ZN(n14377) );
  OAI211_X1 U16341 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14378), .A(n14377), 
        .B(n15060), .ZN(n14383) );
  INV_X1 U16342 ( .A(n14379), .ZN(n14389) );
  OAI21_X1 U16343 ( .B1(n15064), .B2(n8916), .A(n14380), .ZN(n14381) );
  AOI21_X1 U16344 ( .B1(n14389), .B2(n14398), .A(n14381), .ZN(n14382) );
  OAI211_X1 U16345 ( .C1(n14384), .C2(n15057), .A(n14383), .B(n14382), .ZN(
        P1_U3261) );
  NOR2_X1 U16346 ( .A1(n14386), .A2(n14385), .ZN(n14388) );
  XOR2_X1 U16347 ( .A(n14388), .B(n14387), .Z(n14397) );
  NAND2_X1 U16348 ( .A1(n14390), .A2(n14389), .ZN(n14393) );
  NAND2_X1 U16349 ( .A1(n14391), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U16350 ( .A1(n14393), .A2(n14392), .ZN(n14394) );
  XOR2_X1 U16351 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14394), .Z(n14395) );
  AOI22_X1 U16352 ( .A1(n14397), .A2(n15060), .B1(n14400), .B2(n14395), .ZN(
        n14402) );
  INV_X1 U16353 ( .A(n14395), .ZN(n14399) );
  INV_X1 U16354 ( .A(n14991), .ZN(n14963) );
  OR2_X1 U16355 ( .A1(n14714), .A2(n14614), .ZN(n14600) );
  NOR2_X2 U16356 ( .A1(n14709), .A2(n14600), .ZN(n14586) );
  NAND2_X1 U16357 ( .A1(n14572), .A2(n14586), .ZN(n14571) );
  NAND2_X1 U16358 ( .A1(n14404), .A2(n15077), .ZN(n14657) );
  INV_X1 U16359 ( .A(P1_B_REG_SCAN_IN), .ZN(n14405) );
  OR2_X1 U16360 ( .A1(n14776), .A2(n14405), .ZN(n14453) );
  NAND3_X1 U16361 ( .A1(n14643), .A2(n14406), .A3(n14453), .ZN(n14658) );
  NOR2_X1 U16362 ( .A1(n15112), .A2(n14658), .ZN(n14412) );
  NOR2_X1 U16363 ( .A1(n7319), .A2(n15106), .ZN(n14408) );
  AOI211_X1 U16364 ( .C1(n15112), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14412), 
        .B(n14408), .ZN(n14409) );
  OAI21_X1 U16365 ( .B1(n14577), .B2(n14657), .A(n14409), .ZN(P1_U3263) );
  OAI211_X1 U16366 ( .C1(n14660), .C2(n14450), .A(n15077), .B(n14410), .ZN(
        n14659) );
  NOR2_X1 U16367 ( .A1(n14660), .A2(n15106), .ZN(n14411) );
  AOI211_X1 U16368 ( .C1(n15112), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14412), 
        .B(n14411), .ZN(n14413) );
  OAI21_X1 U16369 ( .B1(n14577), .B2(n14659), .A(n14413), .ZN(P1_U3264) );
  OR2_X1 U16370 ( .A1(n14416), .A2(n14642), .ZN(n14417) );
  OR2_X1 U16371 ( .A1(n14951), .A2(n14959), .ZN(n14418) );
  AND2_X1 U16372 ( .A1(n14727), .A2(n14957), .ZN(n14421) );
  OR2_X1 U16373 ( .A1(n14721), .A2(n14627), .ZN(n14423) );
  NAND2_X1 U16374 ( .A1(n14714), .A2(n14584), .ZN(n14425) );
  INV_X1 U16375 ( .A(n14581), .ZN(n14439) );
  NAND2_X1 U16376 ( .A1(n14572), .A2(n14440), .ZN(n14426) );
  NAND2_X1 U16377 ( .A1(n14562), .A2(n14566), .ZN(n14428) );
  INV_X1 U16378 ( .A(n14466), .ZN(n14471) );
  INV_X1 U16379 ( .A(n14497), .ZN(n14495) );
  INV_X1 U16380 ( .A(n14431), .ZN(n14432) );
  INV_X1 U16381 ( .A(n14652), .ZN(n14639) );
  NAND2_X1 U16382 ( .A1(n14951), .A2(n14738), .ZN(n14734) );
  INV_X1 U16383 ( .A(n14644), .ZN(n14942) );
  NAND2_X1 U16384 ( .A1(n14595), .A2(n14437), .ZN(n14582) );
  INV_X1 U16385 ( .A(n14709), .ZN(n14438) );
  INV_X1 U16386 ( .A(n14529), .ZN(n14521) );
  OR2_X1 U16387 ( .A1(n14549), .A2(n14443), .ZN(n14519) );
  NAND3_X1 U16388 ( .A1(n14541), .A2(n14521), .A3(n14519), .ZN(n14520) );
  INV_X1 U16389 ( .A(n14486), .ZN(n14483) );
  OR2_X1 U16390 ( .A1(n15097), .A2(n14488), .ZN(n14662) );
  AOI21_X1 U16391 ( .B1(n14668), .B2(n14662), .A(n15112), .ZN(n14464) );
  INV_X1 U16392 ( .A(n14450), .ZN(n14452) );
  NAND2_X1 U16393 ( .A1(n14472), .A2(n14661), .ZN(n14451) );
  AND2_X1 U16394 ( .A1(n14452), .A2(n14451), .ZN(n14666) );
  NAND2_X1 U16395 ( .A1(n14666), .A2(n15100), .ZN(n14461) );
  NAND2_X1 U16396 ( .A1(n14454), .A2(n14453), .ZN(n14455) );
  OR2_X1 U16397 ( .A1(n15102), .A2(n14455), .ZN(n14663) );
  INV_X1 U16398 ( .A(n14456), .ZN(n14457) );
  OAI22_X1 U16399 ( .A1(n14458), .A2(n14663), .B1(n14457), .B2(n14648), .ZN(
        n14459) );
  AOI21_X1 U16400 ( .B1(n15112), .B2(P1_REG2_REG_29__SCAN_IN), .A(n14459), 
        .ZN(n14460) );
  OAI211_X1 U16401 ( .C1(n14462), .C2(n15106), .A(n14461), .B(n14460), .ZN(
        n14463) );
  NOR2_X1 U16402 ( .A1(n14464), .A2(n14463), .ZN(n14465) );
  OAI21_X1 U16403 ( .B1(n14669), .B2(n14623), .A(n14465), .ZN(P1_U3356) );
  OAI211_X1 U16404 ( .C1(n14673), .C2(n14492), .A(n15077), .B(n14472), .ZN(
        n14671) );
  INV_X1 U16405 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14475) );
  INV_X1 U16406 ( .A(n14473), .ZN(n14474) );
  OAI22_X1 U16407 ( .A1(n15103), .A2(n14475), .B1(n14474), .B2(n14648), .ZN(
        n14476) );
  AOI21_X1 U16408 ( .B1(n14477), .B2(n15074), .A(n14476), .ZN(n14478) );
  OAI21_X1 U16409 ( .B1(n14671), .B2(n14577), .A(n14478), .ZN(n14479) );
  AOI21_X1 U16410 ( .B1(n14670), .B2(n14654), .A(n14479), .ZN(n14480) );
  OAI21_X1 U16411 ( .B1(n14481), .B2(n15112), .A(n14480), .ZN(P1_U3265) );
  OAI21_X1 U16412 ( .B1(n14484), .B2(n14483), .A(n14482), .ZN(n14491) );
  OAI22_X1 U16413 ( .A1(n14489), .A2(n15097), .B1(n15102), .B2(n14488), .ZN(
        n14490) );
  INV_X1 U16414 ( .A(n14509), .ZN(n14494) );
  INV_X1 U16415 ( .A(n14492), .ZN(n14493) );
  OAI211_X1 U16416 ( .C1(n14495), .C2(n14494), .A(n14493), .B(n15077), .ZN(
        n14677) );
  AOI22_X1 U16417 ( .A1(n15112), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14496), 
        .B2(n15099), .ZN(n14499) );
  NAND2_X1 U16418 ( .A1(n14497), .A2(n15074), .ZN(n14498) );
  OAI211_X1 U16419 ( .C1(n14677), .C2(n14577), .A(n14499), .B(n14498), .ZN(
        n14500) );
  AOI21_X1 U16420 ( .B1(n14676), .B2(n15081), .A(n14500), .ZN(n14501) );
  OAI21_X1 U16421 ( .B1(n14680), .B2(n15112), .A(n14501), .ZN(P1_U3266) );
  OAI21_X1 U16422 ( .B1(n14514), .B2(n14503), .A(n14502), .ZN(n14506) );
  AOI222_X1 U16423 ( .A1(n14506), .A2(n14645), .B1(n14505), .B2(n14643), .C1(
        n14504), .C2(n14641), .ZN(n14685) );
  OAI211_X1 U16424 ( .C1(n7320), .C2(n14508), .A(n15077), .B(n14509), .ZN(
        n14682) );
  INV_X1 U16425 ( .A(n14682), .ZN(n14513) );
  AOI22_X1 U16426 ( .A1(n15112), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14510), 
        .B2(n15099), .ZN(n14511) );
  OAI21_X1 U16427 ( .B1(n7320), .B2(n15106), .A(n14511), .ZN(n14512) );
  AOI21_X1 U16428 ( .B1(n14513), .B2(n15080), .A(n14512), .ZN(n14517) );
  XNOR2_X1 U16429 ( .A(n14515), .B(n14514), .ZN(n14681) );
  NAND2_X1 U16430 ( .A1(n14681), .A2(n14654), .ZN(n14516) );
  OAI211_X1 U16431 ( .C1(n14685), .C2(n15112), .A(n14517), .B(n14516), .ZN(
        P1_U3267) );
  AOI211_X1 U16432 ( .C1(n14518), .C2(n14547), .A(n15159), .B(n14508), .ZN(
        n14688) );
  AND2_X1 U16433 ( .A1(n14541), .A2(n14519), .ZN(n14522) );
  OAI21_X1 U16434 ( .B1(n14522), .B2(n14521), .A(n14520), .ZN(n14525) );
  AOI222_X1 U16435 ( .A1(n14525), .A2(n14645), .B1(n14524), .B2(n14643), .C1(
        n14523), .C2(n14641), .ZN(n14690) );
  INV_X1 U16436 ( .A(n14690), .ZN(n14526) );
  AOI21_X1 U16437 ( .B1(n14688), .B2(n14527), .A(n14526), .ZN(n14536) );
  OAI21_X1 U16438 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n14691) );
  INV_X1 U16439 ( .A(n14691), .ZN(n14534) );
  AOI22_X1 U16440 ( .A1(n15112), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n14531), 
        .B2(n15099), .ZN(n14532) );
  OAI21_X1 U16441 ( .B1(n7321), .B2(n15106), .A(n14532), .ZN(n14533) );
  AOI21_X1 U16442 ( .B1(n14534), .B2(n14654), .A(n14533), .ZN(n14535) );
  OAI21_X1 U16443 ( .B1(n14536), .B2(n15112), .A(n14535), .ZN(P1_U3268) );
  XNOR2_X1 U16444 ( .A(n14537), .B(n14544), .ZN(n14692) );
  OAI22_X1 U16445 ( .A1(n14539), .A2(n15097), .B1(n15102), .B2(n14538), .ZN(
        n14546) );
  INV_X1 U16446 ( .A(n14540), .ZN(n14543) );
  INV_X1 U16447 ( .A(n14541), .ZN(n14542) );
  AOI211_X1 U16448 ( .C1(n14544), .C2(n14543), .A(n15145), .B(n14542), .ZN(
        n14545) );
  AOI211_X1 U16449 ( .C1(n15072), .C2(n14692), .A(n14546), .B(n14545), .ZN(
        n14696) );
  OAI211_X1 U16450 ( .C1(n7323), .C2(n7324), .A(n14547), .B(n15077), .ZN(
        n14693) );
  AOI22_X1 U16451 ( .A1(n15112), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14548), 
        .B2(n15099), .ZN(n14551) );
  NAND2_X1 U16452 ( .A1(n14549), .A2(n15074), .ZN(n14550) );
  OAI211_X1 U16453 ( .C1(n14693), .C2(n14577), .A(n14551), .B(n14550), .ZN(
        n14552) );
  AOI21_X1 U16454 ( .B1(n14692), .B2(n15081), .A(n14552), .ZN(n14553) );
  OAI21_X1 U16455 ( .B1(n14696), .B2(n15112), .A(n14553), .ZN(P1_U3269) );
  OAI21_X1 U16456 ( .B1(n14555), .B2(n14427), .A(n14554), .ZN(n14703) );
  AOI21_X1 U16457 ( .B1(n14562), .B2(n14571), .A(n7324), .ZN(n14700) );
  INV_X1 U16458 ( .A(n14700), .ZN(n14560) );
  AOI21_X1 U16459 ( .B1(n14556), .B2(n14427), .A(n6767), .ZN(n14557) );
  OR2_X1 U16460 ( .A1(n14557), .A2(n15145), .ZN(n14702) );
  AOI21_X1 U16461 ( .B1(n15099), .B2(n14558), .A(n14698), .ZN(n14559) );
  OAI211_X1 U16462 ( .C1(n11216), .C2(n14560), .A(n14702), .B(n14559), .ZN(
        n14561) );
  NAND2_X1 U16463 ( .A1(n14561), .A2(n15103), .ZN(n14564) );
  AOI22_X1 U16464 ( .A1(n14562), .A2(n15074), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15112), .ZN(n14563) );
  OAI211_X1 U16465 ( .C1(n14703), .C2(n14623), .A(n14564), .B(n14563), .ZN(
        P1_U3270) );
  XNOR2_X1 U16466 ( .A(n6795), .B(n7161), .ZN(n14567) );
  AOI222_X1 U16467 ( .A1(n14567), .A2(n14645), .B1(n14566), .B2(n14643), .C1(
        n14565), .C2(n14641), .ZN(n14708) );
  OAI21_X1 U16468 ( .B1(n14570), .B2(n14569), .A(n14568), .ZN(n14704) );
  OAI211_X1 U16469 ( .C1(n14572), .C2(n14586), .A(n15077), .B(n14571), .ZN(
        n14705) );
  AOI22_X1 U16470 ( .A1(n15112), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14573), 
        .B2(n15099), .ZN(n14576) );
  NAND2_X1 U16471 ( .A1(n14574), .A2(n15074), .ZN(n14575) );
  OAI211_X1 U16472 ( .C1(n14705), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14578) );
  AOI21_X1 U16473 ( .B1(n14704), .B2(n14654), .A(n14578), .ZN(n14579) );
  OAI21_X1 U16474 ( .B1(n14708), .B2(n15112), .A(n14579), .ZN(P1_U3271) );
  XNOR2_X1 U16475 ( .A(n14580), .B(n14581), .ZN(n14713) );
  XNOR2_X1 U16476 ( .A(n14582), .B(n14581), .ZN(n14583) );
  AOI222_X1 U16477 ( .A1(n14585), .A2(n14643), .B1(n14584), .B2(n14641), .C1(
        n14645), .C2(n14583), .ZN(n14712) );
  INV_X1 U16478 ( .A(n14712), .ZN(n14590) );
  AOI21_X1 U16479 ( .B1(n14709), .B2(n14600), .A(n14586), .ZN(n14710) );
  INV_X1 U16480 ( .A(n14710), .ZN(n14588) );
  OAI22_X1 U16481 ( .A1(n14588), .A2(n11216), .B1(n14587), .B2(n14648), .ZN(
        n14589) );
  OAI21_X1 U16482 ( .B1(n14590), .B2(n14589), .A(n15103), .ZN(n14592) );
  AOI22_X1 U16483 ( .A1(n14709), .A2(n15074), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15112), .ZN(n14591) );
  OAI211_X1 U16484 ( .C1(n14713), .C2(n14623), .A(n14592), .B(n14591), .ZN(
        P1_U3272) );
  OAI21_X1 U16485 ( .B1(n14594), .B2(n7494), .A(n14593), .ZN(n14718) );
  OAI211_X1 U16486 ( .C1(n14597), .C2(n14596), .A(n14595), .B(n14645), .ZN(
        n14599) );
  INV_X1 U16487 ( .A(n14717), .ZN(n14605) );
  INV_X1 U16488 ( .A(n14600), .ZN(n14601) );
  AOI21_X1 U16489 ( .B1(n14714), .B2(n14614), .A(n14601), .ZN(n14715) );
  INV_X1 U16490 ( .A(n14715), .ZN(n14603) );
  OAI22_X1 U16491 ( .A1(n14603), .A2(n11216), .B1(n14602), .B2(n14648), .ZN(
        n14604) );
  OAI21_X1 U16492 ( .B1(n14605), .B2(n14604), .A(n15103), .ZN(n14607) );
  AOI22_X1 U16493 ( .A1(n14714), .A2(n15074), .B1(n15112), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14606) );
  OAI211_X1 U16494 ( .C1(n14718), .C2(n14623), .A(n14607), .B(n14606), .ZN(
        P1_U3273) );
  XNOR2_X1 U16495 ( .A(n14608), .B(n14609), .ZN(n14724) );
  XNOR2_X1 U16496 ( .A(n14610), .B(n14609), .ZN(n14611) );
  AOI22_X1 U16497 ( .A1(n14611), .A2(n14645), .B1(n14641), .B2(n14957), .ZN(
        n14723) );
  INV_X1 U16498 ( .A(n14723), .ZN(n14613) );
  NOR2_X1 U16499 ( .A1(n14612), .A2(n15102), .ZN(n14720) );
  OAI21_X1 U16500 ( .B1(n14613), .B2(n14720), .A(n15103), .ZN(n14622) );
  OR2_X1 U16501 ( .A1(n14631), .A2(n14619), .ZN(n14615) );
  AND3_X1 U16502 ( .A1(n14615), .A2(n14614), .A3(n15077), .ZN(n14719) );
  INV_X1 U16503 ( .A(n14616), .ZN(n14617) );
  AOI22_X1 U16504 ( .A1(n15112), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14617), 
        .B2(n15099), .ZN(n14618) );
  OAI21_X1 U16505 ( .B1(n14619), .B2(n15106), .A(n14618), .ZN(n14620) );
  AOI21_X1 U16506 ( .B1(n14719), .B2(n15080), .A(n14620), .ZN(n14621) );
  OAI211_X1 U16507 ( .C1(n14724), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        P1_U3274) );
  XNOR2_X1 U16508 ( .A(n14624), .B(n14625), .ZN(n14725) );
  XNOR2_X1 U16509 ( .A(n14626), .B(n14625), .ZN(n14629) );
  AOI22_X1 U16510 ( .A1(n14627), .A2(n14643), .B1(n14641), .B2(n14644), .ZN(
        n14628) );
  OAI21_X1 U16511 ( .B1(n14629), .B2(n15145), .A(n14628), .ZN(n14630) );
  AOI21_X1 U16512 ( .B1(n15072), .B2(n14725), .A(n14630), .ZN(n14729) );
  INV_X1 U16513 ( .A(n14743), .ZN(n14632) );
  AOI211_X1 U16514 ( .C1(n14727), .C2(n14632), .A(n15159), .B(n14631), .ZN(
        n14726) );
  NAND2_X1 U16515 ( .A1(n14726), .A2(n15080), .ZN(n14635) );
  AOI22_X1 U16516 ( .A1(n15112), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14633), 
        .B2(n15099), .ZN(n14634) );
  OAI211_X1 U16517 ( .C1(n14636), .C2(n15106), .A(n14635), .B(n14634), .ZN(
        n14637) );
  AOI21_X1 U16518 ( .B1(n14725), .B2(n15081), .A(n14637), .ZN(n14638) );
  OAI21_X1 U16519 ( .B1(n14729), .B2(n15112), .A(n14638), .ZN(P1_U3275) );
  OAI21_X1 U16520 ( .B1(n14640), .B2(n14639), .A(n14735), .ZN(n14646) );
  AOI222_X1 U16521 ( .A1(n14646), .A2(n14645), .B1(n14644), .B2(n14643), .C1(
        n14642), .C2(n14641), .ZN(n15003) );
  AOI211_X1 U16522 ( .C1(n14951), .C2(n14647), .A(n15159), .B(n14742), .ZN(
        n15000) );
  INV_X1 U16523 ( .A(n14951), .ZN(n15002) );
  NOR2_X1 U16524 ( .A1(n15002), .A2(n15106), .ZN(n14650) );
  OAI22_X1 U16525 ( .A1(n15103), .A2(n11749), .B1(n14954), .B2(n14648), .ZN(
        n14649) );
  AOI211_X1 U16526 ( .C1(n15000), .C2(n15080), .A(n14650), .B(n14649), .ZN(
        n14656) );
  OAI21_X1 U16527 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n15006) );
  NAND2_X1 U16528 ( .A1(n15006), .A2(n14654), .ZN(n14655) );
  OAI211_X1 U16529 ( .C1(n15003), .C2(n15112), .A(n14656), .B(n14655), .ZN(
        P1_U3277) );
  OAI211_X1 U16530 ( .C1(n7319), .C2(n15204), .A(n14657), .B(n14658), .ZN(
        n14746) );
  MUX2_X1 U16531 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14746), .S(n15225), .Z(
        P1_U3559) );
  OAI211_X1 U16532 ( .C1(n14660), .C2(n15204), .A(n14659), .B(n14658), .ZN(
        n14747) );
  MUX2_X1 U16533 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14747), .S(n15225), .Z(
        P1_U3558) );
  NAND2_X1 U16534 ( .A1(n14661), .A2(n15156), .ZN(n14664) );
  NAND3_X1 U16535 ( .A1(n14664), .A2(n14663), .A3(n14662), .ZN(n14665) );
  AOI21_X1 U16536 ( .B1(n14666), .B2(n15077), .A(n14665), .ZN(n14667) );
  NAND2_X1 U16537 ( .A1(n14670), .A2(n15208), .ZN(n14672) );
  OAI211_X1 U16538 ( .C1(n14673), .C2(n15204), .A(n14672), .B(n14671), .ZN(
        n14674) );
  INV_X1 U16539 ( .A(n14674), .ZN(n14675) );
  MUX2_X1 U16540 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14748), .S(n15225), .Z(
        P1_U3556) );
  INV_X1 U16541 ( .A(n15197), .ZN(n15185) );
  NAND2_X1 U16542 ( .A1(n14676), .A2(n15185), .ZN(n14678) );
  NAND4_X1 U16543 ( .A1(n14680), .A2(n14679), .A3(n14678), .A4(n14677), .ZN(
        n14749) );
  MUX2_X1 U16544 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14749), .S(n15225), .Z(
        P1_U3555) );
  NAND2_X1 U16545 ( .A1(n14681), .A2(n15208), .ZN(n14683) );
  NAND4_X1 U16546 ( .A1(n14685), .A2(n14684), .A3(n14683), .A4(n14682), .ZN(
        n14750) );
  MUX2_X1 U16547 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14750), .S(n15225), .Z(
        P1_U3554) );
  INV_X1 U16548 ( .A(n14686), .ZN(n14687) );
  NOR2_X1 U16549 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  OAI211_X1 U16550 ( .C1(n15146), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14751) );
  MUX2_X1 U16551 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14751), .S(n15225), .Z(
        P1_U3553) );
  NAND2_X1 U16552 ( .A1(n14692), .A2(n15185), .ZN(n14694) );
  NAND4_X1 U16553 ( .A1(n14696), .A2(n14695), .A3(n14694), .A4(n14693), .ZN(
        n14752) );
  MUX2_X1 U16554 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14752), .S(n15225), .Z(
        P1_U3552) );
  INV_X1 U16555 ( .A(n14697), .ZN(n14699) );
  AOI211_X1 U16556 ( .C1(n14700), .C2(n15077), .A(n14699), .B(n14698), .ZN(
        n14701) );
  OAI211_X1 U16557 ( .C1(n15146), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14753) );
  MUX2_X1 U16558 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14753), .S(n15225), .Z(
        P1_U3551) );
  NAND2_X1 U16559 ( .A1(n14704), .A2(n15208), .ZN(n14706) );
  NAND4_X1 U16560 ( .A1(n14708), .A2(n14707), .A3(n14706), .A4(n14705), .ZN(
        n14754) );
  MUX2_X1 U16561 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14754), .S(n15225), .Z(
        P1_U3550) );
  AOI22_X1 U16562 ( .A1(n14710), .A2(n15077), .B1(n14709), .B2(n15156), .ZN(
        n14711) );
  OAI211_X1 U16563 ( .C1(n15146), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14755) );
  MUX2_X1 U16564 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14755), .S(n15225), .Z(
        P1_U3549) );
  AOI22_X1 U16565 ( .A1(n14715), .A2(n15077), .B1(n14714), .B2(n15156), .ZN(
        n14716) );
  OAI211_X1 U16566 ( .C1(n15146), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14756) );
  MUX2_X1 U16567 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14756), .S(n15225), .Z(
        P1_U3548) );
  AOI211_X1 U16568 ( .C1(n14721), .C2(n15156), .A(n14720), .B(n14719), .ZN(
        n14722) );
  OAI211_X1 U16569 ( .C1(n15146), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        n14757) );
  MUX2_X1 U16570 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14757), .S(n15225), .Z(
        P1_U3547) );
  INV_X1 U16571 ( .A(n14725), .ZN(n14730) );
  AOI21_X1 U16572 ( .B1(n14727), .B2(n15156), .A(n14726), .ZN(n14728) );
  OAI211_X1 U16573 ( .C1(n14730), .C2(n15197), .A(n14729), .B(n14728), .ZN(
        n14758) );
  MUX2_X1 U16574 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14758), .S(n15225), .Z(
        P1_U3546) );
  XNOR2_X1 U16575 ( .A(n14731), .B(n14733), .ZN(n14986) );
  INV_X1 U16576 ( .A(n14732), .ZN(n14737) );
  AOI21_X1 U16577 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(n14736) );
  NOR3_X1 U16578 ( .A1(n14737), .A2(n14736), .A3(n15145), .ZN(n14741) );
  OAI22_X1 U16579 ( .A1(n14739), .A2(n15102), .B1(n14738), .B2(n15097), .ZN(
        n14740) );
  NOR2_X1 U16580 ( .A1(n14741), .A2(n14740), .ZN(n14993) );
  INV_X1 U16581 ( .A(n14742), .ZN(n14744) );
  AOI21_X1 U16582 ( .B1(n14991), .B2(n14744), .A(n14743), .ZN(n14987) );
  AOI22_X1 U16583 ( .A1(n14987), .A2(n15077), .B1(n14991), .B2(n15156), .ZN(
        n14745) );
  OAI211_X1 U16584 ( .C1(n15146), .C2(n14986), .A(n14993), .B(n14745), .ZN(
        n14759) );
  MUX2_X1 U16585 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14759), .S(n15225), .Z(
        P1_U3545) );
  MUX2_X1 U16586 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14746), .S(n15212), .Z(
        P1_U3527) );
  MUX2_X1 U16587 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14747), .S(n15212), .Z(
        P1_U3526) );
  MUX2_X1 U16588 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14748), .S(n15212), .Z(
        P1_U3524) );
  MUX2_X1 U16589 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14749), .S(n15212), .Z(
        P1_U3523) );
  MUX2_X1 U16590 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14750), .S(n15212), .Z(
        P1_U3522) );
  MUX2_X1 U16591 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14751), .S(n15212), .Z(
        P1_U3521) );
  MUX2_X1 U16592 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14752), .S(n15212), .Z(
        P1_U3520) );
  MUX2_X1 U16593 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14753), .S(n15212), .Z(
        P1_U3519) );
  MUX2_X1 U16594 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14754), .S(n15212), .Z(
        P1_U3518) );
  MUX2_X1 U16595 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14755), .S(n15212), .Z(
        P1_U3517) );
  MUX2_X1 U16596 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14756), .S(n15212), .Z(
        P1_U3516) );
  MUX2_X1 U16597 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14757), .S(n15212), .Z(
        P1_U3515) );
  MUX2_X1 U16598 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14758), .S(n15212), .Z(
        P1_U3513) );
  MUX2_X1 U16599 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14759), .S(n15212), .Z(
        P1_U3510) );
  NOR4_X1 U16600 ( .A1(n14761), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14760), .ZN(n14762) );
  AOI21_X1 U16601 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14763), .A(n14762), 
        .ZN(n14764) );
  OAI21_X1 U16602 ( .B1(n14765), .B2(n14775), .A(n14764), .ZN(P1_U3324) );
  OAI222_X1 U16603 ( .A1(n14780), .A2(n14768), .B1(n14767), .B2(P1_U3086), 
        .C1(n14766), .C2(n14772), .ZN(P1_U3326) );
  INV_X1 U16604 ( .A(n14769), .ZN(n14771) );
  OAI222_X1 U16605 ( .A1(P1_U3086), .A2(n10202), .B1(n14780), .B2(n14771), 
        .C1(n14770), .C2(n14777), .ZN(P1_U3327) );
  OAI222_X1 U16606 ( .A1(n14776), .A2(P1_U3086), .B1(n14775), .B2(n14774), 
        .C1(n14773), .C2(n14772), .ZN(P1_U3328) );
  OAI222_X1 U16607 ( .A1(n14781), .A2(P1_U3086), .B1(n14780), .B2(n14779), 
        .C1(n14778), .C2(n14777), .ZN(P1_U3329) );
  MUX2_X1 U16608 ( .A(n15149), .B(n14782), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16609 ( .A(n14783), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16610 ( .A(n14787), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16611 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14788) );
  OAI21_X1 U16612 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14788), 
        .ZN(U28) );
  AOI21_X1 U16613 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14789) );
  OAI21_X1 U16614 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14789), 
        .ZN(U29) );
  AOI21_X1 U16615 ( .B1(n14792), .B2(n14791), .A(n14790), .ZN(SUB_1596_U61) );
  AOI21_X1 U16616 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(SUB_1596_U57) );
  AOI21_X1 U16617 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(SUB_1596_U55) );
  AOI21_X1 U16618 ( .B1(n14801), .B2(n14800), .A(n14799), .ZN(n14802) );
  XOR2_X1 U16619 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14802), .Z(SUB_1596_U54) );
  AOI21_X1 U16620 ( .B1(n14805), .B2(n14804), .A(n14803), .ZN(n14806) );
  XOR2_X1 U16621 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14806), .Z(SUB_1596_U70)
         );
  OAI222_X1 U16622 ( .A1(n15312), .A2(n14810), .B1(n15312), .B2(n14809), .C1(
        n14808), .C2(n14807), .ZN(SUB_1596_U63) );
  AOI22_X1 U16623 ( .A1(n14827), .A2(n14811), .B1(n15516), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14825) );
  OAI21_X1 U16624 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14813), .A(n14812), 
        .ZN(n14818) );
  AOI211_X1 U16625 ( .C1(n14816), .C2(n14815), .A(n15439), .B(n14814), .ZN(
        n14817) );
  AOI21_X1 U16626 ( .B1(n15519), .B2(n14818), .A(n14817), .ZN(n14824) );
  NAND2_X1 U16627 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n6665), .ZN(n14823) );
  OAI221_X1 U16628 ( .B1(n14821), .B2(n14820), .C1(n14821), .C2(n14819), .A(
        n14837), .ZN(n14822) );
  NAND4_X1 U16629 ( .A1(n14825), .A2(n14824), .A3(n14823), .A4(n14822), .ZN(
        P3_U3199) );
  AOI22_X1 U16630 ( .A1(n14827), .A2(n14826), .B1(n15516), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14843) );
  OAI21_X1 U16631 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14836) );
  AOI21_X1 U16632 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(n14834) );
  NOR2_X1 U16633 ( .A1(n14834), .A2(n15439), .ZN(n14835) );
  AOI21_X1 U16634 ( .B1(n15519), .B2(n14836), .A(n14835), .ZN(n14842) );
  NAND4_X1 U16635 ( .A1(n14843), .A2(n14842), .A3(n14841), .A4(n14840), .ZN(
        P3_U3200) );
  XNOR2_X1 U16636 ( .A(n14844), .B(n14845), .ZN(n14871) );
  AND2_X1 U16637 ( .A1(n14847), .A2(n14846), .ZN(n14850) );
  OAI211_X1 U16638 ( .C1(n14850), .C2(n14849), .A(n14848), .B(n15612), .ZN(
        n14853) );
  AOI22_X1 U16639 ( .A1(n14851), .A2(n15607), .B1(n15610), .B2(n15529), .ZN(
        n14852) );
  NAND2_X1 U16640 ( .A1(n14853), .A2(n14852), .ZN(n14869) );
  AOI21_X1 U16641 ( .B1(n14871), .B2(n14864), .A(n14869), .ZN(n14857) );
  AND2_X1 U16642 ( .A1(n14854), .A2(n15583), .ZN(n14870) );
  AOI22_X1 U16643 ( .A1(n14870), .A2(n15577), .B1(n15576), .B2(n14855), .ZN(
        n14856) );
  OAI221_X1 U16644 ( .B1(n15625), .B2(n14857), .C1(n15623), .C2(n8388), .A(
        n14856), .ZN(P3_U3221) );
  XNOR2_X1 U16645 ( .A(n14858), .B(n14859), .ZN(n14874) );
  XOR2_X1 U16646 ( .A(n14860), .B(n14859), .Z(n14861) );
  OAI222_X1 U16647 ( .A1(n15588), .A2(n14863), .B1(n15590), .B2(n14862), .C1(
        n14861), .C2(n15594), .ZN(n14872) );
  AOI21_X1 U16648 ( .B1(n14874), .B2(n14864), .A(n14872), .ZN(n14868) );
  NOR2_X1 U16649 ( .A1(n14865), .A2(n15605), .ZN(n14873) );
  AOI22_X1 U16650 ( .A1(n14873), .A2(n15577), .B1(n15576), .B2(n14866), .ZN(
        n14867) );
  OAI221_X1 U16651 ( .B1(n15625), .B2(n14868), .C1(n15623), .C2(n8374), .A(
        n14867), .ZN(P3_U3222) );
  AOI211_X1 U16652 ( .C1(n14871), .C2(n15669), .A(n14870), .B(n14869), .ZN(
        n14875) );
  AOI22_X1 U16653 ( .A1(n15685), .A2(n14875), .B1(n8389), .B2(n8704), .ZN(
        P3_U3471) );
  AOI211_X1 U16654 ( .C1(n14874), .C2(n15669), .A(n14873), .B(n14872), .ZN(
        n14877) );
  AOI22_X1 U16655 ( .A1(n15685), .A2(n14877), .B1(n8375), .B2(n8704), .ZN(
        P3_U3470) );
  INV_X1 U16656 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U16657 ( .A1(n15672), .A2(n14876), .B1(n14875), .B2(n15670), .ZN(
        P3_U3426) );
  INV_X1 U16658 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14878) );
  AOI22_X1 U16659 ( .A1(n15672), .A2(n14878), .B1(n14877), .B2(n15670), .ZN(
        P3_U3423) );
  XNOR2_X1 U16660 ( .A(n14879), .B(n14888), .ZN(n14883) );
  INV_X1 U16661 ( .A(n14880), .ZN(n14881) );
  AOI21_X1 U16662 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14904) );
  AOI222_X1 U16663 ( .A1(n14889), .A2(n15314), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n6674), .C1(n14884), .C2(n15316), .ZN(n14895) );
  INV_X1 U16664 ( .A(n14885), .ZN(n14886) );
  AOI21_X1 U16665 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14907) );
  INV_X1 U16666 ( .A(n14889), .ZN(n14903) );
  INV_X1 U16667 ( .A(n14890), .ZN(n14891) );
  OAI211_X1 U16668 ( .C1(n14903), .C2(n14892), .A(n14891), .B(n9576), .ZN(
        n14902) );
  INV_X1 U16669 ( .A(n14902), .ZN(n14893) );
  AOI22_X1 U16670 ( .A1(n14907), .A2(n15320), .B1(n15319), .B2(n14893), .ZN(
        n14894) );
  OAI211_X1 U16671 ( .C1(n6674), .C2(n14904), .A(n14895), .B(n14894), .ZN(
        P2_U3251) );
  NAND2_X1 U16672 ( .A1(n14896), .A2(n15370), .ZN(n14898) );
  OAI211_X1 U16673 ( .C1(n14899), .C2(n15409), .A(n14898), .B(n14897), .ZN(
        n14901) );
  NOR2_X1 U16674 ( .A1(n14901), .A2(n14900), .ZN(n14923) );
  AOI22_X1 U16675 ( .A1(n15431), .A2(n14923), .B1(n15286), .B2(n15429), .ZN(
        P2_U3514) );
  OAI21_X1 U16676 ( .B1(n14903), .B2(n15409), .A(n14902), .ZN(n14906) );
  INV_X1 U16677 ( .A(n14904), .ZN(n14905) );
  AOI211_X1 U16678 ( .C1(n14907), .C2(n15370), .A(n14906), .B(n14905), .ZN(
        n14925) );
  AOI22_X1 U16679 ( .A1(n15431), .A2(n14925), .B1(n11844), .B2(n15429), .ZN(
        P2_U3513) );
  INV_X1 U16680 ( .A(n14908), .ZN(n14909) );
  OAI21_X1 U16681 ( .B1(n14910), .B2(n15409), .A(n14909), .ZN(n14913) );
  INV_X1 U16682 ( .A(n14911), .ZN(n14912) );
  AOI211_X1 U16683 ( .C1(n15370), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        n14927) );
  AOI22_X1 U16684 ( .A1(n15431), .A2(n14927), .B1(n11685), .B2(n15429), .ZN(
        P2_U3512) );
  OAI21_X1 U16685 ( .B1(n14916), .B2(n15409), .A(n14915), .ZN(n14920) );
  OAI21_X1 U16686 ( .B1(n14918), .B2(n15412), .A(n14917), .ZN(n14919) );
  AOI211_X1 U16687 ( .C1(n15417), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14929) );
  AOI22_X1 U16688 ( .A1(n15431), .A2(n14929), .B1(n11333), .B2(n15429), .ZN(
        P2_U3511) );
  INV_X1 U16689 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U16690 ( .A1(n15420), .A2(n14923), .B1(n14922), .B2(n15418), .ZN(
        P2_U3475) );
  INV_X1 U16691 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16692 ( .A1(n15420), .A2(n14925), .B1(n14924), .B2(n15418), .ZN(
        P2_U3472) );
  INV_X1 U16693 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14926) );
  AOI22_X1 U16694 ( .A1(n15420), .A2(n14927), .B1(n14926), .B2(n15418), .ZN(
        P2_U3469) );
  INV_X1 U16695 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14928) );
  AOI22_X1 U16696 ( .A1(n15420), .A2(n14929), .B1(n14928), .B2(n15418), .ZN(
        P2_U3466) );
  OAI22_X1 U16697 ( .A1(n14972), .A2(n14930), .B1(n14943), .B2(n14969), .ZN(
        n14937) );
  INV_X1 U16698 ( .A(n14209), .ZN(n14933) );
  OAI21_X1 U16699 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14935) );
  AOI21_X1 U16700 ( .B1(n14935), .B2(n14934), .A(n14976), .ZN(n14936) );
  AOI211_X1 U16701 ( .C1(n14981), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14940) );
  OAI211_X1 U16702 ( .C1(n14985), .C2(n14941), .A(n14940), .B(n14939), .ZN(
        P1_U3215) );
  OAI22_X1 U16703 ( .A1(n14972), .A2(n14943), .B1(n14942), .B2(n14969), .ZN(
        n14950) );
  INV_X1 U16704 ( .A(n14247), .ZN(n14946) );
  OAI21_X1 U16705 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14948) );
  AOI21_X1 U16706 ( .B1(n14948), .B2(n14947), .A(n14976), .ZN(n14949) );
  AOI211_X1 U16707 ( .C1(n14981), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14953) );
  OAI211_X1 U16708 ( .C1(n14985), .C2(n14954), .A(n14953), .B(n14952), .ZN(
        P1_U3226) );
  XNOR2_X1 U16709 ( .A(n14956), .B(n14955), .ZN(n14966) );
  AOI22_X1 U16710 ( .A1(n14960), .A2(n14959), .B1(n14958), .B2(n14957), .ZN(
        n14961) );
  OAI21_X1 U16711 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  AOI21_X1 U16712 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14968) );
  OAI211_X1 U16713 ( .C1(n14985), .C2(n14988), .A(n14968), .B(n14967), .ZN(
        P1_U3228) );
  OAI22_X1 U16714 ( .A1(n14972), .A2(n14971), .B1(n14970), .B2(n14969), .ZN(
        n14980) );
  AOI21_X1 U16715 ( .B1(n14133), .B2(n14974), .A(n14973), .ZN(n14975) );
  INV_X1 U16716 ( .A(n14975), .ZN(n14978) );
  AOI21_X1 U16717 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n14979) );
  AOI211_X1 U16718 ( .C1(n14981), .C2(n15013), .A(n14980), .B(n14979), .ZN(
        n14983) );
  OAI211_X1 U16719 ( .C1(n14985), .C2(n14984), .A(n14983), .B(n14982), .ZN(
        P1_U3236) );
  INV_X1 U16720 ( .A(n14986), .ZN(n14996) );
  INV_X1 U16721 ( .A(n14987), .ZN(n14994) );
  INV_X1 U16722 ( .A(n14988), .ZN(n14989) );
  AOI22_X1 U16723 ( .A1(n14991), .A2(n14990), .B1(n14989), .B2(n15099), .ZN(
        n14992) );
  OAI211_X1 U16724 ( .C1(n11216), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14995) );
  AOI21_X1 U16725 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n14998) );
  AOI22_X1 U16726 ( .A1(n15112), .A2(n14999), .B1(n14998), .B2(n15103), .ZN(
        P1_U3276) );
  INV_X1 U16727 ( .A(n15000), .ZN(n15001) );
  OAI21_X1 U16728 ( .B1(n15002), .B2(n15204), .A(n15001), .ZN(n15005) );
  INV_X1 U16729 ( .A(n15003), .ZN(n15004) );
  AOI211_X1 U16730 ( .C1(n15208), .C2(n15006), .A(n15005), .B(n15004), .ZN(
        n15021) );
  AOI22_X1 U16731 ( .A1(n15225), .A2(n15021), .B1(n15007), .B2(n15223), .ZN(
        P1_U3544) );
  OAI21_X1 U16732 ( .B1(n7312), .B2(n15204), .A(n15008), .ZN(n15010) );
  AOI211_X1 U16733 ( .C1(n15011), .C2(n15208), .A(n15010), .B(n15009), .ZN(
        n15023) );
  AOI22_X1 U16734 ( .A1(n15225), .A2(n15023), .B1(n15012), .B2(n15223), .ZN(
        P1_U3542) );
  NAND2_X1 U16735 ( .A1(n15013), .A2(n15156), .ZN(n15015) );
  OAI211_X1 U16736 ( .C1(n15016), .C2(n15146), .A(n15015), .B(n15014), .ZN(
        n15017) );
  NOR2_X1 U16737 ( .A1(n15018), .A2(n15017), .ZN(n15025) );
  AOI22_X1 U16738 ( .A1(n15225), .A2(n15025), .B1(n15019), .B2(n15223), .ZN(
        P1_U3539) );
  INV_X1 U16739 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16740 ( .A1(n15212), .A2(n15021), .B1(n15020), .B2(n15210), .ZN(
        P1_U3507) );
  INV_X1 U16741 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U16742 ( .A1(n15212), .A2(n15023), .B1(n15022), .B2(n15210), .ZN(
        P1_U3501) );
  INV_X1 U16743 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U16744 ( .A1(n15212), .A2(n15025), .B1(n15024), .B2(n15210), .ZN(
        P1_U3492) );
  AOI21_X1 U16745 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15029) );
  XOR2_X1 U16746 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15029), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16747 ( .B1(n6822), .B2(n15031), .A(n15030), .ZN(n15032) );
  XNOR2_X1 U16748 ( .A(n15032), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U16749 ( .A1(n15037), .A2(n15036), .B1(n15037), .B2(n15035), .C1(
        n15034), .C2(n15033), .ZN(SUB_1596_U67) );
  OAI21_X1 U16750 ( .B1(n15040), .B2(n15039), .A(n15038), .ZN(n15041) );
  XNOR2_X1 U16751 ( .A(n15041), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16752 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15045) );
  XOR2_X1 U16753 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15045), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16754 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15049) );
  XOR2_X1 U16755 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15049), .Z(SUB_1596_U64)
         );
  INV_X1 U16756 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15065) );
  OAI21_X1 U16757 ( .B1(n15052), .B2(n15051), .A(n15050), .ZN(n15061) );
  AOI21_X1 U16758 ( .B1(n15054), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15053), 
        .ZN(n15058) );
  OAI22_X1 U16759 ( .A1(n15058), .A2(n15057), .B1(n15056), .B2(n15055), .ZN(
        n15059) );
  AOI21_X1 U16760 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15063) );
  OAI211_X1 U16761 ( .C1(n15065), .C2(n15064), .A(n15063), .B(n15062), .ZN(
        P1_U3258) );
  XNOR2_X1 U16762 ( .A(n15066), .B(n15068), .ZN(n15184) );
  XOR2_X1 U16763 ( .A(n15068), .B(n15067), .Z(n15069) );
  NOR2_X1 U16764 ( .A1(n15069), .A2(n15145), .ZN(n15070) );
  AOI211_X1 U16765 ( .C1(n15072), .C2(n15184), .A(n15071), .B(n15070), .ZN(
        n15181) );
  AOI222_X1 U16766 ( .A1(n15075), .A2(n15074), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n15112), .C1(n15073), .C2(n15099), .ZN(n15083) );
  OAI211_X1 U16767 ( .C1(n15078), .C2(n15180), .A(n15077), .B(n15076), .ZN(
        n15179) );
  INV_X1 U16768 ( .A(n15179), .ZN(n15079) );
  AOI22_X1 U16769 ( .A1(n15081), .A2(n15184), .B1(n15080), .B2(n15079), .ZN(
        n15082) );
  OAI211_X1 U16770 ( .C1(n15112), .C2(n15181), .A(n15083), .B(n15082), .ZN(
        P1_U3287) );
  INV_X1 U16771 ( .A(n15084), .ZN(n15098) );
  INV_X1 U16772 ( .A(n15085), .ZN(n15088) );
  INV_X1 U16773 ( .A(n15086), .ZN(n15087) );
  AOI21_X1 U16774 ( .B1(n15092), .B2(n15088), .A(n15087), .ZN(n15095) );
  INV_X1 U16775 ( .A(n15095), .ZN(n15162) );
  OR2_X1 U16776 ( .A1(n15107), .A2(n15148), .ZN(n15089) );
  AND2_X1 U16777 ( .A1(n15090), .A2(n15089), .ZN(n15154) );
  XNOR2_X1 U16778 ( .A(n10887), .B(n15154), .ZN(n15093) );
  MUX2_X1 U16779 ( .A(n15093), .B(n15092), .S(n15091), .Z(n15094) );
  OAI222_X1 U16780 ( .A1(n15097), .A2(n15096), .B1(n15198), .B2(n15095), .C1(
        n15094), .C2(n15145), .ZN(n15160) );
  AOI21_X1 U16781 ( .B1(n15098), .B2(n15162), .A(n15160), .ZN(n15111) );
  AOI22_X1 U16782 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n15112), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15099), .ZN(n15110) );
  NAND2_X1 U16783 ( .A1(n15100), .A2(n15154), .ZN(n15105) );
  NOR2_X1 U16784 ( .A1(n15102), .A2(n15101), .ZN(n15155) );
  NAND2_X1 U16785 ( .A1(n15103), .A2(n15155), .ZN(n15104) );
  OAI211_X1 U16786 ( .C1(n15107), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n15108) );
  INV_X1 U16787 ( .A(n15108), .ZN(n15109) );
  OAI211_X1 U16788 ( .C1(n15112), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        P1_U3292) );
  INV_X1 U16789 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U16790 ( .A1(n15143), .A2(n15113), .ZN(P1_U3294) );
  INV_X1 U16791 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15114) );
  NOR2_X1 U16792 ( .A1(n15143), .A2(n15114), .ZN(P1_U3295) );
  INV_X1 U16793 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16794 ( .A1(n15143), .A2(n15115), .ZN(P1_U3296) );
  INV_X1 U16795 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15116) );
  NOR2_X1 U16796 ( .A1(n15143), .A2(n15116), .ZN(P1_U3297) );
  INV_X1 U16797 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U16798 ( .A1(n15143), .A2(n15117), .ZN(P1_U3298) );
  INV_X1 U16799 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U16800 ( .A1(n15143), .A2(n15118), .ZN(P1_U3299) );
  INV_X1 U16801 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15119) );
  NOR2_X1 U16802 ( .A1(n15143), .A2(n15119), .ZN(P1_U3300) );
  INV_X1 U16803 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U16804 ( .A1(n15143), .A2(n15120), .ZN(P1_U3301) );
  INV_X1 U16805 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16806 ( .A1(n15143), .A2(n15121), .ZN(P1_U3302) );
  INV_X1 U16807 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U16808 ( .A1(n15143), .A2(n15122), .ZN(P1_U3303) );
  INV_X1 U16809 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U16810 ( .A1(n15143), .A2(n15123), .ZN(P1_U3304) );
  INV_X1 U16811 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16812 ( .A1(n15143), .A2(n15124), .ZN(P1_U3305) );
  INV_X1 U16813 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15125) );
  NOR2_X1 U16814 ( .A1(n15143), .A2(n15125), .ZN(P1_U3306) );
  INV_X1 U16815 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15126) );
  NOR2_X1 U16816 ( .A1(n15143), .A2(n15126), .ZN(P1_U3307) );
  INV_X1 U16817 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16818 ( .A1(n15143), .A2(n15127), .ZN(P1_U3308) );
  INV_X1 U16819 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15128) );
  NOR2_X1 U16820 ( .A1(n15143), .A2(n15128), .ZN(P1_U3309) );
  INV_X1 U16821 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15129) );
  NOR2_X1 U16822 ( .A1(n15143), .A2(n15129), .ZN(P1_U3310) );
  INV_X1 U16823 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15130) );
  NOR2_X1 U16824 ( .A1(n15143), .A2(n15130), .ZN(P1_U3311) );
  INV_X1 U16825 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15131) );
  NOR2_X1 U16826 ( .A1(n15143), .A2(n15131), .ZN(P1_U3312) );
  INV_X1 U16827 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U16828 ( .A1(n15143), .A2(n15132), .ZN(P1_U3313) );
  INV_X1 U16829 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U16830 ( .A1(n15143), .A2(n15133), .ZN(P1_U3314) );
  INV_X1 U16831 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U16832 ( .A1(n15143), .A2(n15134), .ZN(P1_U3315) );
  INV_X1 U16833 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U16834 ( .A1(n15143), .A2(n15135), .ZN(P1_U3316) );
  INV_X1 U16835 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U16836 ( .A1(n15143), .A2(n15136), .ZN(P1_U3317) );
  INV_X1 U16837 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15137) );
  NOR2_X1 U16838 ( .A1(n15143), .A2(n15137), .ZN(P1_U3318) );
  INV_X1 U16839 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15138) );
  NOR2_X1 U16840 ( .A1(n15143), .A2(n15138), .ZN(P1_U3319) );
  INV_X1 U16841 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15139) );
  NOR2_X1 U16842 ( .A1(n15143), .A2(n15139), .ZN(P1_U3320) );
  INV_X1 U16843 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15140) );
  NOR2_X1 U16844 ( .A1(n15143), .A2(n15140), .ZN(P1_U3321) );
  INV_X1 U16845 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15141) );
  NOR2_X1 U16846 ( .A1(n15143), .A2(n15141), .ZN(P1_U3322) );
  INV_X1 U16847 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15142) );
  NOR2_X1 U16848 ( .A1(n15143), .A2(n15142), .ZN(P1_U3323) );
  AOI21_X1 U16849 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15152) );
  INV_X1 U16850 ( .A(n15147), .ZN(n15151) );
  NOR3_X1 U16851 ( .A1(n15149), .A2(n10570), .A3(n15148), .ZN(n15150) );
  NOR3_X1 U16852 ( .A1(n15152), .A2(n15151), .A3(n15150), .ZN(n15214) );
  INV_X1 U16853 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16854 ( .A1(n15212), .A2(n15214), .B1(n15153), .B2(n15210), .ZN(
        P1_U3459) );
  INV_X1 U16855 ( .A(n15154), .ZN(n15158) );
  AOI21_X1 U16856 ( .B1(n15156), .B2(n10603), .A(n15155), .ZN(n15157) );
  OAI21_X1 U16857 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15161) );
  AOI211_X1 U16858 ( .C1(n15185), .C2(n15162), .A(n15161), .B(n15160), .ZN(
        n15216) );
  INV_X1 U16859 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U16860 ( .A1(n15212), .A2(n15216), .B1(n15163), .B2(n15210), .ZN(
        P1_U3462) );
  OAI21_X1 U16861 ( .B1(n15204), .B2(n15165), .A(n15164), .ZN(n15168) );
  INV_X1 U16862 ( .A(n15166), .ZN(n15167) );
  AOI211_X1 U16863 ( .C1(n15208), .C2(n15169), .A(n15168), .B(n15167), .ZN(
        n15217) );
  INV_X1 U16864 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15170) );
  AOI22_X1 U16865 ( .A1(n15212), .A2(n15217), .B1(n15170), .B2(n15210), .ZN(
        P1_U3465) );
  AOI21_X1 U16866 ( .B1(n15198), .B2(n15197), .A(n15171), .ZN(n15177) );
  INV_X1 U16867 ( .A(n15172), .ZN(n15176) );
  OAI21_X1 U16868 ( .B1(n15174), .B2(n15204), .A(n15173), .ZN(n15175) );
  NOR3_X1 U16869 ( .A1(n15177), .A2(n15176), .A3(n15175), .ZN(n15219) );
  INV_X1 U16870 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U16871 ( .A1(n15212), .A2(n15219), .B1(n15178), .B2(n15210), .ZN(
        P1_U3474) );
  OAI21_X1 U16872 ( .B1(n15180), .B2(n15204), .A(n15179), .ZN(n15183) );
  INV_X1 U16873 ( .A(n15181), .ZN(n15182) );
  AOI211_X1 U16874 ( .C1(n15185), .C2(n15184), .A(n15183), .B(n15182), .ZN(
        n15220) );
  INV_X1 U16875 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U16876 ( .A1(n15212), .A2(n15220), .B1(n15186), .B2(n15210), .ZN(
        P1_U3477) );
  AOI21_X1 U16877 ( .B1(n15198), .B2(n15197), .A(n15187), .ZN(n15190) );
  NOR4_X1 U16878 ( .A1(n15191), .A2(n15190), .A3(n15189), .A4(n15188), .ZN(
        n15221) );
  INV_X1 U16879 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U16880 ( .A1(n15212), .A2(n15221), .B1(n15192), .B2(n15210), .ZN(
        P1_U3480) );
  OAI211_X1 U16881 ( .C1(n15195), .C2(n15204), .A(n15194), .B(n15193), .ZN(
        n15200) );
  AOI21_X1 U16882 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15199) );
  NOR2_X1 U16883 ( .A1(n15200), .A2(n15199), .ZN(n15222) );
  INV_X1 U16884 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15201) );
  AOI22_X1 U16885 ( .A1(n15212), .A2(n15222), .B1(n15201), .B2(n15210), .ZN(
        P1_U3486) );
  OAI211_X1 U16886 ( .C1(n15205), .C2(n15204), .A(n15203), .B(n15202), .ZN(
        n15207) );
  AOI211_X1 U16887 ( .C1(n15209), .C2(n15208), .A(n15207), .B(n15206), .ZN(
        n15224) );
  INV_X1 U16888 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15211) );
  AOI22_X1 U16889 ( .A1(n15212), .A2(n15224), .B1(n15211), .B2(n15210), .ZN(
        P1_U3489) );
  INV_X1 U16890 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15213) );
  AOI22_X1 U16891 ( .A1(n15225), .A2(n15214), .B1(n15213), .B2(n15223), .ZN(
        P1_U3528) );
  INV_X1 U16892 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U16893 ( .A1(n15225), .A2(n15216), .B1(n15215), .B2(n15223), .ZN(
        P1_U3529) );
  AOI22_X1 U16894 ( .A1(n15225), .A2(n15217), .B1(n10349), .B2(n15223), .ZN(
        P1_U3530) );
  AOI22_X1 U16895 ( .A1(n15225), .A2(n15219), .B1(n15218), .B2(n15223), .ZN(
        P1_U3533) );
  AOI22_X1 U16896 ( .A1(n15225), .A2(n15220), .B1(n10469), .B2(n15223), .ZN(
        P1_U3534) );
  AOI22_X1 U16897 ( .A1(n15225), .A2(n15221), .B1(n10471), .B2(n15223), .ZN(
        P1_U3535) );
  AOI22_X1 U16898 ( .A1(n15225), .A2(n15222), .B1(n10473), .B2(n15223), .ZN(
        P1_U3537) );
  AOI22_X1 U16899 ( .A1(n15225), .A2(n15224), .B1(n10474), .B2(n15223), .ZN(
        P1_U3538) );
  NOR2_X1 U16900 ( .A1(n15289), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16901 ( .A1(n15289), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15243) );
  NAND2_X1 U16902 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15229) );
  INV_X1 U16903 ( .A(n15226), .ZN(n15228) );
  AOI211_X1 U16904 ( .C1(n15229), .C2(n15228), .A(n15227), .B(n15298), .ZN(
        n15234) );
  NOR3_X1 U16905 ( .A1(n15232), .A2(n15231), .A3(n15230), .ZN(n15233) );
  NOR2_X1 U16906 ( .A1(n15234), .A2(n15233), .ZN(n15242) );
  NOR2_X1 U16907 ( .A1(n15236), .A2(n15235), .ZN(n15239) );
  INV_X1 U16908 ( .A(n15237), .ZN(n15238) );
  OAI211_X1 U16909 ( .C1(n15240), .C2(n15239), .A(n15307), .B(n15238), .ZN(
        n15241) );
  NAND3_X1 U16910 ( .A1(n15243), .A2(n15242), .A3(n15241), .ZN(P2_U3215) );
  AOI22_X1 U16911 ( .A1(n15289), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15255) );
  AOI211_X1 U16912 ( .C1(n15246), .C2(n15245), .A(n15244), .B(n15298), .ZN(
        n15247) );
  AOI21_X1 U16913 ( .B1(n15305), .B2(n15248), .A(n15247), .ZN(n15254) );
  AOI211_X1 U16914 ( .C1(n15251), .C2(n15250), .A(n15249), .B(n15279), .ZN(
        n15252) );
  INV_X1 U16915 ( .A(n15252), .ZN(n15253) );
  NAND3_X1 U16916 ( .A1(n15255), .A2(n15254), .A3(n15253), .ZN(P2_U3216) );
  OAI21_X1 U16917 ( .B1(n15258), .B2(n15257), .A(n15256), .ZN(n15259) );
  INV_X1 U16918 ( .A(n15259), .ZN(n15270) );
  OAI21_X1 U16919 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15266) );
  INV_X1 U16920 ( .A(n15263), .ZN(n15264) );
  AOI21_X1 U16921 ( .B1(n15266), .B2(n15265), .A(n15264), .ZN(n15269) );
  AOI22_X1 U16922 ( .A1(n15305), .A2(n15267), .B1(n15289), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n15268) );
  OAI211_X1 U16923 ( .C1(n15270), .C2(n15279), .A(n15269), .B(n15268), .ZN(
        P2_U3223) );
  NOR2_X1 U16924 ( .A1(n15272), .A2(n15271), .ZN(n15277) );
  AOI211_X1 U16925 ( .C1(n15275), .C2(n15274), .A(n15298), .B(n15273), .ZN(
        n15276) );
  AOI211_X1 U16926 ( .C1(n15289), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n15277), 
        .B(n15276), .ZN(n15284) );
  AOI211_X1 U16927 ( .C1(n15281), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        n15282) );
  INV_X1 U16928 ( .A(n15282), .ZN(n15283) );
  OAI211_X1 U16929 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9343), .A(n15284), .B(
        n15283), .ZN(P2_U3224) );
  AOI211_X1 U16930 ( .C1(n15287), .C2(n15286), .A(n15285), .B(n15298), .ZN(
        n15288) );
  AOI21_X1 U16931 ( .B1(n15289), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n15288), 
        .ZN(n15296) );
  OAI211_X1 U16932 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15291), .A(n15307), 
        .B(n15290), .ZN(n15294) );
  NAND2_X1 U16933 ( .A1(n15305), .A2(n15292), .ZN(n15293) );
  NAND4_X1 U16934 ( .A1(n15296), .A2(n15295), .A3(n15294), .A4(n15293), .ZN(
        P2_U3229) );
  NOR2_X1 U16935 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15297), .ZN(n15303) );
  AOI211_X1 U16936 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        n15302) );
  AOI211_X1 U16937 ( .C1(n15305), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15311) );
  OAI211_X1 U16938 ( .C1(n15309), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        n15310) );
  OAI211_X1 U16939 ( .C1(n15313), .C2(n15312), .A(n15311), .B(n15310), .ZN(
        P2_U3231) );
  AOI222_X1 U16940 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n6674), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15316), .C1(n15315), .C2(n15314), .ZN(
        n15323) );
  INV_X1 U16941 ( .A(n15317), .ZN(n15318) );
  AOI22_X1 U16942 ( .A1(n15321), .A2(n15320), .B1(n15319), .B2(n15318), .ZN(
        n15322) );
  OAI211_X1 U16943 ( .C1(n6674), .C2(n15324), .A(n15323), .B(n15322), .ZN(
        P2_U3263) );
  INV_X1 U16944 ( .A(n15362), .ZN(n15359) );
  NOR2_X4 U16945 ( .A1(n15325), .A2(n15359), .ZN(n15353) );
  INV_X1 U16946 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U16947 ( .A1(n15353), .A2(n15326), .ZN(P2_U3266) );
  INV_X1 U16948 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15327) );
  NOR2_X1 U16949 ( .A1(n15353), .A2(n15327), .ZN(P2_U3267) );
  INV_X1 U16950 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15328) );
  NOR2_X1 U16951 ( .A1(n15353), .A2(n15328), .ZN(P2_U3268) );
  INV_X1 U16952 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U16953 ( .A1(n15353), .A2(n15329), .ZN(P2_U3269) );
  INV_X1 U16954 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15330) );
  NOR2_X1 U16955 ( .A1(n15353), .A2(n15330), .ZN(P2_U3270) );
  INV_X1 U16956 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U16957 ( .A1(n15353), .A2(n15331), .ZN(P2_U3271) );
  INV_X1 U16958 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U16959 ( .A1(n15353), .A2(n15332), .ZN(P2_U3272) );
  INV_X1 U16960 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16961 ( .A1(n15353), .A2(n15333), .ZN(P2_U3273) );
  INV_X1 U16962 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U16963 ( .A1(n15353), .A2(n15334), .ZN(P2_U3274) );
  INV_X1 U16964 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16965 ( .A1(n15353), .A2(n15335), .ZN(P2_U3275) );
  INV_X1 U16966 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U16967 ( .A1(n15353), .A2(n15336), .ZN(P2_U3276) );
  INV_X1 U16968 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16969 ( .A1(n15353), .A2(n15337), .ZN(P2_U3277) );
  INV_X1 U16970 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U16971 ( .A1(n15353), .A2(n15338), .ZN(P2_U3278) );
  INV_X1 U16972 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16973 ( .A1(n15353), .A2(n15339), .ZN(P2_U3279) );
  INV_X1 U16974 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U16975 ( .A1(n15353), .A2(n15340), .ZN(P2_U3280) );
  INV_X1 U16976 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U16977 ( .A1(n15353), .A2(n15341), .ZN(P2_U3281) );
  INV_X1 U16978 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U16979 ( .A1(n15353), .A2(n15342), .ZN(P2_U3282) );
  INV_X1 U16980 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16981 ( .A1(n15353), .A2(n15343), .ZN(P2_U3283) );
  INV_X1 U16982 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15344) );
  NOR2_X1 U16983 ( .A1(n15353), .A2(n15344), .ZN(P2_U3284) );
  INV_X1 U16984 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15345) );
  NOR2_X1 U16985 ( .A1(n15353), .A2(n15345), .ZN(P2_U3285) );
  INV_X1 U16986 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15346) );
  NOR2_X1 U16987 ( .A1(n15353), .A2(n15346), .ZN(P2_U3286) );
  INV_X1 U16988 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16989 ( .A1(n15353), .A2(n15347), .ZN(P2_U3287) );
  INV_X1 U16990 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U16991 ( .A1(n15353), .A2(n15348), .ZN(P2_U3288) );
  INV_X1 U16992 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16993 ( .A1(n15353), .A2(n15349), .ZN(P2_U3289) );
  INV_X1 U16994 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U16995 ( .A1(n15353), .A2(n15350), .ZN(P2_U3290) );
  INV_X1 U16996 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U16997 ( .A1(n15353), .A2(n15351), .ZN(P2_U3291) );
  INV_X1 U16998 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16999 ( .A1(n15353), .A2(n15352), .ZN(P2_U3292) );
  INV_X1 U17000 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U17001 ( .A1(n15353), .A2(n15354), .ZN(P2_U3293) );
  INV_X1 U17002 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15355) );
  NOR2_X1 U17003 ( .A1(n15353), .A2(n15355), .ZN(P2_U3294) );
  INV_X1 U17004 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15356) );
  NOR2_X1 U17005 ( .A1(n15353), .A2(n15356), .ZN(P2_U3295) );
  INV_X1 U17006 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15358) );
  OAI21_X1 U17007 ( .B1(n15362), .B2(n15358), .A(n15357), .ZN(P2_U3416) );
  INV_X1 U17008 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15360) );
  AOI22_X1 U17009 ( .A1(n15362), .A2(n15361), .B1(n15360), .B2(n15359), .ZN(
        P2_U3417) );
  INV_X1 U17010 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U17011 ( .A1(n15420), .A2(n15364), .B1(n15363), .B2(n15418), .ZN(
        P2_U3430) );
  OAI21_X1 U17012 ( .B1(n15409), .B2(n15366), .A(n15365), .ZN(n15369) );
  INV_X1 U17013 ( .A(n15367), .ZN(n15368) );
  AOI211_X1 U17014 ( .C1(n15371), .C2(n15370), .A(n15369), .B(n15368), .ZN(
        n15422) );
  INV_X1 U17015 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U17016 ( .A1(n15420), .A2(n15422), .B1(n15372), .B2(n15418), .ZN(
        P2_U3433) );
  INV_X1 U17017 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U17018 ( .A1(n15420), .A2(n15374), .B1(n15373), .B2(n15418), .ZN(
        P2_U3436) );
  AOI21_X1 U17019 ( .B1(n15412), .B2(n15401), .A(n15375), .ZN(n15381) );
  INV_X1 U17020 ( .A(n15376), .ZN(n15377) );
  OAI211_X1 U17021 ( .C1(n15379), .C2(n15409), .A(n15378), .B(n15377), .ZN(
        n15380) );
  NOR2_X1 U17022 ( .A1(n15381), .A2(n15380), .ZN(n15424) );
  INV_X1 U17023 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U17024 ( .A1(n15420), .A2(n15424), .B1(n15382), .B2(n15418), .ZN(
        P2_U3439) );
  AOI21_X1 U17025 ( .B1(n15412), .B2(n15401), .A(n15383), .ZN(n15388) );
  OAI211_X1 U17026 ( .C1(n15386), .C2(n15409), .A(n15385), .B(n15384), .ZN(
        n15387) );
  NOR2_X1 U17027 ( .A1(n15388), .A2(n15387), .ZN(n15426) );
  INV_X1 U17028 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U17029 ( .A1(n15420), .A2(n15426), .B1(n15389), .B2(n15418), .ZN(
        P2_U3445) );
  OAI21_X1 U17030 ( .B1(n15391), .B2(n15409), .A(n15390), .ZN(n15392) );
  AOI21_X1 U17031 ( .B1(n15393), .B2(n15417), .A(n15392), .ZN(n15394) );
  INV_X1 U17032 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U17033 ( .A1(n15420), .A2(n15427), .B1(n15396), .B2(n15418), .ZN(
        P2_U3454) );
  INV_X1 U17034 ( .A(n15402), .ZN(n15405) );
  AOI21_X1 U17035 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(n15400) );
  OAI21_X1 U17036 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15404) );
  AOI211_X1 U17037 ( .C1(n15406), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        n15428) );
  INV_X1 U17038 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U17039 ( .A1(n15420), .A2(n15428), .B1(n15407), .B2(n15418), .ZN(
        P2_U3457) );
  OAI21_X1 U17040 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(n15415) );
  OAI21_X1 U17041 ( .B1(n15413), .B2(n15412), .A(n15411), .ZN(n15414) );
  AOI211_X1 U17042 ( .C1(n15417), .C2(n15416), .A(n15415), .B(n15414), .ZN(
        n15430) );
  INV_X1 U17043 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U17044 ( .A1(n15420), .A2(n15430), .B1(n15419), .B2(n15418), .ZN(
        P2_U3463) );
  INV_X1 U17045 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U17046 ( .A1(n15431), .A2(n15422), .B1(n15421), .B2(n15429), .ZN(
        P2_U3500) );
  INV_X1 U17047 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U17048 ( .A1(n15431), .A2(n15424), .B1(n15423), .B2(n15429), .ZN(
        P2_U3502) );
  INV_X1 U17049 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U17050 ( .A1(n15431), .A2(n15426), .B1(n15425), .B2(n15429), .ZN(
        P2_U3504) );
  AOI22_X1 U17051 ( .A1(n15431), .A2(n15427), .B1(n10394), .B2(n15429), .ZN(
        P2_U3507) );
  AOI22_X1 U17052 ( .A1(n15431), .A2(n15428), .B1(n11100), .B2(n15429), .ZN(
        P2_U3508) );
  AOI22_X1 U17053 ( .A1(n15431), .A2(n15430), .B1(n11102), .B2(n15429), .ZN(
        P2_U3510) );
  NOR2_X1 U17054 ( .A1(P3_U3897), .A2(n15516), .ZN(P3_U3150) );
  AOI21_X1 U17055 ( .B1(n15564), .B2(n15433), .A(n15432), .ZN(n15448) );
  INV_X1 U17056 ( .A(n15453), .ZN(n15437) );
  OR2_X1 U17057 ( .A1(n15434), .A2(n15453), .ZN(n15435) );
  AOI22_X1 U17058 ( .A1(n15454), .A2(n15437), .B1(n15436), .B2(n15435), .ZN(
        n15440) );
  OAI22_X1 U17059 ( .A1(n15440), .A2(n15439), .B1(n15438), .B2(n15513), .ZN(
        n15441) );
  AOI211_X1 U17060 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15516), .A(n15442), .B(
        n15441), .ZN(n15447) );
  OAI21_X1 U17061 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15444), .A(n15443), .ZN(
        n15445) );
  NAND2_X1 U17062 ( .A1(n15519), .A2(n15445), .ZN(n15446) );
  OAI211_X1 U17063 ( .C1(n15448), .C2(n15523), .A(n15447), .B(n15446), .ZN(
        P3_U3187) );
  AOI21_X1 U17064 ( .B1(n15451), .B2(n15450), .A(n15449), .ZN(n15467) );
  INV_X1 U17065 ( .A(n15472), .ZN(n15456) );
  NOR3_X1 U17066 ( .A1(n15454), .A2(n15453), .A3(n15452), .ZN(n15455) );
  OAI21_X1 U17067 ( .B1(n15456), .B2(n15455), .A(n15508), .ZN(n15457) );
  OAI21_X1 U17068 ( .B1(n15513), .B2(n15458), .A(n15457), .ZN(n15459) );
  AOI211_X1 U17069 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15516), .A(n15460), .B(
        n15459), .ZN(n15466) );
  OAI21_X1 U17070 ( .B1(n15463), .B2(n15462), .A(n15461), .ZN(n15464) );
  NAND2_X1 U17071 ( .A1(n15464), .A2(n15519), .ZN(n15465) );
  OAI211_X1 U17072 ( .C1(n15467), .C2(n15523), .A(n15466), .B(n15465), .ZN(
        P3_U3188) );
  AOI21_X1 U17073 ( .B1(n11152), .B2(n15469), .A(n15468), .ZN(n15483) );
  AND3_X1 U17074 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n15473) );
  OAI21_X1 U17075 ( .B1(n15489), .B2(n15473), .A(n15508), .ZN(n15474) );
  OAI21_X1 U17076 ( .B1(n15513), .B2(n15475), .A(n15474), .ZN(n15476) );
  AOI211_X1 U17077 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15516), .A(n15477), .B(
        n15476), .ZN(n15482) );
  OAI21_X1 U17078 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15479), .A(n15478), .ZN(
        n15480) );
  NAND2_X1 U17079 ( .A1(n15480), .A2(n15519), .ZN(n15481) );
  OAI211_X1 U17080 ( .C1(n15483), .C2(n15523), .A(n15482), .B(n15481), .ZN(
        P3_U3189) );
  AOI21_X1 U17081 ( .B1(n15486), .B2(n15485), .A(n15484), .ZN(n15502) );
  INV_X1 U17082 ( .A(n15507), .ZN(n15491) );
  NOR3_X1 U17083 ( .A1(n15489), .A2(n15488), .A3(n15487), .ZN(n15490) );
  OAI21_X1 U17084 ( .B1(n15491), .B2(n15490), .A(n15508), .ZN(n15492) );
  OAI21_X1 U17085 ( .B1(n15513), .B2(n15493), .A(n15492), .ZN(n15494) );
  AOI211_X1 U17086 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15516), .A(n15495), .B(
        n15494), .ZN(n15501) );
  OAI21_X1 U17087 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15499) );
  NAND2_X1 U17088 ( .A1(n15499), .A2(n15519), .ZN(n15500) );
  OAI211_X1 U17089 ( .C1(n15502), .C2(n15523), .A(n15501), .B(n15500), .ZN(
        P3_U3190) );
  AOI21_X1 U17090 ( .B1(n11165), .B2(n15504), .A(n15503), .ZN(n15524) );
  AND3_X1 U17091 ( .A1(n15507), .A2(n15506), .A3(n15505), .ZN(n15509) );
  OAI21_X1 U17092 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n15511) );
  OAI21_X1 U17093 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15514) );
  AOI211_X1 U17094 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15516), .A(n15515), .B(
        n15514), .ZN(n15522) );
  OAI21_X1 U17095 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15518), .A(n15517), .ZN(
        n15520) );
  NAND2_X1 U17096 ( .A1(n15520), .A2(n15519), .ZN(n15521) );
  OAI211_X1 U17097 ( .C1(n15524), .C2(n15523), .A(n15522), .B(n15521), .ZN(
        P3_U3191) );
  NAND2_X1 U17098 ( .A1(n15526), .A2(n15525), .ZN(n15527) );
  XNOR2_X1 U17099 ( .A(n15527), .B(n8370), .ZN(n15530) );
  AOI222_X1 U17100 ( .A1(n15612), .A2(n15530), .B1(n15529), .B2(n15607), .C1(
        n15528), .C2(n15610), .ZN(n15665) );
  AOI22_X1 U17101 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15625), .B1(n15576), 
        .B2(n15531), .ZN(n15537) );
  XNOR2_X1 U17102 ( .A(n15533), .B(n15532), .ZN(n15668) );
  NOR2_X1 U17103 ( .A1(n15534), .A2(n15605), .ZN(n15667) );
  AOI22_X1 U17104 ( .A1(n15668), .A2(n15535), .B1(n15577), .B2(n15667), .ZN(
        n15536) );
  OAI211_X1 U17105 ( .C1(n15625), .C2(n15665), .A(n15537), .B(n15536), .ZN(
        P3_U3223) );
  XNOR2_X1 U17106 ( .A(n15538), .B(n15539), .ZN(n15653) );
  XNOR2_X1 U17107 ( .A(n15541), .B(n15540), .ZN(n15545) );
  OAI22_X1 U17108 ( .A1(n15542), .A2(n15588), .B1(n15555), .B2(n15590), .ZN(
        n15543) );
  AOI21_X1 U17109 ( .B1(n15653), .B2(n15599), .A(n15543), .ZN(n15544) );
  OAI21_X1 U17110 ( .B1(n15545), .B2(n15594), .A(n15544), .ZN(n15651) );
  AOI21_X1 U17111 ( .B1(n15602), .B2(n15653), .A(n15651), .ZN(n15550) );
  NOR2_X1 U17112 ( .A1(n15546), .A2(n15605), .ZN(n15652) );
  INV_X1 U17113 ( .A(n15547), .ZN(n15548) );
  AOI22_X1 U17114 ( .A1(n15577), .A2(n15652), .B1(n15576), .B2(n15548), .ZN(
        n15549) );
  OAI221_X1 U17115 ( .B1(n15625), .B2(n15550), .C1(n15623), .C2(n11152), .A(
        n15549), .ZN(P3_U3226) );
  XNOR2_X1 U17116 ( .A(n15551), .B(n15553), .ZN(n15560) );
  INV_X1 U17117 ( .A(n15560), .ZN(n15644) );
  OAI21_X1 U17118 ( .B1(n15554), .B2(n15553), .A(n15552), .ZN(n15558) );
  OAI22_X1 U17119 ( .A1(n15556), .A2(n15590), .B1(n15555), .B2(n15588), .ZN(
        n15557) );
  AOI21_X1 U17120 ( .B1(n15558), .B2(n15612), .A(n15557), .ZN(n15559) );
  OAI21_X1 U17121 ( .B1(n15616), .B2(n15560), .A(n15559), .ZN(n15642) );
  AOI21_X1 U17122 ( .B1(n15602), .B2(n15644), .A(n15642), .ZN(n15565) );
  NOR2_X1 U17123 ( .A1(n15561), .A2(n15605), .ZN(n15643) );
  AOI22_X1 U17124 ( .A1(n15577), .A2(n15643), .B1(n15576), .B2(n15562), .ZN(
        n15563) );
  OAI221_X1 U17125 ( .B1(n15625), .B2(n15565), .C1(n15623), .C2(n15564), .A(
        n15563), .ZN(P3_U3228) );
  XNOR2_X1 U17126 ( .A(n15567), .B(n15566), .ZN(n15640) );
  XNOR2_X1 U17127 ( .A(n15569), .B(n15568), .ZN(n15573) );
  OAI22_X1 U17128 ( .A1(n15589), .A2(n15590), .B1(n15570), .B2(n15588), .ZN(
        n15571) );
  AOI21_X1 U17129 ( .B1(n15640), .B2(n15599), .A(n15571), .ZN(n15572) );
  OAI21_X1 U17130 ( .B1(n15594), .B2(n15573), .A(n15572), .ZN(n15638) );
  AOI21_X1 U17131 ( .B1(n15602), .B2(n15640), .A(n15638), .ZN(n15579) );
  NOR2_X1 U17132 ( .A1(n15574), .A2(n15605), .ZN(n15639) );
  AOI22_X1 U17133 ( .A1(n15577), .A2(n15639), .B1(n15576), .B2(n15575), .ZN(
        n15578) );
  OAI221_X1 U17134 ( .B1(n15625), .B2(n15579), .C1(n15623), .C2(n8268), .A(
        n15578), .ZN(P3_U3229) );
  OAI21_X1 U17135 ( .B1(n15581), .B2(n15593), .A(n15580), .ZN(n15633) );
  INV_X1 U17136 ( .A(n15582), .ZN(n15584) );
  NAND2_X1 U17137 ( .A1(n15584), .A2(n15583), .ZN(n15630) );
  OAI22_X1 U17138 ( .A1(n15618), .A2(n15586), .B1(n15630), .B2(n15585), .ZN(
        n15601) );
  OAI22_X1 U17139 ( .A1(n7689), .A2(n15590), .B1(n15589), .B2(n15588), .ZN(
        n15598) );
  NAND3_X1 U17140 ( .A1(n15591), .A2(n15593), .A3(n15592), .ZN(n15595) );
  AOI21_X1 U17141 ( .B1(n15596), .B2(n15595), .A(n15594), .ZN(n15597) );
  AOI211_X1 U17142 ( .C1(n15599), .C2(n15633), .A(n15598), .B(n15597), .ZN(
        n15600) );
  INV_X1 U17143 ( .A(n15600), .ZN(n15631) );
  AOI211_X1 U17144 ( .C1(n15602), .C2(n15633), .A(n15601), .B(n15631), .ZN(
        n15603) );
  AOI22_X1 U17145 ( .A1(n15625), .A2(n15604), .B1(n15603), .B2(n15623), .ZN(
        P3_U3231) );
  NOR2_X1 U17146 ( .A1(n15606), .A2(n15605), .ZN(n15628) );
  XNOR2_X1 U17147 ( .A(n10413), .B(n15611), .ZN(n15626) );
  AOI22_X1 U17148 ( .A1(n15610), .A2(n15609), .B1(n15608), .B2(n15607), .ZN(
        n15615) );
  NAND2_X1 U17149 ( .A1(n15613), .A2(n15612), .ZN(n15614) );
  OAI211_X1 U17150 ( .C1(n15626), .C2(n15616), .A(n15615), .B(n15614), .ZN(
        n15627) );
  AOI21_X1 U17151 ( .B1(n15628), .B2(n15617), .A(n15627), .ZN(n15624) );
  OAI22_X1 U17152 ( .A1(n15626), .A2(n15620), .B1(n15619), .B2(n15618), .ZN(
        n15621) );
  INV_X1 U17153 ( .A(n15621), .ZN(n15622) );
  OAI221_X1 U17154 ( .B1(n15625), .B2(n15624), .C1(n15623), .C2(n8223), .A(
        n15622), .ZN(P3_U3232) );
  INV_X1 U17155 ( .A(n15626), .ZN(n15629) );
  AOI211_X1 U17156 ( .C1(n15662), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15673) );
  AOI22_X1 U17157 ( .A1(n15672), .A2(n8222), .B1(n15673), .B2(n15670), .ZN(
        P3_U3393) );
  INV_X1 U17158 ( .A(n15630), .ZN(n15632) );
  AOI211_X1 U17159 ( .C1(n15662), .C2(n15633), .A(n15632), .B(n15631), .ZN(
        n15674) );
  AOI22_X1 U17160 ( .A1(n15672), .A2(n8244), .B1(n15674), .B2(n15670), .ZN(
        P3_U3396) );
  INV_X1 U17161 ( .A(n15634), .ZN(n15637) );
  AOI211_X1 U17162 ( .C1(n15637), .C2(n15662), .A(n15636), .B(n15635), .ZN(
        n15675) );
  AOI22_X1 U17163 ( .A1(n15672), .A2(n7002), .B1(n15675), .B2(n15670), .ZN(
        P3_U3399) );
  INV_X1 U17164 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15641) );
  AOI211_X1 U17165 ( .C1(n15640), .C2(n15662), .A(n15639), .B(n15638), .ZN(
        n15677) );
  AOI22_X1 U17166 ( .A1(n15672), .A2(n15641), .B1(n15677), .B2(n15670), .ZN(
        P3_U3402) );
  INV_X1 U17167 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15645) );
  AOI211_X1 U17168 ( .C1(n15644), .C2(n15662), .A(n15643), .B(n15642), .ZN(
        n15679) );
  AOI22_X1 U17169 ( .A1(n15672), .A2(n15645), .B1(n15679), .B2(n15670), .ZN(
        P3_U3405) );
  INV_X1 U17170 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15650) );
  INV_X1 U17171 ( .A(n15646), .ZN(n15648) );
  AOI211_X1 U17172 ( .C1(n15649), .C2(n15662), .A(n15648), .B(n15647), .ZN(
        n15680) );
  AOI22_X1 U17173 ( .A1(n15672), .A2(n15650), .B1(n15680), .B2(n15670), .ZN(
        P3_U3408) );
  INV_X1 U17174 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15654) );
  AOI211_X1 U17175 ( .C1(n15653), .C2(n15662), .A(n15652), .B(n15651), .ZN(
        n15681) );
  AOI22_X1 U17176 ( .A1(n15672), .A2(n15654), .B1(n15681), .B2(n15670), .ZN(
        P3_U3411) );
  INV_X1 U17177 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15659) );
  INV_X1 U17178 ( .A(n15655), .ZN(n15657) );
  AOI211_X1 U17179 ( .C1(n15662), .C2(n15658), .A(n15657), .B(n15656), .ZN(
        n15682) );
  AOI22_X1 U17180 ( .A1(n15672), .A2(n15659), .B1(n15682), .B2(n15670), .ZN(
        P3_U3414) );
  INV_X1 U17181 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15664) );
  AOI211_X1 U17182 ( .C1(n15663), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15683) );
  AOI22_X1 U17183 ( .A1(n15672), .A2(n15664), .B1(n15683), .B2(n15670), .ZN(
        P3_U3417) );
  INV_X1 U17184 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15671) );
  INV_X1 U17185 ( .A(n15665), .ZN(n15666) );
  AOI211_X1 U17186 ( .C1(n15669), .C2(n15668), .A(n15667), .B(n15666), .ZN(
        n15684) );
  AOI22_X1 U17187 ( .A1(n15672), .A2(n15671), .B1(n15684), .B2(n15670), .ZN(
        P3_U3420) );
  AOI22_X1 U17188 ( .A1(n15685), .A2(n15673), .B1(n10685), .B2(n8704), .ZN(
        P3_U3460) );
  AOI22_X1 U17189 ( .A1(n15685), .A2(n15674), .B1(n10750), .B2(n8704), .ZN(
        P3_U3461) );
  AOI22_X1 U17190 ( .A1(n15685), .A2(n15675), .B1(n10770), .B2(n8704), .ZN(
        P3_U3462) );
  AOI22_X1 U17191 ( .A1(n15685), .A2(n15677), .B1(n15676), .B2(n8704), .ZN(
        P3_U3463) );
  AOI22_X1 U17192 ( .A1(n15685), .A2(n15679), .B1(n15678), .B2(n8704), .ZN(
        P3_U3464) );
  AOI22_X1 U17193 ( .A1(n15685), .A2(n15680), .B1(n11145), .B2(n8704), .ZN(
        P3_U3465) );
  AOI22_X1 U17194 ( .A1(n15685), .A2(n15681), .B1(n11151), .B2(n8704), .ZN(
        P3_U3466) );
  AOI22_X1 U17195 ( .A1(n15685), .A2(n15682), .B1(n11158), .B2(n8704), .ZN(
        P3_U3467) );
  AOI22_X1 U17196 ( .A1(n15685), .A2(n15683), .B1(n11164), .B2(n8704), .ZN(
        P3_U3468) );
  AOI22_X1 U17197 ( .A1(n15685), .A2(n15684), .B1(n11171), .B2(n8704), .ZN(
        P3_U3469) );
  AOI21_X1 U17198 ( .B1(n15688), .B2(n15687), .A(n15686), .ZN(SUB_1596_U59) );
  OAI21_X1 U17199 ( .B1(n15691), .B2(n15690), .A(n15689), .ZN(SUB_1596_U58) );
  XOR2_X1 U17200 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15692), .Z(SUB_1596_U53) );
  AOI21_X1 U17201 ( .B1(n15695), .B2(n15694), .A(n15693), .ZN(SUB_1596_U56) );
  OAI21_X1 U17202 ( .B1(n15698), .B2(n15697), .A(n15696), .ZN(n15699) );
  XNOR2_X1 U17203 ( .A(n15699), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17204 ( .B1(n15702), .B2(n15701), .A(n15700), .ZN(SUB_1596_U5) );
  BUF_X1 U7512 ( .A(n10817), .Z(n12726) );
  NAND2_X1 U7728 ( .A1(n14527), .A2(n6670), .ZN(n11216) );
  CLKBUF_X1 U7445 ( .A(n12125), .Z(n12156) );
  CLKBUF_X1 U7486 ( .A(n10818), .Z(n12116) );
  INV_X2 U7530 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n12177) );
  CLKBUF_X1 U7536 ( .A(n12052), .Z(n6671) );
  OAI211_X1 U7747 ( .C1(n10594), .C2(n11914), .A(n6742), .B(n10598), .ZN(
        n10603) );
endmodule

