

module b20_C_AntiSAT_k_256_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738;

  AOI21_X1 U5047 ( .B1(n4911), .B2(n4570), .A(n4910), .ZN(n10306) );
  OR2_X1 U5048 ( .A1(n7227), .A2(n4631), .ZN(n4752) );
  INV_X1 U5049 ( .A(n9795), .ZN(n9941) );
  CLKBUF_X1 U5050 ( .A(n6767), .Z(n8798) );
  BUF_X2 U5052 ( .A(n6299), .Z(n4541) );
  BUF_X1 U5053 ( .A(n6487), .Z(n4547) );
  AND2_X1 U5054 ( .A1(n10188), .A2(n9677), .ZN(n10175) );
  INV_X1 U5055 ( .A(n5454), .ZN(n5639) );
  NAND2_X1 U5056 ( .A1(n6778), .A2(n6585), .ZN(n6277) );
  NAND2_X1 U5057 ( .A1(n8691), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8690) );
  OR2_X1 U5058 ( .A1(n6261), .A2(n9518), .ZN(n6263) );
  INV_X1 U5059 ( .A(n4553), .ZN(n5747) );
  NAND2_X1 U5060 ( .A1(n8441), .A2(n5846), .ZN(n5847) );
  AND2_X1 U5061 ( .A1(n5820), .A2(n9918), .ZN(n5888) );
  OAI22_X2 U5062 ( .A1(n10201), .A2(n5665), .B1(n10209), .B2(n9806), .ZN(
        n10187) );
  INV_X1 U5063 ( .A(n9690), .ZN(n10602) );
  INV_X1 U5064 ( .A(n7313), .ZN(n7513) );
  BUF_X1 U5065 ( .A(n6277), .Z(n8172) );
  NAND2_X1 U5066 ( .A1(n5086), .A2(n5085), .ZN(n9450) );
  NAND2_X1 U5069 ( .A1(n6527), .A2(n6526), .ZN(n8656) );
  INV_X1 U5071 ( .A(n8172), .ZN(n6487) );
  INV_X1 U5072 ( .A(n6112), .ZN(n4544) );
  NAND2_X2 U5073 ( .A1(n10281), .A2(n4686), .ZN(n10263) );
  NAND2_X2 U5074 ( .A1(n10282), .A2(n10287), .ZN(n10281) );
  OR2_X2 U5075 ( .A1(n10069), .A2(n10068), .ZN(n10085) );
  NAND2_X2 U5076 ( .A1(n6678), .A2(n5896), .ZN(n7034) );
  NAND2_X2 U5077 ( .A1(n6680), .A2(n6679), .ZN(n6678) );
  OAI21_X2 U5078 ( .B1(n8930), .B2(n6616), .A(n8233), .ZN(n8921) );
  AOI21_X2 U5079 ( .B1(n4919), .B2(n4571), .A(n4918), .ZN(n10244) );
  BUF_X2 U5080 ( .A(n5420), .Z(n5454) );
  OR2_X1 U5081 ( .A1(n5454), .A2(n6724), .ZN(n5441) );
  AOI21_X2 U5082 ( .B1(n5225), .B2(n5452), .A(n5488), .ZN(n4868) );
  XNOR2_X2 U5083 ( .A(n5226), .B(SI_6_), .ZN(n5488) );
  OAI21_X2 U5084 ( .B1(n5735), .B2(n8423), .A(n4632), .ZN(n10323) );
  NAND2_X2 U5085 ( .A1(n10174), .A2(n9840), .ZN(n10162) );
  AND3_X4 U5086 ( .A1(n4898), .A2(n5402), .A3(n4897), .ZN(n5408) );
  NAND2_X2 U5087 ( .A1(n9635), .A2(n9633), .ZN(n9630) );
  OAI21_X2 U5088 ( .B1(n5667), .B2(n5666), .A(n5294), .ZN(n5679) );
  NAND2_X2 U5089 ( .A1(n4973), .A2(n5289), .ZN(n5667) );
  NAND2_X2 U5090 ( .A1(n8948), .A2(n8955), .ZN(n8947) );
  NOR2_X2 U5091 ( .A1(n8961), .A2(n5011), .ZN(n8948) );
  NAND2_X2 U5092 ( .A1(n5543), .A2(n5542), .ZN(n10486) );
  XNOR2_X2 U5093 ( .A(n5707), .B(n5706), .ZN(n8048) );
  AND2_X2 U5094 ( .A1(n6302), .A2(n6301), .ZN(n7697) );
  XNOR2_X2 U5095 ( .A(n8743), .B(n8748), .ZN(n8733) );
  AND2_X2 U5096 ( .A1(n4757), .A2(n4756), .ZN(n8743) );
  NOR2_X2 U5097 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5419) );
  BUF_X2 U5098 ( .A(n6192), .Z(n8482) );
  INV_X1 U5099 ( .A(n6563), .ZN(n6299) );
  BUF_X4 U5100 ( .A(n5927), .Z(n6110) );
  AOI22_X2 U5101 ( .A1(n10047), .A2(n10046), .B1(n10045), .B2(n10044), .ZN(
        n10066) );
  NOR2_X2 U5102 ( .A1(n10026), .A2(n10025), .ZN(n10047) );
  INV_X1 U5105 ( .A(n6081), .ZN(n6117) );
  AOI21_X2 U5106 ( .B1(n10237), .B2(n10236), .A(n4851), .ZN(n10218) );
  AOI21_X2 U5107 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8615) );
  OAI21_X2 U5108 ( .B1(n8956), .B2(n6614), .A(n8349), .ZN(n8941) );
  AOI21_X2 U5109 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8054), .A(n8050), .ZN(
        n10033) );
  INV_X1 U5110 ( .A(n4544), .ZN(n4545) );
  INV_X2 U5111 ( .A(n4544), .ZN(n4546) );
  XNOR2_X2 U5112 ( .A(n5192), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5195) );
  NAND2_X2 U5113 ( .A1(n10462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5192) );
  XNOR2_X2 U5114 ( .A(n5057), .B(n5056), .ZN(n4985) );
  OAI21_X2 U5115 ( .B1(n10364), .B2(n9967), .A(n5649), .ZN(n10201) );
  AOI21_X2 U5116 ( .B1(n5737), .B2(n5318), .A(n5317), .ZN(n5757) );
  OAI21_X2 U5117 ( .B1(n5350), .B2(n5280), .A(n5279), .ZN(n5634) );
  INV_X2 U5118 ( .A(n4943), .ZN(n5350) );
  NAND2_X2 U5119 ( .A1(n5694), .A2(n5693), .ZN(n10341) );
  XNOR2_X1 U5120 ( .A(n6263), .B(n6262), .ZN(n6798) );
  AOI21_X1 U5121 ( .B1(n9788), .B2(n9838), .A(n9787), .ZN(n9796) );
  OR2_X1 U5122 ( .A1(n9860), .A2(n9859), .ZN(n9923) );
  NOR2_X1 U5123 ( .A1(n7883), .A2(n7884), .ZN(n7959) );
  AND2_X1 U5124 ( .A1(n5050), .A2(n5049), .ZN(n7227) );
  INV_X1 U5126 ( .A(n9698), .ZN(n10557) );
  NAND2_X1 U5127 ( .A1(n9704), .A2(n9808), .ZN(n7188) );
  NAND2_X1 U5128 ( .A1(n8263), .A2(n8259), .ZN(n7075) );
  AND2_X1 U5129 ( .A1(n5037), .A2(n6875), .ZN(n8691) );
  INV_X2 U5130 ( .A(n8671), .ZN(n7324) );
  BUF_X1 U5131 ( .A(n6288), .Z(n8675) );
  INV_X2 U5132 ( .A(n8673), .ZN(n6304) );
  INV_X2 U5133 ( .A(n7140), .ZN(n7503) );
  CLKBUF_X2 U5134 ( .A(n5427), .Z(n4553) );
  NAND2_X1 U5135 ( .A1(n10467), .A2(n10473), .ZN(n5427) );
  BUF_X2 U5136 ( .A(n6270), .Z(n6588) );
  MUX2_X1 U5137 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10475), .S(n6688), .Z(n7488)
         );
  NAND2_X2 U5138 ( .A1(n8482), .A2(n6193), .ZN(n6548) );
  INV_X4 U5139 ( .A(n8402), .ZN(n8392) );
  BUF_X2 U5140 ( .A(n5872), .Z(n4558) );
  OAI21_X1 U5141 ( .B1(n5621), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U5142 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6200) );
  NOR2_X1 U5144 ( .A1(n6179), .A2(n6178), .ZN(n5155) );
  CLKBUF_X1 U5145 ( .A(n6260), .Z(n6261) );
  AND2_X1 U5146 ( .A1(n6260), .A2(n6262), .ZN(n4728) );
  INV_X2 U5147 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9518) );
  INV_X1 U5148 ( .A(n8487), .ZN(n4675) );
  AND2_X1 U5149 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  AOI21_X1 U5150 ( .B1(n4674), .B2(n10451), .A(n4673), .ZN(n4672) );
  OR2_X1 U5151 ( .A1(n10129), .A2(n5733), .ZN(n5735) );
  NOR2_X1 U5152 ( .A1(n9921), .A2(n9938), .ZN(n4955) );
  OR2_X1 U5153 ( .A1(n8791), .A2(n8792), .ZN(n8817) );
  OR2_X1 U5154 ( .A1(n5048), .A2(n8792), .ZN(n8771) );
  OAI211_X1 U5155 ( .C1(n9923), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9924)
         );
  NAND2_X1 U5156 ( .A1(n10175), .A2(n10176), .ZN(n10174) );
  AND2_X1 U5157 ( .A1(n9676), .A2(n9675), .ZN(n10398) );
  AND2_X1 U5158 ( .A1(n8489), .A2(n10453), .ZN(n4673) );
  NAND2_X1 U5159 ( .A1(n5764), .A2(n5763), .ZN(n8489) );
  XNOR2_X1 U5160 ( .A(n8183), .B(n8182), .ZN(n9789) );
  NAND2_X1 U5161 ( .A1(n8166), .A2(n5761), .ZN(n10471) );
  CLKBUF_X1 U5162 ( .A(n10218), .Z(n4687) );
  NAND2_X1 U5163 ( .A1(n4811), .A2(n4810), .ZN(n4809) );
  OR2_X1 U5164 ( .A1(n5760), .A2(SI_29_), .ZN(n5761) );
  INV_X1 U5165 ( .A(n6564), .ZN(n8850) );
  NAND2_X1 U5166 ( .A1(n6530), .A2(n6529), .ZN(n9043) );
  XNOR2_X1 U5167 ( .A(n5741), .B(n5740), .ZN(n8103) );
  NAND2_X1 U5168 ( .A1(n7737), .A2(n5976), .ZN(n7736) );
  AOI21_X1 U5169 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7988), .A(n7985), .ZN(
        n8697) );
  XNOR2_X1 U5170 ( .A(n5721), .B(n5720), .ZN(n8097) );
  XNOR2_X1 U5171 ( .A(n7958), .B(n8666), .ZN(n7883) );
  INV_X1 U5172 ( .A(n8656), .ZN(n8929) );
  NAND2_X1 U5173 ( .A1(n5681), .A2(n5680), .ZN(n10179) );
  NAND2_X1 U5174 ( .A1(n6518), .A2(n6517), .ZN(n8533) );
  NAND2_X1 U5175 ( .A1(n7970), .A2(n9821), .ZN(n8441) );
  NAND2_X1 U5176 ( .A1(n5654), .A2(n5653), .ZN(n10428) );
  AND2_X1 U5177 ( .A1(n10202), .A2(n9681), .ZN(n10217) );
  NAND2_X1 U5178 ( .A1(n5339), .A2(n5338), .ZN(n10364) );
  OAI22_X1 U5179 ( .A1(n6434), .A2(n5005), .B1(n8664), .B2(n8030), .ZN(n5004)
         );
  NAND2_X1 U5180 ( .A1(n6476), .A2(n6475), .ZN(n9444) );
  NAND2_X1 U5181 ( .A1(n5608), .A2(n5607), .ZN(n10454) );
  AOI21_X1 U5182 ( .B1(n7356), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7351), .ZN(
        n7354) );
  NOR2_X1 U5183 ( .A1(n6434), .A2(n5008), .ZN(n5006) );
  NAND2_X1 U5184 ( .A1(n5592), .A2(n5591), .ZN(n9534) );
  NAND2_X1 U5185 ( .A1(n6378), .A2(n6377), .ZN(n7669) );
  NAND2_X1 U5186 ( .A1(n5534), .A2(n5535), .ZN(n5243) );
  NAND2_X1 U5187 ( .A1(n5477), .A2(n4805), .ZN(n9690) );
  NAND2_X1 U5188 ( .A1(n5036), .A2(n6330), .ZN(n7385) );
  NAND2_X1 U5189 ( .A1(n6081), .A2(n5927), .ZN(n5936) );
  NAND2_X1 U5190 ( .A1(n4831), .A2(n6685), .ZN(n6081) );
  NAND2_X1 U5191 ( .A1(n4945), .A2(n5274), .ZN(n4944) );
  INV_X2 U5192 ( .A(n10565), .ZN(n4550) );
  INV_X1 U5193 ( .A(n5884), .ZN(n4831) );
  NAND4_X1 U5194 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n9984)
         );
  NAND4_X1 U5195 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n9986)
         );
  OR2_X1 U5196 ( .A1(n8677), .A2(n6986), .ZN(n8261) );
  NAND2_X1 U5197 ( .A1(n4947), .A2(n4949), .ZN(n4945) );
  OAI211_X1 U5198 ( .C1(n6688), .C2(n4554), .A(n5424), .B(n5423), .ZN(n7140)
         );
  OAI211_X1 U5200 ( .C1(n6563), .C2(n6720), .A(n6265), .B(n6264), .ZN(n8268)
         );
  INV_X1 U5201 ( .A(n5458), .ZN(n5726) );
  INV_X1 U5202 ( .A(n5822), .ZN(n10211) );
  NAND2_X1 U5204 ( .A1(n6711), .A2(n6712), .ZN(n6957) );
  INV_X1 U5205 ( .A(n5195), .ZN(n10467) );
  INV_X1 U5206 ( .A(n5793), .ZN(n8035) );
  XNOR2_X1 U5207 ( .A(n5327), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U5208 ( .A(n5814), .B(n5813), .ZN(n9918) );
  INV_X1 U5209 ( .A(n5196), .ZN(n10473) );
  NAND2_X1 U5210 ( .A1(n9520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U5211 ( .B1(n5812), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5814) );
  OR2_X1 U5212 ( .A1(n6628), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n6637) );
  XNOR2_X1 U5213 ( .A(n6200), .B(n6199), .ZN(n6778) );
  NAND2_X1 U5214 ( .A1(n5193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U5215 ( .A(n5438), .B(n5437), .ZN(n6722) );
  NOR2_X1 U5216 ( .A1(n5118), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4833) );
  XNOR2_X1 U5217 ( .A(n5435), .B(n5434), .ZN(n6721) );
  NAND2_X1 U5218 ( .A1(n4892), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4893) );
  AND4_X1 U5219 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n5183)
         );
  INV_X1 U5220 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6185) );
  INV_X4 U5221 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5222 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5813) );
  INV_X1 U5223 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5486) );
  INV_X1 U5224 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6230) );
  INV_X1 U5225 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6229) );
  INV_X4 U5226 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5227 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6316) );
  NOR2_X1 U5228 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6177) );
  NOR2_X1 U5229 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6173) );
  INV_X1 U5230 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5636) );
  INV_X1 U5231 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8154) );
  INV_X2 U5232 ( .A(n4560), .ZN(n7450) );
  NAND2_X2 U5233 ( .A1(n9631), .A2(n5112), .ZN(n5108) );
  NAND2_X2 U5234 ( .A1(n6086), .A2(n6085), .ZN(n9631) );
  NOR2_X2 U5235 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  INV_X1 U5236 ( .A(n4850), .ZN(n10189) );
  AOI21_X2 U5237 ( .B1(n8397), .B2(n8396), .A(n8395), .ZN(n8403) );
  AOI21_X1 U5238 ( .B1(n5336), .B2(n5286), .A(n4971), .ZN(n4969) );
  AOI22_X2 U5239 ( .A1(n8869), .A2(n6621), .B1(n9474), .B2(n8651), .ZN(n8224)
         );
  INV_X1 U5240 ( .A(n5957), .ZN(n4551) );
  AND2_X4 U5241 ( .A1(n5889), .A2(n5888), .ZN(n5957) );
  INV_X2 U5242 ( .A(n5408), .ZN(n5897) );
  OAI21_X2 U5243 ( .B1(n10147), .B2(n5862), .A(n9848), .ZN(n10131) );
  OAI21_X2 U5244 ( .B1(n10162), .B2(n10160), .A(n5860), .ZN(n10147) );
  INV_X1 U5245 ( .A(n6255), .ZN(n4555) );
  INV_X1 U5246 ( .A(n4555), .ZN(n4556) );
  INV_X1 U5247 ( .A(n4555), .ZN(n4557) );
  NOR2_X2 U5248 ( .A1(n5527), .A2(n7121), .ZN(n5544) );
  OR2_X2 U5249 ( .A1(n5508), .A2(n5507), .ZN(n5527) );
  OAI21_X2 U5250 ( .B1(n5847), .B2(n4855), .A(n4852), .ZN(n10282) );
  AOI211_X2 U5251 ( .C1(n10104), .C2(n10108), .A(n9927), .B(n9926), .ZN(n9928)
         );
  CLKBUF_X2 U5253 ( .A(n9551), .Z(n4561) );
  XNOR2_X2 U5254 ( .A(n5408), .B(n4688), .ZN(n9812) );
  INV_X2 U5255 ( .A(n9987), .ZN(n4688) );
  NAND2_X1 U5256 ( .A1(n8505), .A2(n8951), .ZN(n5135) );
  NOR2_X1 U5257 ( .A1(n5701), .A2(n4935), .ZN(n4934) );
  INV_X1 U5258 ( .A(n4937), .ZN(n4935) );
  NAND2_X1 U5259 ( .A1(n5453), .A2(n5219), .ZN(n5474) );
  INV_X1 U5260 ( .A(n6548), .ZN(n6557) );
  INV_X1 U5261 ( .A(n5130), .ZN(n5128) );
  NAND2_X1 U5262 ( .A1(n4706), .A2(n4606), .ZN(n4704) );
  INV_X1 U5263 ( .A(n5158), .ZN(n4706) );
  AOI21_X1 U5264 ( .B1(n9842), .B2(n9769), .A(n4771), .ZN(n9768) );
  INV_X1 U5265 ( .A(n8279), .ZN(n5060) );
  INV_X1 U5266 ( .A(n8294), .ZN(n5061) );
  INV_X1 U5267 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6327) );
  INV_X1 U5268 ( .A(SI_17_), .ZN(n5270) );
  NOR2_X1 U5269 ( .A1(n5252), .A2(n4962), .ZN(n4961) );
  INV_X1 U5270 ( .A(n5249), .ZN(n4962) );
  AOI21_X1 U5271 ( .B1(n5142), .B2(n5140), .A(n5139), .ZN(n5138) );
  INV_X1 U5272 ( .A(n8623), .ZN(n5139) );
  INV_X1 U5273 ( .A(n5145), .ZN(n5140) );
  MUX2_X1 U5274 ( .A(n8394), .B(n8393), .S(n8392), .Z(n8395) );
  OR2_X1 U5275 ( .A1(n6192), .A2(n6191), .ZN(n6268) );
  NAND2_X1 U5276 ( .A1(n10644), .A2(n6799), .ZN(n6801) );
  NAND2_X1 U5277 ( .A1(n6873), .A2(n6872), .ZN(n6874) );
  NAND2_X1 U5278 ( .A1(n7150), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5051) );
  OAI211_X1 U5279 ( .C1(n4743), .C2(n4741), .A(n4740), .B(n4746), .ZN(n7143)
         );
  INV_X1 U5280 ( .A(n6884), .ZN(n4743) );
  NOR2_X1 U5281 ( .A1(n7471), .A2(n4747), .ZN(n7605) );
  NOR2_X1 U5282 ( .A1(n7228), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U5283 ( .A1(n7677), .A2(n7676), .ZN(n4664) );
  NAND2_X1 U5284 ( .A1(n8732), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4756) );
  INV_X1 U5285 ( .A(n4998), .ZN(n4996) );
  NAND2_X1 U5286 ( .A1(n9501), .A2(n8952), .ZN(n5001) );
  OR2_X1 U5287 ( .A1(n8492), .A2(n8994), .ZN(n8337) );
  INV_X1 U5288 ( .A(n8262), .ZN(n8229) );
  AOI21_X1 U5289 ( .B1(n9620), .B2(n4828), .A(n4607), .ZN(n4827) );
  INV_X1 U5290 ( .A(n6010), .ZN(n4828) );
  INV_X1 U5291 ( .A(n9620), .ZN(n4829) );
  AND2_X1 U5292 ( .A1(n5891), .A2(n6685), .ZN(n4830) );
  INV_X1 U5293 ( .A(n9962), .ZN(n5861) );
  AOI21_X1 U5294 ( .B1(n4913), .B2(n4914), .A(n4621), .ZN(n4912) );
  NOR2_X1 U5295 ( .A1(n5585), .A2(n4916), .ZN(n4913) );
  NAND2_X1 U5296 ( .A1(n5822), .A2(n4549), .ZN(n6122) );
  NAND2_X1 U5297 ( .A1(n5795), .A2(n5785), .ZN(n5889) );
  NOR2_X1 U5298 ( .A1(n5792), .A2(n8035), .ZN(n5785) );
  AND3_X1 U5299 ( .A1(n5636), .A2(n5353), .A3(n5184), .ZN(n5160) );
  INV_X1 U5300 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U5301 ( .A1(n5261), .A2(n5260), .ZN(n5602) );
  AND2_X1 U5302 ( .A1(n5587), .A2(n5258), .ZN(n5259) );
  INV_X1 U5303 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5304 ( .B1(n4586), .B2(n4564), .A(n5518), .ZN(n4967) );
  INV_X1 U5305 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U5306 ( .A1(n4988), .A2(n5218), .ZN(n5453) );
  NAND2_X1 U5307 ( .A1(n8411), .A2(n8229), .ZN(n8402) );
  AOI21_X1 U5308 ( .B1(n5127), .B2(n5132), .A(n5133), .ZN(n5125) );
  NOR2_X1 U5309 ( .A1(n8507), .A2(n8659), .ZN(n5133) );
  NAND2_X1 U5310 ( .A1(n8636), .A2(n5148), .ZN(n8583) );
  AND2_X1 U5311 ( .A1(n8570), .A2(n8571), .ZN(n5148) );
  AOI21_X1 U5312 ( .B1(n8083), .B2(n8082), .A(n4641), .ZN(n8088) );
  NAND2_X1 U5313 ( .A1(n6190), .A2(n6191), .ZN(n6270) );
  INV_X1 U5314 ( .A(n6403), .ZN(n6565) );
  INV_X1 U5315 ( .A(n6267), .ZN(n6255) );
  AND2_X1 U5316 ( .A1(n6191), .A2(n8482), .ZN(n6267) );
  INV_X1 U5317 ( .A(n6191), .ZN(n6193) );
  CLKBUF_X2 U5318 ( .A(n6268), .Z(n6403) );
  AND2_X1 U5319 ( .A1(n7674), .A2(n7673), .ZN(n7808) );
  AND2_X1 U5320 ( .A1(n4733), .A2(n4732), .ZN(n8712) );
  NAND2_X1 U5321 ( .A1(n7988), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U5322 ( .A1(n4731), .A2(n4583), .ZN(n4730) );
  INV_X1 U5323 ( .A(n4660), .ZN(n8747) );
  NAND2_X1 U5324 ( .A1(n8815), .A2(n10648), .ZN(n8813) );
  AND2_X1 U5325 ( .A1(n4737), .A2(n4736), .ZN(n8827) );
  INV_X1 U5326 ( .A(n8816), .ZN(n4736) );
  AND2_X1 U5327 ( .A1(n8372), .A2(n6617), .ZN(n8900) );
  NAND2_X1 U5328 ( .A1(n6169), .A2(n6168), .ZN(n6533) );
  NAND2_X1 U5329 ( .A1(n4657), .A2(n4995), .ZN(n4992) );
  INV_X1 U5330 ( .A(n8947), .ZN(n4657) );
  NAND2_X1 U5331 ( .A1(n5082), .A2(n8997), .ZN(n8996) );
  NAND2_X1 U5332 ( .A1(n6918), .A2(n8392), .ZN(n8993) );
  OR2_X1 U5333 ( .A1(n6918), .A2(n8402), .ZN(n8953) );
  NAND2_X1 U5334 ( .A1(n7653), .A2(n7731), .ZN(n9449) );
  INV_X1 U5335 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6574) );
  AOI21_X1 U5336 ( .B1(n6435), .B2(P2_IR_REG_31__SCAN_IN), .A(n4702), .ZN(
        n4701) );
  NAND2_X1 U5337 ( .A1(n4703), .A2(n6236), .ZN(n4702) );
  INV_X1 U5338 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U5339 ( .A1(n5351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5362) );
  AOI21_X1 U5340 ( .B1(n4934), .B2(n4932), .A(n4612), .ZN(n4931) );
  INV_X1 U5341 ( .A(n4939), .ZN(n4932) );
  AOI21_X1 U5342 ( .B1(n4582), .B2(n4939), .A(n4938), .ZN(n4937) );
  NOR2_X1 U5343 ( .A1(n10346), .A2(n5858), .ZN(n4938) );
  INV_X1 U5344 ( .A(n4920), .ZN(n4918) );
  AND2_X1 U5345 ( .A1(n6121), .A2(n4549), .ZN(n10319) );
  NAND2_X1 U5346 ( .A1(n4834), .A2(n5183), .ZN(n5351) );
  INV_X1 U5347 ( .A(n8655), .ZN(n8919) );
  INV_X1 U5348 ( .A(n8653), .ZN(n8897) );
  INV_X1 U5349 ( .A(n8654), .ZN(n8908) );
  INV_X1 U5350 ( .A(n9903), .ZN(n4803) );
  AOI21_X1 U5351 ( .B1(n4776), .B2(n4779), .A(n4620), .ZN(n4775) );
  NAND2_X1 U5352 ( .A1(n8309), .A2(n4888), .ZN(n4887) );
  AND2_X1 U5353 ( .A1(n8308), .A2(n8392), .ZN(n4888) );
  AOI21_X1 U5354 ( .B1(n9776), .B2(n9774), .A(n9859), .ZN(n4793) );
  OAI21_X1 U5355 ( .B1(n4872), .B2(n4871), .A(n8361), .ZN(n8368) );
  NAND2_X1 U5356 ( .A1(n9848), .A2(n9844), .ZN(n4795) );
  NAND2_X1 U5357 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  INV_X1 U5358 ( .A(n4791), .ZN(n4788) );
  INV_X1 U5359 ( .A(n4789), .ZN(n4787) );
  MUX2_X1 U5360 ( .A(n9773), .B(n9772), .S(n9795), .Z(n4974) );
  AOI21_X1 U5361 ( .B1(n9769), .B2(n4770), .A(n4769), .ZN(n9771) );
  AOI21_X1 U5362 ( .B1(n4793), .B2(n9845), .A(n9795), .ZN(n4789) );
  INV_X1 U5363 ( .A(n4793), .ZN(n4790) );
  NOR2_X1 U5364 ( .A1(n8383), .A2(n8382), .ZN(n4883) );
  INV_X1 U5365 ( .A(n5650), .ZN(n5288) );
  INV_X1 U5366 ( .A(n5147), .ZN(n5144) );
  NAND2_X1 U5367 ( .A1(n6566), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U5368 ( .A1(n6619), .A2(n5034), .ZN(n5031) );
  NAND2_X1 U5369 ( .A1(n6619), .A2(n5030), .ZN(n5029) );
  NAND2_X1 U5370 ( .A1(n4587), .A2(n6618), .ZN(n5030) );
  NAND2_X1 U5371 ( .A1(n8900), .A2(n5032), .ZN(n5025) );
  NOR2_X1 U5372 ( .A1(n5031), .A2(n5035), .ZN(n5027) );
  NOR2_X1 U5373 ( .A1(n8374), .A2(n5077), .ZN(n5076) );
  INV_X1 U5374 ( .A(n8367), .ZN(n5077) );
  OR2_X1 U5375 ( .A1(n8560), .A2(n8952), .ZN(n8358) );
  OR2_X1 U5376 ( .A1(n9062), .A2(n8964), .ZN(n8357) );
  INV_X1 U5377 ( .A(n5020), .ZN(n5017) );
  OR2_X1 U5378 ( .A1(n9444), .A2(n8992), .ZN(n8332) );
  AOI21_X1 U5379 ( .B1(n8294), .B2(n5065), .A(n5063), .ZN(n5062) );
  INV_X1 U5380 ( .A(n8281), .ZN(n5065) );
  OR2_X1 U5381 ( .A1(n8674), .A2(n8268), .ZN(n6290) );
  AND2_X1 U5382 ( .A1(n6622), .A2(n6623), .ZN(n6625) );
  INV_X1 U5383 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9220) );
  INV_X1 U5384 ( .A(n8340), .ZN(n5081) );
  NAND2_X1 U5385 ( .A1(n6622), .A2(n8406), .ZN(n6922) );
  NOR2_X1 U5386 ( .A1(n4825), .A2(n9529), .ZN(n5095) );
  NOR2_X1 U5387 ( .A1(n6024), .A2(n5094), .ZN(n5091) );
  INV_X1 U5388 ( .A(n9529), .ZN(n5094) );
  OR2_X1 U5389 ( .A1(n8479), .A2(n5754), .ZN(n9854) );
  NOR2_X1 U5390 ( .A1(n10326), .A2(n8479), .ZN(n4849) );
  NOR2_X1 U5391 ( .A1(n10443), .A2(n10374), .ZN(n4846) );
  NOR2_X1 U5392 ( .A1(n9743), .A2(n4857), .ZN(n4856) );
  NOR2_X1 U5393 ( .A1(n10625), .A2(n4839), .ZN(n4838) );
  INV_X1 U5394 ( .A(n4840), .ZN(n4839) );
  NAND2_X1 U5395 ( .A1(n7845), .A2(n7852), .ZN(n7844) );
  INV_X1 U5396 ( .A(n9961), .ZN(n5863) );
  AOI21_X1 U5397 ( .B1(n4565), .B2(n4921), .A(n4605), .ZN(n4920) );
  NOR2_X1 U5398 ( .A1(n4923), .A2(n4925), .ZN(n4921) );
  AND2_X1 U5399 ( .A1(n7933), .A2(n9807), .ZN(n6121) );
  NAND2_X1 U5400 ( .A1(n5759), .A2(n5758), .ZN(n8162) );
  NAND2_X1 U5401 ( .A1(n5721), .A2(n5720), .ZN(n5737) );
  INV_X1 U5402 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U5403 ( .A1(n5786), .A2(n5185), .ZN(n5783) );
  AND2_X1 U5404 ( .A1(n5702), .A2(n5304), .ZN(n5691) );
  NOR2_X1 U5405 ( .A1(n5360), .A2(n4952), .ZN(n4951) );
  INV_X1 U5406 ( .A(n5264), .ZN(n4952) );
  AND2_X1 U5407 ( .A1(n5274), .A2(n5273), .ZN(n5619) );
  NAND2_X1 U5408 ( .A1(n4950), .A2(n5269), .ZN(n4949) );
  NAND2_X1 U5409 ( .A1(n4951), .A2(n5265), .ZN(n4950) );
  AOI21_X1 U5410 ( .B1(n4958), .B2(n4960), .A(n5376), .ZN(n4956) );
  NOR2_X1 U5411 ( .A1(n5553), .A2(n4965), .ZN(n4964) );
  INV_X1 U5412 ( .A(n5242), .ZN(n4965) );
  AOI21_X1 U5413 ( .B1(n5138), .B2(n5141), .A(n4574), .ZN(n5136) );
  INV_X1 U5414 ( .A(n5142), .ZN(n5141) );
  OR2_X1 U5415 ( .A1(n8109), .A2(n8108), .ZN(n4708) );
  NAND2_X1 U5416 ( .A1(n8504), .A2(n8994), .ZN(n5134) );
  INV_X1 U5417 ( .A(n5138), .ZN(n4712) );
  AND2_X1 U5418 ( .A1(n5136), .A2(n4715), .ZN(n4714) );
  INV_X1 U5419 ( .A(n8520), .ZN(n4715) );
  NAND2_X1 U5420 ( .A1(n6922), .A2(n4722), .ZN(n7162) );
  INV_X1 U5421 ( .A(n4723), .ZN(n4722) );
  OAI21_X1 U5422 ( .B1(n6924), .B2(n6923), .A(n7364), .ZN(n4723) );
  AND2_X1 U5423 ( .A1(n8513), .A2(n8919), .ZN(n5147) );
  NAND2_X1 U5424 ( .A1(n8605), .A2(n8510), .ZN(n8511) );
  OR2_X1 U5425 ( .A1(n8509), .A2(n8939), .ZN(n8510) );
  NAND2_X1 U5426 ( .A1(n5135), .A2(n4589), .ZN(n5130) );
  INV_X1 U5427 ( .A(n8556), .ZN(n5123) );
  INV_X1 U5428 ( .A(n8613), .ZN(n4719) );
  NAND2_X1 U5429 ( .A1(n5127), .A2(n8556), .ZN(n5124) );
  NAND2_X1 U5430 ( .A1(n4720), .A2(n8613), .ZN(n8612) );
  NAND2_X1 U5431 ( .A1(n4721), .A2(n8503), .ZN(n4720) );
  AND2_X1 U5432 ( .A1(n8172), .A2(n6586), .ZN(n6918) );
  INV_X1 U5433 ( .A(n8087), .ZN(n4709) );
  INV_X1 U5434 ( .A(n8405), .ZN(n4878) );
  MUX2_X1 U5435 ( .A(n8231), .B(n8230), .S(n8229), .Z(n8407) );
  AND4_X1 U5436 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n8247)
         );
  OR2_X1 U5437 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  OR2_X1 U5438 ( .A1(n6268), .A2(n7376), .ZN(n6272) );
  NAND2_X1 U5439 ( .A1(n4738), .A2(n6827), .ZN(n4739) );
  NAND2_X1 U5440 ( .A1(n6801), .A2(n6800), .ZN(n6804) );
  NAND3_X1 U5441 ( .A1(n4739), .A2(P2_REG1_REG_3__SCAN_IN), .A3(n6804), .ZN(
        n6824) );
  NAND2_X1 U5442 ( .A1(n5038), .A2(n6869), .ZN(n5037) );
  INV_X1 U5443 ( .A(n6874), .ZN(n5038) );
  NAND2_X1 U5444 ( .A1(n4751), .A2(n4750), .ZN(n7231) );
  NOR2_X1 U5445 ( .A1(n7227), .A2(n4753), .ZN(n4751) );
  INV_X1 U5446 ( .A(n4754), .ZN(n4750) );
  NAND2_X1 U5447 ( .A1(n4734), .A2(n4600), .ZN(n4976) );
  INV_X1 U5448 ( .A(n4664), .ZN(n7824) );
  OR2_X1 U5449 ( .A1(n7831), .A2(n7830), .ZN(n4733) );
  NAND2_X1 U5450 ( .A1(n4984), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4981) );
  INV_X1 U5451 ( .A(n8717), .ZN(n4984) );
  INV_X1 U5452 ( .A(n8750), .ZN(n4729) );
  INV_X1 U5453 ( .A(n5072), .ZN(n5071) );
  OAI22_X1 U5454 ( .A1(n4563), .A2(n5073), .B1(n8518), .B2(n8887), .ZN(n5072)
         );
  OAI21_X1 U5455 ( .B1(n8895), .B2(n8900), .A(n5032), .ZN(n8885) );
  NOR2_X1 U5456 ( .A1(n8887), .A2(n8953), .ZN(n4685) );
  AOI21_X1 U5457 ( .B1(n6617), .B2(n8366), .A(n8373), .ZN(n5075) );
  AOI21_X1 U5458 ( .B1(n4995), .B2(n4994), .A(n4613), .ZN(n4993) );
  INV_X1 U5459 ( .A(n4999), .ZN(n4994) );
  AND2_X1 U5460 ( .A1(n8362), .A2(n8911), .ZN(n8920) );
  AND2_X1 U5461 ( .A1(n5001), .A2(n5002), .ZN(n4999) );
  NAND2_X1 U5462 ( .A1(n8940), .A2(n5001), .ZN(n4998) );
  AND2_X1 U5463 ( .A1(n8234), .A2(n8233), .ZN(n8931) );
  INV_X1 U5464 ( .A(n8657), .ZN(n8939) );
  INV_X1 U5465 ( .A(n8658), .ZN(n8952) );
  AND2_X1 U5466 ( .A1(n8967), .A2(n8977), .ZN(n5011) );
  NOR2_X1 U5467 ( .A1(n8326), .A2(n5021), .ZN(n5020) );
  INV_X1 U5468 ( .A(n6459), .ZN(n5021) );
  NOR2_X1 U5469 ( .A1(n6612), .A2(n5088), .ZN(n5087) );
  INV_X1 U5470 ( .A(n6610), .ZN(n5088) );
  AND2_X1 U5471 ( .A1(n8329), .A2(n8328), .ZN(n8326) );
  NAND2_X1 U5472 ( .A1(n6155), .A2(n7821), .ZN(n6438) );
  INV_X1 U5473 ( .A(n6427), .ZN(n6155) );
  NOR2_X1 U5474 ( .A1(n7726), .A2(n8665), .ZN(n5009) );
  AND2_X1 U5475 ( .A1(n6608), .A2(n6607), .ZN(n8314) );
  CLKBUF_X1 U5476 ( .A(n7720), .Z(n4658) );
  OR2_X1 U5477 ( .A1(n7479), .A2(n8198), .ZN(n6604) );
  OR2_X1 U5478 ( .A1(n7324), .A2(n7385), .ZN(n8281) );
  NAND2_X1 U5479 ( .A1(n6602), .A2(n8279), .ZN(n7264) );
  AND2_X1 U5480 ( .A1(n6651), .A2(n6650), .ZN(n7338) );
  AND2_X1 U5481 ( .A1(n8996), .A2(n5080), .ZN(n9073) );
  NAND2_X1 U5482 ( .A1(n8996), .A2(n8340), .ZN(n8981) );
  NAND2_X1 U5483 ( .A1(n6451), .A2(n6450), .ZN(n8107) );
  OR2_X1 U5484 ( .A1(n6922), .A2(n8402), .ZN(n7345) );
  AND2_X1 U5485 ( .A1(n6916), .A2(n6915), .ZN(n7050) );
  NAND2_X1 U5486 ( .A1(n6664), .A2(n6663), .ZN(n6903) );
  INV_X1 U5487 ( .A(n6915), .ZN(n6912) );
  INV_X1 U5488 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6199) );
  AND2_X1 U5489 ( .A1(n6639), .A2(n6201), .ZN(n6642) );
  INV_X1 U5490 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6635) );
  OAI21_X1 U5491 ( .B1(n6628), .B2(n5153), .A(n5151), .ZN(n6629) );
  AOI21_X1 U5492 ( .B1(n5152), .B2(n9518), .A(n9518), .ZN(n5151) );
  INV_X1 U5493 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6634) );
  INV_X1 U5494 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6573) );
  AND3_X1 U5495 ( .A1(n4728), .A2(n4727), .A3(n4726), .ZN(n6374) );
  XNOR2_X1 U5496 ( .A(n6341), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7148) );
  INV_X1 U5497 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5056) );
  NOR2_X1 U5498 ( .A1(n9518), .A2(n6794), .ZN(n5057) );
  NOR2_X1 U5499 ( .A1(n4820), .A2(n4813), .ZN(n4812) );
  INV_X1 U5500 ( .A(n4821), .ZN(n4820) );
  INV_X1 U5501 ( .A(n5109), .ZN(n4813) );
  NAND2_X1 U5502 ( .A1(n4826), .A2(n4824), .ZN(n9526) );
  AOI21_X1 U5503 ( .B1(n4827), .B2(n4829), .A(n4825), .ZN(n4824) );
  NAND2_X1 U5504 ( .A1(n5106), .A2(n9630), .ZN(n5111) );
  INV_X1 U5505 ( .A(n5108), .ZN(n5106) );
  NAND2_X1 U5506 ( .A1(n4831), .A2(n4830), .ZN(n5892) );
  NAND2_X1 U5507 ( .A1(n5098), .A2(n6060), .ZN(n5097) );
  NAND2_X1 U5508 ( .A1(n5101), .A2(n5103), .ZN(n5098) );
  AND2_X1 U5509 ( .A1(n9654), .A2(n4823), .ZN(n4821) );
  INV_X1 U5510 ( .A(n6131), .ZN(n6132) );
  AND2_X1 U5511 ( .A1(n10398), .A2(n9929), .ZN(n9933) );
  INV_X1 U5512 ( .A(n7933), .ZN(n9802) );
  INV_X1 U5513 ( .A(n5766), .ZN(n5714) );
  INV_X1 U5514 ( .A(n5695), .ZN(n5729) );
  NAND2_X1 U5515 ( .A1(n5195), .A2(n5196), .ZN(n5425) );
  NAND2_X1 U5516 ( .A1(n10005), .A2(n4689), .ZN(n6711) );
  NAND2_X1 U5517 ( .A1(n4690), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5518 ( .A1(n10035), .A2(n10034), .ZN(n10038) );
  OR2_X1 U5519 ( .A1(n10038), .A2(n10039), .ZN(n10051) );
  NAND2_X1 U5520 ( .A1(n5171), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U5521 ( .A1(n10306), .A2(n5157), .ZN(n5617) );
  NAND2_X1 U5522 ( .A1(n5847), .A2(n4856), .ZN(n10299) );
  NOR2_X1 U5523 ( .A1(n5161), .A2(n4602), .ZN(n4914) );
  NAND2_X1 U5524 ( .A1(n7975), .A2(n5585), .ZN(n4915) );
  INV_X1 U5525 ( .A(n9821), .ZN(n7974) );
  NAND2_X1 U5526 ( .A1(n7922), .A2(n5566), .ZN(n7975) );
  OR2_X1 U5527 ( .A1(n10625), .A2(n9976), .ZN(n5566) );
  NAND2_X1 U5528 ( .A1(n7924), .A2(n7923), .ZN(n7922) );
  NAND2_X1 U5529 ( .A1(n7755), .A2(n5533), .ZN(n7799) );
  OR2_X1 U5530 ( .A1(n4559), .A2(n9978), .ZN(n5533) );
  NAND2_X1 U5531 ( .A1(n4899), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4898) );
  INV_X1 U5532 ( .A(n10319), .ZN(n10308) );
  AOI21_X1 U5533 ( .B1(n4929), .B2(n4931), .A(n4928), .ZN(n4927) );
  NOR2_X1 U5534 ( .A1(n10152), .A2(n5861), .ZN(n4928) );
  INV_X1 U5535 ( .A(n4934), .ZN(n4933) );
  NOR2_X1 U5536 ( .A1(n5690), .A2(n4940), .ZN(n4939) );
  INV_X1 U5537 ( .A(n4941), .ZN(n4940) );
  AND2_X1 U5538 ( .A1(n9770), .A2(n9840), .ZN(n10176) );
  NAND2_X1 U5539 ( .A1(n4942), .A2(n6082), .ZN(n4941) );
  OR2_X1 U5540 ( .A1(n10256), .A2(n5853), .ZN(n5162) );
  NAND2_X1 U5541 ( .A1(n5364), .A2(n5363), .ZN(n10384) );
  INV_X1 U5542 ( .A(n6688), .ZN(n5638) );
  NAND2_X1 U5543 ( .A1(n5865), .A2(n9801), .ZN(n10285) );
  AND2_X1 U5544 ( .A1(n5796), .A2(n5795), .ZN(n6747) );
  NAND2_X1 U5545 ( .A1(n5777), .A2(n5778), .ZN(n5781) );
  XNOR2_X1 U5546 ( .A(n5791), .B(n5790), .ZN(n7937) );
  NAND2_X1 U5547 ( .A1(n5809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5791) );
  AND2_X1 U5548 ( .A1(n5787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U5549 ( .A1(n5789), .A2(n5788), .ZN(n5809) );
  INV_X1 U5550 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5788) );
  INV_X1 U5551 ( .A(n5807), .ZN(n5789) );
  NAND2_X1 U5552 ( .A1(n5160), .A2(n4601), .ZN(n5118) );
  NAND2_X1 U5553 ( .A1(n5287), .A2(n4970), .ZN(n5652) );
  NAND2_X1 U5554 ( .A1(n5160), .A2(n5117), .ZN(n5812) );
  INV_X1 U5555 ( .A(n5351), .ZN(n5117) );
  OAI21_X1 U5556 ( .B1(n5243), .B2(n4960), .A(n4958), .ZN(n5377) );
  XNOR2_X1 U5557 ( .A(n5476), .B(n5475), .ZN(n6324) );
  XNOR2_X1 U5558 ( .A(n8511), .B(n8512), .ZN(n8529) );
  AND2_X1 U5559 ( .A1(n6498), .A2(n6497), .ZN(n8975) );
  AND2_X1 U5560 ( .A1(n7318), .A2(n7317), .ZN(n7320) );
  NAND2_X1 U5561 ( .A1(n6205), .A2(n6204), .ZN(n8630) );
  NAND2_X1 U5562 ( .A1(n6538), .A2(n6537), .ZN(n8654) );
  INV_X1 U5563 ( .A(n7617), .ZN(n5044) );
  NOR2_X1 U5564 ( .A1(n6415), .A2(n7675), .ZN(n7809) );
  OR2_X1 U5565 ( .A1(n7984), .A2(n8010), .ZN(n4983) );
  OR2_X1 U5566 ( .A1(n8724), .A2(n9400), .ZN(n4731) );
  INV_X1 U5567 ( .A(n5042), .ZN(n8744) );
  INV_X1 U5568 ( .A(n8813), .ZN(n8808) );
  OAI21_X1 U5569 ( .B1(n8867), .B2(n8990), .A(n8866), .ZN(n9034) );
  NOR2_X1 U5570 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NOR2_X1 U5571 ( .A1(n8863), .A2(n8953), .ZN(n8865) );
  NAND2_X1 U5572 ( .A1(n4696), .A2(n4693), .ZN(n9037) );
  NOR2_X1 U5573 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  NOR2_X1 U5574 ( .A1(n8897), .A2(n8993), .ZN(n4694) );
  OAI21_X1 U5575 ( .B1(n8896), .B2(n8990), .A(n4666), .ZN(n9044) );
  NOR2_X1 U5576 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  NOR2_X1 U5577 ( .A1(n8919), .A2(n8993), .ZN(n4667) );
  AOI21_X1 U5578 ( .B1(n8912), .B2(n8367), .A(n8366), .ZN(n8901) );
  AND2_X1 U5579 ( .A1(n8859), .A2(n9449), .ZN(n6624) );
  OAI21_X1 U5580 ( .B1(n6435), .B2(n4704), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6241) );
  INV_X1 U5581 ( .A(n5116), .ZN(n5115) );
  INV_X1 U5582 ( .A(n10547), .ZN(n9638) );
  AOI21_X1 U5583 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6974), .A(n6969), .ZN(
        n6972) );
  AOI21_X1 U5584 ( .B1(n7356), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7355), .ZN(
        n7359) );
  INV_X1 U5585 ( .A(n10406), .ZN(n10142) );
  NAND2_X1 U5586 ( .A1(n8489), .A2(n10392), .ZN(n4860) );
  AND2_X1 U5587 ( .A1(n8099), .A2(n5792), .ZN(n6749) );
  AOI21_X1 U5588 ( .B1(n9734), .B2(n9733), .A(n5843), .ZN(n4780) );
  NAND2_X1 U5589 ( .A1(n4588), .A2(n4879), .ZN(n8257) );
  AOI21_X1 U5590 ( .B1(n4881), .B2(n8402), .A(n4880), .ZN(n4879) );
  AND2_X1 U5591 ( .A1(n8243), .A2(n8392), .ZN(n4880) );
  NAND2_X1 U5592 ( .A1(n8250), .A2(n8251), .ZN(n4881) );
  INV_X1 U5593 ( .A(n9738), .ZN(n4781) );
  INV_X1 U5594 ( .A(n4780), .ZN(n4779) );
  AND2_X1 U5595 ( .A1(n4783), .A2(n4777), .ZN(n4776) );
  AND2_X1 U5596 ( .A1(n9737), .A2(n9891), .ZN(n4783) );
  NAND2_X1 U5597 ( .A1(n4780), .A2(n4778), .ZN(n4777) );
  INV_X1 U5598 ( .A(n9733), .ZN(n4778) );
  AND2_X1 U5599 ( .A1(n4801), .A2(n4799), .ZN(n9744) );
  AOI21_X1 U5600 ( .B1(n9749), .B2(n10310), .A(n4800), .ZN(n4799) );
  NOR2_X1 U5601 ( .A1(n4804), .A2(n4803), .ZN(n4802) );
  NAND2_X1 U5602 ( .A1(n4886), .A2(n4885), .ZN(n8319) );
  INV_X1 U5603 ( .A(n8313), .ZN(n4885) );
  OAI211_X1 U5604 ( .C1(n8310), .C2(n8392), .A(n8314), .B(n4887), .ZN(n4886)
         );
  INV_X1 U5605 ( .A(n8319), .ZN(n8317) );
  AND2_X1 U5606 ( .A1(n4865), .A2(n8341), .ZN(n4863) );
  AND2_X1 U5607 ( .A1(n8326), .A2(n8325), .ZN(n4865) );
  NAND2_X1 U5608 ( .A1(n4622), .A2(n8341), .ZN(n4862) );
  NAND2_X1 U5609 ( .A1(n8339), .A2(n4609), .ZN(n4864) );
  AOI21_X1 U5610 ( .B1(n8355), .B2(n4873), .A(n4590), .ZN(n4872) );
  AND2_X1 U5611 ( .A1(n8354), .A2(n8356), .ZN(n4873) );
  NAND2_X1 U5612 ( .A1(n8931), .A2(n4597), .ZN(n4871) );
  NAND2_X1 U5613 ( .A1(n9766), .A2(n9767), .ZN(n4773) );
  NOR2_X1 U5614 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  INV_X1 U5615 ( .A(n9852), .ZN(n4772) );
  INV_X1 U5616 ( .A(n9770), .ZN(n4769) );
  AOI22_X1 U5617 ( .A1(n4789), .A2(n4790), .B1(n4791), .B2(n4792), .ZN(n4784)
         );
  INV_X1 U5618 ( .A(n4794), .ZN(n4792) );
  NAND2_X1 U5619 ( .A1(n4882), .A2(n4884), .ZN(n8387) );
  AND2_X1 U5620 ( .A1(n6886), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5621 ( .A1(n6303), .A2(n6304), .ZN(n8286) );
  NAND2_X1 U5622 ( .A1(n4649), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U5623 ( .A1(n5286), .A2(n5333), .ZN(n4972) );
  INV_X1 U5624 ( .A(n4948), .ZN(n4947) );
  OAI21_X1 U5625 ( .B1(n4949), .B2(n4951), .A(n5619), .ZN(n4948) );
  INV_X1 U5626 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5276) );
  INV_X1 U5627 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5275) );
  NOR2_X1 U5628 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5176) );
  NAND2_X1 U5629 ( .A1(n4699), .A2(n4698), .ZN(n5222) );
  NAND2_X1 U5630 ( .A1(n5330), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4698) );
  OR2_X1 U5631 ( .A1(n5330), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U5632 ( .A1(n4677), .A2(n4676), .ZN(n5220) );
  NAND2_X1 U5633 ( .A1(n5330), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4676) );
  OR2_X1 U5634 ( .A1(n5330), .A2(n4678), .ZN(n4677) );
  OAI21_X1 U5635 ( .B1(n5330), .B2(n5215), .A(n5214), .ZN(n5217) );
  NAND2_X1 U5636 ( .A1(n5330), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5214) );
  INV_X1 U5637 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4768) );
  NAND2_X1 U5638 ( .A1(n5203), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4892) );
  INV_X1 U5639 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5203) );
  NAND2_X1 U5640 ( .A1(n5046), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U5641 ( .A1(n8389), .A2(n8221), .ZN(n8385) );
  NAND2_X1 U5642 ( .A1(n8877), .A2(n8379), .ZN(n5073) );
  NOR2_X1 U5643 ( .A1(n5073), .A2(n5068), .ZN(n5067) );
  INV_X1 U5644 ( .A(n5076), .ZN(n5068) );
  NAND2_X1 U5645 ( .A1(n5009), .A2(n5007), .ZN(n5005) );
  NOR2_X1 U5646 ( .A1(n7669), .A2(n7633), .ZN(n8243) );
  NAND2_X1 U5647 ( .A1(n7637), .A2(n7885), .ZN(n8251) );
  OAI21_X1 U5648 ( .B1(n7207), .B2(n6351), .A(n6350), .ZN(n7407) );
  INV_X1 U5649 ( .A(n7075), .ZN(n8190) );
  OR2_X1 U5650 ( .A1(n6647), .A2(n6662), .ZN(n6900) );
  NAND2_X1 U5651 ( .A1(n7073), .A2(n8263), .ZN(n7056) );
  AND2_X1 U5652 ( .A1(n6895), .A2(n6900), .ZN(n6916) );
  INV_X1 U5653 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6202) );
  INV_X1 U5654 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5655 ( .A1(n4704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4703) );
  NOR2_X1 U5656 ( .A1(n6383), .A2(n6232), .ZN(n6423) );
  INV_X1 U5657 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6231) );
  INV_X1 U5658 ( .A(n4724), .ZN(n4727) );
  AND3_X1 U5659 ( .A1(n4728), .A2(n4727), .A3(n4725), .ZN(n6380) );
  AND2_X1 U5660 ( .A1(n6229), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5661 ( .A1(n9644), .A2(n9643), .ZN(n5104) );
  AND2_X1 U5662 ( .A1(n9557), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U5663 ( .A1(n5105), .A2(n5104), .ZN(n5102) );
  NAND2_X1 U5664 ( .A1(n5669), .A2(n4604), .ZN(n9677) );
  OR2_X1 U5665 ( .A1(n5671), .A2(n5670), .ZN(n5683) );
  NAND2_X1 U5666 ( .A1(n9852), .A2(n9677), .ZN(n9832) );
  OR2_X1 U5667 ( .A1(n10625), .A2(n5565), .ZN(n9737) );
  NOR2_X1 U5668 ( .A1(n4559), .A2(n10486), .ZN(n4840) );
  INV_X1 U5669 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7121) );
  AND2_X1 U5670 ( .A1(n5408), .A2(n7185), .ZN(n4836) );
  INV_X1 U5671 ( .A(n5762), .ZN(n4807) );
  OR2_X1 U5672 ( .A1(n8489), .A2(n5774), .ZN(n9866) );
  AND2_X1 U5673 ( .A1(n4931), .A2(n4591), .ZN(n4930) );
  AND2_X1 U5674 ( .A1(n4933), .A2(n4591), .ZN(n4929) );
  NAND2_X1 U5675 ( .A1(n10289), .A2(n10274), .ZN(n10273) );
  NAND2_X1 U5676 ( .A1(n7490), .A2(n9812), .ZN(n5836) );
  NAND2_X1 U5677 ( .A1(n8166), .A2(n8165), .ZN(n8183) );
  INV_X1 U5678 ( .A(n5704), .ZN(n5308) );
  AND2_X1 U5679 ( .A1(n5736), .A2(n5313), .ZN(n5720) );
  AOI21_X1 U5680 ( .B1(n4959), .B2(n4961), .A(n4617), .ZN(n4958) );
  INV_X1 U5681 ( .A(n4964), .ZN(n4959) );
  INV_X1 U5682 ( .A(n4961), .ZN(n4960) );
  INV_X1 U5683 ( .A(n5501), .ZN(n4968) );
  XNOR2_X1 U5684 ( .A(n5208), .B(SI_1_), .ZN(n5397) );
  XNOR2_X1 U5685 ( .A(n7697), .B(n7162), .ZN(n7159) );
  OR2_X1 U5686 ( .A1(n6477), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U5687 ( .A1(n8088), .A2(n8087), .ZN(n8110) );
  NAND2_X1 U5688 ( .A1(n6165), .A2(n6164), .ZN(n6510) );
  INV_X1 U5689 ( .A(n6501), .ZN(n6165) );
  NAND2_X1 U5690 ( .A1(n7882), .A2(n7881), .ZN(n7958) );
  NAND2_X1 U5691 ( .A1(n7097), .A2(n6928), .ZN(n6929) );
  NOR2_X1 U5692 ( .A1(n8564), .A2(n5146), .ZN(n5145) );
  INV_X1 U5693 ( .A(n8590), .ZN(n5146) );
  AND2_X1 U5694 ( .A1(n5143), .A2(n4629), .ZN(n5142) );
  OR2_X1 U5695 ( .A1(n8564), .A2(n5144), .ZN(n5143) );
  NAND2_X1 U5696 ( .A1(n6159), .A2(n6158), .ZN(n6477) );
  INV_X1 U5697 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6158) );
  INV_X1 U5698 ( .A(n6467), .ZN(n6159) );
  AND2_X1 U5699 ( .A1(n8181), .A2(n8180), .ZN(n8849) );
  AOI21_X1 U5700 ( .B1(n8870), .B2(n6565), .A(n6560), .ZN(n8876) );
  NAND4_X1 U5701 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n8674)
         );
  NAND2_X1 U5702 ( .A1(n6784), .A2(n6785), .ZN(n6842) );
  NAND2_X1 U5703 ( .A1(n4758), .A2(n6789), .ZN(n6822) );
  INV_X1 U5704 ( .A(n4759), .ZN(n4758) );
  INV_X1 U5705 ( .A(n6876), .ZN(n4761) );
  XNOR2_X1 U5706 ( .A(n7605), .B(n7613), .ZN(n7473) );
  XNOR2_X1 U5707 ( .A(n4664), .B(n4663), .ZN(n7678) );
  OR2_X1 U5708 ( .A1(n8723), .A2(n4661), .ZN(n4660) );
  AND2_X1 U5709 ( .A1(n8732), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4661) );
  NOR2_X1 U5710 ( .A1(n8748), .A2(n8743), .ZN(n8745) );
  OR2_X1 U5711 ( .A1(n6903), .A2(n7083), .ZN(n6777) );
  OR2_X1 U5712 ( .A1(n8805), .A2(n4662), .ZN(n8785) );
  NOR2_X1 U5713 ( .A1(n8876), .A2(n8993), .ZN(n6596) );
  INV_X1 U5714 ( .A(n8385), .ZN(n8223) );
  NAND2_X1 U5715 ( .A1(n5026), .A2(n5023), .ZN(n8862) );
  INV_X1 U5716 ( .A(n5024), .ZN(n5023) );
  OAI21_X1 U5717 ( .B1(n5031), .B2(n5025), .A(n5029), .ZN(n5024) );
  NOR2_X1 U5718 ( .A1(n8876), .A2(n8953), .ZN(n4695) );
  NOR2_X1 U5719 ( .A1(n8897), .A2(n8953), .ZN(n4668) );
  NAND2_X1 U5720 ( .A1(n6167), .A2(n6166), .ZN(n6531) );
  NAND2_X1 U5721 ( .A1(n6163), .A2(n6162), .ZN(n6222) );
  INV_X1 U5722 ( .A(n6248), .ZN(n6163) );
  OR2_X1 U5723 ( .A1(n6222), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6501) );
  INV_X1 U5724 ( .A(n5079), .ZN(n5078) );
  AOI21_X1 U5725 ( .B1(n5080), .B2(n8988), .A(n6613), .ZN(n5079) );
  AND2_X1 U5726 ( .A1(n8346), .A2(n8348), .ZN(n8963) );
  OR2_X1 U5727 ( .A1(n8492), .A2(n8660), .ZN(n5012) );
  NOR2_X1 U5728 ( .A1(n9071), .A2(n8994), .ZN(n5013) );
  NOR2_X1 U5729 ( .A1(n8962), .A2(n8963), .ZN(n8961) );
  INV_X1 U5730 ( .A(n5014), .ZN(n8973) );
  NAND2_X1 U5731 ( .A1(n6161), .A2(n6160), .ZN(n6492) );
  INV_X1 U5732 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6160) );
  INV_X1 U5733 ( .A(n6490), .ZN(n6161) );
  OR2_X1 U5734 ( .A1(n6492), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6248) );
  AOI21_X1 U5735 ( .B1(n8208), .B2(n5019), .A(n4608), .ZN(n5018) );
  INV_X1 U5736 ( .A(n6471), .ZN(n5019) );
  NAND2_X1 U5737 ( .A1(n6157), .A2(n6156), .ZN(n6452) );
  INV_X1 U5738 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6156) );
  INV_X1 U5739 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6153) );
  OR2_X1 U5740 ( .A1(n6368), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U5741 ( .A1(n6603), .A2(n8244), .ZN(n7457) );
  OR2_X1 U5742 ( .A1(n6344), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U5743 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
  AND2_X1 U5744 ( .A1(n8173), .A2(n8172), .ZN(n8226) );
  OR2_X1 U5745 ( .A1(n8849), .A2(n8848), .ZN(n9457) );
  NAND2_X1 U5746 ( .A1(n6509), .A2(n6508), .ZN(n8604) );
  INV_X1 U5747 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U5748 ( .A1(n5084), .A2(n5083), .ZN(n6187) );
  AND2_X1 U5749 ( .A1(n4567), .A2(n6202), .ZN(n5083) );
  AND2_X2 U5750 ( .A1(n5156), .A2(n5155), .ZN(n5084) );
  INV_X1 U5751 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U5752 ( .A1(n6423), .A2(n6233), .ZN(n6435) );
  INV_X1 U5753 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6233) );
  INV_X1 U5754 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6461) );
  NOR2_X1 U5755 ( .A1(n9644), .A2(n9643), .ZN(n5105) );
  INV_X1 U5756 ( .A(n5104), .ZN(n5103) );
  INV_X1 U5757 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5507) );
  AOI21_X1 U5758 ( .B1(n5113), .B2(n5110), .A(n4610), .ZN(n5109) );
  INV_X1 U5759 ( .A(n4581), .ZN(n5110) );
  AND2_X1 U5760 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5478) );
  INV_X1 U5761 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U5762 ( .A1(n6029), .A2(n5091), .ZN(n5090) );
  OR2_X1 U5763 ( .A1(n5095), .A2(n5093), .ZN(n5092) );
  NAND2_X1 U5764 ( .A1(n9526), .A2(n9529), .ZN(n6030) );
  OR2_X1 U5765 ( .A1(n7038), .A2(n10458), .ZN(n6131) );
  NAND2_X1 U5766 ( .A1(n9939), .A2(n9938), .ZN(n4953) );
  NAND2_X1 U5767 ( .A1(n6695), .A2(n6694), .ZN(n6709) );
  AOI21_X1 U5768 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6996), .A(n6995), .ZN(
        n6999) );
  AOI21_X1 U5769 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10017), .A(n10011), .ZN(
        n7119) );
  AOI21_X1 U5770 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8054), .A(n8053), .ZN(
        n10024) );
  AND2_X1 U5771 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  NOR2_X1 U5772 ( .A1(n4908), .A2(n4904), .ZN(n4902) );
  NOR2_X1 U5773 ( .A1(n10208), .A2(n10194), .ZN(n10178) );
  INV_X1 U5774 ( .A(n9832), .ZN(n10190) );
  OAI21_X1 U5775 ( .B1(n10218), .B2(n9861), .A(n9851), .ZN(n4850) );
  NAND2_X1 U5776 ( .A1(n5170), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5671) );
  INV_X1 U5777 ( .A(n5656), .ZN(n5170) );
  AND2_X1 U5778 ( .A1(n10289), .A2(n4842), .ZN(n10221) );
  NOR2_X1 U5779 ( .A1(n10364), .A2(n4844), .ZN(n4842) );
  OR2_X1 U5780 ( .A1(n5644), .A2(n9613), .ZN(n5656) );
  OR2_X1 U5781 ( .A1(n5626), .A2(n9648), .ZN(n5642) );
  NAND2_X1 U5782 ( .A1(n5169), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5644) );
  INV_X1 U5783 ( .A(n5642), .ZN(n5169) );
  NAND2_X1 U5784 ( .A1(n10289), .A2(n4846), .ZN(n10250) );
  OR2_X1 U5785 ( .A1(n5611), .A2(n5365), .ZN(n5624) );
  NAND2_X1 U5786 ( .A1(n5168), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5626) );
  INV_X1 U5787 ( .A(n5624), .ZN(n5168) );
  AND2_X1 U5788 ( .A1(n10268), .A2(n10260), .ZN(n4686) );
  NOR2_X1 U5789 ( .A1(n10287), .A2(n4924), .ZN(n4923) );
  AND2_X1 U5790 ( .A1(n10307), .A2(n10293), .ZN(n10289) );
  AND2_X1 U5791 ( .A1(n9900), .A2(n10260), .ZN(n10287) );
  AOI21_X1 U5792 ( .B1(n5851), .B2(n4854), .A(n4853), .ZN(n4852) );
  INV_X1 U5793 ( .A(n5851), .ZN(n4855) );
  INV_X1 U5794 ( .A(n4856), .ZN(n4854) );
  OR2_X1 U5795 ( .A1(n8452), .A2(n9534), .ZN(n10309) );
  OR2_X1 U5796 ( .A1(n5575), .A2(n5574), .ZN(n5577) );
  INV_X1 U5797 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9623) );
  OR2_X1 U5798 ( .A1(n5577), .A2(n9623), .ZN(n5594) );
  OR2_X1 U5799 ( .A1(n10503), .A2(n5582), .ZN(n9739) );
  AND2_X1 U5800 ( .A1(n9739), .A2(n9893), .ZN(n9821) );
  AND2_X1 U5801 ( .A1(n7857), .A2(n4575), .ZN(n8453) );
  AND2_X1 U5802 ( .A1(n5544), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5803 ( .A1(n7857), .A2(n4838), .ZN(n7976) );
  OR2_X1 U5804 ( .A1(n10486), .A2(n9977), .ZN(n5552) );
  NAND2_X1 U5805 ( .A1(n7857), .A2(n10618), .ZN(n7801) );
  NAND2_X1 U5806 ( .A1(n7844), .A2(n5165), .ZN(n7757) );
  NAND2_X1 U5807 ( .A1(n7757), .A2(n7756), .ZN(n7755) );
  AND2_X1 U5808 ( .A1(n7856), .A2(n10525), .ZN(n7857) );
  AND2_X1 U5809 ( .A1(n9713), .A2(n7850), .ZN(n9711) );
  NAND2_X1 U5810 ( .A1(n10211), .A2(n5888), .ZN(n5883) );
  AOI21_X1 U5811 ( .B1(n6324), .B2(n5337), .A(n4806), .ZN(n4805) );
  NOR2_X1 U5812 ( .A1(n6688), .A2(n6963), .ZN(n4806) );
  NAND2_X1 U5813 ( .A1(n10602), .A2(n4580), .ZN(n7594) );
  NAND2_X1 U5814 ( .A1(n4835), .A2(n4836), .ZN(n7290) );
  AND2_X1 U5815 ( .A1(n7450), .A2(n7503), .ZN(n4835) );
  INV_X1 U5816 ( .A(n9959), .ZN(n5755) );
  AND2_X1 U5817 ( .A1(n9866), .A2(n9913), .ZN(n9838) );
  AND2_X1 U5818 ( .A1(n10369), .A2(n9968), .ZN(n5647) );
  AND2_X1 U5819 ( .A1(n9906), .A2(n9869), .ZN(n10236) );
  AND2_X1 U5820 ( .A1(n9905), .A2(n9760), .ZN(n10246) );
  AND2_X1 U5821 ( .A1(n10245), .A2(n9753), .ZN(n10268) );
  INV_X1 U5822 ( .A(n4912), .ZN(n4910) );
  INV_X1 U5823 ( .A(n7975), .ZN(n4911) );
  INV_X1 U5824 ( .A(n10617), .ZN(n10626) );
  NOR2_X1 U5825 ( .A1(n6858), .A2(n6857), .ZN(n7261) );
  XNOR2_X1 U5826 ( .A(n8162), .B(n8163), .ZN(n5760) );
  NAND2_X1 U5827 ( .A1(n5760), .A2(SI_29_), .ZN(n8166) );
  AND2_X1 U5828 ( .A1(n5758), .A2(n5322), .ZN(n5756) );
  NAND2_X1 U5829 ( .A1(n5325), .A2(n10461), .ZN(n4900) );
  NAND2_X1 U5830 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U5831 ( .A(n5784), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5793) );
  AND2_X1 U5832 ( .A1(n5299), .A2(n5298), .ZN(n5678) );
  XNOR2_X1 U5833 ( .A(n5667), .B(n5666), .ZN(n7931) );
  INV_X1 U5834 ( .A(SI_20_), .ZN(n5333) );
  INV_X1 U5835 ( .A(n4946), .ZN(n5620) );
  AOI21_X1 U5836 ( .B1(n5602), .B2(n4951), .A(n4949), .ZN(n4946) );
  OAI21_X1 U5837 ( .B1(n5602), .B2(n5265), .A(n5264), .ZN(n5361) );
  NAND2_X1 U5838 ( .A1(n4963), .A2(n5249), .ZN(n5568) );
  NAND2_X1 U5839 ( .A1(n5243), .A2(n4964), .ZN(n4963) );
  NAND2_X1 U5840 ( .A1(n5243), .A2(n5242), .ZN(n5554) );
  NAND2_X1 U5841 ( .A1(n5231), .A2(n5230), .ZN(n5502) );
  NOR2_X1 U5842 ( .A1(n4870), .A2(n4585), .ZN(n5489) );
  NOR2_X1 U5843 ( .A1(n8139), .A2(n10730), .ZN(n8141) );
  NAND2_X1 U5844 ( .A1(n7422), .A2(n7421), .ZN(n7429) );
  NAND2_X1 U5845 ( .A1(n4716), .A2(n5136), .ZN(n8521) );
  NAND2_X1 U5846 ( .A1(n4716), .A2(n4714), .ZN(n8545) );
  NAND2_X1 U5847 ( .A1(n4707), .A2(n4708), .ZN(n8494) );
  NAND2_X1 U5848 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  NAND2_X1 U5849 ( .A1(n8612), .A2(n5134), .ZN(n8538) );
  AOI21_X1 U5850 ( .B1(n4714), .B2(n4712), .A(n4711), .ZN(n4710) );
  INV_X1 U5851 ( .A(n4714), .ZN(n4713) );
  INV_X1 U5852 ( .A(n8544), .ZN(n4711) );
  NAND2_X1 U5853 ( .A1(n6554), .A2(n6553), .ZN(n8552) );
  NAND2_X1 U5854 ( .A1(n6926), .A2(n6928), .ZN(n7099) );
  OAI21_X1 U5855 ( .B1(n8612), .B2(n5126), .A(n5125), .ZN(n8555) );
  NAND2_X1 U5856 ( .A1(n6500), .A2(n6499), .ZN(n8560) );
  NAND2_X1 U5857 ( .A1(n8022), .A2(n5149), .ZN(n8083) );
  OR2_X1 U5858 ( .A1(n8023), .A2(n8028), .ZN(n5149) );
  AOI21_X1 U5859 ( .B1(n8589), .B2(n8590), .A(n5147), .ZN(n8563) );
  AND4_X1 U5860 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n7282)
         );
  NAND2_X1 U5861 ( .A1(n6207), .A2(n6206), .ZN(n8594) );
  AND2_X1 U5862 ( .A1(n7161), .A2(n7160), .ZN(n7167) );
  AND2_X1 U5863 ( .A1(n7050), .A2(n6917), .ZN(n8639) );
  NAND2_X1 U5864 ( .A1(n7636), .A2(n5150), .ZN(n7882) );
  AND2_X1 U5865 ( .A1(n7638), .A2(n7635), .ZN(n5150) );
  AND2_X1 U5866 ( .A1(n7636), .A2(n7635), .ZN(n7639) );
  NAND2_X1 U5867 ( .A1(n5129), .A2(n5130), .ZN(n8597) );
  NAND2_X1 U5868 ( .A1(n8612), .A2(n5131), .ZN(n5129) );
  OAI21_X1 U5869 ( .B1(n8615), .B2(n4718), .A(n4717), .ZN(n8607) );
  NAND2_X1 U5870 ( .A1(n5121), .A2(n8503), .ZN(n4718) );
  NAND2_X1 U5871 ( .A1(n5121), .A2(n4573), .ZN(n4717) );
  NAND2_X1 U5872 ( .A1(n8607), .A2(n8606), .ZN(n8605) );
  INV_X1 U5873 ( .A(n8664), .ZN(n7965) );
  NAND2_X1 U5874 ( .A1(n7962), .A2(n8023), .ZN(n8022) );
  NAND2_X1 U5875 ( .A1(n5137), .A2(n5142), .ZN(n8622) );
  NAND2_X1 U5876 ( .A1(n8589), .A2(n5145), .ZN(n5137) );
  NAND2_X1 U5877 ( .A1(n6914), .A2(n9018), .ZN(n8629) );
  NAND2_X1 U5878 ( .A1(n4707), .A2(n4640), .ZN(n8636) );
  AND2_X1 U5879 ( .A1(n4707), .A2(n4579), .ZN(n8638) );
  INV_X1 U5880 ( .A(n8632), .ZN(n8635) );
  OAI21_X1 U5881 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(n4874) );
  OR2_X1 U5882 ( .A1(n8404), .A2(n6896), .ZN(n4876) );
  XNOR2_X1 U5883 ( .A(n6576), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8411) );
  AND2_X1 U5884 ( .A1(n8181), .A2(n6593), .ZN(n8186) );
  NAND2_X1 U5885 ( .A1(n6198), .A2(n6197), .ZN(n8653) );
  INV_X1 U5886 ( .A(n7282), .ZN(n8672) );
  CLKBUF_X1 U5887 ( .A(n8674), .Z(n4669) );
  OR2_X1 U5888 ( .A1(n6548), .A2(n7375), .ZN(n6274) );
  OR2_X2 U5889 ( .A1(n6777), .A2(P2_U3151), .ZN(n8676) );
  AND2_X1 U5890 ( .A1(n4739), .A2(n6804), .ZN(n6825) );
  NAND2_X1 U5891 ( .A1(n4745), .A2(n6885), .ZN(n4744) );
  NOR2_X1 U5892 ( .A1(n7227), .A2(n4754), .ZN(n7152) );
  AND2_X1 U5893 ( .A1(n4653), .A2(n4978), .ZN(n7216) );
  OAI21_X1 U5894 ( .B1(n7219), .B2(n7218), .A(n4749), .ZN(n7471) );
  AND2_X1 U5895 ( .A1(n7217), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4977) );
  INV_X1 U5896 ( .A(n5045), .ZN(n7618) );
  NAND2_X1 U5897 ( .A1(n4976), .A2(n4975), .ZN(n7677) );
  INV_X1 U5898 ( .A(n7609), .ZN(n4975) );
  INV_X1 U5899 ( .A(n4976), .ZN(n7610) );
  NOR2_X1 U5900 ( .A1(n7810), .A2(n7809), .ZN(n7813) );
  INV_X1 U5901 ( .A(n4733), .ZN(n7983) );
  NOR2_X1 U5902 ( .A1(n7987), .A2(n7986), .ZN(n8698) );
  INV_X1 U5903 ( .A(n8715), .ZN(n4982) );
  OAI21_X1 U5904 ( .B1(n7987), .B2(n5054), .A(n5053), .ZN(n8731) );
  NAND2_X1 U5905 ( .A1(n5055), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5054) );
  INV_X1 U5906 ( .A(n8700), .ZN(n5055) );
  XNOR2_X1 U5907 ( .A(n4660), .B(n4659), .ZN(n8724) );
  OR2_X1 U5908 ( .A1(n8733), .A2(n9270), .ZN(n5042) );
  INV_X1 U5909 ( .A(n8745), .ZN(n5041) );
  INV_X1 U5910 ( .A(n4730), .ZN(n8751) );
  OAI21_X1 U5911 ( .B1(n5040), .B2(n8733), .A(n5039), .ZN(n8769) );
  NAND2_X1 U5912 ( .A1(n5043), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U5913 ( .A1(n8745), .A2(n5043), .ZN(n5039) );
  INV_X1 U5914 ( .A(n8746), .ZN(n5043) );
  NAND2_X1 U5915 ( .A1(n6833), .A2(n6782), .ZN(n8841) );
  NOR2_X1 U5916 ( .A1(n8827), .A2(n4735), .ZN(n8830) );
  NOR2_X1 U5917 ( .A1(n8833), .A2(n8814), .ZN(n4735) );
  INV_X1 U5918 ( .A(n5069), .ZN(n8878) );
  AOI21_X1 U5919 ( .B1(n5074), .B2(n4563), .A(n5070), .ZN(n5069) );
  INV_X1 U5920 ( .A(n8379), .ZN(n5070) );
  OAI21_X1 U5921 ( .B1(n8886), .B2(n8990), .A(n4683), .ZN(n9039) );
  NOR2_X1 U5922 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  NOR2_X1 U5923 ( .A1(n8908), .A2(n8993), .ZN(n4684) );
  NAND2_X1 U5924 ( .A1(n5074), .A2(n5075), .ZN(n8889) );
  NAND2_X1 U5925 ( .A1(n4992), .A2(n4993), .ZN(n8917) );
  NAND2_X1 U5926 ( .A1(n4997), .A2(n4998), .ZN(n8927) );
  NAND2_X1 U5927 ( .A1(n8947), .A2(n4999), .ZN(n4997) );
  NAND2_X1 U5928 ( .A1(n8947), .A2(n5002), .ZN(n8937) );
  NAND2_X1 U5929 ( .A1(n6216), .A2(n6215), .ZN(n9062) );
  NAND2_X1 U5930 ( .A1(n5022), .A2(n6471), .ZN(n9011) );
  NAND2_X1 U5931 ( .A1(n6460), .A2(n5020), .ZN(n5022) );
  AND2_X1 U5932 ( .A1(n8326), .A2(n8324), .ZN(n5085) );
  NAND2_X1 U5933 ( .A1(n6460), .A2(n6459), .ZN(n8001) );
  NAND2_X1 U5934 ( .A1(n6611), .A2(n6610), .ZN(n8039) );
  NAND2_X1 U5935 ( .A1(n6437), .A2(n6436), .ZN(n8318) );
  INV_X1 U5936 ( .A(n9023), .ZN(n9002) );
  NOR2_X2 U5937 ( .A1(n9000), .A2(n7654), .ZN(n9004) );
  OAI21_X1 U5938 ( .B1(n4658), .B2(n5009), .A(n5007), .ZN(n7903) );
  NAND2_X1 U5939 ( .A1(n7264), .A2(n8281), .ZN(n7210) );
  NAND2_X1 U5940 ( .A1(n6324), .A2(n4541), .ZN(n5036) );
  OR2_X1 U5941 ( .A1(n6913), .A2(n6912), .ZN(n9018) );
  INV_X1 U5942 ( .A(n9018), .ZN(n8999) );
  INV_X1 U5943 ( .A(n8226), .ZN(n9459) );
  NOR2_X1 U5944 ( .A1(n9034), .A2(n5163), .ZN(n9471) );
  INV_X1 U5945 ( .A(n8630), .ZN(n9481) );
  NOR2_X1 U5946 ( .A1(n9039), .A2(n4682), .ZN(n9478) );
  AND2_X1 U5947 ( .A1(n9040), .A2(n9449), .ZN(n4682) );
  NOR2_X1 U5948 ( .A1(n9044), .A2(n4596), .ZN(n9482) );
  INV_X1 U5949 ( .A(n8594), .ZN(n9489) );
  INV_X1 U5950 ( .A(n8533), .ZN(n9493) );
  INV_X1 U5951 ( .A(n8604), .ZN(n9497) );
  INV_X1 U5952 ( .A(n8560), .ZN(n9501) );
  OR2_X1 U5953 ( .A1(n9075), .A2(n9074), .ZN(n9510) );
  INV_X1 U5954 ( .A(n8580), .ZN(n9515) );
  INV_X1 U5955 ( .A(n8107), .ZN(n8118) );
  NAND2_X1 U5956 ( .A1(n6644), .A2(n6643), .ZN(n6899) );
  AND2_X1 U5957 ( .A1(n6903), .A2(n6909), .ZN(n6915) );
  INV_X1 U5958 ( .A(n6642), .ZN(n8102) );
  OR2_X1 U5959 ( .A1(n6629), .A2(n6634), .ZN(n6630) );
  INV_X1 U5960 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7942) );
  INV_X1 U5961 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9186) );
  INV_X1 U5962 ( .A(n8411), .ZN(n7932) );
  INV_X1 U5963 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U5964 ( .A1(n6628), .A2(n6579), .ZN(n8262) );
  INV_X1 U5965 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9185) );
  INV_X1 U5966 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6237) );
  INV_X1 U5967 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7331) );
  INV_X1 U5968 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7303) );
  INV_X1 U5969 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7177) );
  INV_X1 U5970 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7181) );
  XNOR2_X1 U5971 ( .A(n6462), .B(n6461), .ZN(n8732) );
  INV_X1 U5972 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6893) );
  INV_X1 U5973 ( .A(n7829), .ZN(n7988) );
  INV_X1 U5974 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9274) );
  INV_X1 U5975 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9151) );
  INV_X1 U5976 ( .A(n4985), .ZN(n6768) );
  NAND2_X1 U5977 ( .A1(n4819), .A2(n4818), .ZN(n8472) );
  AOI21_X1 U5978 ( .B1(n4821), .B2(n4816), .A(n4647), .ZN(n4818) );
  NAND2_X1 U5979 ( .A1(n4814), .A2(n4812), .ZN(n4819) );
  NOR2_X1 U5980 ( .A1(n8471), .A2(n4647), .ZN(n5114) );
  OR2_X1 U5981 ( .A1(n5762), .A2(n6723), .ZN(n5442) );
  INV_X1 U5982 ( .A(n5099), .ZN(n9556) );
  AOI21_X1 U5983 ( .B1(n9646), .B2(n5100), .A(n5103), .ZN(n5099) );
  INV_X1 U5984 ( .A(n5105), .ZN(n5100) );
  AND2_X1 U5985 ( .A1(n6128), .A2(n10527), .ZN(n6129) );
  NAND2_X1 U5986 ( .A1(n5332), .A2(n5331), .ZN(n10326) );
  NAND2_X1 U5987 ( .A1(n5932), .A2(n5931), .ZN(n7308) );
  INV_X1 U5988 ( .A(n7306), .ZN(n5931) );
  INV_X1 U5989 ( .A(n4665), .ZN(n9566) );
  CLKBUF_X1 U5990 ( .A(n5096), .Z(n4665) );
  NAND2_X1 U5991 ( .A1(n9619), .A2(n9620), .ZN(n9618) );
  NAND2_X1 U5992 ( .A1(n10499), .A2(n6010), .ZN(n9619) );
  NAND2_X1 U5993 ( .A1(n6083), .A2(n6080), .ZN(n9635) );
  CLKBUF_X1 U5994 ( .A(n10493), .Z(n10494) );
  NAND2_X1 U5995 ( .A1(n10480), .A2(n4808), .ZN(n10512) );
  AND2_X1 U5996 ( .A1(n4809), .A2(n10511), .ZN(n4808) );
  CLKBUF_X1 U5997 ( .A(n10502), .Z(n10515) );
  OR2_X1 U5998 ( .A1(n5420), .A2(n6719), .ZN(n5424) );
  OR2_X1 U5999 ( .A1(n6720), .A2(n5762), .ZN(n5423) );
  NAND2_X1 U6000 ( .A1(n5359), .A2(n5358), .ZN(n10374) );
  INV_X1 U6001 ( .A(n10492), .ZN(n10541) );
  AND2_X1 U6002 ( .A1(n4822), .A2(n4823), .ZN(n9655) );
  INV_X1 U6003 ( .A(n10535), .ZN(n10527) );
  NAND2_X1 U6004 ( .A1(n6132), .A2(n6124), .ZN(n10535) );
  NAND2_X1 U6005 ( .A1(n6137), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10547) );
  INV_X1 U6006 ( .A(n9933), .ZN(n9943) );
  NAND2_X1 U6007 ( .A1(n5753), .A2(n5752), .ZN(n9960) );
  NAND2_X1 U6008 ( .A1(n5719), .A2(n5718), .ZN(n9962) );
  NAND2_X1 U6009 ( .A1(n5700), .A2(n5699), .ZN(n9963) );
  NAND2_X1 U6010 ( .A1(n5689), .A2(n5688), .ZN(n9964) );
  NAND2_X1 U6011 ( .A1(n5695), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5417) );
  OR2_X1 U6012 ( .A1(n5458), .A2(n7242), .ZN(n5414) );
  AOI21_X1 U6013 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n4690), .A(n10001), .ZN(
        n6708) );
  INV_X1 U6014 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9412) );
  AOI21_X1 U6015 ( .B1(n6959), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6958), .ZN(
        n6962) );
  NAND2_X1 U6016 ( .A1(n7003), .A2(n4679), .ZN(n7007) );
  OR2_X1 U6017 ( .A1(n7004), .A2(n7005), .ZN(n4679) );
  NAND2_X1 U6018 ( .A1(n7007), .A2(n7006), .ZN(n7108) );
  AOI21_X1 U6019 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10017), .A(n7111), .ZN(
        n7112) );
  AOI21_X1 U6020 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7395), .A(n7389), .ZN(
        n7392) );
  AOI21_X1 U6021 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7871), .A(n7866), .ZN(
        n7869) );
  AOI21_X1 U6022 ( .B1(n7871), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7870), .ZN(
        n7873) );
  AND2_X1 U6023 ( .A1(n6944), .A2(n6697), .ZN(n10093) );
  NOR2_X1 U6024 ( .A1(n10102), .A2(n10308), .ZN(n10315) );
  AND2_X1 U6025 ( .A1(n10137), .A2(n4576), .ZN(n10101) );
  NAND2_X1 U6026 ( .A1(n9836), .A2(n4904), .ZN(n4903) );
  NOR2_X1 U6027 ( .A1(n10116), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U6028 ( .A1(n4901), .A2(n4905), .ZN(n10324) );
  AND2_X1 U6029 ( .A1(n10116), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U6030 ( .A1(n5735), .A2(n4902), .ZN(n4901) );
  NAND2_X1 U6031 ( .A1(n8423), .A2(n4909), .ZN(n4906) );
  NAND2_X1 U6032 ( .A1(n5847), .A2(n9894), .ZN(n8063) );
  NAND2_X1 U6033 ( .A1(n4915), .A2(n4914), .ZN(n8067) );
  NAND2_X1 U6034 ( .A1(n5382), .A2(n5381), .ZN(n8456) );
  AND2_X1 U6035 ( .A1(n4915), .A2(n4917), .ZN(n8449) );
  OR2_X1 U6036 ( .A1(n5830), .A2(n10211), .ZN(n10275) );
  INV_X1 U6037 ( .A(n10275), .ZN(n10548) );
  INV_X1 U6038 ( .A(n8491), .ZN(n4674) );
  NAND2_X1 U6039 ( .A1(n5735), .A2(n5734), .ZN(n8418) );
  OAI21_X1 U6040 ( .B1(n10187), .B2(n4933), .A(n4931), .ZN(n10145) );
  NAND2_X1 U6041 ( .A1(n4936), .A2(n4937), .ZN(n10159) );
  NAND2_X1 U6042 ( .A1(n10187), .A2(n4939), .ZN(n4936) );
  OAI21_X1 U6043 ( .B1(n10187), .B2(n4582), .A(n4941), .ZN(n10173) );
  AND2_X1 U6044 ( .A1(n10449), .A2(n10626), .ZN(n10453) );
  NAND2_X1 U6045 ( .A1(n6685), .A2(n6674), .ZN(n10458) );
  AND2_X1 U6046 ( .A1(n5190), .A2(n5191), .ZN(n5119) );
  INV_X1 U6047 ( .A(n5323), .ZN(n5120) );
  INV_X1 U6048 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5191) );
  CLKBUF_X1 U6049 ( .A(n5870), .Z(n5871) );
  XNOR2_X1 U6050 ( .A(n5757), .B(n5756), .ZN(n8159) );
  INV_X1 U6051 ( .A(n5777), .ZN(n5780) );
  INV_X1 U6052 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7939) );
  INV_X1 U6053 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U6054 ( .A1(n5809), .A2(n5808), .ZN(n7933) );
  XNOR2_X1 U6055 ( .A(n5811), .B(n5810), .ZN(n9807) );
  INV_X1 U6056 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9174) );
  INV_X1 U6057 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7333) );
  INV_X1 U6058 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7176) );
  INV_X1 U6059 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7180) );
  INV_X1 U6060 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9295) );
  AND2_X1 U6061 ( .A1(n5541), .A2(n5555), .ZN(n7356) );
  INV_X1 U6062 ( .A(n6324), .ZN(n6731) );
  XNOR2_X1 U6063 ( .A(n5421), .B(n5422), .ZN(n6720) );
  XNOR2_X1 U6064 ( .A(n5399), .B(n5398), .ZN(n6727) );
  INV_X1 U6065 ( .A(n4987), .ZN(n4986) );
  INV_X1 U6066 ( .A(n4983), .ZN(n8714) );
  AND2_X1 U6067 ( .A1(n8821), .A2(n4652), .ZN(n4765) );
  OAI21_X1 U6068 ( .B1(n4614), .B2(n4764), .A(n8833), .ZN(n4763) );
  OAI21_X1 U6069 ( .B1(n9463), .B2(n4671), .A(n6673), .ZN(P2_U3488) );
  OAI21_X1 U6070 ( .B1(n9475), .B2(n4671), .A(n4648), .ZN(P2_U3486) );
  NAND2_X1 U6071 ( .A1(n4671), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n4670) );
  OAI21_X1 U6072 ( .B1(n9475), .B2(n10685), .A(n4680), .ZN(P2_U3454) );
  AOI21_X1 U6073 ( .B1(n8518), .B2(n9467), .A(n4681), .ZN(n4680) );
  NOR2_X1 U6074 ( .A1(n10683), .A2(n9476), .ZN(n4681) );
  NAND2_X1 U6075 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  AOI21_X1 U6076 ( .B1(n8488), .B2(n10643), .A(n4858), .ZN(n8490) );
  NAND2_X1 U6077 ( .A1(n4860), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U6078 ( .A1(n10641), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4859) );
  OR2_X1 U6079 ( .A1(n8594), .A2(n8919), .ZN(n8363) );
  INV_X1 U6080 ( .A(n7151), .ZN(n5049) );
  INV_X2 U6081 ( .A(n5762), .ZN(n5337) );
  INV_X1 U6082 ( .A(n6722), .ZN(n4690) );
  NOR2_X1 U6083 ( .A1(n9567), .A2(n6071), .ZN(n4562) );
  AND2_X1 U6084 ( .A1(n5075), .A2(n8378), .ZN(n4563) );
  NAND2_X1 U6085 ( .A1(n5516), .A2(n5519), .ZN(n4564) );
  NAND2_X1 U6086 ( .A1(n10384), .A2(n9971), .ZN(n4565) );
  AND2_X1 U6087 ( .A1(n5829), .A2(n4849), .ZN(n4566) );
  INV_X1 U6088 ( .A(n9836), .ZN(n8423) );
  AND4_X1 U6089 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n5154), .ZN(n4567)
         );
  OR2_X1 U6090 ( .A1(n9859), .A2(n9941), .ZN(n4568) );
  AND4_X1 U6091 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5486), .ZN(n4569)
         );
  AND2_X1 U6092 ( .A1(n4914), .A2(n5600), .ZN(n4570) );
  INV_X1 U6093 ( .A(n8665), .ZN(n8028) );
  AND2_X1 U6094 ( .A1(n4565), .A2(n5631), .ZN(n4571) );
  AND2_X1 U6095 ( .A1(n5185), .A2(n5186), .ZN(n4572) );
  OR2_X1 U6096 ( .A1(n5124), .A2(n4719), .ZN(n4573) );
  AND2_X1 U6097 ( .A1(n8516), .A2(n8897), .ZN(n4574) );
  AND2_X1 U6098 ( .A1(n4838), .A2(n4837), .ZN(n4575) );
  AND2_X1 U6099 ( .A1(n4566), .A2(n4848), .ZN(n4576) );
  AND2_X1 U6100 ( .A1(n7426), .A2(n7421), .ZN(n4577) );
  INV_X1 U6101 ( .A(n6024), .ZN(n4825) );
  INV_X1 U6102 ( .A(n9579), .ZN(n4816) );
  OR3_X1 U6103 ( .A1(n6435), .A2(n5158), .A3(P2_IR_REG_16__SCAN_IN), .ZN(n4578) );
  INV_X1 U6104 ( .A(n5734), .ZN(n4904) );
  NAND2_X1 U6105 ( .A1(n7857), .A2(n4840), .ZN(n4841) );
  INV_X1 U6106 ( .A(n8518), .ZN(n9477) );
  NAND2_X1 U6107 ( .A1(n6541), .A2(n6540), .ZN(n8518) );
  AND2_X1 U6108 ( .A1(n4708), .A2(n4645), .ZN(n4579) );
  NAND2_X1 U6109 ( .A1(n6884), .A2(n4651), .ZN(n4745) );
  OAI211_X1 U6110 ( .C1(n6688), .C2(n6722), .A(n5442), .B(n5441), .ZN(n9551)
         );
  AND4_X1 U6111 ( .A1(n7513), .A2(n4836), .A3(n7503), .A4(n7450), .ZN(n4580)
         );
  NAND2_X1 U6112 ( .A1(n6089), .A2(n6088), .ZN(n4581) );
  NAND2_X1 U6113 ( .A1(n5323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NOR2_X1 U6114 ( .A1(n4942), .A2(n6082), .ZN(n4582) );
  OR2_X1 U6115 ( .A1(n8748), .A2(n8747), .ZN(n4583) );
  INV_X1 U6116 ( .A(n9894), .ZN(n4857) );
  AND2_X1 U6117 ( .A1(n5111), .A2(n4581), .ZN(n4584) );
  NOR2_X1 U6118 ( .A1(n5224), .A2(n5223), .ZN(n4585) );
  AND2_X1 U6119 ( .A1(n4968), .A2(n5230), .ZN(n4586) );
  INV_X1 U6120 ( .A(n9840), .ZN(n4771) );
  NAND2_X1 U6121 ( .A1(n8630), .A2(n8653), .ZN(n4587) );
  OR2_X1 U6122 ( .A1(n7637), .A2(n7885), .ZN(n4588) );
  NAND2_X1 U6123 ( .A1(n5623), .A2(n5622), .ZN(n10443) );
  AND2_X1 U6124 ( .A1(n8536), .A2(n8977), .ZN(n4589) );
  INV_X1 U6125 ( .A(n9746), .ZN(n4853) );
  INV_X1 U6126 ( .A(n8668), .ZN(n7633) );
  AND2_X1 U6127 ( .A1(n8359), .A2(n8392), .ZN(n4590) );
  OR2_X1 U6128 ( .A1(n10411), .A2(n9962), .ZN(n4591) );
  NAND2_X1 U6129 ( .A1(n5669), .A2(n5668), .ZN(n10194) );
  INV_X1 U6130 ( .A(n10194), .ZN(n4942) );
  INV_X1 U6131 ( .A(n8285), .ZN(n5063) );
  OR2_X1 U6132 ( .A1(n9851), .A2(n9795), .ZN(n4592) );
  AND2_X1 U6133 ( .A1(n5891), .A2(n5957), .ZN(n4593) );
  NOR2_X1 U6134 ( .A1(n8811), .A2(n8832), .ZN(n4594) );
  OR2_X1 U6135 ( .A1(n8533), .A2(n8656), .ZN(n4595) );
  NOR2_X1 U6136 ( .A1(n8980), .A2(n5081), .ZN(n5080) );
  AND2_X1 U6137 ( .A1(n9045), .A2(n9449), .ZN(n4596) );
  OR2_X1 U6138 ( .A1(n8360), .A2(n8402), .ZN(n4597) );
  NAND2_X1 U6139 ( .A1(n5743), .A2(n5742), .ZN(n8479) );
  NAND2_X1 U6140 ( .A1(n5558), .A2(n5557), .ZN(n10625) );
  AND2_X1 U6141 ( .A1(n8332), .A2(n8331), .ZN(n9010) );
  NOR2_X1 U6142 ( .A1(n8109), .A2(n4709), .ZN(n4598) );
  OR2_X1 U6143 ( .A1(n8342), .A2(n8402), .ZN(n4599) );
  OR2_X1 U6144 ( .A1(n7613), .A2(n7605), .ZN(n4600) );
  NOR2_X1 U6145 ( .A1(n4996), .A2(n8931), .ZN(n4995) );
  INV_X1 U6146 ( .A(n6869), .ZN(n8684) );
  AND2_X1 U6147 ( .A1(n6329), .A2(n6340), .ZN(n6869) );
  INV_X1 U6149 ( .A(n5889), .ZN(n4832) );
  AND2_X1 U6150 ( .A1(n5813), .A2(n5355), .ZN(n4601) );
  INV_X1 U6151 ( .A(n5132), .ZN(n5131) );
  NAND2_X1 U6152 ( .A1(n5135), .A2(n5134), .ZN(n5132) );
  NOR2_X1 U6153 ( .A1(n8456), .A2(n9974), .ZN(n4602) );
  AND2_X1 U6154 ( .A1(n10190), .A2(n4592), .ZN(n4603) );
  AND2_X1 U6155 ( .A1(n9965), .A2(n5668), .ZN(n4604) );
  INV_X1 U6156 ( .A(n5631), .ZN(n4925) );
  INV_X1 U6157 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4726) );
  AND2_X1 U6158 ( .A1(n10274), .A2(n5852), .ZN(n4605) );
  AND2_X1 U6159 ( .A1(n6235), .A2(n4705), .ZN(n4606) );
  INV_X1 U6160 ( .A(n5600), .ZN(n4916) );
  AND2_X1 U6161 ( .A1(n6017), .A2(n6016), .ZN(n4607) );
  AND2_X1 U6162 ( .A1(n9444), .A2(n8661), .ZN(n4608) );
  INV_X1 U6163 ( .A(n5008), .ZN(n5007) );
  NOR2_X1 U6164 ( .A1(n5010), .A2(n8028), .ZN(n5008) );
  INV_X1 U6165 ( .A(n5035), .ZN(n5032) );
  NOR2_X1 U6166 ( .A1(n9043), .A2(n8654), .ZN(n5035) );
  INV_X1 U6167 ( .A(n5034), .ZN(n5033) );
  NAND2_X1 U6168 ( .A1(n9481), .A2(n8897), .ZN(n5034) );
  NAND2_X1 U6169 ( .A1(n8330), .A2(n9010), .ZN(n4609) );
  INV_X1 U6170 ( .A(n5153), .ZN(n5152) );
  OAI21_X1 U6171 ( .B1(n5154), .B2(n9518), .A(n6666), .ZN(n5153) );
  NOR2_X1 U6172 ( .A1(n6095), .A2(n6094), .ZN(n4610) );
  OR2_X1 U6173 ( .A1(n5351), .A2(n5118), .ZN(n4611) );
  INV_X1 U6174 ( .A(n4844), .ZN(n4843) );
  NAND2_X1 U6175 ( .A1(n4846), .A2(n4845), .ZN(n4844) );
  INV_X1 U6176 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U6177 ( .A1(n10341), .A2(n9963), .ZN(n4612) );
  NOR2_X1 U6178 ( .A1(n8604), .A2(n8657), .ZN(n4613) );
  AND2_X1 U6179 ( .A1(n8808), .A2(n8814), .ZN(n4614) );
  NAND2_X1 U6180 ( .A1(n5325), .A2(n5186), .ZN(n4615) );
  NOR2_X1 U6181 ( .A1(n6071), .A2(n9568), .ZN(n4616) );
  INV_X1 U6182 ( .A(n5127), .ZN(n5126) );
  NOR2_X1 U6183 ( .A1(n8598), .A2(n5128), .ZN(n5127) );
  AND2_X1 U6184 ( .A1(n5251), .A2(SI_12_), .ZN(n4617) );
  NAND2_X1 U6185 ( .A1(n8508), .A2(n8952), .ZN(n4618) );
  INV_X1 U6186 ( .A(n9859), .ZN(n9775) );
  AND2_X1 U6187 ( .A1(n10406), .A2(n5863), .ZN(n9859) );
  AND2_X1 U6188 ( .A1(n7093), .A2(n7089), .ZN(n4619) );
  OR2_X1 U6189 ( .A1(n4782), .A2(n4781), .ZN(n4620) );
  AND2_X1 U6190 ( .A1(n8358), .A2(n8360), .ZN(n8940) );
  AND2_X1 U6191 ( .A1(n9534), .A2(n9973), .ZN(n4621) );
  INV_X1 U6192 ( .A(n5122), .ZN(n5121) );
  OAI21_X1 U6193 ( .B1(n5125), .B2(n5123), .A(n4618), .ZN(n5122) );
  NAND2_X1 U6194 ( .A1(n4864), .A2(n4866), .ZN(n4622) );
  OR2_X1 U6195 ( .A1(n6277), .A2(n4985), .ZN(n4623) );
  OR2_X1 U6196 ( .A1(n10607), .A2(n9980), .ZN(n4624) );
  AND2_X1 U6197 ( .A1(n9038), .A2(n9449), .ZN(n4625) );
  OR2_X1 U6198 ( .A1(n7613), .A2(n7612), .ZN(n4626) );
  AND2_X1 U6199 ( .A1(n4993), .A2(n4595), .ZN(n4627) );
  NAND2_X1 U6200 ( .A1(n6688), .A2(n5330), .ZN(n5762) );
  OR2_X1 U6201 ( .A1(n9743), .A2(n9741), .ZN(n4628) );
  OR2_X1 U6202 ( .A1(n8515), .A2(n8654), .ZN(n4629) );
  AND2_X1 U6203 ( .A1(n6366), .A2(n8668), .ZN(n4630) );
  OR2_X1 U6204 ( .A1(n7230), .A2(n4753), .ZN(n4631) );
  AND2_X1 U6205 ( .A1(n4907), .A2(n4903), .ZN(n4632) );
  OR2_X1 U6206 ( .A1(n9493), .A2(n8929), .ZN(n4633) );
  NAND2_X1 U6207 ( .A1(n8580), .A2(n9015), .ZN(n4634) );
  AND2_X1 U6208 ( .A1(n4572), .A2(n5190), .ZN(n4635) );
  AND2_X1 U6209 ( .A1(n4862), .A2(n4599), .ZN(n4636) );
  INV_X1 U6210 ( .A(n9604), .ZN(n5113) );
  NAND2_X1 U6211 ( .A1(n9791), .A2(n9790), .ZN(n10108) );
  INV_X1 U6212 ( .A(n10108), .ZN(n4848) );
  NAND2_X1 U6213 ( .A1(n8088), .A2(n4598), .ZN(n4707) );
  INV_X1 U6214 ( .A(n7162), .ZN(n8517) );
  NAND2_X1 U6215 ( .A1(n5641), .A2(n5640), .ZN(n10369) );
  INV_X1 U6216 ( .A(n10369), .ZN(n4845) );
  XNOR2_X1 U6217 ( .A(n5779), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5795) );
  INV_X1 U6218 ( .A(n6029), .ZN(n5093) );
  INV_X1 U6219 ( .A(n10260), .ZN(n4804) );
  INV_X1 U6220 ( .A(n9869), .ZN(n4851) );
  AND2_X1 U6221 ( .A1(n4922), .A2(n4565), .ZN(n4637) );
  AND2_X1 U6222 ( .A1(n6384), .A2(n6383), .ZN(n7613) );
  INV_X1 U6223 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U6224 ( .A1(n5782), .A2(n5781), .ZN(n5792) );
  OR2_X1 U6225 ( .A1(n9477), .A2(n9442), .ZN(n4638) );
  NAND2_X1 U6226 ( .A1(n8436), .A2(n5754), .ZN(n4909) );
  INV_X1 U6227 ( .A(n4909), .ZN(n4908) );
  OR2_X1 U6228 ( .A1(n10384), .A2(n5618), .ZN(n9900) );
  INV_X1 U6229 ( .A(n9900), .ZN(n4800) );
  NOR2_X1 U6230 ( .A1(n8698), .A2(n8699), .ZN(n4639) );
  AND2_X1 U6231 ( .A1(n4579), .A2(n8637), .ZN(n4640) );
  INV_X1 U6232 ( .A(n8995), .ZN(n5082) );
  NAND2_X1 U6233 ( .A1(n10289), .A2(n4843), .ZN(n4847) );
  AND2_X1 U6234 ( .A1(n8085), .A2(n8664), .ZN(n4641) );
  AND2_X1 U6235 ( .A1(n5042), .A2(n5041), .ZN(n4642) );
  AND2_X1 U6236 ( .A1(n4983), .A2(n4982), .ZN(n4643) );
  OR2_X1 U6237 ( .A1(n6435), .A2(n5158), .ZN(n4644) );
  NAND2_X1 U6238 ( .A1(n8495), .A2(n8642), .ZN(n4645) );
  INV_X1 U6239 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U6240 ( .A1(n5086), .A2(n8324), .ZN(n4646) );
  AND2_X1 U6241 ( .A1(n6106), .A2(n6105), .ZN(n4647) );
  AND2_X1 U6242 ( .A1(n4638), .A2(n4670), .ZN(n4648) );
  NAND2_X1 U6243 ( .A1(n5617), .A2(n4923), .ZN(n4922) );
  OR2_X1 U6244 ( .A1(n5288), .A2(SI_21_), .ZN(n4649) );
  INV_X1 U6245 ( .A(n8748), .ZN(n4659) );
  NAND2_X1 U6246 ( .A1(n6640), .A2(n6642), .ZN(n6647) );
  OAI21_X1 U6247 ( .B1(n6647), .B2(P2_D_REG_0__SCAN_IN), .A(n6646), .ZN(n6924)
         );
  INV_X2 U6248 ( .A(n10685), .ZN(n10683) );
  NAND2_X1 U6249 ( .A1(n6637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U6250 ( .A1(n7320), .A2(n7319), .ZN(n7422) );
  OR2_X1 U6251 ( .A1(n9802), .A2(n9938), .ZN(n9795) );
  INV_X1 U6252 ( .A(n5161), .ZN(n4917) );
  INV_X1 U6253 ( .A(n7726), .ZN(n5010) );
  AND2_X2 U6254 ( .A1(n7338), .A2(n6670), .ZN(n9456) );
  INV_X1 U6255 ( .A(n9456), .ZN(n4671) );
  AND2_X1 U6256 ( .A1(n6584), .A2(n6583), .ZN(n8990) );
  INV_X1 U6257 ( .A(n8990), .ZN(n9017) );
  AND2_X2 U6258 ( .A1(n7261), .A2(n10459), .ZN(n10643) );
  NAND2_X1 U6259 ( .A1(n5573), .A2(n5572), .ZN(n10503) );
  INV_X1 U6260 ( .A(n10503), .ZN(n4837) );
  NAND2_X1 U6261 ( .A1(n4619), .A2(n7090), .ZN(n7161) );
  AND2_X1 U6262 ( .A1(n4744), .A2(n6886), .ZN(n4650) );
  INV_X1 U6263 ( .A(n7697), .ZN(n6303) );
  AND2_X1 U6264 ( .A1(n6885), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U6265 ( .A1(n4762), .A2(n4761), .ZN(n5052) );
  INV_X1 U6266 ( .A(n4745), .ZN(n8686) );
  OR2_X1 U6267 ( .A1(n10657), .A2(n10693), .ZN(n4652) );
  AND2_X1 U6268 ( .A1(n7219), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4653) );
  NOR2_X1 U6269 ( .A1(n6852), .A2(n4986), .ZN(n4654) );
  NAND2_X1 U6270 ( .A1(n6577), .A2(n6582), .ZN(n8406) );
  NAND2_X1 U6271 ( .A1(n5046), .A2(n6789), .ZN(n4655) );
  NAND2_X1 U6272 ( .A1(n4691), .A2(n6274), .ZN(n6280) );
  INV_X1 U6273 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4896) );
  INV_X1 U6274 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4678) );
  INV_X1 U6275 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4700) );
  INV_X1 U6276 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n4748) );
  XNOR2_X1 U6277 ( .A(n7808), .B(n7825), .ZN(n7675) );
  INV_X1 U6278 ( .A(n7825), .ZN(n4663) );
  XNOR2_X1 U6279 ( .A(n8712), .B(n8713), .ZN(n7984) );
  XNOR2_X1 U6280 ( .A(n8697), .B(n8713), .ZN(n7987) );
  NAND2_X1 U6281 ( .A1(n4656), .A2(n9762), .ZN(n9765) );
  NAND3_X1 U6282 ( .A1(n9761), .A2(n9760), .A3(n9869), .ZN(n4656) );
  OAI21_X1 U6283 ( .B1(n9781), .B2(n9864), .A(n9857), .ZN(n9780) );
  NAND2_X1 U6284 ( .A1(n4796), .A2(n4955), .ZN(n4954) );
  MUX2_X1 U6285 ( .A(n9745), .B(n9744), .S(n9941), .Z(n9751) );
  NAND2_X1 U6286 ( .A1(n5384), .A2(n5228), .ZN(n5231) );
  OAI21_X1 U6287 ( .B1(n9799), .B2(n9798), .A(n9931), .ZN(n4798) );
  OAI21_X1 U6288 ( .B1(n9742), .B2(n4628), .A(n4802), .ZN(n4801) );
  NAND2_X1 U6289 ( .A1(n6604), .A2(n4588), .ZN(n7570) );
  AOI21_X2 U6290 ( .B1(n8995), .B2(n5080), .A(n5078), .ZN(n8960) );
  NAND2_X1 U6291 ( .A1(n6609), .A2(n6608), .ZN(n7946) );
  NAND2_X1 U6292 ( .A1(n8407), .A2(n6896), .ZN(n4875) );
  NAND2_X1 U6293 ( .A1(n6602), .A2(n5059), .ZN(n5064) );
  NAND2_X1 U6294 ( .A1(n4992), .A2(n4627), .ZN(n5000) );
  OAI21_X1 U6295 ( .B1(n5014), .B2(n5013), .A(n5012), .ZN(n8962) );
  AOI22_X1 U6296 ( .A1(n8862), .A2(n6561), .B1(n8651), .B2(n8552), .ZN(n6572)
         );
  INV_X1 U6297 ( .A(n6280), .ZN(n6288) );
  INV_X1 U6298 ( .A(n5003), .ZN(n7943) );
  AOI21_X2 U6299 ( .B1(n9489), .B2(n8919), .A(n6528), .ZN(n8895) );
  NAND2_X1 U6300 ( .A1(n6410), .A2(n6409), .ZN(n7720) );
  NAND2_X1 U6301 ( .A1(n7075), .A2(n7072), .ZN(n7071) );
  NAND2_X1 U6302 ( .A1(n7071), .A2(n6289), .ZN(n7058) );
  NAND2_X1 U6303 ( .A1(n7406), .A2(n6366), .ZN(n7455) );
  NAND2_X1 U6304 ( .A1(n6379), .A2(n4990), .ZN(n7480) );
  NAND2_X1 U6305 ( .A1(n6365), .A2(n6364), .ZN(n7406) );
  INV_X1 U6306 ( .A(n5225), .ZN(n4869) );
  AOI21_X1 U6307 ( .B1(n5602), .B2(n4947), .A(n4944), .ZN(n4943) );
  OAI21_X1 U6308 ( .B1(n4867), .B2(n4585), .A(n5227), .ZN(n5384) );
  INV_X1 U6309 ( .A(n5084), .ZN(n6580) );
  NAND2_X1 U6310 ( .A1(n7128), .A2(n6305), .ZN(n7065) );
  NAND2_X1 U6311 ( .A1(n7771), .A2(n4624), .ZN(n7845) );
  INV_X1 U6312 ( .A(n9812), .ZN(n5833) );
  NAND2_X1 U6313 ( .A1(n4675), .A2(n4672), .ZN(P1_U3519) );
  NAND2_X1 U6314 ( .A1(n5000), .A2(n4633), .ZN(n8906) );
  OAI21_X1 U6315 ( .B1(n6842), .B2(n7375), .A(n6785), .ZN(n10661) );
  NAND2_X1 U6316 ( .A1(n4755), .A2(n4626), .ZN(n5045) );
  NOR2_X2 U6317 ( .A1(n8771), .A2(n6495), .ZN(n8791) );
  NAND2_X1 U6318 ( .A1(n10660), .A2(n6786), .ZN(n6788) );
  AOI21_X2 U6319 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7472), .A(n7461), .ZN(
        n7612) );
  NOR2_X1 U6320 ( .A1(n8784), .A2(n8783), .ZN(n4662) );
  AND2_X1 U6321 ( .A1(n8784), .A2(n8783), .ZN(n8805) );
  INV_X1 U6322 ( .A(n7606), .ZN(n4734) );
  NAND2_X1 U6323 ( .A1(n8715), .A2(n4984), .ZN(n4980) );
  NOR2_X1 U6324 ( .A1(n7826), .A2(n7827), .ZN(n7831) );
  NAND3_X1 U6325 ( .A1(n9527), .A2(n6030), .A3(n5093), .ZN(n9662) );
  AOI21_X2 U6326 ( .B1(n5108), .B2(n5109), .A(n4816), .ZN(n4815) );
  OAI21_X2 U6327 ( .B1(n7034), .B2(n7036), .A(n7033), .ZN(n5904) );
  NAND2_X2 U6328 ( .A1(n7537), .A2(n5964), .ZN(n5971) );
  NAND2_X1 U6329 ( .A1(n9653), .A2(n5114), .ZN(n8474) );
  NAND2_X1 U6330 ( .A1(n5015), .A2(n5018), .ZN(n8989) );
  OAI21_X1 U6331 ( .B1(n6598), .B2(n8990), .A(n6597), .ZN(n8854) );
  NAND2_X4 U6332 ( .A1(n5870), .A2(n4558), .ZN(n6688) );
  NAND2_X1 U6333 ( .A1(n4822), .A2(n4821), .ZN(n9653) );
  INV_X1 U6334 ( .A(n8474), .ZN(n6146) );
  NAND2_X1 U6335 ( .A1(n6460), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U6336 ( .A1(n4807), .A2(n6275), .ZN(n4897) );
  NOR2_X2 U6337 ( .A1(n8854), .A2(n6624), .ZN(n9463) );
  AND3_X1 U6338 ( .A1(n6273), .A2(n6271), .A3(n6272), .ZN(n4691) );
  XNOR2_X2 U6339 ( .A(n6186), .B(n6185), .ZN(n6191) );
  INV_X1 U6340 ( .A(n4728), .ZN(n6297) );
  AND2_X2 U6341 ( .A1(n4727), .A2(n4728), .ZN(n5156) );
  NOR2_X1 U6342 ( .A1(n9794), .A2(n9793), .ZN(n4797) );
  NAND2_X1 U6343 ( .A1(n4954), .A2(n4953), .ZN(n9947) );
  NAND2_X1 U6344 ( .A1(n4957), .A2(n4956), .ZN(n5586) );
  OR2_X2 U6345 ( .A1(n10406), .A2(n5863), .ZN(n9847) );
  AND2_X1 U6346 ( .A1(n9776), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6347 ( .A1(n9922), .A2(n9942), .ZN(n4796) );
  NAND2_X1 U6348 ( .A1(n4785), .A2(n4784), .ZN(n9781) );
  INV_X1 U6349 ( .A(n5156), .ZN(n6352) );
  NAND2_X1 U6350 ( .A1(n8036), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U6351 ( .A1(n7736), .A2(n5980), .ZN(n5985) );
  NAND2_X1 U6352 ( .A1(n9595), .A2(n9596), .ZN(n9594) );
  OAI21_X1 U6353 ( .B1(n6023), .B2(n5092), .A(n5090), .ZN(n5089) );
  NAND2_X2 U6354 ( .A1(n6009), .A2(n10495), .ZN(n10499) );
  AOI21_X2 U6355 ( .B1(n5936), .B2(n7488), .A(n4593), .ZN(n5895) );
  OR2_X2 U6356 ( .A1(n5107), .A2(n5108), .ZN(n4814) );
  NAND2_X1 U6357 ( .A1(n10662), .A2(n10661), .ZN(n10660) );
  NAND2_X1 U6358 ( .A1(n5045), .A2(n5044), .ZN(n7674) );
  NAND2_X1 U6359 ( .A1(n5052), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U6360 ( .A1(n8690), .A2(n6875), .ZN(n4762) );
  NAND2_X1 U6361 ( .A1(n4760), .A2(n6790), .ZN(n6873) );
  INV_X1 U6362 ( .A(n8731), .ZN(n4757) );
  OAI22_X2 U6363 ( .A1(n4752), .A2(n4754), .B1(n7230), .B2(n7229), .ZN(n7461)
         );
  INV_X1 U6364 ( .A(n6788), .ZN(n5047) );
  INV_X1 U6365 ( .A(n7614), .ZN(n4755) );
  NAND2_X1 U6366 ( .A1(n8699), .A2(n5055), .ZN(n5053) );
  NAND2_X1 U6367 ( .A1(n4692), .A2(n4634), .ZN(n5014) );
  NAND2_X1 U6368 ( .A1(n8989), .A2(n8988), .ZN(n4692) );
  NAND2_X1 U6369 ( .A1(n6445), .A2(n6444), .ZN(n8036) );
  NAND2_X1 U6370 ( .A1(n7057), .A2(n6290), .ZN(n7130) );
  NAND2_X1 U6371 ( .A1(n8486), .A2(n8485), .ZN(n8488) );
  NAND2_X1 U6372 ( .A1(n5838), .A2(n9879), .ZN(n7529) );
  NAND2_X1 U6373 ( .A1(n7749), .A2(n9882), .ZN(n5840) );
  NAND2_X1 U6374 ( .A1(n7058), .A2(n8274), .ZN(n7057) );
  NAND2_X1 U6375 ( .A1(n4991), .A2(n7458), .ZN(n4990) );
  NAND2_X1 U6376 ( .A1(n6280), .A2(n7079), .ZN(n8259) );
  XNOR2_X1 U6377 ( .A(n8875), .B(n6620), .ZN(n4697) );
  NAND2_X1 U6378 ( .A1(n4697), .A2(n9017), .ZN(n4696) );
  INV_X1 U6379 ( .A(n4834), .ZN(n5378) );
  AND2_X2 U6380 ( .A1(n4569), .A2(n5178), .ZN(n4834) );
  NAND2_X1 U6381 ( .A1(n7137), .A2(n5915), .ZN(n9547) );
  NAND4_X1 U6382 ( .A1(n5904), .A2(n5914), .A3(n5915), .A4(n5903), .ZN(n7137)
         );
  OAI21_X2 U6383 ( .B1(n10499), .B2(n4829), .A(n4827), .ZN(n6023) );
  NAND2_X2 U6384 ( .A1(n9594), .A2(n6048), .ZN(n9646) );
  NAND2_X1 U6385 ( .A1(n5362), .A2(n5352), .ZN(n5621) );
  AOI21_X2 U6386 ( .B1(n5096), .B2(n4562), .A(n4616), .ZN(n6083) );
  NAND2_X1 U6387 ( .A1(n4817), .A2(n4815), .ZN(n4822) );
  AOI21_X1 U6388 ( .B1(n8655), .B2(n8594), .A(n8906), .ZN(n6528) );
  NAND2_X1 U6389 ( .A1(n6339), .A2(n6338), .ZN(n7207) );
  NOR2_X1 U6390 ( .A1(n9037), .A2(n4625), .ZN(n9475) );
  AOI21_X1 U6391 ( .B1(n7720), .B2(n5006), .A(n5004), .ZN(n5003) );
  OAI21_X1 U6392 ( .B1(n8885), .B2(n5033), .A(n4587), .ZN(n5028) );
  INV_X1 U6393 ( .A(n5028), .ZN(n8875) );
  NOR2_X1 U6394 ( .A1(n8400), .A2(n4878), .ZN(n4877) );
  NOR2_X1 U6395 ( .A1(n8385), .A2(n4883), .ZN(n4882) );
  XNOR2_X1 U6396 ( .A(n4874), .B(n6622), .ZN(n8414) );
  AOI21_X1 U6397 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8405) );
  NOR2_X2 U6398 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6260) );
  INV_X1 U6399 ( .A(n4701), .ZN(n6243) );
  OAI21_X1 U6400 ( .B1(n8589), .B2(n4713), .A(n4710), .ZN(n8548) );
  NAND2_X1 U6401 ( .A1(n8589), .A2(n5138), .ZN(n4716) );
  INV_X1 U6402 ( .A(n8615), .ZN(n4721) );
  NAND2_X1 U6403 ( .A1(n7275), .A2(n7274), .ZN(n7277) );
  NAND3_X1 U6404 ( .A1(n7161), .A2(n7166), .A3(n7160), .ZN(n7275) );
  NAND4_X1 U6405 ( .A1(n6316), .A2(n6327), .A3(n6172), .A4(n6171), .ZN(n4724)
         );
  INV_X1 U6406 ( .A(n4731), .ZN(n8749) );
  NAND2_X1 U6407 ( .A1(n4730), .A2(n4729), .ZN(n8782) );
  INV_X1 U6408 ( .A(n4737), .ZN(n8815) );
  OR2_X1 U6409 ( .A1(n8804), .A2(n8805), .ZN(n4737) );
  NOR2_X1 U6410 ( .A1(n8785), .A2(n9440), .ZN(n8804) );
  INV_X1 U6411 ( .A(n6801), .ZN(n4738) );
  NAND2_X1 U6412 ( .A1(n6887), .A2(n6886), .ZN(n4740) );
  NAND2_X1 U6413 ( .A1(n6885), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U6414 ( .A1(n6884), .A2(n6885), .ZN(n8688) );
  OR2_X1 U6415 ( .A1(n7148), .A2(n7213), .ZN(n4746) );
  NAND3_X1 U6416 ( .A1(n4978), .A2(n7219), .A3(n4977), .ZN(n4749) );
  NAND2_X1 U6417 ( .A1(n4985), .A2(n6795), .ZN(n6796) );
  NOR2_X1 U6418 ( .A1(n5050), .A2(n5049), .ZN(n4754) );
  NAND2_X1 U6419 ( .A1(n4759), .A2(n6789), .ZN(n4760) );
  NAND3_X1 U6420 ( .A1(n4766), .A2(n4765), .A3(n4763), .ZN(P2_U3200) );
  OAI21_X1 U6421 ( .B1(n8811), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8807), .ZN(
        n4764) );
  OAI21_X1 U6422 ( .B1(n4594), .B2(n4767), .A(n8828), .ZN(n4766) );
  OAI21_X1 U6423 ( .B1(n8813), .B2(n8814), .A(n8812), .ZN(n4767) );
  NAND2_X1 U6424 ( .A1(n8154), .A2(n4768), .ZN(n4895) );
  NAND2_X1 U6425 ( .A1(n4773), .A2(n4603), .ZN(n9769) );
  NAND2_X1 U6426 ( .A1(n4774), .A2(n4775), .ZN(n9740) );
  NAND2_X1 U6427 ( .A1(n9735), .A2(n4776), .ZN(n4774) );
  INV_X1 U6428 ( .A(n9893), .ZN(n4782) );
  NAND2_X1 U6429 ( .A1(n4974), .A2(n4786), .ZN(n4785) );
  AOI21_X1 U6430 ( .B1(n4794), .B2(n9774), .A(n4568), .ZN(n4791) );
  NOR2_X2 U6431 ( .A1(n4798), .A2(n4797), .ZN(n9922) );
  NAND2_X1 U6432 ( .A1(n4809), .A2(n5986), .ZN(n10481) );
  NAND2_X1 U6433 ( .A1(n5116), .A2(n4809), .ZN(n5999) );
  NAND2_X1 U6434 ( .A1(n5115), .A2(n4809), .ZN(n10480) );
  INV_X1 U6435 ( .A(n5984), .ZN(n4810) );
  INV_X1 U6436 ( .A(n5985), .ZN(n4811) );
  NAND2_X1 U6437 ( .A1(n4814), .A2(n5109), .ZN(n9578) );
  NAND2_X1 U6438 ( .A1(n5107), .A2(n5109), .ZN(n4817) );
  NAND2_X1 U6439 ( .A1(n6101), .A2(n6100), .ZN(n4823) );
  NAND2_X1 U6440 ( .A1(n10499), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U6441 ( .A1(n5914), .A2(n5915), .ZN(n7135) );
  NAND2_X1 U6442 ( .A1(n5904), .A2(n5903), .ZN(n7136) );
  XNOR2_X2 U6443 ( .A(n5329), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5872) );
  AND3_X2 U6444 ( .A1(n4834), .A2(n5183), .A3(n4833), .ZN(n5786) );
  NAND2_X1 U6445 ( .A1(n4836), .A2(n7503), .ZN(n7200) );
  INV_X1 U6446 ( .A(n4841), .ZN(n7800) );
  INV_X1 U6447 ( .A(n4847), .ZN(n10231) );
  NAND2_X1 U6448 ( .A1(n10137), .A2(n4566), .ZN(n10109) );
  NAND2_X1 U6449 ( .A1(n10137), .A2(n8436), .ZN(n10121) );
  AND2_X1 U6450 ( .A1(n10137), .A2(n4849), .ZN(n10120) );
  OAI21_X2 U6451 ( .B1(n7529), .B2(n9815), .A(n9884), .ZN(n7749) );
  NAND2_X1 U6452 ( .A1(n5786), .A2(n4635), .ZN(n5193) );
  NAND2_X1 U6453 ( .A1(n5786), .A2(n4572), .ZN(n5323) );
  AOI21_X2 U6454 ( .B1(n5877), .B2(n10285), .A(n5876), .ZN(n8486) );
  NAND3_X1 U6455 ( .A1(n8327), .A2(n4863), .A3(n8339), .ZN(n4861) );
  NAND2_X1 U6456 ( .A1(n4861), .A2(n4636), .ZN(n8343) );
  INV_X1 U6457 ( .A(n8338), .ZN(n4866) );
  OAI21_X1 U6458 ( .B1(n5453), .B2(n4869), .A(n4868), .ZN(n4867) );
  AND2_X1 U6459 ( .A1(n5474), .A2(n5225), .ZN(n4870) );
  AND2_X2 U6460 ( .A1(n8387), .A2(n8386), .ZN(n8391) );
  NAND3_X1 U6461 ( .A1(n8381), .A2(n8380), .A3(n8877), .ZN(n4884) );
  NAND2_X1 U6462 ( .A1(n4895), .A2(n10100), .ZN(n4894) );
  NAND3_X1 U6463 ( .A1(n4891), .A2(n4890), .A3(n4889), .ZN(n5208) );
  NAND3_X1 U6464 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n4892), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4889) );
  NAND3_X1 U6465 ( .A1(n4895), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n10100), .ZN(
        n4890) );
  NAND3_X1 U6466 ( .A1(n4894), .A2(n4893), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4891) );
  AND2_X2 U6467 ( .A1(n4894), .A2(n4893), .ZN(n5204) );
  INV_X1 U6468 ( .A(n5420), .ZN(n4899) );
  OAI21_X2 U6469 ( .B1(n5783), .B2(n4615), .A(n4900), .ZN(n5328) );
  NAND3_X1 U6470 ( .A1(n10323), .A2(n10622), .A3(n10324), .ZN(n10329) );
  INV_X1 U6471 ( .A(n5617), .ZN(n4919) );
  NAND2_X1 U6472 ( .A1(n5617), .A2(n5616), .ZN(n10288) );
  INV_X1 U6473 ( .A(n4922), .ZN(n10388) );
  INV_X1 U6474 ( .A(n5616), .ZN(n4924) );
  NAND2_X1 U6475 ( .A1(n10187), .A2(n4930), .ZN(n4926) );
  NAND2_X1 U6476 ( .A1(n4926), .A2(n4927), .ZN(n10129) );
  NAND2_X2 U6477 ( .A1(n6688), .A2(n8171), .ZN(n5420) );
  NAND2_X1 U6478 ( .A1(n5243), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U6479 ( .A1(n5231), .A2(n4586), .ZN(n5517) );
  OAI21_X2 U6480 ( .B1(n5231), .B2(n4564), .A(n4966), .ZN(n5534) );
  OAI21_X1 U6481 ( .B1(n5336), .B2(n5333), .A(n5286), .ZN(n4970) );
  NAND2_X1 U6482 ( .A1(n5287), .A2(n4969), .ZN(n4973) );
  NAND2_X1 U6483 ( .A1(n4978), .A2(n7219), .ZN(n7144) );
  NAND2_X1 U6484 ( .A1(n4979), .A2(n7151), .ZN(n4978) );
  INV_X1 U6485 ( .A(n7143), .ZN(n4979) );
  OAI21_X1 U6486 ( .B1(n4981), .B2(n7984), .A(n4980), .ZN(n8723) );
  NAND2_X1 U6487 ( .A1(n4985), .A2(n6783), .ZN(n6784) );
  XNOR2_X1 U6488 ( .A(n6769), .B(n4985), .ZN(n6849) );
  AOI21_X1 U6489 ( .B1(n10650), .B2(n4985), .A(n6853), .ZN(n4987) );
  NAND2_X1 U6490 ( .A1(n5440), .A2(n5216), .ZN(n4988) );
  NAND2_X1 U6491 ( .A1(n4989), .A2(n5213), .ZN(n5440) );
  NAND2_X1 U6492 ( .A1(n5422), .A2(n5421), .ZN(n4989) );
  NAND2_X1 U6493 ( .A1(n7406), .A2(n4630), .ZN(n4991) );
  NAND2_X1 U6494 ( .A1(n7480), .A2(n6395), .ZN(n6397) );
  OR2_X1 U6495 ( .A1(n9062), .A2(n8659), .ZN(n5002) );
  NOR2_X1 U6496 ( .A1(n5017), .A2(n9010), .ZN(n5016) );
  NAND2_X1 U6497 ( .A1(n8895), .A2(n5027), .ZN(n5026) );
  INV_X2 U6498 ( .A(n5204), .ZN(n8171) );
  NOR2_X2 U6499 ( .A1(n7462), .A2(n6390), .ZN(n7614) );
  NAND2_X1 U6500 ( .A1(n5047), .A2(n6827), .ZN(n5046) );
  NOR2_X1 U6501 ( .A1(n8770), .A2(n8797), .ZN(n8792) );
  AND2_X1 U6502 ( .A1(n8770), .A2(n8797), .ZN(n5048) );
  NAND2_X1 U6503 ( .A1(n5058), .A2(n8189), .ZN(n6601) );
  XNOR2_X1 U6504 ( .A(n5058), .B(n7129), .ZN(n7703) );
  NAND2_X1 U6505 ( .A1(n6600), .A2(n8267), .ZN(n5058) );
  NOR2_X1 U6506 ( .A1(n5061), .A2(n5060), .ZN(n5059) );
  NAND2_X1 U6507 ( .A1(n5064), .A2(n5062), .ZN(n7405) );
  NAND2_X1 U6508 ( .A1(n8912), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U6509 ( .A1(n5066), .A2(n5071), .ZN(n8869) );
  NAND2_X1 U6510 ( .A1(n8912), .A2(n5076), .ZN(n5074) );
  NAND2_X1 U6511 ( .A1(n5084), .A2(n4567), .ZN(n6201) );
  NAND2_X1 U6512 ( .A1(n6611), .A2(n5087), .ZN(n5086) );
  OAI21_X2 U6513 ( .B1(n7457), .B2(n8243), .A(n8250), .ZN(n7479) );
  INV_X1 U6514 ( .A(n5089), .ZN(n9663) );
  OR2_X2 U6515 ( .A1(n6023), .A2(n6024), .ZN(n9527) );
  AOI21_X2 U6516 ( .B1(n9646), .B2(n5101), .A(n5097), .ZN(n5096) );
  NAND2_X1 U6517 ( .A1(n9630), .A2(n5113), .ZN(n5107) );
  INV_X1 U6518 ( .A(n5111), .ZN(n9538) );
  NAND2_X1 U6519 ( .A1(n9630), .A2(n9631), .ZN(n9537) );
  INV_X1 U6520 ( .A(n9539), .ZN(n5112) );
  NAND2_X1 U6521 ( .A1(n5986), .A2(n5989), .ZN(n5116) );
  NAND2_X1 U6522 ( .A1(n5120), .A2(n5119), .ZN(n10462) );
  INV_X1 U6523 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6524 ( .A1(n7422), .A2(n4577), .ZN(n7560) );
  NAND3_X1 U6525 ( .A1(n5156), .A2(n5155), .A3(n6573), .ZN(n6577) );
  NAND3_X1 U6526 ( .A1(n6926), .A2(n6928), .A3(n6927), .ZN(n7097) );
  NAND2_X1 U6527 ( .A1(n5833), .A2(n7487), .ZN(n7486) );
  OR2_X1 U6528 ( .A1(n4556), .A2(n6254), .ZN(n6258) );
  NAND4_X1 U6529 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n8677)
         );
  XNOR2_X1 U6530 ( .A(n6632), .B(n6635), .ZN(n6641) );
  INV_X1 U6531 ( .A(n10563), .ZN(n10241) );
  NAND2_X1 U6532 ( .A1(n7862), .A2(n5824), .ZN(n10560) );
  AND2_X2 U6533 ( .A1(n7261), .A2(n7260), .ZN(n10449) );
  OR2_X1 U6534 ( .A1(n10310), .A2(n5849), .ZN(n5157) );
  NAND3_X1 U6535 ( .A1(n6461), .A2(n6446), .A3(n6234), .ZN(n5158) );
  OR2_X1 U6536 ( .A1(n10225), .A2(n5856), .ZN(n5159) );
  NOR2_X1 U6537 ( .A1(n5584), .A2(n8448), .ZN(n5161) );
  INV_X1 U6538 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5215) );
  INV_X1 U6539 ( .A(n9807), .ZN(n5820) );
  INV_X1 U6540 ( .A(n9667), .ZN(n7846) );
  AND2_X1 U6541 ( .A1(n9033), .A2(n9449), .ZN(n5163) );
  INV_X1 U6542 ( .A(n6727), .ZN(n5400) );
  INV_X1 U6543 ( .A(n6622), .ZN(n6898) );
  INV_X1 U6544 ( .A(n8822), .ZN(n6767) );
  INV_X1 U6545 ( .A(n10178), .ZN(n10193) );
  INV_X1 U6546 ( .A(n6927), .ZN(n7100) );
  AND2_X1 U6547 ( .A1(n9468), .A2(n9028), .ZN(n5164) );
  INV_X1 U6548 ( .A(n8298), .ZN(n6364) );
  OR2_X1 U6549 ( .A1(n7950), .A2(n9979), .ZN(n5165) );
  INV_X1 U6550 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5174) );
  INV_X1 U6551 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6172) );
  INV_X1 U6552 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5187) );
  NOR2_X1 U6553 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5185) );
  INV_X1 U6554 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5179) );
  INV_X1 U6555 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7821) );
  NOR2_X1 U6556 ( .A1(n8186), .A2(n8848), .ZN(n6595) );
  AND2_X1 U6557 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  INV_X1 U6558 ( .A(SI_26_), .ZN(n5310) );
  INV_X1 U6559 ( .A(SI_23_), .ZN(n5295) );
  INV_X1 U6560 ( .A(SI_19_), .ZN(n5281) );
  INV_X1 U6561 ( .A(SI_16_), .ZN(n9273) );
  NOR2_X1 U6562 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5177) );
  INV_X1 U6563 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6162) );
  INV_X1 U6564 ( .A(n8641), .ZN(n8624) );
  XNOR2_X1 U6565 ( .A(n6203), .B(n6202), .ZN(n6585) );
  NOR2_X1 U6566 ( .A1(n8887), .A2(n8993), .ZN(n8864) );
  NOR2_X1 U6567 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  AND2_X1 U6568 ( .A1(n6922), .A2(n8392), .ZN(n6904) );
  NAND2_X1 U6569 ( .A1(n6631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6632) );
  INV_X1 U6570 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6446) );
  INV_X1 U6571 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5365) );
  INV_X1 U6573 ( .A(n9960), .ZN(n5754) );
  AND2_X1 U6574 ( .A1(n9802), .A2(n5820), .ZN(n9932) );
  NAND2_X1 U6575 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6576 ( .A1(n10178), .A2(n10346), .ZN(n10180) );
  NAND2_X1 U6577 ( .A1(n8076), .A2(n5848), .ZN(n5600) );
  INV_X1 U6578 ( .A(n10625), .ZN(n5828) );
  AND2_X1 U6579 ( .A1(n9891), .A2(n9736), .ZN(n9820) );
  INV_X1 U6580 ( .A(n7203), .ZN(n7196) );
  INV_X1 U6581 ( .A(n5738), .ZN(n5317) );
  INV_X1 U6582 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5355) );
  OAI21_X1 U6583 ( .B1(n7162), .B2(n7344), .A(n8261), .ZN(n6927) );
  NAND2_X1 U6584 ( .A1(n7050), .A2(n6920), .ZN(n8641) );
  AND2_X1 U6585 ( .A1(n6781), .A2(n6780), .ZN(n8837) );
  INV_X1 U6586 ( .A(n6585), .ZN(n8822) );
  INV_X1 U6587 ( .A(n8652), .ZN(n8887) );
  INV_X1 U6588 ( .A(n8977), .ZN(n8951) );
  INV_X1 U6589 ( .A(n8660), .ZN(n8994) );
  OR2_X1 U6590 ( .A1(n6901), .A2(n9454), .ZN(n6913) );
  OR2_X1 U6591 ( .A1(n6904), .A2(n6667), .ZN(n7340) );
  OR2_X1 U6592 ( .A1(n6649), .A2(n6899), .ZN(n6651) );
  INV_X1 U6593 ( .A(n8666), .ZN(n7960) );
  NOR2_X1 U6594 ( .A1(n6645), .A2(n8102), .ZN(n6663) );
  XNOR2_X1 U6595 ( .A(n6665), .B(n6666), .ZN(n6814) );
  INV_X1 U6596 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U6597 ( .A1(n6132), .A2(n9949), .ZN(n10492) );
  INV_X1 U6598 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10015) );
  INV_X1 U6599 ( .A(n7124), .ZN(n7252) );
  INV_X1 U6600 ( .A(n10563), .ZN(n5878) );
  AND2_X1 U6601 ( .A1(n9779), .A2(n9778), .ZN(n10116) );
  NOR2_X1 U6602 ( .A1(n7780), .A2(n10607), .ZN(n7856) );
  AOI21_X1 U6603 ( .B1(n6747), .B2(n5818), .A(n6749), .ZN(n6856) );
  OR2_X1 U6604 ( .A1(n5420), .A2(n8098), .ZN(n5722) );
  OR2_X1 U6605 ( .A1(n10443), .A2(n5852), .ZN(n10245) );
  NOR2_X1 U6606 ( .A1(n10309), .A2(n10454), .ZN(n10307) );
  INV_X1 U6607 ( .A(n9820), .ZN(n7798) );
  NAND2_X1 U6608 ( .A1(n6122), .A2(n6121), .ZN(n10617) );
  NAND2_X1 U6609 ( .A1(n9703), .A2(n9809), .ZN(n7203) );
  INV_X1 U6610 ( .A(n10285), .ZN(n10302) );
  INV_X1 U6611 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5790) );
  OR2_X1 U6612 ( .A1(n5569), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5590) );
  INV_X1 U6613 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10461) );
  AOI21_X1 U6614 ( .B1(n7961), .B2(n7960), .A(n7959), .ZN(n7962) );
  NAND2_X1 U6615 ( .A1(n7084), .A2(n8413), .ZN(n8645) );
  AOI21_X1 U6616 ( .B1(n8954), .B2(n6565), .A(n6220), .ZN(n8964) );
  INV_X1 U6617 ( .A(n8837), .ZN(n10650) );
  INV_X1 U6618 ( .A(n10657), .ZN(n8839) );
  INV_X1 U6619 ( .A(n8953), .ZN(n9014) );
  INV_X1 U6620 ( .A(n9022), .ZN(n9020) );
  INV_X1 U6621 ( .A(n8194), .ZN(n7266) );
  NOR2_X1 U6622 ( .A1(n9456), .A2(n6671), .ZN(n6672) );
  NOR2_X1 U6623 ( .A1(n4671), .A2(n9454), .ZN(n9028) );
  NOR2_X1 U6624 ( .A1(n7340), .A2(n6669), .ZN(n6670) );
  NAND2_X1 U6625 ( .A1(n10685), .A2(n9464), .ZN(n9465) );
  INV_X1 U6626 ( .A(n9443), .ZN(n9454) );
  AND2_X1 U6627 ( .A1(n7932), .A2(n8262), .ZN(n9443) );
  INV_X1 U6628 ( .A(n6647), .ZN(n6755) );
  INV_X1 U6629 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6262) );
  OAI21_X1 U6630 ( .B1(n6131), .B2(n6130), .A(n10270), .ZN(n10502) );
  INV_X1 U6631 ( .A(n10090), .ZN(n10087) );
  INV_X1 U6632 ( .A(n10093), .ZN(n10037) );
  AND2_X1 U6633 ( .A1(n6691), .A2(n6689), .ZN(n6944) );
  INV_X1 U6634 ( .A(n10089), .ZN(n10072) );
  INV_X1 U6635 ( .A(n10270), .ZN(n10551) );
  OR2_X1 U6636 ( .A1(n10458), .A2(n6854), .ZN(n10270) );
  AND2_X1 U6637 ( .A1(n10643), .A2(n10626), .ZN(n10392) );
  INV_X1 U6638 ( .A(n9838), .ZN(n5775) );
  OR2_X1 U6639 ( .A1(n7796), .A2(n10478), .ZN(n7837) );
  NAND2_X1 U6640 ( .A1(n7776), .A2(n10629), .ZN(n10622) );
  AND2_X1 U6641 ( .A1(n7937), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6674) );
  AND2_X1 U6642 ( .A1(n8099), .A2(n8035), .ZN(n5816) );
  AND2_X1 U6643 ( .A1(n5571), .A2(n5590), .ZN(n7709) );
  INV_X1 U6644 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5471) );
  AND2_X1 U6645 ( .A1(n5204), .A2(P1_U3086), .ZN(n7936) );
  INV_X1 U6646 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8129) );
  NOR2_X1 U6647 ( .A1(n8137), .A2(n10727), .ZN(n8138) );
  INV_X1 U6648 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10710) );
  INV_X1 U6649 ( .A(n8645), .ZN(n8524) );
  AND2_X1 U6650 ( .A1(n6935), .A2(n6934), .ZN(n8632) );
  NAND2_X1 U6651 ( .A1(n6552), .A2(n6551), .ZN(n8652) );
  INV_X1 U6652 ( .A(n8975), .ZN(n9015) );
  INV_X1 U6653 ( .A(n8247), .ZN(n8669) );
  NAND2_X1 U6654 ( .A1(n6833), .A2(n6806), .ZN(n8806) );
  OR2_X1 U6655 ( .A1(P2_U3150), .A2(n6766), .ZN(n10657) );
  INV_X1 U6656 ( .A(n9020), .ZN(n9000) );
  AND2_X1 U6657 ( .A1(n7343), .A2(n9018), .ZN(n9022) );
  INV_X1 U6658 ( .A(n9004), .ZN(n9026) );
  NOR2_X1 U6659 ( .A1(n5164), .A2(n6672), .ZN(n6673) );
  INV_X1 U6660 ( .A(n9028), .ZN(n9442) );
  INV_X1 U6661 ( .A(n8552), .ZN(n9474) );
  INV_X1 U6662 ( .A(n9467), .ZN(n9514) );
  AND2_X1 U6663 ( .A1(n7052), .A2(n7051), .ZN(n10685) );
  NOR2_X1 U6664 ( .A1(n6912), .A2(n6755), .ZN(n7010) );
  INV_X1 U6665 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U6666 ( .A1(n6146), .A2(n6129), .ZN(n6144) );
  INV_X1 U6667 ( .A(n10443), .ZN(n10274) );
  INV_X1 U6668 ( .A(n8456), .ZN(n9629) );
  INV_X1 U6669 ( .A(n10502), .ZN(n10543) );
  NAND2_X1 U6670 ( .A1(n5202), .A2(n5201), .ZN(n9959) );
  NAND2_X1 U6671 ( .A1(n6944), .A2(n4558), .ZN(n10090) );
  INV_X1 U6672 ( .A(n10278), .ZN(n10556) );
  AND2_X1 U6673 ( .A1(n10267), .A2(n10266), .ZN(n10378) );
  INV_X1 U6674 ( .A(n10241), .ZN(n10553) );
  OR2_X1 U6675 ( .A1(n10553), .A2(n5883), .ZN(n7862) );
  INV_X1 U6676 ( .A(n10560), .ZN(n10259) );
  AND2_X1 U6677 ( .A1(n5830), .A2(n10270), .ZN(n10563) );
  NAND2_X1 U6678 ( .A1(n10643), .A2(n10622), .ZN(n10381) );
  INV_X1 U6679 ( .A(n10643), .ZN(n10641) );
  INV_X1 U6680 ( .A(n10453), .ZN(n10425) );
  NAND2_X1 U6681 ( .A1(n10449), .A2(n10622), .ZN(n10447) );
  AND2_X1 U6682 ( .A1(n10614), .A2(n10613), .ZN(n10639) );
  INV_X1 U6683 ( .A(n10449), .ZN(n10634) );
  AOI21_X1 U6684 ( .B1(n6747), .B2(n5817), .A(n5816), .ZN(n10459) );
  INV_X1 U6685 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8098) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7790) );
  INV_X1 U6687 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7305) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9293) );
  INV_X2 U6689 ( .A(n7936), .ZN(n10472) );
  INV_X1 U6690 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10729) );
  INV_X1 U6691 ( .A(n8676), .ZN(P2_U3893) );
  INV_X1 U6692 ( .A(n9985), .ZN(P1_U3973) );
  NAND2_X1 U6693 ( .A1(n5478), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5493) );
  INV_X1 U6694 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6695 ( .A1(n5494), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6696 ( .A1(n5559), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5575) );
  INV_X1 U6697 ( .A(n5594), .ZN(n5166) );
  NAND2_X1 U6698 ( .A1(n5166), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5609) );
  INV_X1 U6699 ( .A(n5609), .ZN(n5167) );
  NAND2_X1 U6700 ( .A1(n5167), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5611) );
  INV_X1 U6701 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9613) );
  INV_X1 U6702 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5670) );
  INV_X1 U6703 ( .A(n5683), .ZN(n5171) );
  INV_X1 U6704 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5711) );
  INV_X1 U6705 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5710) );
  OR3_X2 U6706 ( .A1(n5712), .A2(n5711), .A3(n5710), .ZN(n5724) );
  INV_X1 U6707 ( .A(n5724), .ZN(n5172) );
  NAND2_X1 U6708 ( .A1(n5172), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5745) );
  INV_X1 U6709 ( .A(n5745), .ZN(n5173) );
  NAND2_X1 U6710 ( .A1(n5173), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5827) );
  XNOR2_X1 U6711 ( .A(n5827), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U6712 ( .A1(n5419), .A2(n5177), .ZN(n5385) );
  INV_X1 U6713 ( .A(n5385), .ZN(n5178) );
  NOR2_X1 U6714 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5182) );
  NOR2_X1 U6715 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5181) );
  NOR2_X1 U6716 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5180) );
  INV_X1 U6717 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6718 ( .A1(n5778), .A2(n5187), .ZN(n5324) );
  INV_X1 U6719 ( .A(n5324), .ZN(n5189) );
  NOR2_X1 U6720 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5188) );
  XNOR2_X2 U6721 ( .A(n5194), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6722 ( .A1(n10122), .A2(n5714), .ZN(n5202) );
  INV_X1 U6723 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5199) );
  NAND2_X2 U6724 ( .A1(n5195), .A2(n10473), .ZN(n5458) );
  AND2_X4 U6725 ( .A1(n10467), .A2(n5196), .ZN(n5695) );
  NAND2_X1 U6726 ( .A1(n5695), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6727 ( .A1(n5747), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5197) );
  OAI211_X1 U6728 ( .C1(n5199), .C2(n5458), .A(n5198), .B(n5197), .ZN(n5200)
         );
  INV_X1 U6729 ( .A(n5200), .ZN(n5201) );
  INV_X1 U6730 ( .A(n5397), .ZN(n5207) );
  AND2_X1 U6731 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6732 ( .A1(n5204), .A2(n5205), .ZN(n5411) );
  NAND3_X1 U6733 ( .A1(n8171), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5206) );
  NAND2_X1 U6734 ( .A1(n5411), .A2(n5206), .ZN(n5396) );
  NAND2_X1 U6735 ( .A1(n5207), .A2(n5396), .ZN(n5210) );
  NAND2_X1 U6736 ( .A1(n5208), .A2(SI_1_), .ZN(n5209) );
  NAND2_X1 U6737 ( .A1(n5210), .A2(n5209), .ZN(n5422) );
  INV_X1 U6738 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6718) );
  INV_X1 U6739 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6719) );
  MUX2_X1 U6740 ( .A(n6718), .B(n6719), .S(n5204), .Z(n5211) );
  XNOR2_X1 U6741 ( .A(n5211), .B(SI_2_), .ZN(n5421) );
  INV_X1 U6742 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6743 ( .A1(n5212), .A2(SI_2_), .ZN(n5213) );
  BUF_X8 U6744 ( .A(n5204), .Z(n5330) );
  XNOR2_X1 U6745 ( .A(n5217), .B(SI_3_), .ZN(n5439) );
  INV_X1 U6746 ( .A(n5439), .ZN(n5216) );
  NAND2_X1 U6747 ( .A1(n5217), .A2(SI_3_), .ZN(n5218) );
  XNOR2_X1 U6748 ( .A(n5220), .B(SI_4_), .ZN(n5452) );
  INV_X1 U6749 ( .A(n5452), .ZN(n5219) );
  NAND2_X1 U6750 ( .A1(n5220), .A2(SI_4_), .ZN(n5473) );
  NAND2_X1 U6751 ( .A1(n5222), .A2(SI_5_), .ZN(n5221) );
  AND2_X1 U6752 ( .A1(n5473), .A2(n5221), .ZN(n5225) );
  INV_X1 U6753 ( .A(n5221), .ZN(n5224) );
  XNOR2_X1 U6754 ( .A(n5222), .B(SI_5_), .ZN(n5475) );
  INV_X1 U6755 ( .A(n5475), .ZN(n5223) );
  MUX2_X1 U6756 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5330), .Z(n5226) );
  NAND2_X1 U6757 ( .A1(n5226), .A2(SI_6_), .ZN(n5227) );
  MUX2_X1 U6758 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5330), .Z(n5229) );
  XNOR2_X1 U6759 ( .A(n5229), .B(SI_7_), .ZN(n5383) );
  INV_X1 U6760 ( .A(n5383), .ZN(n5228) );
  NAND2_X1 U6761 ( .A1(n5229), .A2(SI_7_), .ZN(n5230) );
  INV_X1 U6762 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6745) );
  INV_X1 U6763 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5232) );
  MUX2_X1 U6764 ( .A(n6745), .B(n5232), .S(n5330), .Z(n5233) );
  INV_X1 U6765 ( .A(SI_8_), .ZN(n9422) );
  NAND2_X1 U6766 ( .A1(n5233), .A2(n9422), .ZN(n5516) );
  INV_X1 U6767 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6768 ( .A1(n5234), .A2(SI_8_), .ZN(n5235) );
  NAND2_X1 U6769 ( .A1(n5516), .A2(n5235), .ZN(n5501) );
  INV_X1 U6770 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6752) );
  MUX2_X1 U6771 ( .A(n9151), .B(n6752), .S(n5330), .Z(n5237) );
  INV_X1 U6772 ( .A(SI_9_), .ZN(n5236) );
  NAND2_X1 U6773 ( .A1(n5237), .A2(n5236), .ZN(n5519) );
  INV_X1 U6774 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6775 ( .A1(n5238), .A2(SI_9_), .ZN(n5518) );
  INV_X1 U6776 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5239) );
  MUX2_X1 U6777 ( .A(n9274), .B(n5239), .S(n5330), .Z(n5240) );
  XNOR2_X1 U6778 ( .A(n5240), .B(SI_10_), .ZN(n5535) );
  INV_X1 U6779 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6780 ( .A1(n5241), .A2(SI_10_), .ZN(n5242) );
  INV_X1 U6781 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5244) );
  MUX2_X1 U6782 ( .A(n5244), .B(n9293), .S(n5330), .Z(n5246) );
  INV_X1 U6783 ( .A(SI_11_), .ZN(n5245) );
  NAND2_X1 U6784 ( .A1(n5246), .A2(n5245), .ZN(n5249) );
  INV_X1 U6785 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6786 ( .A1(n5247), .A2(SI_11_), .ZN(n5248) );
  NAND2_X1 U6787 ( .A1(n5249), .A2(n5248), .ZN(n5553) );
  MUX2_X1 U6788 ( .A(n6893), .B(n9295), .S(n5330), .Z(n5250) );
  XNOR2_X1 U6789 ( .A(n5250), .B(SI_12_), .ZN(n5567) );
  INV_X1 U6790 ( .A(n5567), .ZN(n5252) );
  INV_X1 U6791 ( .A(n5250), .ZN(n5251) );
  MUX2_X1 U6792 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5330), .Z(n5253) );
  XNOR2_X1 U6793 ( .A(n5253), .B(SI_13_), .ZN(n5376) );
  NAND2_X1 U6794 ( .A1(n5253), .A2(SI_13_), .ZN(n5587) );
  MUX2_X1 U6795 ( .A(n7181), .B(n7180), .S(n5330), .Z(n5255) );
  INV_X1 U6796 ( .A(SI_14_), .ZN(n5254) );
  NAND2_X1 U6797 ( .A1(n5255), .A2(n5254), .ZN(n5260) );
  INV_X1 U6798 ( .A(n5255), .ZN(n5256) );
  NAND2_X1 U6799 ( .A1(n5256), .A2(SI_14_), .ZN(n5257) );
  NAND2_X1 U6800 ( .A1(n5260), .A2(n5257), .ZN(n5588) );
  INV_X1 U6801 ( .A(n5588), .ZN(n5258) );
  NAND2_X1 U6802 ( .A1(n5586), .A2(n5259), .ZN(n5261) );
  MUX2_X1 U6803 ( .A(n7177), .B(n7176), .S(n5330), .Z(n5262) );
  XNOR2_X1 U6804 ( .A(n5262), .B(SI_15_), .ZN(n5601) );
  INV_X1 U6805 ( .A(n5601), .ZN(n5265) );
  INV_X1 U6806 ( .A(n5262), .ZN(n5263) );
  NAND2_X1 U6807 ( .A1(n5263), .A2(SI_15_), .ZN(n5264) );
  MUX2_X1 U6808 ( .A(n7303), .B(n7305), .S(n5330), .Z(n5266) );
  NAND2_X1 U6809 ( .A1(n5266), .A2(n9273), .ZN(n5269) );
  INV_X1 U6810 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6811 ( .A1(n5267), .A2(SI_16_), .ZN(n5268) );
  NAND2_X1 U6812 ( .A1(n5269), .A2(n5268), .ZN(n5360) );
  MUX2_X1 U6813 ( .A(n7331), .B(n7333), .S(n5330), .Z(n5271) );
  NAND2_X1 U6814 ( .A1(n5271), .A2(n5270), .ZN(n5274) );
  INV_X1 U6815 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6816 ( .A1(n5272), .A2(SI_17_), .ZN(n5273) );
  MUX2_X1 U6817 ( .A(n5276), .B(n5275), .S(n5330), .Z(n5277) );
  XNOR2_X1 U6818 ( .A(n5277), .B(SI_18_), .ZN(n5349) );
  INV_X1 U6819 ( .A(n5349), .ZN(n5280) );
  INV_X1 U6820 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6821 ( .A1(n5278), .A2(SI_18_), .ZN(n5279) );
  MUX2_X1 U6822 ( .A(n9185), .B(n9174), .S(n5330), .Z(n5282) );
  NAND2_X1 U6823 ( .A1(n5282), .A2(n5281), .ZN(n5285) );
  INV_X1 U6824 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6825 ( .A1(n5283), .A2(SI_19_), .ZN(n5284) );
  NAND2_X1 U6826 ( .A1(n5285), .A2(n5284), .ZN(n5633) );
  OAI21_X2 U6827 ( .B1(n5634), .B2(n5633), .A(n5285), .ZN(n5336) );
  MUX2_X1 U6828 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5204), .Z(n5334) );
  INV_X1 U6829 ( .A(n5334), .ZN(n5286) );
  NAND2_X1 U6830 ( .A1(n5336), .A2(n5333), .ZN(n5287) );
  MUX2_X1 U6831 ( .A(n9264), .B(n7790), .S(n5330), .Z(n5650) );
  NAND2_X1 U6832 ( .A1(n5288), .A2(SI_21_), .ZN(n5289) );
  MUX2_X1 U6833 ( .A(n9186), .B(n7935), .S(n5204), .Z(n5291) );
  INV_X1 U6834 ( .A(SI_22_), .ZN(n5290) );
  NAND2_X1 U6835 ( .A1(n5291), .A2(n5290), .ZN(n5294) );
  INV_X1 U6836 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6837 ( .A1(n5292), .A2(SI_22_), .ZN(n5293) );
  NAND2_X1 U6838 ( .A1(n5294), .A2(n5293), .ZN(n5666) );
  MUX2_X1 U6839 ( .A(n7942), .B(n7939), .S(n5330), .Z(n5296) );
  NAND2_X1 U6840 ( .A1(n5296), .A2(n5295), .ZN(n5299) );
  INV_X1 U6841 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6842 ( .A1(n5297), .A2(SI_23_), .ZN(n5298) );
  NAND2_X1 U6843 ( .A1(n5679), .A2(n5678), .ZN(n5300) );
  NAND2_X1 U6844 ( .A1(n5300), .A2(n5299), .ZN(n5692) );
  INV_X1 U6845 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8469) );
  INV_X1 U6846 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8034) );
  MUX2_X1 U6847 ( .A(n8469), .B(n8034), .S(n5330), .Z(n5302) );
  INV_X1 U6848 ( .A(SI_24_), .ZN(n5301) );
  NAND2_X1 U6849 ( .A1(n5302), .A2(n5301), .ZN(n5702) );
  INV_X1 U6850 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U6851 ( .A1(n5303), .A2(SI_24_), .ZN(n5304) );
  NAND2_X1 U6852 ( .A1(n5692), .A2(n5691), .ZN(n5703) );
  INV_X1 U6853 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8415) );
  INV_X1 U6854 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8049) );
  MUX2_X1 U6855 ( .A(n8415), .B(n8049), .S(n5204), .Z(n5306) );
  INV_X1 U6856 ( .A(SI_25_), .ZN(n5305) );
  NAND2_X1 U6857 ( .A1(n5306), .A2(n5305), .ZN(n5705) );
  AND2_X1 U6858 ( .A1(n5702), .A2(n5705), .ZN(n5309) );
  INV_X1 U6859 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6860 ( .A1(n5307), .A2(SI_25_), .ZN(n5704) );
  AOI21_X2 U6861 ( .B1(n5703), .B2(n5309), .A(n5308), .ZN(n5721) );
  MUX2_X1 U6862 ( .A(n8100), .B(n8098), .S(n5330), .Z(n5311) );
  NAND2_X1 U6863 ( .A1(n5311), .A2(n5310), .ZN(n5736) );
  INV_X1 U6864 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6865 ( .A1(n5312), .A2(SI_26_), .ZN(n5313) );
  INV_X1 U6866 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6539) );
  INV_X1 U6867 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8158) );
  MUX2_X1 U6868 ( .A(n6539), .B(n8158), .S(n5204), .Z(n5315) );
  INV_X1 U6869 ( .A(SI_27_), .ZN(n5314) );
  NAND2_X1 U6870 ( .A1(n5315), .A2(n5314), .ZN(n5739) );
  AND2_X1 U6871 ( .A1(n5736), .A2(n5739), .ZN(n5318) );
  INV_X1 U6872 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6873 ( .A1(n5316), .A2(SI_27_), .ZN(n5738) );
  INV_X1 U6874 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8122) );
  INV_X1 U6875 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8161) );
  MUX2_X1 U6876 ( .A(n8122), .B(n8161), .S(n5330), .Z(n5320) );
  INV_X1 U6877 ( .A(SI_28_), .ZN(n5319) );
  NAND2_X1 U6878 ( .A1(n5320), .A2(n5319), .ZN(n5758) );
  INV_X1 U6879 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6880 ( .A1(n5321), .A2(SI_28_), .ZN(n5322) );
  NAND2_X1 U6881 ( .A1(n5324), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6882 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5326) );
  NAND2_X1 U6883 ( .A1(n5328), .A2(n5326), .ZN(n5327) );
  INV_X1 U6884 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6885 ( .A1(n8159), .A2(n5337), .ZN(n5332) );
  OR2_X1 U6886 ( .A1(n5420), .A2(n8161), .ZN(n5331) );
  INV_X1 U6887 ( .A(n10326), .ZN(n10124) );
  XNOR2_X1 U6888 ( .A(n5334), .B(n5333), .ZN(n5335) );
  XNOR2_X1 U6889 ( .A(n5336), .B(n5335), .ZN(n7694) );
  NAND2_X1 U6890 ( .A1(n7694), .A2(n5337), .ZN(n5339) );
  INV_X1 U6891 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7651) );
  OR2_X1 U6892 ( .A1(n5454), .A2(n7651), .ZN(n5338) );
  NAND2_X1 U6893 ( .A1(n5644), .A2(n9613), .ZN(n5340) );
  AND2_X1 U6894 ( .A1(n5656), .A2(n5340), .ZN(n10222) );
  NAND2_X1 U6895 ( .A1(n10222), .A2(n5714), .ZN(n5345) );
  INV_X1 U6896 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U6897 ( .A1(n5695), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6898 ( .A1(n5726), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5341) );
  OAI211_X1 U6899 ( .C1(n4552), .C2(n10432), .A(n5342), .B(n5341), .ZN(n5343)
         );
  INV_X1 U6900 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U6901 ( .A1(n5345), .A2(n5344), .ZN(n9967) );
  NAND2_X1 U6902 ( .A1(n5626), .A2(n9648), .ZN(n5346) );
  NAND2_X1 U6903 ( .A1(n5642), .A2(n5346), .ZN(n10252) );
  AOI22_X1 U6904 ( .A1(n5695), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5747), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6905 ( .A1(n5726), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6906 ( .C1(n10252), .C2(n5766), .A(n5348), .B(n5347), .ZN(n9969)
         );
  XNOR2_X1 U6907 ( .A(n5350), .B(n5349), .ZN(n7334) );
  NAND2_X1 U6908 ( .A1(n7334), .A2(n5337), .ZN(n5359) );
  NAND2_X1 U6909 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n5352) );
  INV_X1 U6910 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5353) );
  INV_X1 U6911 ( .A(n5356), .ZN(n5354) );
  NAND2_X1 U6912 ( .A1(n5354), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6913 ( .A1(n5356), .A2(n5355), .ZN(n5635) );
  AND2_X1 U6914 ( .A1(n5357), .A2(n5635), .ZN(n10075) );
  AOI22_X1 U6915 ( .A1(n5639), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5638), .B2(
        n10075), .ZN(n5358) );
  XNOR2_X1 U6916 ( .A(n5361), .B(n5360), .ZN(n7302) );
  NAND2_X1 U6917 ( .A1(n7302), .A2(n5337), .ZN(n5364) );
  XNOR2_X1 U6918 ( .A(n5362), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U6919 ( .A1(n5639), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5638), .B2(
        n10049), .ZN(n5363) );
  NAND2_X1 U6920 ( .A1(n5747), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6921 ( .A1(n5611), .A2(n5365), .ZN(n5366) );
  AND2_X1 U6922 ( .A1(n5624), .A2(n5366), .ZN(n10291) );
  NAND2_X1 U6923 ( .A1(n5714), .A2(n10291), .ZN(n5369) );
  INV_X1 U6924 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10044) );
  OR2_X1 U6925 ( .A1(n5729), .A2(n10044), .ZN(n5368) );
  INV_X1 U6926 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10029) );
  OR2_X1 U6927 ( .A1(n5458), .A2(n10029), .ZN(n5367) );
  NAND4_X1 U6928 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n9971)
         );
  NAND2_X1 U6929 ( .A1(n5747), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6930 ( .A1(n5695), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6931 ( .A1(n5577), .A2(n9623), .ZN(n5371) );
  NAND2_X1 U6932 ( .A1(n5594), .A2(n5371), .ZN(n9622) );
  OR2_X1 U6933 ( .A1(n5766), .A2(n9622), .ZN(n5373) );
  INV_X1 U6934 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8451) );
  OR2_X1 U6935 ( .A1(n5458), .A2(n8451), .ZN(n5372) );
  NAND4_X1 U6936 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n9974)
         );
  XNOR2_X1 U6937 ( .A(n5377), .B(n5376), .ZN(n6940) );
  NAND2_X1 U6938 ( .A1(n6940), .A2(n5337), .ZN(n5382) );
  NOR2_X1 U6939 ( .A1(n5378), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5537) );
  NOR2_X1 U6940 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5379) );
  NAND2_X1 U6941 ( .A1(n5537), .A2(n5379), .ZN(n5569) );
  NAND2_X1 U6942 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6943 ( .A(n5380), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7871) );
  AOI22_X1 U6944 ( .A1(n5639), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5638), .B2(
        n7871), .ZN(n5381) );
  XNOR2_X1 U6945 ( .A(n5384), .B(n5383), .ZN(n6739) );
  NAND2_X1 U6946 ( .A1(n6739), .A2(n5337), .ZN(n5390) );
  OR2_X1 U6947 ( .A1(n5385), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5470) );
  INV_X1 U6948 ( .A(n5470), .ZN(n5386) );
  NAND2_X1 U6949 ( .A1(n5386), .A2(n5471), .ZN(n5485) );
  INV_X1 U6950 ( .A(n5485), .ZN(n5387) );
  NAND2_X1 U6951 ( .A1(n5387), .A2(n5486), .ZN(n5503) );
  NAND2_X1 U6952 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5388) );
  XNOR2_X1 U6953 ( .A(n5388), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7115) );
  AOI22_X1 U6954 ( .A1(n5639), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5638), .B2(
        n7115), .ZN(n5389) );
  NAND2_X1 U6955 ( .A1(n5390), .A2(n5389), .ZN(n10607) );
  NAND2_X1 U6956 ( .A1(n5747), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6957 ( .A1(n5695), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6958 ( .A1(n5494), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6959 ( .A1(n5508), .A2(n5391), .ZN(n7783) );
  OR2_X1 U6960 ( .A1(n5766), .A2(n7783), .ZN(n5393) );
  INV_X1 U6961 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7779) );
  OR2_X1 U6962 ( .A1(n5458), .A2(n7779), .ZN(n5392) );
  NAND4_X1 U6963 ( .A1(n5395), .A2(n5394), .A3(n5393), .A4(n5392), .ZN(n9980)
         );
  XNOR2_X1 U6964 ( .A(n5397), .B(n5396), .ZN(n6275) );
  INV_X1 U6965 ( .A(n6275), .ZN(n6726) );
  INV_X1 U6966 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6725) );
  INV_X1 U6967 ( .A(n6688), .ZN(n5401) );
  INV_X1 U6968 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6969 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5398) );
  NAND2_X1 U6970 ( .A1(n5695), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5407) );
  INV_X1 U6971 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7042) );
  OR2_X1 U6972 ( .A1(n5425), .A2(n7042), .ZN(n5406) );
  INV_X1 U6973 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7494) );
  OR2_X1 U6974 ( .A1(n5458), .A2(n7494), .ZN(n5405) );
  INV_X1 U6975 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5403) );
  OR2_X1 U6976 ( .A1(n4553), .A2(n5403), .ZN(n5404) );
  NAND4_X2 U6977 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n9987)
         );
  INV_X1 U6978 ( .A(SI_0_), .ZN(n5410) );
  INV_X1 U6979 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5409) );
  OAI21_X1 U6980 ( .B1(n8171), .B2(n5410), .A(n5409), .ZN(n5412) );
  AND2_X1 U6981 ( .A1(n5412), .A2(n5411), .ZN(n10475) );
  INV_X1 U6982 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7297) );
  OR2_X1 U6983 ( .A1(n5425), .A2(n7297), .ZN(n5416) );
  INV_X1 U6984 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6985 ( .A1(n5427), .A2(n5413), .ZN(n5415) );
  INV_X1 U6986 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7242) );
  NAND4_X2 U6987 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n5891)
         );
  NAND2_X1 U6988 ( .A1(n7488), .A2(n5891), .ZN(n7487) );
  NAND2_X1 U6989 ( .A1(n5408), .A2(n4688), .ZN(n5418) );
  NAND2_X1 U6990 ( .A1(n7486), .A2(n5418), .ZN(n7189) );
  OR2_X1 U6991 ( .A1(n5419), .A2(n10461), .ZN(n5435) );
  INV_X1 U6992 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6993 ( .A1(n5695), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5431) );
  INV_X1 U6994 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7502) );
  OR2_X1 U6995 ( .A1(n5425), .A2(n7502), .ZN(n5430) );
  INV_X1 U6996 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7501) );
  OR2_X1 U6997 ( .A1(n5458), .A2(n7501), .ZN(n5429) );
  INV_X1 U6998 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5426) );
  OR2_X1 U6999 ( .A1(n4552), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U7000 ( .A1(n7503), .A2(n9986), .ZN(n9704) );
  INV_X1 U7001 ( .A(n9986), .ZN(n5432) );
  NAND2_X1 U7002 ( .A1(n5432), .A2(n7140), .ZN(n9808) );
  NAND2_X1 U7003 ( .A1(n7189), .A2(n7188), .ZN(n7191) );
  NAND2_X1 U7004 ( .A1(n7503), .A2(n5432), .ZN(n5433) );
  NAND2_X1 U7005 ( .A1(n7191), .A2(n5433), .ZN(n7204) );
  NAND2_X1 U7006 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  NAND2_X1 U7007 ( .A1(n5436), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5438) );
  INV_X1 U7008 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U7009 ( .A(n5440), .B(n5439), .ZN(n6300) );
  INV_X1 U7010 ( .A(n6300), .ZN(n6723) );
  INV_X1 U7011 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U7012 ( .A1(n5695), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7013 ( .A1(n5726), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5446) );
  OR2_X1 U7014 ( .A1(n5766), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5445) );
  INV_X1 U7015 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5443) );
  OR2_X1 U7016 ( .A1(n4552), .A2(n5443), .ZN(n5444) );
  NAND2_X1 U7017 ( .A1(n7450), .A2(n9984), .ZN(n9703) );
  INV_X1 U7018 ( .A(n9984), .ZN(n5448) );
  NAND2_X1 U7019 ( .A1(n5448), .A2(n4561), .ZN(n9809) );
  NAND2_X1 U7020 ( .A1(n7204), .A2(n7203), .ZN(n7202) );
  NAND2_X1 U7021 ( .A1(n7450), .A2(n5448), .ZN(n5449) );
  NAND2_X1 U7022 ( .A1(n7202), .A2(n5449), .ZN(n7293) );
  NAND2_X1 U7023 ( .A1(n5385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  INV_X1 U7024 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5450) );
  XNOR2_X1 U7025 ( .A(n5451), .B(n5450), .ZN(n6952) );
  XNOR2_X1 U7026 ( .A(n5453), .B(n5452), .ZN(n6313) );
  INV_X1 U7027 ( .A(n6313), .ZN(n6728) );
  OR2_X1 U7028 ( .A1(n5762), .A2(n6728), .ZN(n5456) );
  INV_X1 U7029 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6729) );
  OR2_X1 U7030 ( .A1(n5454), .A2(n6729), .ZN(n5455) );
  OAI211_X1 U7031 ( .C1(n6688), .C2(n6952), .A(n5456), .B(n5455), .ZN(n7313)
         );
  NAND2_X1 U7032 ( .A1(n5695), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5467) );
  INV_X1 U7033 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5457) );
  OR2_X1 U7034 ( .A1(n5458), .A2(n5457), .ZN(n5466) );
  INV_X1 U7035 ( .A(n5478), .ZN(n5462) );
  INV_X1 U7036 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5460) );
  INV_X1 U7037 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7038 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U7039 ( .A1(n5462), .A2(n5461), .ZN(n7510) );
  OR2_X1 U7040 ( .A1(n5766), .A2(n7510), .ZN(n5465) );
  INV_X1 U7041 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5463) );
  OR2_X1 U7042 ( .A1(n4552), .A2(n5463), .ZN(n5464) );
  NAND4_X1 U7043 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n9983)
         );
  NAND2_X1 U7044 ( .A1(n7513), .A2(n9983), .ZN(n9876) );
  INV_X1 U7045 ( .A(n9983), .ZN(n5468) );
  NAND2_X1 U7046 ( .A1(n5468), .A2(n7313), .ZN(n9879) );
  AND2_X1 U7047 ( .A1(n9876), .A2(n9879), .ZN(n9813) );
  INV_X1 U7048 ( .A(n9813), .ZN(n7292) );
  NAND2_X1 U7049 ( .A1(n7293), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U7050 ( .A1(n7513), .A2(n5468), .ZN(n5469) );
  NAND2_X1 U7051 ( .A1(n7291), .A2(n5469), .ZN(n7526) );
  NAND2_X1 U7052 ( .A1(n5470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5472) );
  XNOR2_X1 U7053 ( .A(n5472), .B(n5471), .ZN(n6963) );
  NAND2_X1 U7054 ( .A1(n5474), .A2(n5473), .ZN(n5476) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6730) );
  OR2_X1 U7056 ( .A1(n5454), .A2(n6730), .ZN(n5477) );
  NAND2_X1 U7057 ( .A1(n5747), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7058 ( .A1(n5695), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5482) );
  OAI21_X1 U7059 ( .B1(n5478), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5493), .ZN(
        n7586) );
  OR2_X1 U7060 ( .A1(n5766), .A2(n7586), .ZN(n5481) );
  INV_X1 U7061 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5479) );
  OR2_X1 U7062 ( .A1(n5458), .A2(n5479), .ZN(n5480) );
  NAND4_X1 U7063 ( .A1(n5483), .A2(n5482), .A3(n5481), .A4(n5480), .ZN(n9982)
         );
  NAND2_X1 U7064 ( .A1(n10602), .A2(n9982), .ZN(n9884) );
  INV_X1 U7065 ( .A(n9982), .ZN(n9688) );
  NAND2_X1 U7066 ( .A1(n9688), .A2(n9690), .ZN(n9880) );
  NAND2_X1 U7067 ( .A1(n9884), .A2(n9880), .ZN(n9815) );
  NAND2_X1 U7068 ( .A1(n7526), .A2(n9815), .ZN(n7525) );
  NAND2_X1 U7069 ( .A1(n10602), .A2(n9688), .ZN(n5484) );
  NAND2_X1 U7070 ( .A1(n7525), .A2(n5484), .ZN(n7592) );
  NAND2_X1 U7071 ( .A1(n5485), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U7072 ( .A(n5487), .B(n5486), .ZN(n7004) );
  XNOR2_X1 U7073 ( .A(n5489), .B(n5488), .ZN(n6732) );
  NAND2_X1 U7074 ( .A1(n5337), .A2(n6732), .ZN(n5491) );
  INV_X1 U7075 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6733) );
  OR2_X1 U7076 ( .A1(n5454), .A2(n6733), .ZN(n5490) );
  OAI211_X1 U7077 ( .C1(n6688), .C2(n7004), .A(n5491), .B(n5490), .ZN(n9698)
         );
  NAND2_X1 U7078 ( .A1(n5695), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7079 ( .A1(n5747), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5498) );
  AND2_X1 U7080 ( .A1(n5493), .A2(n5492), .ZN(n5495) );
  OR2_X1 U7081 ( .A1(n5495), .A2(n5494), .ZN(n10550) );
  OR2_X1 U7082 ( .A1(n5766), .A2(n10550), .ZN(n5497) );
  INV_X1 U7083 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7005) );
  OR2_X1 U7084 ( .A1(n5458), .A2(n7005), .ZN(n5496) );
  NAND4_X1 U7085 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n9981)
         );
  NAND2_X1 U7086 ( .A1(n10557), .A2(n9981), .ZN(n9706) );
  INV_X1 U7087 ( .A(n9981), .ZN(n9693) );
  NAND2_X1 U7088 ( .A1(n9693), .A2(n9698), .ZN(n9882) );
  NAND2_X1 U7089 ( .A1(n9706), .A2(n9882), .ZN(n7595) );
  NAND2_X1 U7090 ( .A1(n7592), .A2(n7595), .ZN(n7591) );
  NAND2_X1 U7091 ( .A1(n10557), .A2(n9693), .ZN(n5500) );
  NAND2_X1 U7092 ( .A1(n7591), .A2(n5500), .ZN(n7769) );
  INV_X1 U7093 ( .A(n9980), .ZN(n7849) );
  OR2_X1 U7094 ( .A1(n7849), .A2(n10607), .ZN(n9713) );
  NAND2_X1 U7095 ( .A1(n10607), .A2(n7849), .ZN(n7850) );
  INV_X1 U7096 ( .A(n9711), .ZN(n7768) );
  NAND2_X1 U7097 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  XNOR2_X1 U7098 ( .A(n5502), .B(n5501), .ZN(n6743) );
  NAND2_X1 U7099 ( .A1(n6743), .A2(n5337), .ZN(n5506) );
  OAI21_X1 U7100 ( .B1(n5503), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5504) );
  XNOR2_X1 U7101 ( .A(n5504), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10017) );
  AOI22_X1 U7102 ( .A1(n5639), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5638), .B2(
        n10017), .ZN(n5505) );
  NAND2_X1 U7103 ( .A1(n5506), .A2(n5505), .ZN(n7950) );
  NAND2_X1 U7104 ( .A1(n5695), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7105 ( .A1(n5726), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7106 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  NAND2_X1 U7107 ( .A1(n5527), .A2(n5509), .ZN(n10530) );
  OR2_X1 U7108 ( .A1(n5766), .A2(n10530), .ZN(n5512) );
  INV_X1 U7109 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5510) );
  OR2_X1 U7110 ( .A1(n4553), .A2(n5510), .ZN(n5511) );
  NAND4_X1 U7111 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n9979)
         );
  INV_X1 U7112 ( .A(n9979), .ZN(n5515) );
  OR2_X1 U7113 ( .A1(n7950), .A2(n5515), .ZN(n9714) );
  NAND2_X1 U7114 ( .A1(n7950), .A2(n5515), .ZN(n9722) );
  NAND2_X1 U7115 ( .A1(n9714), .A2(n9722), .ZN(n7852) );
  NAND2_X1 U7116 ( .A1(n5517), .A2(n5516), .ZN(n5521) );
  AND2_X1 U7117 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  XNOR2_X1 U7118 ( .A(n5521), .B(n5520), .ZN(n6750) );
  NAND2_X1 U7119 ( .A1(n6750), .A2(n5337), .ZN(n5526) );
  NAND2_X1 U7120 ( .A1(n5378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5522) );
  MUX2_X1 U7121 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5522), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5524) );
  INV_X1 U7122 ( .A(n5537), .ZN(n5523) );
  NAND2_X1 U7123 ( .A1(n5524), .A2(n5523), .ZN(n7124) );
  AOI22_X1 U7124 ( .A1(n5639), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5638), .B2(
        n7252), .ZN(n5525) );
  NAND2_X1 U7125 ( .A1(n5526), .A2(n5525), .ZN(n7763) );
  NAND2_X1 U7126 ( .A1(n5726), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7127 ( .A1(n5747), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5531) );
  INV_X1 U7128 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7117) );
  OR2_X1 U7129 ( .A1(n5729), .A2(n7117), .ZN(n5530) );
  AND2_X1 U7130 ( .A1(n5527), .A2(n7121), .ZN(n5528) );
  OR2_X1 U7131 ( .A1(n5528), .A2(n5544), .ZN(n7760) );
  OR2_X1 U7132 ( .A1(n5766), .A2(n7760), .ZN(n5529) );
  NAND4_X1 U7133 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n9978)
         );
  INV_X1 U7134 ( .A(n9978), .ZN(n7847) );
  OR2_X1 U7135 ( .A1(n7763), .A2(n7847), .ZN(n9733) );
  NAND2_X1 U7136 ( .A1(n4559), .A2(n7847), .ZN(n9732) );
  NAND2_X1 U7137 ( .A1(n9733), .A2(n9732), .ZN(n7756) );
  INV_X1 U7138 ( .A(n5534), .ZN(n5536) );
  XNOR2_X1 U7139 ( .A(n5536), .B(n5535), .ZN(n6753) );
  NAND2_X1 U7140 ( .A1(n6753), .A2(n5337), .ZN(n5543) );
  OR2_X1 U7141 ( .A1(n5537), .A2(n10461), .ZN(n5540) );
  INV_X1 U7142 ( .A(n5540), .ZN(n5538) );
  NAND2_X1 U7143 ( .A1(n5538), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5541) );
  INV_X1 U7144 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7145 ( .A1(n5540), .A2(n5539), .ZN(n5555) );
  AOI22_X1 U7146 ( .A1(n5639), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5638), .B2(
        n7356), .ZN(n5542) );
  NAND2_X1 U7147 ( .A1(n5695), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7148 ( .A1(n5726), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5549) );
  NOR2_X1 U7149 ( .A1(n5544), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5545) );
  OR2_X1 U7150 ( .A1(n5559), .A2(n5545), .ZN(n10488) );
  OR2_X1 U7151 ( .A1(n5766), .A2(n10488), .ZN(n5548) );
  INV_X1 U7152 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5546) );
  OR2_X1 U7153 ( .A1(n4553), .A2(n5546), .ZN(n5547) );
  NAND4_X1 U7154 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n9977)
         );
  INV_X1 U7155 ( .A(n9977), .ZN(n5551) );
  OR2_X1 U7156 ( .A1(n10486), .A2(n5551), .ZN(n9891) );
  NAND2_X1 U7157 ( .A1(n10486), .A2(n5551), .ZN(n9736) );
  NAND2_X1 U7158 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  NAND2_X1 U7159 ( .A1(n7797), .A2(n5552), .ZN(n7924) );
  XNOR2_X1 U7160 ( .A(n5554), .B(n5553), .ZN(n6817) );
  NAND2_X1 U7161 ( .A1(n6817), .A2(n5337), .ZN(n5558) );
  NAND2_X1 U7162 ( .A1(n5555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5556) );
  XNOR2_X1 U7163 ( .A(n5556), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7395) );
  AOI22_X1 U7164 ( .A1(n5639), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5638), .B2(
        n7395), .ZN(n5557) );
  NAND2_X1 U7165 ( .A1(n5695), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7166 ( .A1(n5747), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5563) );
  OR2_X1 U7167 ( .A1(n5559), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7168 ( .A1(n5575), .A2(n5560), .ZN(n10517) );
  OR2_X1 U7169 ( .A1(n5766), .A2(n10517), .ZN(n5562) );
  INV_X1 U7170 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7926) );
  OR2_X1 U7171 ( .A1(n5458), .A2(n7926), .ZN(n5561) );
  NAND4_X1 U7172 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n9976)
         );
  INV_X1 U7173 ( .A(n9976), .ZN(n5565) );
  NAND2_X1 U7174 ( .A1(n10625), .A2(n5565), .ZN(n9738) );
  NAND2_X1 U7175 ( .A1(n9737), .A2(n9738), .ZN(n7923) );
  XNOR2_X1 U7176 ( .A(n5568), .B(n5567), .ZN(n6892) );
  NAND2_X1 U7177 ( .A1(n6892), .A2(n5337), .ZN(n5573) );
  NAND2_X1 U7178 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  MUX2_X1 U7179 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5570), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5571) );
  AOI22_X1 U7180 ( .A1(n5639), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5638), .B2(
        n7709), .ZN(n5572) );
  NAND2_X1 U7181 ( .A1(n5747), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7182 ( .A1(n5695), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7183 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  NAND2_X1 U7184 ( .A1(n5577), .A2(n5576), .ZN(n10505) );
  OR2_X1 U7185 ( .A1(n5766), .A2(n10505), .ZN(n5579) );
  INV_X1 U7186 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7977) );
  OR2_X1 U7187 ( .A1(n5458), .A2(n7977), .ZN(n5578) );
  NAND4_X1 U7188 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n9975)
         );
  INV_X1 U7189 ( .A(n9975), .ZN(n5582) );
  NAND2_X1 U7190 ( .A1(n10503), .A2(n5582), .ZN(n9893) );
  INV_X1 U7191 ( .A(n9974), .ZN(n5583) );
  OR2_X1 U7192 ( .A1(n8456), .A2(n5583), .ZN(n9897) );
  NAND2_X1 U7193 ( .A1(n8456), .A2(n5583), .ZN(n9894) );
  NAND2_X1 U7194 ( .A1(n9897), .A2(n9894), .ZN(n9823) );
  AND2_X1 U7195 ( .A1(n7974), .A2(n9823), .ZN(n5585) );
  INV_X1 U7196 ( .A(n9823), .ZN(n5584) );
  OR2_X1 U7197 ( .A1(n10503), .A2(n9975), .ZN(n8448) );
  NAND2_X1 U7198 ( .A1(n5586), .A2(n5587), .ZN(n5589) );
  XNOR2_X1 U7199 ( .A(n5589), .B(n5588), .ZN(n7179) );
  NAND2_X1 U7200 ( .A1(n7179), .A2(n5337), .ZN(n5592) );
  OAI21_X1 U7201 ( .B1(n5590), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5604) );
  XNOR2_X1 U7202 ( .A(n5604), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8054) );
  AOI22_X1 U7203 ( .A1(n5639), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5638), .B2(
        n8054), .ZN(n5591) );
  INV_X1 U7204 ( .A(n9534), .ZN(n8076) );
  NAND2_X1 U7205 ( .A1(n5747), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7206 ( .A1(n5695), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5598) );
  INV_X1 U7207 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7208 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  NAND2_X1 U7209 ( .A1(n5609), .A2(n5595), .ZN(n9532) );
  OR2_X1 U7210 ( .A1(n5766), .A2(n9532), .ZN(n5597) );
  INV_X1 U7211 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8068) );
  OR2_X1 U7212 ( .A1(n5458), .A2(n8068), .ZN(n5596) );
  NAND4_X1 U7213 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n9973)
         );
  INV_X1 U7214 ( .A(n9973), .ZN(n5848) );
  XNOR2_X1 U7215 ( .A(n5602), .B(n5601), .ZN(n7175) );
  NAND2_X1 U7216 ( .A1(n7175), .A2(n5337), .ZN(n5608) );
  INV_X1 U7217 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7218 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U7219 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  XNOR2_X1 U7220 ( .A(n5606), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8057) );
  AOI22_X1 U7221 ( .A1(n5639), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5638), .B2(
        n8057), .ZN(n5607) );
  INV_X1 U7222 ( .A(n10454), .ZN(n10310) );
  NAND2_X1 U7223 ( .A1(n5747), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7224 ( .A1(n5726), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5614) );
  INV_X1 U7225 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8055) );
  OR2_X1 U7226 ( .A1(n5729), .A2(n8055), .ZN(n5613) );
  INV_X1 U7227 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U7228 ( .A1(n5609), .A2(n9668), .ZN(n5610) );
  NAND2_X1 U7229 ( .A1(n5611), .A2(n5610), .ZN(n10297) );
  OR2_X1 U7230 ( .A1(n5766), .A2(n10297), .ZN(n5612) );
  NAND4_X1 U7231 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n9972)
         );
  INV_X1 U7232 ( .A(n9972), .ZN(n5849) );
  NAND2_X1 U7233 ( .A1(n10310), .A2(n5849), .ZN(n5616) );
  INV_X1 U7234 ( .A(n9971), .ZN(n5618) );
  NAND2_X1 U7235 ( .A1(n10384), .A2(n5618), .ZN(n10260) );
  XNOR2_X1 U7236 ( .A(n5620), .B(n5619), .ZN(n7330) );
  NAND2_X1 U7237 ( .A1(n7330), .A2(n5337), .ZN(n5623) );
  XNOR2_X1 U7238 ( .A(n5621), .B(n5353), .ZN(n10064) );
  AOI22_X1 U7239 ( .A1(n5639), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5638), .B2(
        n10064), .ZN(n5622) );
  INV_X1 U7240 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U7241 ( .A1(n5624), .A2(n9600), .ZN(n5625) );
  NAND2_X1 U7242 ( .A1(n5626), .A2(n5625), .ZN(n10271) );
  OR2_X1 U7243 ( .A1(n10271), .A2(n5766), .ZN(n5630) );
  NAND2_X1 U7244 ( .A1(n5747), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7245 ( .A1(n5695), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5628) );
  INV_X1 U7246 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10272) );
  OR2_X1 U7247 ( .A1(n5458), .A2(n10272), .ZN(n5627) );
  NAND4_X1 U7248 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n9970)
         );
  NAND2_X1 U7249 ( .A1(n10443), .A2(n9970), .ZN(n5631) );
  INV_X1 U7250 ( .A(n9970), .ZN(n5852) );
  OAI21_X1 U7251 ( .B1(n9969), .B2(n10374), .A(n10244), .ZN(n5632) );
  INV_X1 U7252 ( .A(n10374), .ZN(n10256) );
  INV_X1 U7253 ( .A(n9969), .ZN(n5853) );
  NAND2_X1 U7254 ( .A1(n5632), .A2(n5162), .ZN(n10228) );
  XNOR2_X1 U7255 ( .A(n5634), .B(n5633), .ZN(n7548) );
  NAND2_X1 U7256 ( .A1(n7548), .A2(n5337), .ZN(n5641) );
  NAND2_X1 U7257 ( .A1(n5635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U7258 ( .A(n5637), .B(n5636), .ZN(n5822) );
  AOI22_X1 U7259 ( .A1(n5639), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5638), .B2(
        n10211), .ZN(n5640) );
  INV_X1 U7260 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10233) );
  INV_X1 U7261 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U7262 ( .A1(n5642), .A2(n9559), .ZN(n5643) );
  NAND2_X1 U7263 ( .A1(n5644), .A2(n5643), .ZN(n10232) );
  OR2_X1 U7264 ( .A1(n10232), .A2(n5766), .ZN(n5646) );
  AOI22_X1 U7265 ( .A1(n5695), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5747), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5645) );
  OAI211_X1 U7266 ( .C1(n5458), .C2(n10233), .A(n5646), .B(n5645), .ZN(n9968)
         );
  INV_X1 U7267 ( .A(n9968), .ZN(n5855) );
  NAND2_X1 U7268 ( .A1(n4845), .A2(n5855), .ZN(n5648) );
  AOI21_X2 U7269 ( .B1(n10228), .B2(n5648), .A(n5647), .ZN(n10215) );
  INV_X1 U7270 ( .A(n10364), .ZN(n10225) );
  INV_X1 U7271 ( .A(n9967), .ZN(n5856) );
  NAND2_X1 U7272 ( .A1(n10215), .A2(n5159), .ZN(n5649) );
  XNOR2_X1 U7273 ( .A(n5650), .B(SI_21_), .ZN(n5651) );
  XNOR2_X1 U7274 ( .A(n5652), .B(n5651), .ZN(n7789) );
  NAND2_X1 U7275 ( .A1(n7789), .A2(n5337), .ZN(n5654) );
  OR2_X1 U7276 ( .A1(n5454), .A2(n7790), .ZN(n5653) );
  INV_X1 U7277 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7278 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  NAND2_X1 U7279 ( .A1(n5671), .A2(n5657), .ZN(n10210) );
  OR2_X1 U7280 ( .A1(n10210), .A2(n5766), .ZN(n5664) );
  INV_X1 U7281 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7282 ( .A1(n5695), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5660) );
  INV_X1 U7283 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5658) );
  OR2_X1 U7284 ( .A1(n4553), .A2(n5658), .ZN(n5659) );
  OAI211_X1 U7285 ( .C1(n5661), .C2(n5458), .A(n5660), .B(n5659), .ZN(n5662)
         );
  INV_X1 U7286 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7287 ( .A1(n5664), .A2(n5663), .ZN(n9966) );
  NOR2_X1 U7288 ( .A1(n10428), .A2(n9966), .ZN(n5665) );
  INV_X1 U7289 ( .A(n10428), .ZN(n10209) );
  INV_X1 U7290 ( .A(n9966), .ZN(n9806) );
  NAND2_X1 U7291 ( .A1(n7931), .A2(n5337), .ZN(n5669) );
  OR2_X1 U7292 ( .A1(n5420), .A2(n7935), .ZN(n5668) );
  NAND2_X1 U7293 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  AND2_X1 U7294 ( .A1(n5683), .A2(n5672), .ZN(n10195) );
  NAND2_X1 U7295 ( .A1(n10195), .A2(n5714), .ZN(n5677) );
  INV_X1 U7296 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U7297 ( .A1(n5747), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5674) );
  INV_X1 U7298 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9162) );
  OR2_X1 U7299 ( .A1(n5458), .A2(n9162), .ZN(n5673) );
  OAI211_X1 U7300 ( .C1(n5729), .C2(n10354), .A(n5674), .B(n5673), .ZN(n5675)
         );
  INV_X1 U7301 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U7302 ( .A1(n5677), .A2(n5676), .ZN(n9965) );
  INV_X1 U7303 ( .A(n9965), .ZN(n6082) );
  XNOR2_X1 U7304 ( .A(n5679), .B(n5678), .ZN(n7940) );
  NAND2_X1 U7305 ( .A1(n7940), .A2(n5337), .ZN(n5681) );
  OR2_X1 U7306 ( .A1(n5420), .A2(n7939), .ZN(n5680) );
  INV_X1 U7307 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7308 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  NAND2_X1 U7309 ( .A1(n5712), .A2(n5684), .ZN(n9541) );
  OR2_X1 U7310 ( .A1(n9541), .A2(n5766), .ZN(n5689) );
  INV_X1 U7311 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U7312 ( .A1(n5747), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7313 ( .A1(n5726), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5685) );
  OAI211_X1 U7314 ( .C1(n5729), .C2(n10349), .A(n5686), .B(n5685), .ZN(n5687)
         );
  INV_X1 U7315 ( .A(n5687), .ZN(n5688) );
  NOR2_X1 U7316 ( .A1(n10179), .A2(n9964), .ZN(n5690) );
  INV_X1 U7317 ( .A(n10179), .ZN(n10346) );
  INV_X1 U7318 ( .A(n9964), .ZN(n5858) );
  XNOR2_X1 U7319 ( .A(n5692), .B(n5691), .ZN(n8033) );
  NAND2_X1 U7320 ( .A1(n8033), .A2(n5337), .ZN(n5694) );
  OR2_X1 U7321 ( .A1(n5420), .A2(n8034), .ZN(n5693) );
  INV_X1 U7322 ( .A(n10341), .ZN(n10170) );
  XNOR2_X1 U7323 ( .A(n5712), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U7324 ( .A1(n10167), .A2(n5714), .ZN(n5700) );
  INV_X1 U7325 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U7326 ( .A1(n5726), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7327 ( .A1(n5695), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7328 ( .C1(n4552), .C2(n10415), .A(n5697), .B(n5696), .ZN(n5698)
         );
  INV_X1 U7329 ( .A(n5698), .ZN(n5699) );
  INV_X1 U7330 ( .A(n9963), .ZN(n5859) );
  NOR2_X1 U7331 ( .A1(n10170), .A2(n5859), .ZN(n5701) );
  NAND2_X1 U7332 ( .A1(n5703), .A2(n5702), .ZN(n5707) );
  AND2_X1 U7333 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  NAND2_X1 U7334 ( .A1(n8048), .A2(n5337), .ZN(n5709) );
  OR2_X1 U7335 ( .A1(n5420), .A2(n8049), .ZN(n5708) );
  NAND2_X2 U7336 ( .A1(n5709), .A2(n5708), .ZN(n10411) );
  OAI21_X1 U7337 ( .B1(n5712), .B2(n5711), .A(n5710), .ZN(n5713) );
  AND2_X1 U7338 ( .A1(n5713), .A2(n5724), .ZN(n10153) );
  NAND2_X1 U7339 ( .A1(n10153), .A2(n5714), .ZN(n5719) );
  INV_X1 U7340 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U7341 ( .A1(n5726), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7342 ( .A1(n5695), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5715) );
  OAI211_X1 U7343 ( .C1(n4553), .C2(n9329), .A(n5716), .B(n5715), .ZN(n5717)
         );
  INV_X1 U7344 ( .A(n5717), .ZN(n5718) );
  INV_X1 U7345 ( .A(n10411), .ZN(n10152) );
  NAND2_X1 U7346 ( .A1(n8097), .A2(n5337), .ZN(n5723) );
  NAND2_X2 U7347 ( .A1(n5723), .A2(n5722), .ZN(n10406) );
  INV_X1 U7348 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U7349 ( .A1(n5724), .A2(n9658), .ZN(n5725) );
  NAND2_X1 U7350 ( .A1(n5745), .A2(n5725), .ZN(n10138) );
  OR2_X1 U7351 ( .A1(n10138), .A2(n5766), .ZN(n5732) );
  INV_X1 U7352 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U7353 ( .A1(n5747), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7354 ( .A1(n5726), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5727) );
  OAI211_X1 U7355 ( .C1(n5729), .C2(n10332), .A(n5728), .B(n5727), .ZN(n5730)
         );
  INV_X1 U7356 ( .A(n5730), .ZN(n5731) );
  NAND2_X2 U7357 ( .A1(n5732), .A2(n5731), .ZN(n9961) );
  NOR2_X1 U7358 ( .A1(n10142), .A2(n5863), .ZN(n5733) );
  NAND2_X1 U7359 ( .A1(n10142), .A2(n5863), .ZN(n5734) );
  NAND2_X1 U7360 ( .A1(n5737), .A2(n5736), .ZN(n5741) );
  AND2_X1 U7361 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  NAND2_X1 U7362 ( .A1(n8103), .A2(n5337), .ZN(n5743) );
  OR2_X1 U7363 ( .A1(n5420), .A2(n8158), .ZN(n5742) );
  INV_X1 U7364 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7365 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NAND2_X1 U7366 ( .A1(n5827), .A2(n5746), .ZN(n8433) );
  OR2_X1 U7367 ( .A1(n8433), .A2(n5766), .ZN(n5753) );
  INV_X1 U7368 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7369 ( .A1(n5747), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7370 ( .A1(n5695), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5748) );
  OAI211_X1 U7371 ( .C1(n5750), .C2(n5458), .A(n5749), .B(n5748), .ZN(n5751)
         );
  INV_X1 U7372 ( .A(n5751), .ZN(n5752) );
  NAND2_X1 U7373 ( .A1(n8479), .A2(n5754), .ZN(n9777) );
  NAND2_X1 U7374 ( .A1(n9854), .A2(n9777), .ZN(n9836) );
  INV_X1 U7375 ( .A(n8479), .ZN(n8436) );
  NOR2_X1 U7376 ( .A1(n10326), .A2(n5755), .ZN(n9863) );
  INV_X1 U7377 ( .A(n9863), .ZN(n9779) );
  NAND2_X1 U7378 ( .A1(n10326), .A2(n5755), .ZN(n9778) );
  OAI21_X1 U7379 ( .B1(n5755), .B2(n10124), .A(n10323), .ZN(n5776) );
  NAND2_X1 U7380 ( .A1(n5757), .A2(n5756), .ZN(n5759) );
  MUX2_X1 U7381 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8171), .Z(n8163) );
  OR2_X1 U7382 ( .A1(n10471), .A2(n5762), .ZN(n5764) );
  INV_X1 U7383 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10474) );
  OR2_X1 U7384 ( .A1(n5420), .A2(n10474), .ZN(n5763) );
  INV_X1 U7385 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5765) );
  OR2_X1 U7386 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  OR2_X1 U7387 ( .A1(n5827), .A2(n5767), .ZN(n5773) );
  INV_X1 U7388 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7389 ( .A1(n5695), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5770) );
  INV_X1 U7390 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5768) );
  OR2_X1 U7391 ( .A1(n4552), .A2(n5768), .ZN(n5769) );
  OAI211_X1 U7392 ( .C1(n5825), .C2(n5458), .A(n5770), .B(n5769), .ZN(n5771)
         );
  INV_X1 U7393 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7394 ( .A1(n5773), .A2(n5772), .ZN(n9958) );
  INV_X1 U7395 ( .A(n9958), .ZN(n5774) );
  NAND2_X1 U7396 ( .A1(n8489), .A2(n5774), .ZN(n9913) );
  XNOR2_X2 U7397 ( .A(n5776), .B(n5775), .ZN(n8491) );
  NAND2_X1 U7398 ( .A1(n5780), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7399 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5784) );
  INV_X1 U7400 ( .A(n5786), .ZN(n5787) );
  INV_X1 U7401 ( .A(n10458), .ZN(n5815) );
  NAND2_X1 U7402 ( .A1(n5792), .A2(P1_B_REG_SCAN_IN), .ZN(n5794) );
  MUX2_X1 U7403 ( .A(n5794), .B(P1_B_REG_SCAN_IN), .S(n5793), .Z(n5796) );
  NOR4_X1 U7404 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5805) );
  NOR4_X1 U7405 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5804) );
  INV_X1 U7406 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10564) );
  INV_X1 U7407 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10594) );
  INV_X1 U7408 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10586) );
  INV_X1 U7409 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U7410 ( .A1(n10564), .A2(n10594), .A3(n10586), .A4(n10592), .ZN(
        n5802) );
  NOR4_X1 U7411 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5800) );
  NOR4_X1 U7412 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5799) );
  NOR4_X1 U7413 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5798) );
  NOR4_X1 U7414 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5797) );
  NAND4_X1 U7415 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n5801)
         );
  NOR4_X1 U7416 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5802), .A4(n5801), .ZN(n5803) );
  NAND3_X1 U7417 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n5806) );
  NAND2_X1 U7418 ( .A1(n6747), .A2(n5806), .ZN(n6120) );
  NAND2_X1 U7419 ( .A1(n5807), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7420 ( .A1(n4611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7421 ( .A1(n9932), .A2(n6122), .ZN(n6134) );
  NAND3_X1 U7422 ( .A1(n5815), .A2(n6120), .A3(n6134), .ZN(n6857) );
  INV_X1 U7423 ( .A(n6857), .ZN(n5819) );
  INV_X1 U7424 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5817) );
  INV_X1 U7425 ( .A(n5795), .ZN(n8099) );
  INV_X1 U7426 ( .A(n10459), .ZN(n7260) );
  INV_X1 U7427 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5818) );
  NAND3_X1 U7428 ( .A1(n5819), .A2(n7260), .A3(n6856), .ZN(n5830) );
  NAND2_X1 U7429 ( .A1(n10319), .A2(n10211), .ZN(n6854) );
  INV_X1 U7430 ( .A(n6122), .ZN(n9949) );
  NAND2_X1 U7431 ( .A1(n9949), .A2(n9932), .ZN(n5821) );
  INV_X1 U7432 ( .A(n6121), .ZN(n6861) );
  NAND2_X1 U7433 ( .A1(n5821), .A2(n6861), .ZN(n7239) );
  NAND2_X1 U7434 ( .A1(n9938), .A2(n9802), .ZN(n5886) );
  AND2_X1 U7435 ( .A1(n6122), .A2(n5886), .ZN(n5823) );
  OR2_X1 U7436 ( .A1(n7239), .A2(n5823), .ZN(n7776) );
  OR2_X1 U7437 ( .A1(n10553), .A2(n7776), .ZN(n5824) );
  OR2_X1 U7438 ( .A1(n6861), .A2(n4549), .ZN(n6130) );
  NOR2_X2 U7439 ( .A1(n10563), .A2(n6130), .ZN(n10278) );
  NAND2_X1 U7440 ( .A1(n10551), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5826) );
  OAI22_X1 U7441 ( .A1(n5827), .A2(n5826), .B1(n5825), .B2(n5878), .ZN(n5832)
         );
  INV_X1 U7442 ( .A(n8489), .ZN(n5829) );
  INV_X1 U7443 ( .A(n7488), .ZN(n7185) );
  OR2_X1 U7444 ( .A1(n7594), .A2(n9698), .ZN(n7780) );
  INV_X1 U7445 ( .A(n7950), .ZN(n10525) );
  INV_X1 U7446 ( .A(n4559), .ZN(n10618) );
  NAND2_X1 U7447 ( .A1(n8453), .A2(n9629), .ZN(n8452) );
  INV_X1 U7448 ( .A(n10384), .ZN(n10293) );
  NAND2_X1 U7449 ( .A1(n10209), .A2(n10221), .ZN(n10208) );
  NOR2_X1 U7450 ( .A1(n10180), .A2(n10341), .ZN(n10166) );
  NAND2_X1 U7451 ( .A1(n10166), .A2(n10152), .ZN(n10151) );
  NOR2_X2 U7452 ( .A1(n10151), .A2(n10406), .ZN(n10137) );
  OAI211_X1 U7453 ( .C1(n5829), .C2(n10120), .A(n10109), .B(n10319), .ZN(n8485) );
  NOR2_X1 U7454 ( .A1(n8485), .A2(n10275), .ZN(n5831) );
  AOI211_X1 U7455 ( .C1(n10278), .C2(n8489), .A(n5832), .B(n5831), .ZN(n5881)
         );
  NAND2_X1 U7456 ( .A1(n10194), .A2(n6082), .ZN(n9852) );
  OR2_X1 U7457 ( .A1(n10428), .A2(n9806), .ZN(n9762) );
  OR2_X1 U7458 ( .A1(n10364), .A2(n5856), .ZN(n10202) );
  NAND2_X1 U7459 ( .A1(n9762), .A2(n10202), .ZN(n9861) );
  INV_X1 U7460 ( .A(n5891), .ZN(n5834) );
  AND2_X1 U7461 ( .A1(n5834), .A2(n7488), .ZN(n7490) );
  NAND2_X1 U7462 ( .A1(n4688), .A2(n5897), .ZN(n5835) );
  NAND2_X1 U7463 ( .A1(n5836), .A2(n5835), .ZN(n9701) );
  NAND2_X1 U7464 ( .A1(n9701), .A2(n9704), .ZN(n5837) );
  NAND2_X1 U7465 ( .A1(n5837), .A2(n9808), .ZN(n9684) );
  NAND2_X1 U7466 ( .A1(n9684), .A2(n7196), .ZN(n7195) );
  NAND2_X1 U7467 ( .A1(n7195), .A2(n9809), .ZN(n7286) );
  NAND2_X1 U7468 ( .A1(n7286), .A2(n9876), .ZN(n5838) );
  NAND2_X1 U7469 ( .A1(n9733), .A2(n9714), .ZN(n9720) );
  NAND2_X1 U7470 ( .A1(n9713), .A2(n9706), .ZN(n5839) );
  NOR2_X1 U7471 ( .A1(n9720), .A2(n5839), .ZN(n9886) );
  NAND2_X1 U7472 ( .A1(n5840), .A2(n9886), .ZN(n7792) );
  AND2_X1 U7473 ( .A1(n9722), .A2(n7850), .ZN(n7751) );
  OR2_X1 U7474 ( .A1(n9720), .A2(n7751), .ZN(n5841) );
  AND2_X1 U7475 ( .A1(n5841), .A2(n9732), .ZN(n9887) );
  NAND2_X1 U7476 ( .A1(n7792), .A2(n9887), .ZN(n5842) );
  NAND2_X1 U7477 ( .A1(n5842), .A2(n9820), .ZN(n7916) );
  INV_X1 U7478 ( .A(n9736), .ZN(n5843) );
  NOR2_X1 U7479 ( .A1(n7923), .A2(n5843), .ZN(n5844) );
  NAND2_X1 U7480 ( .A1(n7916), .A2(n5844), .ZN(n7920) );
  NAND2_X1 U7481 ( .A1(n7920), .A2(n9737), .ZN(n7970) );
  INV_X1 U7482 ( .A(n9739), .ZN(n5845) );
  NOR2_X1 U7483 ( .A1(n9823), .A2(n5845), .ZN(n5846) );
  OR2_X1 U7484 ( .A1(n9534), .A2(n5848), .ZN(n10298) );
  NAND2_X1 U7485 ( .A1(n9534), .A2(n5848), .ZN(n9731) );
  NAND2_X1 U7486 ( .A1(n10298), .A2(n9731), .ZN(n9743) );
  OR2_X1 U7487 ( .A1(n10454), .A2(n5849), .ZN(n9899) );
  NAND2_X1 U7488 ( .A1(n10454), .A2(n5849), .ZN(n9746) );
  NAND2_X1 U7489 ( .A1(n9899), .A2(n9746), .ZN(n10305) );
  INV_X1 U7490 ( .A(n10298), .ZN(n5850) );
  NOR2_X1 U7491 ( .A1(n10305), .A2(n5850), .ZN(n5851) );
  NAND2_X1 U7492 ( .A1(n10443), .A2(n5852), .ZN(n9753) );
  OR2_X1 U7493 ( .A1(n10374), .A2(n5853), .ZN(n9905) );
  NAND2_X1 U7494 ( .A1(n10374), .A2(n5853), .ZN(n9760) );
  NAND3_X1 U7495 ( .A1(n10263), .A2(n10246), .A3(n10245), .ZN(n5854) );
  NAND2_X1 U7496 ( .A1(n5854), .A2(n9760), .ZN(n10237) );
  OR2_X1 U7497 ( .A1(n10369), .A2(n5855), .ZN(n9906) );
  NAND2_X1 U7498 ( .A1(n10369), .A2(n5855), .ZN(n9869) );
  NAND2_X1 U7499 ( .A1(n10428), .A2(n9806), .ZN(n9763) );
  NAND2_X1 U7500 ( .A1(n10364), .A2(n5856), .ZN(n9681) );
  NAND2_X1 U7501 ( .A1(n9763), .A2(n9681), .ZN(n5857) );
  NAND2_X1 U7502 ( .A1(n5857), .A2(n9762), .ZN(n9851) );
  NAND2_X1 U7503 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  OR2_X1 U7504 ( .A1(n10179), .A2(n5858), .ZN(n9770) );
  NAND2_X1 U7505 ( .A1(n10179), .A2(n5858), .ZN(n9840) );
  NOR2_X1 U7506 ( .A1(n10341), .A2(n5859), .ZN(n9844) );
  INV_X1 U7507 ( .A(n9844), .ZN(n5860) );
  NAND2_X1 U7508 ( .A1(n10341), .A2(n5859), .ZN(n9841) );
  NAND2_X1 U7509 ( .A1(n5860), .A2(n9841), .ZN(n10160) );
  OR2_X1 U7510 ( .A1(n10411), .A2(n5861), .ZN(n9805) );
  INV_X1 U7511 ( .A(n9805), .ZN(n5862) );
  NAND2_X1 U7512 ( .A1(n10411), .A2(n5861), .ZN(n9848) );
  NAND2_X1 U7513 ( .A1(n9847), .A2(n9775), .ZN(n10128) );
  INV_X1 U7514 ( .A(n10128), .ZN(n10132) );
  NAND2_X1 U7515 ( .A1(n10131), .A2(n10132), .ZN(n10130) );
  NAND2_X1 U7516 ( .A1(n10130), .A2(n9775), .ZN(n8422) );
  NAND2_X1 U7517 ( .A1(n8422), .A2(n8423), .ZN(n8421) );
  NAND2_X1 U7518 ( .A1(n8421), .A2(n9777), .ZN(n10115) );
  NAND2_X1 U7519 ( .A1(n10115), .A2(n10116), .ZN(n10114) );
  NAND2_X1 U7520 ( .A1(n10114), .A2(n9778), .ZN(n5864) );
  XNOR2_X1 U7521 ( .A(n5864), .B(n9838), .ZN(n5877) );
  OR2_X1 U7522 ( .A1(n7933), .A2(n9938), .ZN(n5865) );
  OR2_X1 U7523 ( .A1(n9807), .A2(n4549), .ZN(n9801) );
  NAND2_X1 U7524 ( .A1(n5695), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5869) );
  INV_X1 U7525 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7526 ( .A1(n5458), .A2(n5866), .ZN(n5868) );
  INV_X1 U7527 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10400) );
  OR2_X1 U7528 ( .A1(n4553), .A2(n10400), .ZN(n5867) );
  AND3_X1 U7529 ( .A1(n5869), .A2(n5868), .A3(n5867), .ZN(n9804) );
  AND2_X2 U7530 ( .A1(n5871), .A2(n9932), .ZN(n9667) );
  INV_X1 U7531 ( .A(P1_B_REG_SCAN_IN), .ZN(n5873) );
  OR2_X1 U7532 ( .A1(n4558), .A2(n5873), .ZN(n5874) );
  NAND2_X1 U7533 ( .A1(n9667), .A2(n5874), .ZN(n10103) );
  INV_X1 U7534 ( .A(n5871), .ZN(n6682) );
  NAND2_X1 U7535 ( .A1(n6682), .A2(n9932), .ZN(n7848) );
  INV_X2 U7536 ( .A(n7848), .ZN(n9666) );
  NAND2_X1 U7537 ( .A1(n9959), .A2(n9666), .ZN(n5875) );
  OAI21_X1 U7538 ( .B1(n9804), .B2(n10103), .A(n5875), .ZN(n5876) );
  INV_X1 U7539 ( .A(n8486), .ZN(n5879) );
  OAI21_X1 U7540 ( .B1(n8491), .B2(n10259), .A(n5882), .ZN(P1_U3356) );
  OAI21_X1 U7541 ( .B1(n6122), .B2(n9802), .A(n5883), .ZN(n5884) );
  INV_X1 U7542 ( .A(n5888), .ZN(n5885) );
  AND2_X1 U7543 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7544 ( .A1(n5889), .A2(n5887), .ZN(n5927) );
  NAND2_X1 U7545 ( .A1(n4832), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7546 ( .A1(n5895), .A2(n5890), .ZN(n6680) );
  INV_X1 U7547 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7548 ( .A1(n7488), .A2(n5957), .ZN(n5893) );
  OAI211_X1 U7549 ( .C1(n6685), .C2(n5894), .A(n5893), .B(n5892), .ZN(n6679)
         );
  INV_X2 U7550 ( .A(n6110), .ZN(n6074) );
  NAND2_X1 U7551 ( .A1(n5895), .A2(n6074), .ZN(n5896) );
  NAND2_X1 U7552 ( .A1(n5897), .A2(n5936), .ZN(n5899) );
  NAND2_X1 U7553 ( .A1(n9987), .A2(n5957), .ZN(n5898) );
  NAND2_X1 U7554 ( .A1(n5899), .A2(n5898), .ZN(n5900) );
  XNOR2_X2 U7555 ( .A(n5900), .B(n6110), .ZN(n7036) );
  NAND2_X1 U7556 ( .A1(n5897), .A2(n5957), .ZN(n5902) );
  NAND2_X1 U7557 ( .A1(n9987), .A2(n4543), .ZN(n5901) );
  NAND2_X1 U7558 ( .A1(n5902), .A2(n5901), .ZN(n7033) );
  NAND2_X1 U7559 ( .A1(n7034), .A2(n7036), .ZN(n5903) );
  NAND2_X1 U7560 ( .A1(n7140), .A2(n5936), .ZN(n5906) );
  NAND2_X1 U7561 ( .A1(n9986), .A2(n5957), .ZN(n5905) );
  NAND2_X1 U7562 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  XNOR2_X1 U7563 ( .A(n5907), .B(n6074), .ZN(n5910) );
  NAND2_X1 U7564 ( .A1(n7140), .A2(n5957), .ZN(n5909) );
  NAND2_X1 U7565 ( .A1(n9986), .A2(n4543), .ZN(n5908) );
  AND2_X1 U7566 ( .A1(n5909), .A2(n5908), .ZN(n5911) );
  NAND2_X1 U7567 ( .A1(n5910), .A2(n5911), .ZN(n5915) );
  INV_X1 U7568 ( .A(n5910), .ZN(n5913) );
  INV_X1 U7569 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7570 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  NAND2_X1 U7571 ( .A1(n9984), .A2(n5957), .ZN(n5917) );
  NAND2_X1 U7572 ( .A1(n4561), .A2(n5936), .ZN(n5916) );
  NAND2_X1 U7573 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  XNOR2_X1 U7574 ( .A(n5918), .B(n6074), .ZN(n5923) );
  NAND2_X1 U7575 ( .A1(n4561), .A2(n5957), .ZN(n5920) );
  NAND2_X1 U7576 ( .A1(n9984), .A2(n4543), .ZN(n5919) );
  NAND2_X1 U7577 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  XNOR2_X1 U7578 ( .A(n5923), .B(n5921), .ZN(n9548) );
  NAND2_X1 U7579 ( .A1(n9547), .A2(n9548), .ZN(n9546) );
  INV_X1 U7580 ( .A(n5921), .ZN(n5922) );
  NAND2_X1 U7581 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U7582 ( .A1(n9546), .A2(n5924), .ZN(n7307) );
  INV_X1 U7583 ( .A(n7307), .ZN(n5932) );
  NAND2_X1 U7584 ( .A1(n7313), .A2(n4545), .ZN(n5926) );
  NAND2_X1 U7585 ( .A1(n9983), .A2(n5957), .ZN(n5925) );
  NAND2_X1 U7586 ( .A1(n5926), .A2(n5925), .ZN(n5928) );
  XNOR2_X1 U7587 ( .A(n5928), .B(n6115), .ZN(n5934) );
  NAND2_X1 U7588 ( .A1(n7313), .A2(n5957), .ZN(n5930) );
  NAND2_X1 U7589 ( .A1(n9983), .A2(n4543), .ZN(n5929) );
  NAND2_X1 U7590 ( .A1(n5930), .A2(n5929), .ZN(n5933) );
  XNOR2_X1 U7591 ( .A(n5934), .B(n5933), .ZN(n7306) );
  NAND2_X1 U7592 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  NAND2_X1 U7593 ( .A1(n7308), .A2(n5935), .ZN(n7580) );
  NAND2_X1 U7594 ( .A1(n9690), .A2(n4546), .ZN(n5938) );
  NAND2_X1 U7595 ( .A1(n9982), .A2(n5957), .ZN(n5937) );
  NAND2_X1 U7596 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  XNOR2_X1 U7597 ( .A(n5939), .B(n6074), .ZN(n5951) );
  NAND2_X1 U7598 ( .A1(n9690), .A2(n5957), .ZN(n5941) );
  NAND2_X1 U7599 ( .A1(n9982), .A2(n4543), .ZN(n5940) );
  AND2_X1 U7600 ( .A1(n5941), .A2(n5940), .ZN(n7582) );
  NAND2_X1 U7601 ( .A1(n5951), .A2(n7582), .ZN(n5942) );
  NAND2_X1 U7602 ( .A1(n7580), .A2(n5942), .ZN(n5955) );
  NAND2_X1 U7603 ( .A1(n9698), .A2(n4546), .ZN(n5944) );
  NAND2_X1 U7604 ( .A1(n9981), .A2(n5957), .ZN(n5943) );
  NAND2_X1 U7605 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  XNOR2_X1 U7606 ( .A(n5945), .B(n6074), .ZN(n5946) );
  AOI22_X1 U7607 ( .A1(n9698), .A2(n5957), .B1(n9981), .B2(n4543), .ZN(n5947)
         );
  NAND2_X1 U7608 ( .A1(n5946), .A2(n5947), .ZN(n5956) );
  INV_X1 U7609 ( .A(n5946), .ZN(n5949) );
  INV_X1 U7610 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7611 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7612 ( .A1(n5956), .A2(n5950), .ZN(n10533) );
  INV_X1 U7613 ( .A(n5951), .ZN(n7579) );
  INV_X1 U7614 ( .A(n7582), .ZN(n5952) );
  AND2_X1 U7615 ( .A1(n7579), .A2(n5952), .ZN(n5953) );
  NOR2_X1 U7616 ( .A1(n10533), .A2(n5953), .ZN(n5954) );
  NAND2_X1 U7617 ( .A1(n5955), .A2(n5954), .ZN(n10536) );
  NAND2_X1 U7618 ( .A1(n10536), .A2(n5956), .ZN(n7538) );
  NAND2_X1 U7619 ( .A1(n10607), .A2(n4546), .ZN(n5959) );
  NAND2_X1 U7620 ( .A1(n9980), .A2(n5957), .ZN(n5958) );
  NAND2_X1 U7621 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  XNOR2_X1 U7622 ( .A(n5960), .B(n6110), .ZN(n5961) );
  AOI22_X1 U7623 ( .A1(n10607), .A2(n5957), .B1(n4543), .B2(n9980), .ZN(n5962)
         );
  XNOR2_X1 U7624 ( .A(n5961), .B(n5962), .ZN(n7539) );
  NAND2_X1 U7625 ( .A1(n7538), .A2(n7539), .ZN(n7537) );
  INV_X1 U7626 ( .A(n5961), .ZN(n5963) );
  NAND2_X1 U7627 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  NAND2_X1 U7628 ( .A1(n7950), .A2(n4546), .ZN(n5966) );
  NAND2_X1 U7629 ( .A1(n9979), .A2(n5957), .ZN(n5965) );
  NAND2_X1 U7630 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7631 ( .A(n5967), .B(n6110), .ZN(n5969) );
  XNOR2_X2 U7632 ( .A(n5971), .B(n5969), .ZN(n10519) );
  AND2_X1 U7633 ( .A1(n9979), .A2(n4543), .ZN(n5968) );
  AOI21_X1 U7634 ( .B1(n7950), .B2(n5957), .A(n5968), .ZN(n10520) );
  NAND2_X2 U7635 ( .A1(n10519), .A2(n10520), .ZN(n7737) );
  INV_X1 U7636 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7637 ( .A1(n5971), .A2(n5970), .ZN(n7739) );
  NAND2_X1 U7638 ( .A1(n4559), .A2(n4546), .ZN(n5973) );
  NAND2_X1 U7639 ( .A1(n9978), .A2(n5957), .ZN(n5972) );
  NAND2_X1 U7640 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  XNOR2_X1 U7641 ( .A(n5974), .B(n6115), .ZN(n5979) );
  AND2_X1 U7642 ( .A1(n9978), .A2(n4543), .ZN(n5975) );
  AOI21_X1 U7643 ( .B1(n4559), .B2(n5957), .A(n5975), .ZN(n5977) );
  XNOR2_X1 U7644 ( .A(n5979), .B(n5977), .ZN(n7738) );
  AND2_X1 U7645 ( .A1(n7739), .A2(n7738), .ZN(n5976) );
  INV_X1 U7646 ( .A(n5977), .ZN(n5978) );
  NAND2_X1 U7647 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND2_X1 U7648 ( .A1(n10486), .A2(n4546), .ZN(n5982) );
  NAND2_X1 U7649 ( .A1(n9977), .A2(n5957), .ZN(n5981) );
  NAND2_X1 U7650 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  XNOR2_X1 U7651 ( .A(n5983), .B(n6115), .ZN(n5984) );
  NAND2_X1 U7652 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7653 ( .A1(n10486), .A2(n5957), .ZN(n5988) );
  NAND2_X1 U7654 ( .A1(n9977), .A2(n4543), .ZN(n5987) );
  NAND2_X1 U7655 ( .A1(n5988), .A2(n5987), .ZN(n10482) );
  INV_X1 U7656 ( .A(n10482), .ZN(n5989) );
  NAND2_X1 U7657 ( .A1(n10625), .A2(n4546), .ZN(n5991) );
  NAND2_X1 U7658 ( .A1(n9976), .A2(n5957), .ZN(n5990) );
  NAND2_X1 U7659 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  XNOR2_X1 U7660 ( .A(n5992), .B(n6074), .ZN(n5994) );
  AND2_X1 U7661 ( .A1(n9976), .A2(n4543), .ZN(n5993) );
  AOI21_X1 U7662 ( .B1(n10625), .B2(n5957), .A(n5993), .ZN(n5995) );
  NAND2_X1 U7663 ( .A1(n5994), .A2(n5995), .ZN(n10497) );
  INV_X1 U7664 ( .A(n5994), .ZN(n5997) );
  INV_X1 U7665 ( .A(n5995), .ZN(n5996) );
  NAND2_X1 U7666 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  AND2_X1 U7667 ( .A1(n10497), .A2(n5998), .ZN(n10510) );
  NAND2_X1 U7668 ( .A1(n5999), .A2(n10510), .ZN(n10493) );
  NAND2_X1 U7669 ( .A1(n10493), .A2(n10497), .ZN(n6009) );
  NAND2_X1 U7670 ( .A1(n10503), .A2(n4546), .ZN(n6001) );
  NAND2_X1 U7671 ( .A1(n9975), .A2(n5957), .ZN(n6000) );
  NAND2_X1 U7672 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  XNOR2_X1 U7673 ( .A(n6002), .B(n6074), .ZN(n6004) );
  AND2_X1 U7674 ( .A1(n9975), .A2(n4543), .ZN(n6003) );
  AOI21_X1 U7675 ( .B1(n10503), .B2(n5957), .A(n6003), .ZN(n6005) );
  NAND2_X1 U7676 ( .A1(n6004), .A2(n6005), .ZN(n6010) );
  INV_X1 U7677 ( .A(n6004), .ZN(n6007) );
  INV_X1 U7678 ( .A(n6005), .ZN(n6006) );
  NAND2_X1 U7679 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  AND2_X1 U7680 ( .A1(n6010), .A2(n6008), .ZN(n10495) );
  NAND2_X1 U7681 ( .A1(n8456), .A2(n4546), .ZN(n6012) );
  NAND2_X1 U7682 ( .A1(n9974), .A2(n5957), .ZN(n6011) );
  NAND2_X1 U7683 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  XNOR2_X1 U7684 ( .A(n6013), .B(n6110), .ZN(n6015) );
  AND2_X1 U7685 ( .A1(n9974), .A2(n4543), .ZN(n6014) );
  AOI21_X1 U7686 ( .B1(n8456), .B2(n5957), .A(n6014), .ZN(n6016) );
  XNOR2_X1 U7687 ( .A(n6015), .B(n6016), .ZN(n9620) );
  INV_X1 U7688 ( .A(n6015), .ZN(n6017) );
  NAND2_X1 U7689 ( .A1(n9534), .A2(n4546), .ZN(n6019) );
  NAND2_X1 U7690 ( .A1(n9973), .A2(n5957), .ZN(n6018) );
  NAND2_X1 U7691 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  XNOR2_X1 U7692 ( .A(n6020), .B(n6074), .ZN(n6024) );
  NAND2_X1 U7693 ( .A1(n9534), .A2(n5957), .ZN(n6022) );
  NAND2_X1 U7694 ( .A1(n9973), .A2(n4543), .ZN(n6021) );
  NAND2_X1 U7695 ( .A1(n6022), .A2(n6021), .ZN(n9529) );
  NAND2_X1 U7696 ( .A1(n10454), .A2(n4546), .ZN(n6026) );
  NAND2_X1 U7697 ( .A1(n9972), .A2(n5957), .ZN(n6025) );
  NAND2_X1 U7698 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7699 ( .A(n6027), .B(n6115), .ZN(n6029) );
  AND2_X1 U7700 ( .A1(n9972), .A2(n4543), .ZN(n6028) );
  AOI21_X1 U7701 ( .B1(n10454), .B2(n5957), .A(n6028), .ZN(n9664) );
  NAND2_X1 U7702 ( .A1(n9663), .A2(n9664), .ZN(n6031) );
  NAND2_X1 U7703 ( .A1(n6031), .A2(n9662), .ZN(n9586) );
  NAND2_X1 U7704 ( .A1(n10384), .A2(n4546), .ZN(n6033) );
  NAND2_X1 U7705 ( .A1(n9971), .A2(n5957), .ZN(n6032) );
  NAND2_X1 U7706 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  XNOR2_X1 U7707 ( .A(n6034), .B(n6110), .ZN(n6037) );
  NAND2_X1 U7708 ( .A1(n10384), .A2(n5957), .ZN(n6036) );
  NAND2_X1 U7709 ( .A1(n9971), .A2(n4543), .ZN(n6035) );
  NAND2_X1 U7710 ( .A1(n6036), .A2(n6035), .ZN(n6038) );
  NAND2_X1 U7711 ( .A1(n6037), .A2(n6038), .ZN(n9588) );
  NAND2_X1 U7712 ( .A1(n9586), .A2(n9588), .ZN(n9585) );
  INV_X1 U7713 ( .A(n6037), .ZN(n6040) );
  INV_X1 U7714 ( .A(n6038), .ZN(n6039) );
  NAND2_X1 U7715 ( .A1(n6040), .A2(n6039), .ZN(n9587) );
  NAND2_X1 U7716 ( .A1(n9585), .A2(n9587), .ZN(n9595) );
  NAND2_X1 U7717 ( .A1(n10443), .A2(n6112), .ZN(n6042) );
  NAND2_X1 U7718 ( .A1(n9970), .A2(n5957), .ZN(n6041) );
  NAND2_X1 U7719 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  XNOR2_X1 U7720 ( .A(n6043), .B(n6115), .ZN(n6045) );
  AND2_X1 U7721 ( .A1(n9970), .A2(n4543), .ZN(n6044) );
  AOI21_X1 U7722 ( .B1(n10443), .B2(n5957), .A(n6044), .ZN(n6046) );
  XNOR2_X1 U7723 ( .A(n6045), .B(n6046), .ZN(n9596) );
  INV_X1 U7724 ( .A(n6045), .ZN(n6047) );
  NAND2_X1 U7725 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U7726 ( .A1(n10374), .A2(n6112), .ZN(n6050) );
  NAND2_X1 U7727 ( .A1(n9969), .A2(n5957), .ZN(n6049) );
  NAND2_X1 U7728 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7729 ( .A(n6051), .B(n6074), .ZN(n9644) );
  AND2_X1 U7730 ( .A1(n9969), .A2(n4543), .ZN(n6052) );
  AOI21_X1 U7731 ( .B1(n10374), .B2(n5957), .A(n6052), .ZN(n9643) );
  NAND2_X1 U7732 ( .A1(n10369), .A2(n4546), .ZN(n6054) );
  NAND2_X1 U7733 ( .A1(n9968), .A2(n5957), .ZN(n6053) );
  NAND2_X1 U7734 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7735 ( .A(n6055), .B(n6110), .ZN(n6057) );
  AND2_X1 U7736 ( .A1(n9968), .A2(n4543), .ZN(n6056) );
  AOI21_X1 U7737 ( .B1(n10369), .B2(n5957), .A(n6056), .ZN(n6058) );
  XNOR2_X1 U7738 ( .A(n6057), .B(n6058), .ZN(n9557) );
  INV_X1 U7739 ( .A(n6057), .ZN(n6059) );
  NAND2_X1 U7740 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7741 ( .A1(n10364), .A2(n6112), .ZN(n6062) );
  NAND2_X1 U7742 ( .A1(n9967), .A2(n5957), .ZN(n6061) );
  NAND2_X1 U7743 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  XNOR2_X1 U7744 ( .A(n6063), .B(n6074), .ZN(n9610) );
  AND2_X1 U7745 ( .A1(n9967), .A2(n4543), .ZN(n6064) );
  AOI21_X1 U7746 ( .B1(n10364), .B2(n5957), .A(n6064), .ZN(n9609) );
  AND2_X1 U7747 ( .A1(n9610), .A2(n9609), .ZN(n9567) );
  NAND2_X1 U7748 ( .A1(n10428), .A2(n4546), .ZN(n6066) );
  NAND2_X1 U7749 ( .A1(n9966), .A2(n5957), .ZN(n6065) );
  NAND2_X1 U7750 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  XNOR2_X1 U7751 ( .A(n6067), .B(n6074), .ZN(n6076) );
  AND2_X1 U7752 ( .A1(n9966), .A2(n4543), .ZN(n6068) );
  AOI21_X1 U7753 ( .B1(n10428), .B2(n5957), .A(n6068), .ZN(n6077) );
  NAND2_X1 U7754 ( .A1(n6076), .A2(n6077), .ZN(n9564) );
  INV_X1 U7755 ( .A(n9564), .ZN(n6071) );
  INV_X1 U7756 ( .A(n9610), .ZN(n6070) );
  INV_X1 U7757 ( .A(n9609), .ZN(n6069) );
  NAND2_X1 U7758 ( .A1(n6070), .A2(n6069), .ZN(n9568) );
  NAND2_X1 U7759 ( .A1(n10194), .A2(n6112), .ZN(n6073) );
  NAND2_X1 U7760 ( .A1(n9965), .A2(n5957), .ZN(n6072) );
  NAND2_X1 U7761 ( .A1(n6073), .A2(n6072), .ZN(n6075) );
  XNOR2_X1 U7762 ( .A(n6075), .B(n6074), .ZN(n6084) );
  INV_X1 U7763 ( .A(n6076), .ZN(n6079) );
  INV_X1 U7764 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7765 ( .A1(n6079), .A2(n6078), .ZN(n9565) );
  AND2_X1 U7766 ( .A1(n6084), .A2(n9565), .ZN(n6080) );
  OAI22_X1 U7767 ( .A1(n4942), .A2(n4551), .B1(n6082), .B2(n6081), .ZN(n9633)
         );
  NAND2_X1 U7768 ( .A1(n6083), .A2(n9565), .ZN(n6086) );
  INV_X1 U7769 ( .A(n6084), .ZN(n6085) );
  AOI22_X1 U7770 ( .A1(n10179), .A2(n4546), .B1(n5957), .B2(n9964), .ZN(n6087)
         );
  XNOR2_X1 U7771 ( .A(n6087), .B(n6115), .ZN(n6089) );
  AOI22_X1 U7772 ( .A1(n10179), .A2(n5957), .B1(n4543), .B2(n9964), .ZN(n6088)
         );
  XNOR2_X1 U7773 ( .A(n6089), .B(n6088), .ZN(n9539) );
  AOI22_X1 U7774 ( .A1(n10341), .A2(n5957), .B1(n4543), .B2(n9963), .ZN(n6093)
         );
  NAND2_X1 U7775 ( .A1(n10341), .A2(n4546), .ZN(n6091) );
  NAND2_X1 U7776 ( .A1(n9963), .A2(n5957), .ZN(n6090) );
  NAND2_X1 U7777 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7778 ( .A(n6092), .B(n6110), .ZN(n6095) );
  XOR2_X1 U7779 ( .A(n6093), .B(n6095), .Z(n9604) );
  INV_X1 U7780 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7781 ( .A1(n10411), .A2(n4546), .ZN(n6097) );
  NAND2_X1 U7782 ( .A1(n9962), .A2(n5957), .ZN(n6096) );
  NAND2_X1 U7783 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  XNOR2_X1 U7784 ( .A(n6098), .B(n6115), .ZN(n6099) );
  AOI22_X1 U7785 ( .A1(n10411), .A2(n5957), .B1(n4543), .B2(n9962), .ZN(n6100)
         );
  XNOR2_X1 U7786 ( .A(n6099), .B(n6100), .ZN(n9579) );
  INV_X1 U7787 ( .A(n6099), .ZN(n6101) );
  AOI22_X1 U7788 ( .A1(n10406), .A2(n5957), .B1(n4543), .B2(n9961), .ZN(n6104)
         );
  AOI22_X1 U7789 ( .A1(n10406), .A2(n6112), .B1(n5957), .B2(n9961), .ZN(n6102)
         );
  XNOR2_X1 U7790 ( .A(n6102), .B(n6110), .ZN(n6103) );
  XOR2_X1 U7791 ( .A(n6104), .B(n6103), .Z(n9654) );
  INV_X1 U7792 ( .A(n6103), .ZN(n6106) );
  INV_X1 U7793 ( .A(n6104), .ZN(n6105) );
  AND2_X1 U7794 ( .A1(n9960), .A2(n4543), .ZN(n6107) );
  AOI21_X1 U7795 ( .B1(n8479), .B2(n5957), .A(n6107), .ZN(n6125) );
  NAND2_X1 U7796 ( .A1(n8479), .A2(n4546), .ZN(n6109) );
  NAND2_X1 U7797 ( .A1(n9960), .A2(n5957), .ZN(n6108) );
  NAND2_X1 U7798 ( .A1(n6109), .A2(n6108), .ZN(n6111) );
  XNOR2_X1 U7799 ( .A(n6111), .B(n6110), .ZN(n6127) );
  XOR2_X1 U7800 ( .A(n6125), .B(n6127), .Z(n8471) );
  NAND2_X1 U7801 ( .A1(n10326), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7802 ( .A1(n9959), .A2(n5957), .ZN(n6113) );
  NAND2_X1 U7803 ( .A1(n6114), .A2(n6113), .ZN(n6116) );
  XNOR2_X1 U7804 ( .A(n6116), .B(n6115), .ZN(n6119) );
  AOI22_X1 U7805 ( .A1(n10326), .A2(n5957), .B1(n4543), .B2(n9959), .ZN(n6118)
         );
  XNOR2_X1 U7806 ( .A(n6119), .B(n6118), .ZN(n6128) );
  INV_X1 U7807 ( .A(n6128), .ZN(n6140) );
  NAND3_X1 U7808 ( .A1(n6856), .A2(n10459), .A3(n6120), .ZN(n7038) );
  INV_X1 U7809 ( .A(n9932), .ZN(n6123) );
  AND2_X1 U7810 ( .A1(n10617), .A2(n6123), .ZN(n6124) );
  INV_X1 U7811 ( .A(n6125), .ZN(n6126) );
  OR2_X1 U7812 ( .A1(n6127), .A2(n6126), .ZN(n6139) );
  NAND3_X1 U7813 ( .A1(n6140), .A2(n10527), .A3(n6139), .ZN(n6145) );
  AOI22_X1 U7814 ( .A1(n9960), .A2(n9666), .B1(n9667), .B2(n9958), .ZN(n10117)
         );
  INV_X1 U7815 ( .A(n4549), .ZN(n9936) );
  NAND2_X1 U7816 ( .A1(n7038), .A2(n9936), .ZN(n6133) );
  NAND3_X1 U7817 ( .A1(n6133), .A2(n7937), .A3(n6685), .ZN(n6136) );
  NAND2_X1 U7818 ( .A1(n7038), .A2(n10617), .ZN(n6135) );
  NAND2_X1 U7819 ( .A1(n6135), .A2(n6134), .ZN(n7037) );
  OR2_X1 U7820 ( .A1(n6136), .A2(n7037), .ZN(n6137) );
  AOI22_X1 U7821 ( .A1(n10122), .A2(n9638), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6138) );
  OAI21_X1 U7822 ( .B1(n10117), .B2(n10492), .A(n6138), .ZN(n6142) );
  NOR3_X1 U7823 ( .A1(n6140), .A2(n10535), .A3(n6139), .ZN(n6141) );
  AOI211_X1 U7824 ( .C1(n10326), .C2(n10515), .A(n6142), .B(n6141), .ZN(n6143)
         );
  OAI211_X1 U7825 ( .C1(n6146), .C2(n6145), .A(n6144), .B(n6143), .ZN(P1_U3220) );
  INV_X1 U7826 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6148) );
  INV_X1 U7827 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7828 ( .A1(n6148), .A2(n6147), .ZN(n6331) );
  INV_X1 U7829 ( .A(n6331), .ZN(n6150) );
  INV_X1 U7830 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7831 ( .A1(n6150), .A2(n6149), .ZN(n6344) );
  INV_X1 U7832 ( .A(n6357), .ZN(n6152) );
  INV_X1 U7833 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7834 ( .A1(n6152), .A2(n6151), .ZN(n6368) );
  INV_X1 U7835 ( .A(n6388), .ZN(n6154) );
  NAND2_X1 U7836 ( .A1(n6154), .A2(n6153), .ZN(n6401) );
  OR2_X2 U7837 ( .A1(n6401), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6411) );
  OR2_X2 U7838 ( .A1(n6411), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6427) );
  INV_X1 U7839 ( .A(n6438), .ZN(n6157) );
  OR2_X2 U7840 ( .A1(n6452), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6467) );
  INV_X1 U7841 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6164) );
  OR2_X2 U7842 ( .A1(n6510), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6519) );
  OR2_X2 U7843 ( .A1(n6519), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6521) );
  INV_X1 U7844 ( .A(n6521), .ZN(n6167) );
  INV_X1 U7845 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6166) );
  INV_X1 U7846 ( .A(n6531), .ZN(n6169) );
  INV_X1 U7847 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6168) );
  OR2_X2 U7848 ( .A1(n6533), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U7849 ( .A1(n6533), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7850 ( .A1(n6544), .A2(n6170), .ZN(n8890) );
  INV_X1 U7851 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6171) );
  NOR2_X1 U7852 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6176) );
  NOR2_X1 U7853 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6175) );
  NOR2_X1 U7854 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6174) );
  NAND4_X1 U7855 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n6179)
         );
  NAND4_X1 U7856 ( .A1(n6177), .A2(n6230), .A3(n6229), .A4(n4726), .ZN(n6178)
         );
  NOR2_X1 U7857 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n6182) );
  NOR2_X1 U7858 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n6181) );
  NOR2_X1 U7859 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6180) );
  INV_X1 U7860 ( .A(n6187), .ZN(n6184) );
  NOR2_X1 U7861 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6183) );
  NAND2_X1 U7862 ( .A1(n6184), .A2(n6183), .ZN(n9520) );
  NAND2_X1 U7863 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n6188) );
  NAND2_X1 U7864 ( .A1(n6200), .A2(n6188), .ZN(n6189) );
  XNOR2_X2 U7865 ( .A(n6189), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6192) );
  INV_X1 U7866 ( .A(n6192), .ZN(n6190) );
  NAND2_X1 U7867 ( .A1(n8890), .A2(n6565), .ZN(n6198) );
  INV_X1 U7868 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9479) );
  INV_X2 U7869 ( .A(n6270), .ZN(n6566) );
  NAND2_X1 U7870 ( .A1(n6566), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7871 ( .A1(n6557), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7872 ( .C1(n4557), .C2(n9479), .A(n6195), .B(n6194), .ZN(n6196)
         );
  INV_X1 U7873 ( .A(n6196), .ZN(n6197) );
  NAND2_X1 U7874 ( .A1(n6201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7875 ( .A1(n6277), .A2(n8171), .ZN(n6563) );
  NAND2_X1 U7876 ( .A1(n8097), .A2(n4541), .ZN(n6205) );
  NAND2_X4 U7877 ( .A1(n6277), .A2(n5330), .ZN(n6276) );
  OR2_X1 U7878 ( .A1(n6276), .A2(n8100), .ZN(n6204) );
  NAND2_X1 U7879 ( .A1(n8033), .A2(n4541), .ZN(n6207) );
  OR2_X1 U7880 ( .A1(n6276), .A2(n8469), .ZN(n6206) );
  NAND2_X1 U7881 ( .A1(n6521), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7882 ( .A1(n6531), .A2(n6208), .ZN(n8910) );
  NAND2_X1 U7883 ( .A1(n8910), .A2(n6565), .ZN(n6214) );
  INV_X1 U7884 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6211) );
  BUF_X4 U7885 ( .A(n6267), .Z(n8174) );
  NAND2_X1 U7886 ( .A1(n8174), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7887 ( .A1(n6566), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6209) );
  OAI211_X1 U7888 ( .C1(n6569), .C2(n6211), .A(n6210), .B(n6209), .ZN(n6212)
         );
  INV_X1 U7889 ( .A(n6212), .ZN(n6213) );
  NAND2_X1 U7890 ( .A1(n6214), .A2(n6213), .ZN(n8655) );
  NAND2_X1 U7891 ( .A1(n7694), .A2(n4541), .ZN(n6216) );
  INV_X1 U7892 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7695) );
  OR2_X1 U7893 ( .A1(n6276), .A2(n7695), .ZN(n6215) );
  NAND2_X1 U7894 ( .A1(n6222), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7895 ( .A1(n6501), .A2(n6217), .ZN(n8954) );
  INV_X1 U7896 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U7897 ( .A1(n6557), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7898 ( .A1(n8174), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7899 ( .C1(n6588), .C2(n9175), .A(n6219), .B(n6218), .ZN(n6220)
         );
  INV_X1 U7900 ( .A(n8964), .ZN(n8659) );
  NAND2_X1 U7901 ( .A1(n6248), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7902 ( .A1(n6222), .A2(n6221), .ZN(n8968) );
  NAND2_X1 U7903 ( .A1(n8968), .A2(n6565), .ZN(n6228) );
  INV_X1 U7904 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7905 ( .A1(n6566), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7906 ( .A1(n8174), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6223) );
  OAI211_X1 U7907 ( .C1(n6225), .C2(n6569), .A(n6224), .B(n6223), .ZN(n6226)
         );
  INV_X1 U7908 ( .A(n6226), .ZN(n6227) );
  NAND2_X1 U7909 ( .A1(n6228), .A2(n6227), .ZN(n8977) );
  NAND2_X1 U7910 ( .A1(n7548), .A2(n4541), .ZN(n6240) );
  NAND2_X1 U7911 ( .A1(n6380), .A2(n6230), .ZN(n6383) );
  NAND2_X1 U7912 ( .A1(n9220), .A2(n6231), .ZN(n6232) );
  NAND2_X1 U7913 ( .A1(n6243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  XNOR2_X1 U7914 ( .A(n6238), .B(n6237), .ZN(n6622) );
  INV_X2 U7915 ( .A(n6276), .ZN(n6486) );
  AOI22_X1 U7916 ( .A1(n6898), .A2(n4547), .B1(n6486), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7917 ( .A1(n6240), .A2(n6239), .ZN(n8967) );
  NAND2_X1 U7918 ( .A1(n7334), .A2(n4541), .ZN(n6246) );
  INV_X1 U7919 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U7920 ( .A1(n6242), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6244) );
  AND2_X1 U7921 ( .A1(n6244), .A2(n6243), .ZN(n8833) );
  AOI22_X1 U7922 ( .A1(n8833), .A2(n4547), .B1(n6486), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7923 ( .A1(n6246), .A2(n6245), .ZN(n8492) );
  NAND2_X1 U7924 ( .A1(n6492), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7925 ( .A1(n6248), .A2(n6247), .ZN(n8983) );
  NAND2_X1 U7926 ( .A1(n8983), .A2(n6565), .ZN(n6253) );
  INV_X1 U7927 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U7928 ( .A1(n6566), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7929 ( .A1(n8174), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6249) );
  OAI211_X1 U7930 ( .C1(n8832), .C2(n6569), .A(n6250), .B(n6249), .ZN(n6251)
         );
  INV_X1 U7931 ( .A(n6251), .ZN(n6252) );
  NAND2_X1 U7932 ( .A1(n6253), .A2(n6252), .ZN(n8660) );
  INV_X1 U7933 ( .A(n8492), .ZN(n9071) );
  INV_X1 U7934 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7371) );
  OR2_X1 U7935 ( .A1(n6548), .A2(n7371), .ZN(n6259) );
  INV_X1 U7936 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6254) );
  INV_X1 U7937 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6939) );
  OR2_X1 U7938 ( .A1(n6403), .A2(n6939), .ZN(n6257) );
  OR2_X1 U7939 ( .A1(n6276), .A2(n6718), .ZN(n6265) );
  OR2_X1 U7940 ( .A1(n8172), .A2(n4548), .ZN(n6264) );
  NAND2_X1 U7941 ( .A1(n8674), .A2(n8268), .ZN(n6266) );
  AND2_X2 U7942 ( .A1(n6290), .A2(n6266), .ZN(n8274) );
  NAND2_X1 U7943 ( .A1(n6267), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6273) );
  INV_X1 U7944 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7376) );
  INV_X1 U7945 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6269) );
  INV_X1 U7946 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7375) );
  OR2_X1 U7947 ( .A1(n6563), .A2(n6275), .ZN(n6279) );
  OR2_X1 U7948 ( .A1(n6276), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6278) );
  AND3_X2 U7949 ( .A1(n6279), .A2(n6278), .A3(n4623), .ZN(n7378) );
  NAND2_X2 U7950 ( .A1(n6288), .A2(n7378), .ZN(n8263) );
  NAND2_X1 U7951 ( .A1(n8174), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6286) );
  INV_X1 U7952 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6281) );
  OR2_X1 U7953 ( .A1(n6588), .A2(n6281), .ZN(n6285) );
  INV_X1 U7954 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6990) );
  OR2_X1 U7955 ( .A1(n6403), .A2(n6990), .ZN(n6284) );
  INV_X1 U7956 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6282) );
  OR2_X1 U7957 ( .A1(n6548), .A2(n6282), .ZN(n6283) );
  NAND2_X1 U7958 ( .A1(n8171), .A2(SI_0_), .ZN(n6287) );
  XNOR2_X1 U7959 ( .A(n6287), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9525) );
  MUX2_X1 U7960 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9525), .S(n8172), .Z(n7344) );
  NAND2_X1 U7961 ( .A1(n8677), .A2(n7344), .ZN(n7072) );
  INV_X1 U7962 ( .A(n7378), .ZN(n7079) );
  NAND2_X1 U7963 ( .A1(n7079), .A2(n8675), .ZN(n6289) );
  INV_X1 U7964 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6291) );
  OR2_X1 U7965 ( .A1(n6588), .A2(n6291), .ZN(n6296) );
  NAND2_X1 U7966 ( .A1(n8174), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6295) );
  OR2_X1 U7967 ( .A1(n6403), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6294) );
  INV_X1 U7968 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6292) );
  OR2_X1 U7969 ( .A1(n6548), .A2(n6292), .ZN(n6293) );
  NAND4_X2 U7970 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n8673)
         );
  NAND2_X1 U7971 ( .A1(n6297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6298) );
  XNOR2_X1 U7972 ( .A(n6298), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7973 ( .A1(n6486), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6487), .B2(
        n6827), .ZN(n6302) );
  NAND2_X1 U7974 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NAND2_X1 U7975 ( .A1(n7697), .A2(n8673), .ZN(n8278) );
  AND2_X1 U7976 ( .A1(n8286), .A2(n8278), .ZN(n8189) );
  INV_X1 U7977 ( .A(n8189), .ZN(n7129) );
  NAND2_X1 U7978 ( .A1(n7130), .A2(n7129), .ZN(n7128) );
  NAND2_X1 U7979 ( .A1(n6304), .A2(n7697), .ZN(n6305) );
  NAND2_X1 U7980 ( .A1(n6566), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6312) );
  INV_X1 U7981 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7982 ( .A1(n4557), .A2(n6306), .ZN(n6311) );
  NAND2_X1 U7983 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6307) );
  AND2_X1 U7984 ( .A1(n6331), .A2(n6307), .ZN(n7897) );
  OR2_X1 U7985 ( .A1(n6403), .A2(n7897), .ZN(n6310) );
  INV_X1 U7986 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6308) );
  OR2_X1 U7987 ( .A1(n6548), .A2(n6308), .ZN(n6309) );
  NAND2_X1 U7988 ( .A1(n6313), .A2(n4541), .ZN(n6320) );
  OR2_X1 U7989 ( .A1(n6297), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7990 ( .A1(n6315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6314) );
  MUX2_X1 U7991 ( .A(n6314), .B(P2_IR_REG_31__SCAN_IN), .S(n6316), .Z(n6318)
         );
  INV_X1 U7992 ( .A(n6315), .ZN(n6317) );
  NAND2_X1 U7993 ( .A1(n6317), .A2(n6316), .ZN(n6326) );
  NAND2_X1 U7994 ( .A1(n6318), .A2(n6326), .ZN(n6880) );
  INV_X1 U7995 ( .A(n6880), .ZN(n6866) );
  AOI22_X1 U7996 ( .A1(n6486), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n4547), .B2(
        n6866), .ZN(n6319) );
  NAND2_X1 U7997 ( .A1(n6320), .A2(n6319), .ZN(n7895) );
  NAND2_X1 U7998 ( .A1(n8672), .A2(n7895), .ZN(n6321) );
  NAND2_X1 U7999 ( .A1(n7065), .A2(n6321), .ZN(n6323) );
  OR2_X1 U8000 ( .A1(n8672), .A2(n7895), .ZN(n6322) );
  NAND2_X1 U8001 ( .A1(n6323), .A2(n6322), .ZN(n7265) );
  NAND2_X1 U8002 ( .A1(n6326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6325) );
  MUX2_X1 U8003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6325), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6329) );
  INV_X1 U8004 ( .A(n6326), .ZN(n6328) );
  NAND2_X1 U8005 ( .A1(n6328), .A2(n6327), .ZN(n6340) );
  AOI22_X1 U8006 ( .A1(n6486), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n4547), .B2(
        n6869), .ZN(n6330) );
  NAND2_X1 U8007 ( .A1(n8174), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6337) );
  OR2_X1 U8008 ( .A1(n6588), .A2(n8687), .ZN(n6336) );
  NAND2_X1 U8009 ( .A1(n6331), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6332) );
  AND2_X1 U8010 ( .A1(n6344), .A2(n6332), .ZN(n7383) );
  OR2_X1 U8011 ( .A1(n6403), .A2(n7383), .ZN(n6335) );
  BUF_X1 U8012 ( .A(n6548), .Z(n6569) );
  INV_X1 U8013 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6333) );
  OR2_X1 U8014 ( .A1(n6569), .A2(n6333), .ZN(n6334) );
  NAND4_X1 U8015 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n8671)
         );
  NAND2_X1 U8016 ( .A1(n7385), .A2(n7324), .ZN(n7209) );
  AND2_X1 U8017 ( .A1(n8281), .A2(n7209), .ZN(n8194) );
  NAND2_X1 U8018 ( .A1(n7265), .A2(n7266), .ZN(n6339) );
  OR2_X1 U8019 ( .A1(n7385), .A2(n8671), .ZN(n6338) );
  NAND2_X1 U8020 ( .A1(n6732), .A2(n4541), .ZN(n6343) );
  NAND2_X1 U8021 ( .A1(n6340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  AOI22_X1 U8022 ( .A1(n6486), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4547), .B2(
        n7148), .ZN(n6342) );
  NAND2_X1 U8023 ( .A1(n6343), .A2(n6342), .ZN(n7660) );
  NAND2_X1 U8024 ( .A1(n8174), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6349) );
  INV_X1 U8025 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7657) );
  OR2_X1 U8026 ( .A1(n6548), .A2(n7657), .ZN(n6348) );
  NAND2_X1 U8027 ( .A1(n6344), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6345) );
  AND2_X1 U8028 ( .A1(n6357), .A2(n6345), .ZN(n7658) );
  OR2_X1 U8029 ( .A1(n6403), .A2(n7658), .ZN(n6347) );
  OR2_X1 U8030 ( .A1(n6588), .A2(n7213), .ZN(n6346) );
  NAND4_X1 U8031 ( .A1(n6349), .A2(n6348), .A3(n6347), .A4(n6346), .ZN(n8670)
         );
  NOR2_X1 U8032 ( .A1(n7660), .A2(n8670), .ZN(n6351) );
  NAND2_X1 U8033 ( .A1(n7660), .A2(n8670), .ZN(n6350) );
  INV_X1 U8034 ( .A(n7407), .ZN(n6365) );
  NAND2_X1 U8035 ( .A1(n6739), .A2(n4541), .ZN(n6355) );
  NAND2_X1 U8036 ( .A1(n6352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6353) );
  XNOR2_X1 U8037 ( .A(n6353), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7151) );
  AOI22_X1 U8038 ( .A1(n6486), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4547), .B2(
        n7151), .ZN(n6354) );
  NAND2_X1 U8039 ( .A1(n6355), .A2(n6354), .ZN(n8248) );
  NAND2_X1 U8040 ( .A1(n6566), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6362) );
  INV_X1 U8041 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6356) );
  OR2_X1 U8042 ( .A1(n4557), .A2(n6356), .ZN(n6361) );
  OR2_X1 U8043 ( .A1(n6548), .A2(n4753), .ZN(n6360) );
  NAND2_X1 U8044 ( .A1(n6357), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6358) );
  AND2_X1 U8045 ( .A1(n6368), .A2(n6358), .ZN(n7550) );
  OR2_X1 U8046 ( .A1(n6403), .A2(n7550), .ZN(n6359) );
  OR2_X1 U8047 ( .A1(n8248), .A2(n8669), .ZN(n6366) );
  NAND2_X1 U8048 ( .A1(n8248), .A2(n8669), .ZN(n6363) );
  NAND2_X1 U8049 ( .A1(n6366), .A2(n6363), .ZN(n8298) );
  NAND2_X1 U8050 ( .A1(n6566), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6373) );
  INV_X1 U8051 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6367) );
  OR2_X1 U8052 ( .A1(n4557), .A2(n6367), .ZN(n6372) );
  NAND2_X1 U8053 ( .A1(n6368), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6369) );
  AND2_X1 U8054 ( .A1(n6388), .A2(n6369), .ZN(n7667) );
  OR2_X1 U8055 ( .A1(n6403), .A2(n7667), .ZN(n6371) );
  INV_X1 U8056 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7666) );
  OR2_X1 U8057 ( .A1(n6569), .A2(n7666), .ZN(n6370) );
  NAND4_X1 U8058 ( .A1(n6373), .A2(n6372), .A3(n6371), .A4(n6370), .ZN(n8668)
         );
  NAND2_X1 U8059 ( .A1(n6743), .A2(n4541), .ZN(n6378) );
  NOR2_X1 U8060 ( .A1(n6374), .A2(n9518), .ZN(n6375) );
  MUX2_X1 U8061 ( .A(n9518), .B(n6375), .S(P2_IR_REG_8__SCAN_IN), .Z(n6376) );
  NOR2_X1 U8062 ( .A1(n6376), .A2(n6380), .ZN(n7228) );
  AOI22_X1 U8063 ( .A1(n6486), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4547), .B2(
        n7228), .ZN(n6377) );
  INV_X1 U8064 ( .A(n7669), .ZN(n7458) );
  NAND2_X1 U8065 ( .A1(n7455), .A2(n7633), .ZN(n6379) );
  NAND2_X1 U8066 ( .A1(n6750), .A2(n4541), .ZN(n6386) );
  NOR2_X1 U8067 ( .A1(n6380), .A2(n9518), .ZN(n6381) );
  MUX2_X1 U8068 ( .A(n9518), .B(n6381), .S(P2_IR_REG_9__SCAN_IN), .Z(n6382) );
  INV_X1 U8069 ( .A(n6382), .ZN(n6384) );
  AOI22_X1 U8070 ( .A1(n6486), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4547), .B2(
        n7613), .ZN(n6385) );
  NAND2_X1 U8071 ( .A1(n6386), .A2(n6385), .ZN(n7637) );
  NAND2_X1 U8072 ( .A1(n8174), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6394) );
  INV_X1 U8073 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6387) );
  OR2_X1 U8074 ( .A1(n6588), .A2(n6387), .ZN(n6393) );
  NAND2_X1 U8075 ( .A1(n6388), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6389) );
  AND2_X1 U8076 ( .A1(n6401), .A2(n6389), .ZN(n7640) );
  OR2_X1 U8077 ( .A1(n6403), .A2(n7640), .ZN(n6392) );
  INV_X1 U8078 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6390) );
  OR2_X1 U8079 ( .A1(n6548), .A2(n6390), .ZN(n6391) );
  NAND4_X1 U8080 ( .A1(n6394), .A2(n6393), .A3(n6392), .A4(n6391), .ZN(n8667)
         );
  NAND2_X1 U8081 ( .A1(n7637), .A2(n8667), .ZN(n6395) );
  OR2_X1 U8082 ( .A1(n7637), .A2(n8667), .ZN(n6396) );
  NAND2_X1 U8083 ( .A1(n6397), .A2(n6396), .ZN(n7571) );
  NAND2_X1 U8084 ( .A1(n6753), .A2(n4541), .ZN(n6400) );
  NAND2_X1 U8085 ( .A1(n6383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6398) );
  XNOR2_X1 U8086 ( .A(n6398), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7627) );
  AOI22_X1 U8087 ( .A1(n6486), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4547), .B2(
        n7627), .ZN(n6399) );
  NAND2_X1 U8088 ( .A1(n6400), .A2(n6399), .ZN(n7891) );
  NAND2_X1 U8089 ( .A1(n8174), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6407) );
  INV_X1 U8090 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7607) );
  OR2_X1 U8091 ( .A1(n6588), .A2(n7607), .ZN(n6406) );
  NAND2_X1 U8092 ( .A1(n6401), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6402) );
  AND2_X1 U8093 ( .A1(n6411), .A2(n6402), .ZN(n7889) );
  OR2_X1 U8094 ( .A1(n6403), .A2(n7889), .ZN(n6405) );
  INV_X1 U8095 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7615) );
  OR2_X1 U8096 ( .A1(n6548), .A2(n7615), .ZN(n6404) );
  NAND4_X1 U8097 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n8666)
         );
  NAND2_X1 U8098 ( .A1(n7891), .A2(n8666), .ZN(n6408) );
  NAND2_X1 U8099 ( .A1(n7571), .A2(n6408), .ZN(n6410) );
  OR2_X1 U8100 ( .A1(n7891), .A2(n8666), .ZN(n6409) );
  NAND2_X1 U8101 ( .A1(n6411), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U8102 ( .A1(n6427), .A2(n6412), .ZN(n7967) );
  NAND2_X1 U8103 ( .A1(n6565), .A2(n7967), .ZN(n6419) );
  INV_X1 U8104 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6413) );
  OR2_X1 U8105 ( .A1(n4557), .A2(n6413), .ZN(n6418) );
  INV_X1 U8106 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6414) );
  OR2_X1 U8107 ( .A1(n6588), .A2(n6414), .ZN(n6417) );
  INV_X1 U8108 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6415) );
  OR2_X1 U8109 ( .A1(n6569), .A2(n6415), .ZN(n6416) );
  NAND4_X1 U8110 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n8665)
         );
  NAND2_X1 U8111 ( .A1(n6817), .A2(n4541), .ZN(n6422) );
  OAI21_X1 U8112 ( .B1(n6383), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6420) );
  XNOR2_X1 U8113 ( .A(n6420), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7825) );
  AOI22_X1 U8114 ( .A1(n6486), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4547), .B2(
        n7825), .ZN(n6421) );
  NAND2_X1 U8115 ( .A1(n6422), .A2(n6421), .ZN(n7726) );
  NAND2_X1 U8116 ( .A1(n6892), .A2(n4541), .ZN(n6426) );
  OR2_X1 U8117 ( .A1(n6423), .A2(n9518), .ZN(n6424) );
  XNOR2_X1 U8118 ( .A(n6424), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7829) );
  AOI22_X1 U8119 ( .A1(n6486), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7829), .B2(
        n4547), .ZN(n6425) );
  NAND2_X1 U8120 ( .A1(n6426), .A2(n6425), .ZN(n8030) );
  NAND2_X1 U8121 ( .A1(n6427), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8122 ( .A1(n6438), .A2(n6428), .ZN(n8024) );
  NAND2_X1 U8123 ( .A1(n6565), .A2(n8024), .ZN(n6433) );
  INV_X1 U8124 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7828) );
  OR2_X1 U8125 ( .A1(n6588), .A2(n7828), .ZN(n6432) );
  INV_X1 U8126 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6429) );
  OR2_X1 U8127 ( .A1(n4557), .A2(n6429), .ZN(n6431) );
  INV_X1 U8128 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7811) );
  OR2_X1 U8129 ( .A1(n6548), .A2(n7811), .ZN(n6430) );
  NAND4_X1 U8130 ( .A1(n6433), .A2(n6432), .A3(n6431), .A4(n6430), .ZN(n8664)
         );
  AND2_X1 U8131 ( .A1(n8030), .A2(n8664), .ZN(n6434) );
  NAND2_X1 U8132 ( .A1(n6940), .A2(n4541), .ZN(n6437) );
  NAND2_X1 U8133 ( .A1(n6435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U8134 ( .A(n6447), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8713) );
  AOI22_X1 U8135 ( .A1(n8713), .A2(n4547), .B1(n6486), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8136 ( .A1(n6438), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8137 ( .A1(n6452), .A2(n6439), .ZN(n8093) );
  NAND2_X1 U8138 ( .A1(n8093), .A2(n6565), .ZN(n6443) );
  INV_X1 U8139 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9402) );
  OR2_X1 U8140 ( .A1(n4557), .A2(n9402), .ZN(n6442) );
  INV_X1 U8141 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7986) );
  OR2_X1 U8142 ( .A1(n6548), .A2(n7986), .ZN(n6441) );
  INV_X1 U8143 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8010) );
  OR2_X1 U8144 ( .A1(n6588), .A2(n8010), .ZN(n6440) );
  NAND4_X1 U8145 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n8663)
         );
  XNOR2_X1 U8146 ( .A(n8318), .B(n8663), .ZN(n8205) );
  INV_X1 U8147 ( .A(n8205), .ZN(n7945) );
  NAND2_X1 U8148 ( .A1(n7943), .A2(n7945), .ZN(n6445) );
  NOR2_X1 U8149 ( .A1(n8318), .A2(n8663), .ZN(n8316) );
  INV_X1 U8150 ( .A(n8316), .ZN(n6444) );
  NAND2_X1 U8151 ( .A1(n7179), .A2(n4541), .ZN(n6451) );
  NAND2_X1 U8152 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  NAND2_X1 U8153 ( .A1(n6448), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6462) );
  OAI22_X1 U8154 ( .A1(n8732), .A2(n8172), .B1(n6276), .B2(n7181), .ZN(n6449)
         );
  INV_X1 U8155 ( .A(n6449), .ZN(n6450) );
  INV_X1 U8156 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U8157 ( .A1(n6452), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U8158 ( .A1(n6467), .A2(n6453), .ZN(n8115) );
  NAND2_X1 U8159 ( .A1(n8115), .A2(n6565), .ZN(n6457) );
  INV_X1 U8160 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8046) );
  OR2_X1 U8161 ( .A1(n4557), .A2(n8046), .ZN(n6455) );
  INV_X1 U8162 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8701) );
  OR2_X1 U8163 ( .A1(n6588), .A2(n8701), .ZN(n6454) );
  AND2_X1 U8164 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  OAI211_X1 U8165 ( .C1(n6569), .C2(n8702), .A(n6457), .B(n6456), .ZN(n8662)
         );
  NAND2_X1 U8166 ( .A1(n8107), .A2(n8662), .ZN(n6458) );
  OR2_X1 U8167 ( .A1(n8107), .A2(n8662), .ZN(n6459) );
  NAND2_X1 U8168 ( .A1(n7175), .A2(n4541), .ZN(n6466) );
  NAND2_X1 U8169 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U8170 ( .A1(n6463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6464) );
  XNOR2_X1 U8171 ( .A(n6464), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8748) );
  AOI22_X1 U8172 ( .A1(n8748), .A2(n4547), .B1(n6486), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8173 ( .A1(n6466), .A2(n6465), .ZN(n8634) );
  INV_X1 U8174 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U8175 ( .A1(n6467), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8176 ( .A1(n6477), .A2(n6468), .ZN(n8644) );
  NAND2_X1 U8177 ( .A1(n8644), .A2(n6565), .ZN(n6470) );
  AOI22_X1 U8178 ( .A1(n6566), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n8174), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n6469) );
  OAI211_X1 U8179 ( .C1(n6548), .C2(n9270), .A(n6470), .B(n6469), .ZN(n9013)
         );
  INV_X1 U8180 ( .A(n9013), .ZN(n8575) );
  OR2_X1 U8181 ( .A1(n8634), .A2(n8575), .ZN(n8329) );
  NAND2_X1 U8182 ( .A1(n8634), .A2(n8575), .ZN(n8328) );
  NAND2_X1 U8183 ( .A1(n8634), .A2(n9013), .ZN(n6471) );
  NAND2_X1 U8184 ( .A1(n7302), .A2(n4541), .ZN(n6476) );
  NAND2_X1 U8185 ( .A1(n4644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6472) );
  MUX2_X1 U8186 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6472), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6473) );
  NAND2_X1 U8187 ( .A1(n6473), .A2(n4578), .ZN(n8772) );
  OAI22_X1 U8188 ( .A1(n8772), .A2(n8172), .B1(n6276), .B2(n7303), .ZN(n6474)
         );
  INV_X1 U8189 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8190 ( .A1(n6477), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8191 ( .A1(n6490), .A2(n6478), .ZN(n9009) );
  NAND2_X1 U8192 ( .A1(n9009), .A2(n6565), .ZN(n6484) );
  INV_X1 U8193 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8194 ( .A1(n6566), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8195 ( .A1(n6557), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6479) );
  OAI211_X1 U8196 ( .C1(n4557), .C2(n6481), .A(n6480), .B(n6479), .ZN(n6482)
         );
  INV_X1 U8197 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8198 ( .A1(n6484), .A2(n6483), .ZN(n8661) );
  INV_X1 U8199 ( .A(n8661), .ZN(n8992) );
  NAND2_X1 U8200 ( .A1(n9444), .A2(n8992), .ZN(n8331) );
  INV_X1 U8201 ( .A(n9010), .ZN(n8208) );
  NAND2_X1 U8202 ( .A1(n7330), .A2(n4541), .ZN(n6489) );
  NAND2_X1 U8203 ( .A1(n4578), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6485) );
  XNOR2_X1 U8204 ( .A(n6485), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8797) );
  AOI22_X1 U8205 ( .A1(n8797), .A2(n4547), .B1(n6486), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8206 ( .A1(n6489), .A2(n6488), .ZN(n8580) );
  NAND2_X1 U8207 ( .A1(n6490), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8208 ( .A1(n6492), .A2(n6491), .ZN(n8998) );
  NAND2_X1 U8209 ( .A1(n8998), .A2(n6565), .ZN(n6498) );
  INV_X1 U8210 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8211 ( .A1(n8174), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6494) );
  INV_X1 U8212 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9440) );
  OR2_X1 U8213 ( .A1(n6588), .A2(n9440), .ZN(n6493) );
  OAI211_X1 U8214 ( .C1(n6495), .C2(n6548), .A(n6494), .B(n6493), .ZN(n6496)
         );
  INV_X1 U8215 ( .A(n6496), .ZN(n6497) );
  OR2_X1 U8216 ( .A1(n8580), .A2(n8975), .ZN(n8336) );
  NAND2_X1 U8217 ( .A1(n8580), .A2(n8975), .ZN(n8340) );
  NAND2_X1 U8218 ( .A1(n8336), .A2(n8340), .ZN(n8988) );
  OR2_X1 U8219 ( .A1(n8967), .A2(n8951), .ZN(n8346) );
  AND2_X1 U8220 ( .A1(n8967), .A2(n8951), .ZN(n8241) );
  INV_X1 U8221 ( .A(n8241), .ZN(n8348) );
  NAND2_X1 U8222 ( .A1(n9062), .A2(n8964), .ZN(n8349) );
  NAND2_X1 U8223 ( .A1(n8357), .A2(n8349), .ZN(n8955) );
  NAND2_X1 U8224 ( .A1(n7789), .A2(n4541), .ZN(n6500) );
  OR2_X1 U8225 ( .A1(n6276), .A2(n9264), .ZN(n6499) );
  NAND2_X1 U8226 ( .A1(n6501), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8227 ( .A1(n6510), .A2(n6502), .ZN(n8942) );
  NAND2_X1 U8228 ( .A1(n8942), .A2(n6565), .ZN(n6507) );
  INV_X1 U8229 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U8230 ( .A1(n6557), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8231 ( .A1(n8174), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6503) );
  OAI211_X1 U8232 ( .C1(n6588), .C2(n9279), .A(n6504), .B(n6503), .ZN(n6505)
         );
  INV_X1 U8233 ( .A(n6505), .ZN(n6506) );
  NAND2_X1 U8234 ( .A1(n6507), .A2(n6506), .ZN(n8658) );
  NAND2_X1 U8235 ( .A1(n8560), .A2(n8952), .ZN(n8360) );
  NAND2_X1 U8236 ( .A1(n7931), .A2(n4541), .ZN(n6509) );
  OR2_X1 U8237 ( .A1(n6276), .A2(n9186), .ZN(n6508) );
  NAND2_X1 U8238 ( .A1(n6510), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U8239 ( .A1(n6519), .A2(n6511), .ZN(n8932) );
  NAND2_X1 U8240 ( .A1(n8932), .A2(n6565), .ZN(n6516) );
  INV_X1 U8241 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U8242 ( .A1(n6557), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8243 ( .A1(n8174), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6512) );
  OAI211_X1 U8244 ( .C1(n6270), .C2(n9409), .A(n6513), .B(n6512), .ZN(n6514)
         );
  INV_X1 U8245 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U8246 ( .A1(n6516), .A2(n6515), .ZN(n8657) );
  OR2_X1 U8247 ( .A1(n8604), .A2(n8939), .ZN(n8234) );
  NAND2_X1 U8248 ( .A1(n8604), .A2(n8939), .ZN(n8233) );
  NAND2_X1 U8249 ( .A1(n7940), .A2(n4541), .ZN(n6518) );
  OR2_X1 U8250 ( .A1(n6276), .A2(n7942), .ZN(n6517) );
  NAND2_X1 U8251 ( .A1(n6519), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8252 ( .A1(n6521), .A2(n6520), .ZN(n8922) );
  NAND2_X1 U8253 ( .A1(n8922), .A2(n6565), .ZN(n6527) );
  INV_X1 U8254 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8255 ( .A1(n6566), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8256 ( .A1(n8174), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8257 ( .C1(n6524), .C2(n6548), .A(n6523), .B(n6522), .ZN(n6525)
         );
  INV_X1 U8258 ( .A(n6525), .ZN(n6526) );
  NAND2_X1 U8259 ( .A1(n8048), .A2(n4541), .ZN(n6530) );
  OR2_X1 U8260 ( .A1(n6276), .A2(n8415), .ZN(n6529) );
  NAND2_X1 U8261 ( .A1(n6531), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8262 ( .A1(n6533), .A2(n6532), .ZN(n8899) );
  NAND2_X1 U8263 ( .A1(n8899), .A2(n6565), .ZN(n6538) );
  INV_X1 U8264 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U8265 ( .A1(n6566), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8266 ( .A1(n6557), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6534) );
  OAI211_X1 U8267 ( .C1(n4557), .C2(n9483), .A(n6535), .B(n6534), .ZN(n6536)
         );
  INV_X1 U8268 ( .A(n6536), .ZN(n6537) );
  OR2_X1 U8269 ( .A1(n9043), .A2(n8908), .ZN(n8372) );
  NAND2_X1 U8270 ( .A1(n9043), .A2(n8908), .ZN(n6617) );
  NAND2_X1 U8271 ( .A1(n8103), .A2(n4541), .ZN(n6541) );
  OR2_X1 U8272 ( .A1(n6276), .A2(n6539), .ZN(n6540) );
  INV_X1 U8273 ( .A(n6544), .ZN(n6543) );
  INV_X1 U8274 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8275 ( .A1(n6543), .A2(n6542), .ZN(n6555) );
  NAND2_X1 U8276 ( .A1(n6544), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8277 ( .A1(n6555), .A2(n6545), .ZN(n8879) );
  NAND2_X1 U8278 ( .A1(n8879), .A2(n6565), .ZN(n6552) );
  INV_X1 U8279 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8280 ( .A1(n8174), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8281 ( .A1(n6566), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6546) );
  OAI211_X1 U8282 ( .C1(n6549), .C2(n6548), .A(n6547), .B(n6546), .ZN(n6550)
         );
  INV_X1 U8283 ( .A(n6550), .ZN(n6551) );
  NAND2_X1 U8284 ( .A1(n8518), .A2(n8652), .ZN(n6618) );
  OR2_X1 U8285 ( .A1(n8518), .A2(n8652), .ZN(n6619) );
  INV_X1 U8286 ( .A(n6619), .ZN(n8383) );
  NAND2_X1 U8287 ( .A1(n8159), .A2(n4541), .ZN(n6554) );
  OR2_X1 U8288 ( .A1(n6276), .A2(n8122), .ZN(n6553) );
  OR2_X2 U8289 ( .A1(n6555), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U8290 ( .A1(n6555), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8291 ( .A1(n6564), .A2(n6556), .ZN(n8870) );
  INV_X1 U8292 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U8293 ( .A1(n6566), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8294 ( .A1(n6557), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6558) );
  OAI211_X1 U8295 ( .C1(n4557), .C2(n9472), .A(n6559), .B(n6558), .ZN(n6560)
         );
  NAND2_X1 U8296 ( .A1(n9474), .A2(n8876), .ZN(n6561) );
  INV_X1 U8297 ( .A(n8876), .ZN(n8651) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8483) );
  OR2_X1 U8299 ( .A1(n6276), .A2(n8483), .ZN(n6562) );
  OAI21_X2 U8300 ( .B1(n10471), .B2(n6563), .A(n6562), .ZN(n9468) );
  NAND2_X1 U8301 ( .A1(n8850), .A2(n6565), .ZN(n8181) );
  INV_X1 U8302 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U8303 ( .A1(n6566), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8304 ( .A1(n8174), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U8305 ( .C1(n8857), .C2(n6569), .A(n6568), .B(n6567), .ZN(n6570)
         );
  INV_X1 U8306 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U8307 ( .A1(n8181), .A2(n6571), .ZN(n8650) );
  INV_X1 U8308 ( .A(n8650), .ZN(n8863) );
  OR2_X1 U8309 ( .A1(n9468), .A2(n8863), .ZN(n8389) );
  NAND2_X1 U8310 ( .A1(n9468), .A2(n8863), .ZN(n8221) );
  XNOR2_X1 U8311 ( .A(n6572), .B(n8223), .ZN(n6598) );
  INV_X1 U8312 ( .A(n6577), .ZN(n6575) );
  NAND2_X1 U8313 ( .A1(n6575), .A2(n6574), .ZN(n6628) );
  NAND2_X1 U8314 ( .A1(n6628), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6576) );
  OR2_X1 U8315 ( .A1(n6622), .A2(n7932), .ZN(n6584) );
  NAND2_X1 U8316 ( .A1(n6577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6578) );
  MUX2_X1 U8317 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6578), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6579) );
  NAND2_X1 U8318 ( .A1(n6580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U8319 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6581), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6582) );
  INV_X1 U8320 ( .A(n8406), .ZN(n6896) );
  NAND2_X1 U8321 ( .A1(n8229), .A2(n6896), .ZN(n6583) );
  INV_X1 U8322 ( .A(n6778), .ZN(n8408) );
  NAND2_X1 U8323 ( .A1(n8408), .A2(n8822), .ZN(n6586) );
  INV_X1 U8324 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8325 ( .A1(n8174), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6590) );
  INV_X1 U8326 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6587) );
  OR2_X1 U8327 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  OAI211_X1 U8328 ( .C1(n6591), .C2(n6569), .A(n6590), .B(n6589), .ZN(n6592)
         );
  INV_X1 U8329 ( .A(n6592), .ZN(n6593) );
  NAND2_X1 U8330 ( .A1(n8172), .A2(P2_B_REG_SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8331 ( .A1(n9014), .A2(n6594), .ZN(n8848) );
  INV_X1 U8332 ( .A(n7344), .ZN(n6986) );
  INV_X1 U8333 ( .A(n8261), .ZN(n6599) );
  NAND2_X1 U8334 ( .A1(n8190), .A2(n6599), .ZN(n7073) );
  INV_X1 U8335 ( .A(n8274), .ZN(n8187) );
  NAND2_X1 U8336 ( .A1(n7056), .A2(n8187), .ZN(n6600) );
  INV_X1 U8337 ( .A(n8268), .ZN(n7366) );
  OR2_X1 U8338 ( .A1(n7366), .A2(n4669), .ZN(n8267) );
  NAND2_X1 U8339 ( .A1(n6601), .A2(n8286), .ZN(n7067) );
  OR2_X1 U8340 ( .A1(n7895), .A2(n7282), .ZN(n8287) );
  NAND2_X1 U8341 ( .A1(n7067), .A2(n8287), .ZN(n6602) );
  NAND2_X1 U8342 ( .A1(n7895), .A2(n7282), .ZN(n8279) );
  INV_X1 U8343 ( .A(n8670), .ZN(n7431) );
  NAND2_X1 U8344 ( .A1(n7660), .A2(n7431), .ZN(n8282) );
  AND2_X1 U8345 ( .A1(n8282), .A2(n7209), .ZN(n8294) );
  OR2_X1 U8346 ( .A1(n7660), .A2(n7431), .ZN(n8285) );
  NAND2_X1 U8347 ( .A1(n7405), .A2(n8298), .ZN(n6603) );
  OR2_X1 U8348 ( .A1(n8248), .A2(n8247), .ZN(n8244) );
  NAND2_X1 U8349 ( .A1(n7669), .A2(n7633), .ZN(n8250) );
  INV_X1 U8350 ( .A(n8667), .ZN(n7885) );
  NAND2_X1 U8351 ( .A1(n4588), .A2(n8251), .ZN(n8198) );
  OR2_X1 U8352 ( .A1(n7891), .A2(n7960), .ZN(n8304) );
  INV_X1 U8353 ( .A(n8304), .ZN(n6605) );
  OR2_X2 U8354 ( .A1(n7570), .A2(n6605), .ZN(n7718) );
  NAND2_X1 U8355 ( .A1(n7726), .A2(n8028), .ZN(n8306) );
  NAND2_X1 U8356 ( .A1(n7891), .A2(n7960), .ZN(n8252) );
  AND2_X1 U8357 ( .A1(n8306), .A2(n8252), .ZN(n8303) );
  NAND2_X1 U8358 ( .A1(n7718), .A2(n8303), .ZN(n6606) );
  OR2_X1 U8359 ( .A1(n7726), .A2(n8028), .ZN(n8308) );
  NAND2_X1 U8360 ( .A1(n6606), .A2(n8308), .ZN(n7905) );
  NOR2_X1 U8361 ( .A1(n8030), .A2(n7965), .ZN(n8311) );
  INV_X1 U8362 ( .A(n8311), .ZN(n6608) );
  AND2_X1 U8363 ( .A1(n8030), .A2(n7965), .ZN(n8312) );
  INV_X1 U8364 ( .A(n8312), .ZN(n6607) );
  NAND2_X1 U8365 ( .A1(n7905), .A2(n8314), .ZN(n6609) );
  NAND2_X1 U8366 ( .A1(n7946), .A2(n8205), .ZN(n6611) );
  INV_X1 U8367 ( .A(n8663), .ZN(n8113) );
  OR2_X1 U8368 ( .A1(n8318), .A2(n8113), .ZN(n6610) );
  INV_X1 U8369 ( .A(n8662), .ZN(n8642) );
  OR2_X1 U8370 ( .A1(n8107), .A2(n8642), .ZN(n8323) );
  INV_X1 U8371 ( .A(n8323), .ZN(n6612) );
  NAND2_X1 U8372 ( .A1(n8107), .A2(n8642), .ZN(n8324) );
  NAND2_X1 U8373 ( .A1(n9450), .A2(n8329), .ZN(n9008) );
  NAND2_X1 U8374 ( .A1(n9008), .A2(n9010), .ZN(n9007) );
  NAND2_X1 U8375 ( .A1(n9007), .A2(n8332), .ZN(n8995) );
  NAND2_X1 U8376 ( .A1(n8492), .A2(n8994), .ZN(n8341) );
  NAND2_X1 U8377 ( .A1(n8337), .A2(n8341), .ZN(n8980) );
  INV_X1 U8378 ( .A(n8337), .ZN(n6613) );
  AOI21_X1 U8379 ( .B1(n8960), .B2(n8346), .A(n8241), .ZN(n8956) );
  INV_X1 U8380 ( .A(n8357), .ZN(n6614) );
  INV_X1 U8381 ( .A(n8360), .ZN(n6615) );
  OAI21_X1 U8382 ( .B1(n8941), .B2(n6615), .A(n8358), .ZN(n8930) );
  INV_X1 U8383 ( .A(n8234), .ZN(n6616) );
  OR2_X1 U8384 ( .A1(n8533), .A2(n8929), .ZN(n8362) );
  NAND2_X1 U8385 ( .A1(n8921), .A2(n8362), .ZN(n8912) );
  AND2_X1 U8386 ( .A1(n8594), .A2(n8919), .ZN(n8364) );
  INV_X1 U8387 ( .A(n8364), .ZN(n8213) );
  NAND2_X1 U8388 ( .A1(n8533), .A2(n8929), .ZN(n8911) );
  AND2_X1 U8389 ( .A1(n8213), .A2(n8911), .ZN(n8367) );
  INV_X1 U8390 ( .A(n8363), .ZN(n8366) );
  INV_X1 U8391 ( .A(n6617), .ZN(n8374) );
  OR2_X1 U8392 ( .A1(n8630), .A2(n8897), .ZN(n8378) );
  NAND2_X1 U8393 ( .A1(n8630), .A2(n8897), .ZN(n8379) );
  NAND2_X1 U8394 ( .A1(n6619), .A2(n6618), .ZN(n8877) );
  INV_X1 U8395 ( .A(n8877), .ZN(n6620) );
  XNOR2_X1 U8396 ( .A(n8552), .B(n8876), .ZN(n8868) );
  INV_X1 U8397 ( .A(n8868), .ZN(n6621) );
  XNOR2_X1 U8398 ( .A(n8224), .B(n8223), .ZN(n8859) );
  NAND2_X1 U8399 ( .A1(n8229), .A2(n8406), .ZN(n7364) );
  NAND2_X1 U8400 ( .A1(n7932), .A2(n7364), .ZN(n6623) );
  NAND2_X1 U8401 ( .A1(n7345), .A2(n6625), .ZN(n7653) );
  NAND2_X1 U8402 ( .A1(n6898), .A2(n8406), .ZN(n6901) );
  OR2_X1 U8403 ( .A1(n6901), .A2(n8411), .ZN(n7731) );
  INV_X1 U8404 ( .A(n6625), .ZN(n6626) );
  OR2_X1 U8405 ( .A1(n6626), .A2(n8406), .ZN(n6627) );
  NAND2_X1 U8406 ( .A1(n6627), .A2(n8402), .ZN(n6649) );
  NAND2_X1 U8407 ( .A1(n6629), .A2(n6634), .ZN(n6631) );
  NAND2_X1 U8408 ( .A1(n6631), .A2(n6630), .ZN(n6645) );
  XNOR2_X1 U8409 ( .A(n6645), .B(P2_B_REG_SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8410 ( .A1(n6633), .A2(n6641), .ZN(n6640) );
  NAND3_X1 U8411 ( .A1(n6635), .A2(n6634), .A3(n6666), .ZN(n6636) );
  OAI21_X1 U8412 ( .B1(n6637), .B2(n6636), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6638) );
  MUX2_X1 U8413 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6638), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6639) );
  OR2_X1 U8414 ( .A1(n6647), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8415 ( .A1(n6641), .A2(n8102), .ZN(n6643) );
  NAND2_X1 U8416 ( .A1(n6645), .A2(n8102), .ZN(n6646) );
  INV_X1 U8417 ( .A(n6924), .ZN(n6648) );
  NAND2_X1 U8418 ( .A1(n6649), .A2(n6648), .ZN(n6650) );
  NOR2_X1 U8419 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n6655) );
  NOR4_X1 U8420 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6654) );
  NOR4_X1 U8421 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6653) );
  NOR4_X1 U8422 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6652) );
  NAND4_X1 U8423 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(n6661)
         );
  NOR4_X1 U8424 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6659) );
  NOR4_X1 U8425 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6658) );
  NOR4_X1 U8426 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6657) );
  NOR4_X1 U8427 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6656) );
  NAND4_X1 U8428 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6660)
         );
  NOR2_X1 U8429 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  INV_X1 U8430 ( .A(n6641), .ZN(n6664) );
  AND2_X1 U8431 ( .A1(n6814), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8432 ( .A1(n6900), .A2(n6915), .ZN(n6667) );
  AND2_X1 U8433 ( .A1(n6899), .A2(n6924), .ZN(n6895) );
  INV_X1 U8434 ( .A(n6895), .ZN(n6668) );
  NAND2_X1 U8435 ( .A1(n6668), .A2(n6913), .ZN(n6669) );
  INV_X1 U8436 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6671) );
  INV_X1 U8437 ( .A(n6674), .ZN(n6675) );
  OR2_X2 U8438 ( .A1(n6685), .A2(n6675), .ZN(n9985) );
  INV_X1 U8439 ( .A(n6814), .ZN(n7083) );
  NAND2_X1 U8440 ( .A1(n6903), .A2(n8402), .ZN(n6676) );
  NAND2_X1 U8441 ( .A1(n6676), .A2(n6814), .ZN(n6833) );
  NAND2_X1 U8442 ( .A1(n6833), .A2(n8172), .ZN(n6677) );
  NAND2_X1 U8443 ( .A1(n6677), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  OAI21_X1 U8444 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n7301) );
  AND2_X1 U8445 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9992) );
  INV_X1 U8446 ( .A(n4558), .ZN(n9948) );
  MUX2_X1 U8447 ( .A(n7301), .B(n9992), .S(n9948), .Z(n6683) );
  AOI21_X1 U8448 ( .B1(n9948), .B2(n7242), .A(n5871), .ZN(n6942) );
  OAI21_X1 U8449 ( .B1(n6942), .B2(P1_IR_REG_0__SCAN_IN), .A(P1_U3973), .ZN(
        n6681) );
  AOI21_X1 U8450 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6717) );
  INV_X1 U8451 ( .A(n7937), .ZN(n6684) );
  OR2_X1 U8452 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  AND2_X1 U8453 ( .A1(n6686), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8454 ( .A1(n9932), .A2(n7937), .ZN(n6687) );
  AND2_X1 U8455 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U8456 ( .A1(n6944), .A2(n5871), .ZN(n10089) );
  NOR2_X1 U8457 ( .A1(n10089), .A2(n4554), .ZN(n6704) );
  INV_X1 U8458 ( .A(n6689), .ZN(n6690) );
  NAND2_X1 U8459 ( .A1(n6691), .A2(n6690), .ZN(n10099) );
  INV_X1 U8460 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6692) );
  OAI22_X1 U8461 ( .A1(n10099), .A2(n6692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7502), .ZN(n6703) );
  INV_X1 U8462 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7192) );
  MUX2_X1 U8463 ( .A(n7192), .B(P1_REG1_REG_2__SCAN_IN), .S(n4554), .Z(n6695)
         );
  INV_X1 U8464 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10636) );
  MUX2_X1 U8465 ( .A(n10636), .B(P1_REG1_REG_1__SCAN_IN), .S(n6727), .Z(n9990)
         );
  AND2_X1 U8466 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9989) );
  NAND2_X1 U8467 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  NAND2_X1 U8468 ( .A1(n5400), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8469 ( .A1(n9988), .A2(n6693), .ZN(n6694) );
  OAI21_X1 U8470 ( .B1(n6695), .B2(n6694), .A(n6709), .ZN(n6701) );
  MUX2_X1 U8471 ( .A(n7501), .B(P1_REG2_REG_2__SCAN_IN), .S(n4554), .Z(n6699)
         );
  MUX2_X1 U8472 ( .A(n7494), .B(P1_REG2_REG_1__SCAN_IN), .S(n6727), .Z(n9993)
         );
  NAND2_X1 U8473 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  NAND2_X1 U8474 ( .A1(n5400), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8475 ( .A1(n9991), .A2(n6696), .ZN(n6698) );
  NOR2_X1 U8476 ( .A1(n5871), .A2(n4558), .ZN(n6697) );
  NAND2_X1 U8477 ( .A1(n6699), .A2(n6698), .ZN(n6705) );
  OAI211_X1 U8478 ( .C1(n6699), .C2(n6698), .A(n10093), .B(n6705), .ZN(n6700)
         );
  OAI21_X1 U8479 ( .B1(n10090), .B2(n6701), .A(n6700), .ZN(n6702) );
  OR4_X1 U8480 ( .A1(n6717), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(P1_U3245)
         );
  OAI21_X1 U8481 ( .B1(n7501), .B2(n4554), .A(n6705), .ZN(n10003) );
  INV_X1 U8482 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6706) );
  MUX2_X1 U8483 ( .A(n6706), .B(P1_REG2_REG_3__SCAN_IN), .S(n6722), .Z(n10004)
         );
  AND2_X1 U8484 ( .A1(n10003), .A2(n10004), .ZN(n10001) );
  XOR2_X1 U8485 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6952), .Z(n6707) );
  NOR2_X1 U8486 ( .A1(n6708), .A2(n6707), .ZN(n6953) );
  AOI211_X1 U8487 ( .C1(n6708), .C2(n6707), .A(n6953), .B(n10037), .ZN(n6716)
         );
  NAND2_X1 U8488 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7310) );
  OAI21_X1 U8489 ( .B1(n10099), .B2(n9412), .A(n7310), .ZN(n6715) );
  INV_X1 U8490 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9397) );
  MUX2_X1 U8491 ( .A(n9397), .B(P1_REG1_REG_4__SCAN_IN), .S(n6952), .Z(n6712)
         );
  INV_X1 U8492 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U8493 ( .B1(n7192), .B2(n4554), .A(n6709), .ZN(n10006) );
  MUX2_X1 U8494 ( .A(n6710), .B(P1_REG1_REG_3__SCAN_IN), .S(n6722), .Z(n10007)
         );
  NAND2_X1 U8495 ( .A1(n10006), .A2(n10007), .ZN(n10005) );
  OAI211_X1 U8496 ( .C1(n6712), .C2(n6711), .A(n10087), .B(n6957), .ZN(n6713)
         );
  OAI21_X1 U8497 ( .B1(n10089), .B2(n6952), .A(n6713), .ZN(n6714) );
  OR4_X1 U8498 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(P1_U3247)
         );
  AND2_X1 U8499 ( .A1(n8171), .A2(P2_U3151), .ZN(n8119) );
  INV_X2 U8500 ( .A(n8119), .ZN(n9524) );
  NOR2_X1 U8501 ( .A1(n8171), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9522) );
  INV_X2 U8502 ( .A(n9522), .ZN(n8484) );
  OAI222_X1 U8503 ( .A1(P2_U3151), .A2(n6768), .B1(n9524), .B2(n6726), .C1(
        n4896), .C2(n8484), .ZN(P2_U3294) );
  OAI222_X1 U8504 ( .A1(n4548), .A2(P2_U3151), .B1(n9524), .B2(n6720), .C1(
        n6718), .C2(n8484), .ZN(P2_U3293) );
  INV_X1 U8505 ( .A(n6827), .ZN(n6800) );
  OAI222_X1 U8506 ( .A1(n6800), .A2(P2_U3151), .B1(n9524), .B2(n6723), .C1(
        n5215), .C2(n8484), .ZN(P2_U3292) );
  AND2_X1 U8507 ( .A1(n8171), .A2(P1_U3086), .ZN(n10464) );
  INV_X2 U8508 ( .A(n10464), .ZN(n10470) );
  OAI222_X1 U8509 ( .A1(P1_U3086), .A2(n4554), .B1(n10472), .B2(n6720), .C1(
        n6719), .C2(n10470), .ZN(P1_U3353) );
  OAI222_X1 U8510 ( .A1(n10470), .A2(n6724), .B1(n10472), .B2(n6723), .C1(
        P1_U3086), .C2(n6722), .ZN(P1_U3352) );
  OAI222_X1 U8511 ( .A1(P1_U3086), .A2(n6727), .B1(n10472), .B2(n6726), .C1(
        n6725), .C2(n10470), .ZN(P1_U3354) );
  OAI222_X1 U8512 ( .A1(n6880), .A2(P2_U3151), .B1(n9524), .B2(n6728), .C1(
        n4678), .C2(n8484), .ZN(P2_U3291) );
  OAI222_X1 U8513 ( .A1(n10470), .A2(n6729), .B1(n10472), .B2(n6728), .C1(
        P1_U3086), .C2(n6952), .ZN(P1_U3351) );
  OAI222_X1 U8514 ( .A1(n10470), .A2(n6730), .B1(n10472), .B2(n6731), .C1(
        P1_U3086), .C2(n6963), .ZN(P1_U3350) );
  OAI222_X1 U8515 ( .A1(n8684), .A2(P2_U3151), .B1(n9524), .B2(n6731), .C1(
        n4700), .C2(n8484), .ZN(P2_U3290) );
  INV_X1 U8516 ( .A(n6732), .ZN(n6735) );
  OAI222_X1 U8517 ( .A1(n10470), .A2(n6733), .B1(n10472), .B2(n6735), .C1(
        P1_U3086), .C2(n7004), .ZN(P1_U3349) );
  INV_X1 U8518 ( .A(n7148), .ZN(n7150) );
  INV_X1 U8519 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6734) );
  OAI222_X1 U8520 ( .A1(n7150), .A2(P2_U3151), .B1(n9524), .B2(n6735), .C1(
        n6734), .C2(n8484), .ZN(P2_U3289) );
  INV_X1 U8521 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6738) );
  INV_X1 U8522 ( .A(n6899), .ZN(n6736) );
  NAND2_X1 U8523 ( .A1(n6736), .A2(n6915), .ZN(n6737) );
  OAI21_X1 U8524 ( .B1(n6915), .B2(n6738), .A(n6737), .ZN(P2_U3377) );
  INV_X1 U8525 ( .A(n6739), .ZN(n6741) );
  INV_X1 U8526 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6740) );
  OAI222_X1 U8527 ( .A1(n5049), .A2(P2_U3151), .B1(n9524), .B2(n6741), .C1(
        n6740), .C2(n8484), .ZN(P2_U3288) );
  INV_X1 U8528 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6742) );
  INV_X1 U8529 ( .A(n7115), .ZN(n7109) );
  OAI222_X1 U8530 ( .A1(n10470), .A2(n6742), .B1(n10472), .B2(n6741), .C1(
        P1_U3086), .C2(n7109), .ZN(P1_U3348) );
  INV_X1 U8531 ( .A(n6743), .ZN(n6746) );
  AOI22_X1 U8532 ( .A1(n10017), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10464), .ZN(n6744) );
  OAI21_X1 U8533 ( .B1(n6746), .B2(n10472), .A(n6744), .ZN(P1_U3347) );
  INV_X1 U8534 ( .A(n7228), .ZN(n7472) );
  OAI222_X1 U8535 ( .A1(n7472), .A2(P2_U3151), .B1(n9524), .B2(n6746), .C1(
        n6745), .C2(n8484), .ZN(P2_U3287) );
  OR2_X1 U8536 ( .A1(n10458), .A2(n6747), .ZN(n10565) );
  NAND2_X1 U8537 ( .A1(n10565), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6748) );
  OAI21_X1 U8538 ( .B1(n10565), .B2(n6749), .A(n6748), .ZN(P1_U3440) );
  INV_X1 U8539 ( .A(n7613), .ZN(n7620) );
  INV_X1 U8540 ( .A(n6750), .ZN(n6751) );
  OAI222_X1 U8541 ( .A1(P2_U3151), .A2(n7620), .B1(n9524), .B2(n6751), .C1(
        n9151), .C2(n8484), .ZN(P2_U3286) );
  OAI222_X1 U8542 ( .A1(n10470), .A2(n6752), .B1(n10472), .B2(n6751), .C1(
        n7124), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8543 ( .A(n6753), .ZN(n6759) );
  AOI22_X1 U8544 ( .A1(n7356), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10464), .ZN(n6754) );
  OAI21_X1 U8545 ( .B1(n6759), .B2(n10472), .A(n6754), .ZN(P1_U3345) );
  INV_X1 U8546 ( .A(n10099), .ZN(n10055) );
  NOR2_X1 U8547 ( .A1(n10055), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8548 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6756) );
  NOR2_X1 U8549 ( .A1(n7010), .A2(n6756), .ZN(P2_U3247) );
  INV_X1 U8550 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6757) );
  NOR2_X1 U8551 ( .A1(n7010), .A2(n6757), .ZN(P2_U3249) );
  INV_X1 U8552 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6758) );
  NOR2_X1 U8553 ( .A1(n7010), .A2(n6758), .ZN(P2_U3258) );
  INV_X1 U8554 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9228) );
  NOR2_X1 U8555 ( .A1(n7010), .A2(n9228), .ZN(P2_U3259) );
  INV_X1 U8556 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9140) );
  NOR2_X1 U8557 ( .A1(n7010), .A2(n9140), .ZN(P2_U3260) );
  INV_X1 U8558 ( .A(n7627), .ZN(n7680) );
  OAI222_X1 U8559 ( .A1(P2_U3151), .A2(n7680), .B1(n9524), .B2(n6759), .C1(
        n9274), .C2(n8484), .ZN(P2_U3285) );
  INV_X1 U8560 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8561 ( .A1(n5695), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6763) );
  INV_X1 U8562 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6760) );
  OR2_X1 U8563 ( .A1(n5458), .A2(n6760), .ZN(n6762) );
  INV_X1 U8564 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10396) );
  OR2_X1 U8565 ( .A1(n4552), .A2(n10396), .ZN(n6761) );
  AND3_X1 U8566 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n10104) );
  INV_X1 U8567 ( .A(n10104), .ZN(n9929) );
  NAND2_X1 U8568 ( .A1(n9929), .A2(P1_U3973), .ZN(n6764) );
  OAI21_X1 U8569 ( .B1(P1_U3973), .B2(n6765), .A(n6764), .ZN(P1_U3585) );
  INV_X1 U8570 ( .A(n6777), .ZN(n6766) );
  MUX2_X1 U8571 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8798), .Z(n6773) );
  INV_X1 U8572 ( .A(n6773), .ZN(n6774) );
  INV_X1 U8573 ( .A(n4548), .ZN(n10649) );
  MUX2_X1 U8574 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6767), .Z(n6771) );
  INV_X1 U8575 ( .A(n6771), .ZN(n6772) );
  MUX2_X1 U8576 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6767), .Z(n6769) );
  MUX2_X1 U8577 ( .A(n6282), .B(n6281), .S(n6767), .Z(n6835) );
  NAND2_X1 U8578 ( .A1(n6835), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8579 ( .A1(n6849), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U8580 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  NAND2_X1 U8581 ( .A1(n6847), .A2(n6770), .ZN(n10653) );
  XNOR2_X1 U8582 ( .A(n6771), .B(n10649), .ZN(n10654) );
  NAND2_X1 U8583 ( .A1(n10653), .A2(n10654), .ZN(n10651) );
  OAI21_X1 U8584 ( .B1(n10649), .B2(n6772), .A(n10651), .ZN(n6820) );
  XNOR2_X1 U8585 ( .A(n6773), .B(n6800), .ZN(n6821) );
  NOR2_X1 U8586 ( .A1(n6820), .A2(n6821), .ZN(n6819) );
  AOI21_X1 U8587 ( .B1(n6827), .B2(n6774), .A(n6819), .ZN(n6776) );
  MUX2_X1 U8588 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8798), .Z(n6863) );
  XNOR2_X1 U8589 ( .A(n6863), .B(n6866), .ZN(n6775) );
  NAND2_X1 U8590 ( .A1(n6776), .A2(n6775), .ZN(n6864) );
  NOR2_X2 U8591 ( .A1(n8676), .A2(n8408), .ZN(n10652) );
  OAI211_X1 U8592 ( .C1(n6776), .C2(n6775), .A(n6864), .B(n10652), .ZN(n6811)
         );
  OR2_X1 U8593 ( .A1(n6778), .A2(P2_U3151), .ZN(n8120) );
  OR2_X1 U8594 ( .A1(n6777), .A2(n8120), .ZN(n6781) );
  NOR2_X1 U8595 ( .A1(n8798), .A2(P2_U3151), .ZN(n8104) );
  AND2_X1 U8596 ( .A1(n8104), .A2(n6778), .ZN(n6779) );
  NAND2_X1 U8597 ( .A1(n6833), .A2(n6779), .ZN(n6780) );
  NOR2_X1 U8598 ( .A1(n8120), .A2(n8798), .ZN(n6782) );
  XNOR2_X1 U8599 ( .A(n6798), .B(n7371), .ZN(n10662) );
  INV_X1 U8600 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8601 ( .A1(n6794), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8602 ( .A1(n6261), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8603 ( .A1(n4548), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8604 ( .A1(n6788), .A2(n6800), .ZN(n6789) );
  INV_X1 U8605 ( .A(n6789), .ZN(n6787) );
  MUX2_X1 U8606 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6308), .S(n6880), .Z(n6790)
         );
  NOR2_X1 U8607 ( .A1(n6787), .A2(n6790), .ZN(n6792) );
  INV_X1 U8608 ( .A(n6873), .ZN(n6791) );
  AOI21_X1 U8609 ( .B1(n6792), .B2(n6822), .A(n6791), .ZN(n6793) );
  NAND2_X1 U8610 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7169) );
  OAI21_X1 U8611 ( .B1(n8841), .B2(n6793), .A(n7169), .ZN(n6809) );
  XNOR2_X1 U8612 ( .A(n4548), .B(n7063), .ZN(n10646) );
  NAND2_X1 U8613 ( .A1(n6794), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U8614 ( .A1(n6261), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8615 ( .A1(n6796), .A2(n6797), .ZN(n6846) );
  OR2_X1 U8616 ( .A1(n6846), .A2(n6269), .ZN(n6844) );
  NAND2_X1 U8617 ( .A1(n6844), .A2(n6797), .ZN(n10645) );
  NAND2_X1 U8618 ( .A1(n10646), .A2(n10645), .ZN(n10644) );
  NAND2_X1 U8619 ( .A1(n4548), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8620 ( .A1(n6824), .A2(n6804), .ZN(n6802) );
  INV_X1 U8621 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7069) );
  MUX2_X1 U8622 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7069), .S(n6880), .Z(n6803)
         );
  NAND2_X1 U8623 ( .A1(n6802), .A2(n6803), .ZN(n6882) );
  INV_X1 U8624 ( .A(n6803), .ZN(n6805) );
  NAND3_X1 U8625 ( .A1(n6824), .A2(n6805), .A3(n6804), .ZN(n6807) );
  NOR2_X1 U8626 ( .A1(n8120), .A2(n8822), .ZN(n6806) );
  AOI21_X1 U8627 ( .B1(n6882), .B2(n6807), .A(n8806), .ZN(n6808) );
  AOI211_X1 U8628 ( .C1(n6866), .C2(n10650), .A(n6809), .B(n6808), .ZN(n6810)
         );
  OAI211_X1 U8629 ( .C1(n10657), .C2(n8129), .A(n6811), .B(n6810), .ZN(
        P2_U3186) );
  INV_X1 U8630 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8631 ( .A1(n5891), .A2(P1_U3973), .ZN(n6812) );
  OAI21_X1 U8632 ( .B1(P1_U3973), .B2(n6813), .A(n6812), .ZN(P1_U3554) );
  NAND4_X1 U8633 ( .A1(n8102), .A2(P2_STATE_REG_SCAN_IN), .A3(n6645), .A4(
        n6814), .ZN(n6815) );
  OAI21_X1 U8634 ( .B1(n7010), .B2(P2_D_REG_0__SCAN_IN), .A(n6815), .ZN(n6816)
         );
  INV_X1 U8635 ( .A(n6816), .ZN(P2_U3376) );
  INV_X1 U8636 ( .A(n6817), .ZN(n6841) );
  AOI22_X1 U8637 ( .A1(n7825), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9522), .ZN(n6818) );
  OAI21_X1 U8638 ( .B1(n6841), .B2(n9524), .A(n6818), .ZN(P2_U3284) );
  AOI21_X1 U8639 ( .B1(n6821), .B2(n6820), .A(n6819), .ZN(n6832) );
  INV_X1 U8640 ( .A(n10652), .ZN(n8846) );
  INV_X1 U8641 ( .A(n6822), .ZN(n6823) );
  AOI21_X1 U8642 ( .B1(n6292), .B2(n4655), .A(n6823), .ZN(n6829) );
  INV_X1 U8643 ( .A(n8806), .ZN(n10648) );
  OAI21_X1 U8644 ( .B1(n6825), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6824), .ZN(
        n6826) );
  AOI22_X1 U8645 ( .A1(n10650), .A2(n6827), .B1(n10648), .B2(n6826), .ZN(n6828) );
  NAND2_X1 U8646 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7085) );
  OAI211_X1 U8647 ( .C1(n6829), .C2(n8841), .A(n6828), .B(n7085), .ZN(n6830)
         );
  AOI21_X1 U8648 ( .B1(n8839), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6830), .ZN(
        n6831) );
  OAI21_X1 U8649 ( .B1(n6832), .B2(n8846), .A(n6831), .ZN(P2_U3185) );
  INV_X1 U8650 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6840) );
  INV_X1 U8651 ( .A(n6833), .ZN(n6834) );
  OAI21_X1 U8652 ( .B1(n6834), .B2(n8120), .A(n8846), .ZN(n6837) );
  OAI21_X1 U8653 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6835), .A(n6848), .ZN(n6836) );
  NAND2_X1 U8654 ( .A1(n6837), .A2(n6836), .ZN(n6839) );
  AOI22_X1 U8655 ( .A1(n10650), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6838) );
  OAI211_X1 U8656 ( .C1(n6840), .C2(n10657), .A(n6839), .B(n6838), .ZN(
        P2_U3182) );
  INV_X1 U8657 ( .A(n7395), .ZN(n7357) );
  OAI222_X1 U8658 ( .A1(n10470), .A2(n9293), .B1(n10472), .B2(n6841), .C1(
        P1_U3086), .C2(n7357), .ZN(P1_U3344) );
  INV_X1 U8659 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10690) );
  XNOR2_X1 U8660 ( .A(n6842), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6843) );
  OAI22_X1 U8661 ( .A1(n8841), .A2(n6843), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7376), .ZN(n6853) );
  INV_X1 U8662 ( .A(n6844), .ZN(n6845) );
  AOI21_X1 U8663 ( .B1(n6269), .B2(n6846), .A(n6845), .ZN(n6851) );
  OAI211_X1 U8664 ( .C1(n6849), .C2(n6848), .A(n10652), .B(n6847), .ZN(n6850)
         );
  OAI21_X1 U8665 ( .B1(n6851), .B2(n8806), .A(n6850), .ZN(n6852) );
  OAI21_X1 U8666 ( .B1(n10690), .B2(n10657), .A(n4654), .ZN(P2_U3183) );
  INV_X1 U8667 ( .A(n6854), .ZN(n6855) );
  OR2_X1 U8668 ( .A1(n6856), .A2(n6855), .ZN(n6858) );
  INV_X1 U8669 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U8670 ( .A1(n9941), .A2(n4549), .ZN(n10629) );
  NAND2_X1 U8671 ( .A1(n7185), .A2(n5891), .ZN(n9871) );
  INV_X1 U8672 ( .A(n7490), .ZN(n6859) );
  NAND2_X1 U8673 ( .A1(n9871), .A2(n6859), .ZN(n9811) );
  OAI21_X1 U8674 ( .B1(n10622), .B2(n10285), .A(n9811), .ZN(n6860) );
  NOR2_X1 U8675 ( .A1(n4688), .A2(n7846), .ZN(n7240) );
  INV_X1 U8676 ( .A(n7240), .ZN(n7296) );
  OAI211_X1 U8677 ( .C1(n6861), .C2(n7185), .A(n6860), .B(n7296), .ZN(n7262)
         );
  NAND2_X1 U8678 ( .A1(n7262), .A2(n10643), .ZN(n6862) );
  OAI21_X1 U8679 ( .B1(n10643), .B2(n6945), .A(n6862), .ZN(P1_U3522) );
  MUX2_X1 U8680 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8798), .Z(n7145) );
  XNOR2_X1 U8681 ( .A(n7145), .B(n7150), .ZN(n6871) );
  MUX2_X1 U8682 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8798), .Z(n6867) );
  INV_X1 U8683 ( .A(n6867), .ZN(n6868) );
  INV_X1 U8684 ( .A(n6863), .ZN(n6865) );
  OAI21_X1 U8685 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n8680) );
  XNOR2_X1 U8686 ( .A(n6867), .B(n6869), .ZN(n8679) );
  NAND2_X1 U8687 ( .A1(n8680), .A2(n8679), .ZN(n8678) );
  OAI21_X1 U8688 ( .B1(n6869), .B2(n6868), .A(n8678), .ZN(n6870) );
  NOR2_X1 U8689 ( .A1(n6870), .A2(n6871), .ZN(n7146) );
  AOI21_X1 U8690 ( .B1(n6871), .B2(n6870), .A(n7146), .ZN(n6891) );
  NAND2_X1 U8691 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7321) );
  OAI21_X1 U8692 ( .B1(n8837), .B2(n7150), .A(n7321), .ZN(n6879) );
  NAND2_X1 U8693 ( .A1(n6880), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U8694 ( .A1(n6874), .A2(n8684), .ZN(n6875) );
  XNOR2_X1 U8695 ( .A(n7148), .B(n7657), .ZN(n6876) );
  NAND3_X1 U8696 ( .A1(n8690), .A2(n6876), .A3(n6875), .ZN(n6877) );
  AOI21_X1 U8697 ( .B1(n5052), .B2(n6877), .A(n8841), .ZN(n6878) );
  AOI211_X1 U8698 ( .C1(n8839), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6879), .B(
        n6878), .ZN(n6890) );
  NAND2_X1 U8699 ( .A1(n6880), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8700 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  NAND2_X1 U8701 ( .A1(n6883), .A2(n8684), .ZN(n6885) );
  OR2_X1 U8702 ( .A1(n6883), .A2(n8684), .ZN(n6884) );
  INV_X1 U8703 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8687) );
  INV_X1 U8704 ( .A(n6885), .ZN(n6887) );
  XNOR2_X1 U8705 ( .A(n7148), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6886) );
  NOR3_X1 U8706 ( .A1(n8686), .A2(n6887), .A3(n6886), .ZN(n6888) );
  OAI21_X1 U8707 ( .B1(n4650), .B2(n6888), .A(n10648), .ZN(n6889) );
  OAI211_X1 U8708 ( .C1(n6891), .C2(n8846), .A(n6890), .B(n6889), .ZN(P2_U3188) );
  INV_X1 U8709 ( .A(n6892), .ZN(n6894) );
  INV_X1 U8710 ( .A(n7709), .ZN(n7401) );
  OAI222_X1 U8711 ( .A1(n10470), .A2(n9295), .B1(n10472), .B2(n6894), .C1(
        n7401), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U8712 ( .A1(P2_U3151), .A2(n7988), .B1(n9524), .B2(n6894), .C1(
        n6893), .C2(n8484), .ZN(P2_U3283) );
  NAND2_X1 U8713 ( .A1(n8262), .A2(n6896), .ZN(n6923) );
  NOR2_X1 U8714 ( .A1(n7932), .A2(n6923), .ZN(n6897) );
  NAND2_X1 U8715 ( .A1(n6898), .A2(n6897), .ZN(n7046) );
  NOR2_X1 U8716 ( .A1(n6899), .A2(n6924), .ZN(n7339) );
  NAND2_X1 U8717 ( .A1(n7339), .A2(n6900), .ZN(n6910) );
  NAND2_X1 U8718 ( .A1(n6901), .A2(n9443), .ZN(n8905) );
  AND2_X1 U8719 ( .A1(n8402), .A2(n9454), .ZN(n6902) );
  NAND2_X1 U8720 ( .A1(n7046), .A2(n6902), .ZN(n6931) );
  NAND2_X1 U8721 ( .A1(n8905), .A2(n6931), .ZN(n7049) );
  INV_X1 U8722 ( .A(n6903), .ZN(n6905) );
  AOI211_X1 U8723 ( .C1(n6910), .C2(n7049), .A(n6905), .B(n6904), .ZN(n6906)
         );
  OAI21_X1 U8724 ( .B1(n6916), .B2(n7046), .A(n6906), .ZN(n6908) );
  NOR2_X1 U8725 ( .A1(n7345), .A2(n6912), .ZN(n8409) );
  INV_X1 U8726 ( .A(n6916), .ZN(n6907) );
  AOI22_X1 U8727 ( .A1(n6908), .A2(P2_STATE_REG_SCAN_IN), .B1(n8409), .B2(
        n6907), .ZN(n7084) );
  AND2_X1 U8728 ( .A1(n7084), .A2(n6909), .ZN(n7102) );
  INV_X1 U8729 ( .A(n6910), .ZN(n6911) );
  AND2_X1 U8730 ( .A1(n6911), .A2(n6915), .ZN(n7048) );
  NAND2_X1 U8731 ( .A1(n7048), .A2(n9443), .ZN(n6914) );
  NOR2_X1 U8732 ( .A1(n7345), .A2(n6918), .ZN(n6917) );
  INV_X1 U8733 ( .A(n8639), .ZN(n8627) );
  INV_X1 U8734 ( .A(n6918), .ZN(n6919) );
  NOR2_X1 U8735 ( .A1(n7345), .A2(n6919), .ZN(n6920) );
  OAI22_X1 U8736 ( .A1(n8627), .A2(n6304), .B1(n8675), .B2(n8641), .ZN(n6921)
         );
  AOI21_X1 U8737 ( .B1(n8268), .B2(n8629), .A(n6921), .ZN(n6938) );
  XNOR2_X1 U8738 ( .A(n7162), .B(n8268), .ZN(n7088) );
  XNOR2_X1 U8739 ( .A(n7088), .B(n4669), .ZN(n6930) );
  XNOR2_X1 U8740 ( .A(n7162), .B(n7378), .ZN(n6925) );
  OR2_X1 U8741 ( .A1(n6925), .A2(n8675), .ZN(n6926) );
  NAND2_X1 U8742 ( .A1(n6925), .A2(n8675), .ZN(n6928) );
  NAND2_X1 U8743 ( .A1(n6929), .A2(n6930), .ZN(n7090) );
  OAI21_X1 U8744 ( .B1(n6930), .B2(n6929), .A(n7090), .ZN(n6936) );
  INV_X1 U8745 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U8746 ( .A1(n7048), .A2(n6932), .ZN(n6935) );
  INV_X1 U8747 ( .A(n7046), .ZN(n6933) );
  NAND2_X1 U8748 ( .A1(n7050), .A2(n6933), .ZN(n6934) );
  NAND2_X1 U8749 ( .A1(n6936), .A2(n8635), .ZN(n6937) );
  OAI211_X1 U8750 ( .C1(n7102), .C2(n6939), .A(n6938), .B(n6937), .ZN(P2_U3177) );
  INV_X1 U8751 ( .A(n6940), .ZN(n6991) );
  AOI22_X1 U8752 ( .A1(n8713), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9522), .ZN(n6941) );
  OAI21_X1 U8753 ( .B1(n6991), .B2(n9524), .A(n6941), .ZN(P2_U3282) );
  OAI21_X1 U8754 ( .B1(n9948), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6942), .ZN(
        n6943) );
  MUX2_X1 U8755 ( .A(n6943), .B(n6942), .S(P1_IR_REG_0__SCAN_IN), .Z(n6951) );
  INV_X1 U8756 ( .A(n6944), .ZN(n6950) );
  NAND3_X1 U8757 ( .A1(n10087), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6945), .ZN(
        n6949) );
  INV_X1 U8758 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6946) );
  OAI22_X1 U8759 ( .A1(n10099), .A2(n6946), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7297), .ZN(n6947) );
  INV_X1 U8760 ( .A(n6947), .ZN(n6948) );
  OAI211_X1 U8761 ( .C1(n6951), .C2(n6950), .A(n6949), .B(n6948), .ZN(P1_U3243) );
  INV_X1 U8762 ( .A(n6952), .ZN(n6959) );
  AOI21_X1 U8763 ( .B1(n6959), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6953), .ZN(
        n6956) );
  MUX2_X1 U8764 ( .A(n5479), .B(P1_REG2_REG_5__SCAN_IN), .S(n6963), .Z(n6954)
         );
  INV_X1 U8765 ( .A(n6954), .ZN(n6955) );
  NOR2_X1 U8766 ( .A1(n6956), .A2(n6955), .ZN(n6969) );
  AOI211_X1 U8767 ( .C1(n6956), .C2(n6955), .A(n6969), .B(n10037), .ZN(n6968)
         );
  INV_X1 U8768 ( .A(n6957), .ZN(n6958) );
  INV_X1 U8769 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6960) );
  MUX2_X1 U8770 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6960), .S(n6963), .Z(n6961)
         );
  NOR2_X1 U8771 ( .A1(n6962), .A2(n6961), .ZN(n6973) );
  AOI211_X1 U8772 ( .C1(n6962), .C2(n6961), .A(n6973), .B(n10090), .ZN(n6967)
         );
  INV_X1 U8773 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6965) );
  INV_X1 U8774 ( .A(n6963), .ZN(n6974) );
  NAND2_X1 U8775 ( .A1(n10072), .A2(n6974), .ZN(n6964) );
  NAND2_X1 U8776 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7584) );
  OAI211_X1 U8777 ( .C1(n6965), .C2(n10099), .A(n6964), .B(n7584), .ZN(n6966)
         );
  OR3_X1 U8778 ( .A1(n6968), .A2(n6967), .A3(n6966), .ZN(P1_U3248) );
  MUX2_X1 U8779 ( .A(n7005), .B(P1_REG2_REG_6__SCAN_IN), .S(n7004), .Z(n6970)
         );
  INV_X1 U8780 ( .A(n6970), .ZN(n6971) );
  NOR2_X1 U8781 ( .A1(n6972), .A2(n6971), .ZN(n7002) );
  AOI211_X1 U8782 ( .C1(n6972), .C2(n6971), .A(n10037), .B(n7002), .ZN(n6981)
         );
  AOI21_X1 U8783 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6974), .A(n6973), .ZN(
        n6977) );
  INV_X1 U8784 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U8785 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6975), .S(n7004), .Z(n6976)
         );
  NOR2_X1 U8786 ( .A1(n6977), .A2(n6976), .ZN(n6995) );
  AOI211_X1 U8787 ( .C1(n6977), .C2(n6976), .A(n10090), .B(n6995), .ZN(n6980)
         );
  INV_X1 U8788 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8132) );
  INV_X1 U8789 ( .A(n7004), .ZN(n6996) );
  NAND2_X1 U8790 ( .A1(n10072), .A2(n6996), .ZN(n6978) );
  NAND2_X1 U8791 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10538) );
  OAI211_X1 U8792 ( .C1(n8132), .C2(n10099), .A(n6978), .B(n10538), .ZN(n6979)
         );
  OR3_X1 U8793 ( .A1(n6981), .A2(n6980), .A3(n6979), .ZN(P1_U3249) );
  NAND2_X1 U8794 ( .A1(n6986), .A2(n8677), .ZN(n8258) );
  AND2_X1 U8795 ( .A1(n8258), .A2(n8261), .ZN(n8188) );
  INV_X1 U8796 ( .A(n8188), .ZN(n6988) );
  OAI21_X1 U8797 ( .B1(n9449), .B2(n9017), .A(n6988), .ZN(n6984) );
  NOR2_X1 U8798 ( .A1(n8675), .A2(n8953), .ZN(n7348) );
  AND2_X1 U8799 ( .A1(n7344), .A2(n9443), .ZN(n6982) );
  NOR2_X1 U8800 ( .A1(n7348), .A2(n6982), .ZN(n6983) );
  NAND2_X1 U8801 ( .A1(n6984), .A2(n6983), .ZN(n7053) );
  NAND2_X1 U8802 ( .A1(n7053), .A2(n9456), .ZN(n6985) );
  OAI21_X1 U8803 ( .B1(n9456), .B2(n6281), .A(n6985), .ZN(P2_U3459) );
  INV_X1 U8804 ( .A(n8629), .ZN(n8648) );
  OAI22_X1 U8805 ( .A1(n8648), .A2(n6986), .B1(n8627), .B2(n8675), .ZN(n6987)
         );
  AOI21_X1 U8806 ( .B1(n6988), .B2(n8635), .A(n6987), .ZN(n6989) );
  OAI21_X1 U8807 ( .B1(n7102), .B2(n6990), .A(n6989), .ZN(P2_U3172) );
  INV_X1 U8808 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6992) );
  INV_X1 U8809 ( .A(n7871), .ZN(n7705) );
  OAI222_X1 U8810 ( .A1(n10470), .A2(n6992), .B1(n10472), .B2(n6991), .C1(
        P1_U3086), .C2(n7705), .ZN(P1_U3342) );
  INV_X1 U8811 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6994) );
  INV_X1 U8812 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U8813 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9199), .ZN(n7542) );
  INV_X1 U8814 ( .A(n7542), .ZN(n6993) );
  OAI21_X1 U8815 ( .B1(n10099), .B2(n6994), .A(n6993), .ZN(n7001) );
  INV_X1 U8816 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6997) );
  MUX2_X1 U8817 ( .A(n6997), .B(P1_REG1_REG_7__SCAN_IN), .S(n7115), .Z(n6998)
         );
  NOR2_X1 U8818 ( .A1(n6999), .A2(n6998), .ZN(n7114) );
  AOI211_X1 U8819 ( .C1(n6999), .C2(n6998), .A(n10090), .B(n7114), .ZN(n7000)
         );
  AOI211_X1 U8820 ( .C1(n10072), .C2(n7115), .A(n7001), .B(n7000), .ZN(n7009)
         );
  INV_X1 U8821 ( .A(n7002), .ZN(n7003) );
  MUX2_X1 U8822 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7779), .S(n7115), .Z(n7006)
         );
  OAI211_X1 U8823 ( .C1(n7007), .C2(n7006), .A(n7108), .B(n10093), .ZN(n7008)
         );
  NAND2_X1 U8824 ( .A1(n7009), .A2(n7008), .ZN(P1_U3250) );
  CLKBUF_X2 U8825 ( .A(n7010), .Z(n7032) );
  INV_X1 U8826 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U8827 ( .A1(n7032), .A2(n7011), .ZN(P2_U3251) );
  INV_X1 U8828 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U8829 ( .A1(n7032), .A2(n7012), .ZN(P2_U3250) );
  INV_X1 U8830 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9396) );
  NOR2_X1 U8831 ( .A1(n7032), .A2(n9396), .ZN(P2_U3237) );
  INV_X1 U8832 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U8833 ( .A1(n7032), .A2(n7013), .ZN(P2_U3257) );
  INV_X1 U8834 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n7014) );
  NOR2_X1 U8835 ( .A1(n7032), .A2(n7014), .ZN(P2_U3263) );
  INV_X1 U8836 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9218) );
  NOR2_X1 U8837 ( .A1(n7032), .A2(n9218), .ZN(P2_U3262) );
  INV_X1 U8838 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n7015) );
  NOR2_X1 U8839 ( .A1(n7032), .A2(n7015), .ZN(P2_U3261) );
  INV_X1 U8840 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n7016) );
  NOR2_X1 U8841 ( .A1(n7032), .A2(n7016), .ZN(P2_U3243) );
  INV_X1 U8842 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n7017) );
  NOR2_X1 U8843 ( .A1(n7032), .A2(n7017), .ZN(P2_U3235) );
  INV_X1 U8844 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7018) );
  NOR2_X1 U8845 ( .A1(n7032), .A2(n7018), .ZN(P2_U3242) );
  INV_X1 U8846 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n7019) );
  NOR2_X1 U8847 ( .A1(n7032), .A2(n7019), .ZN(P2_U3239) );
  INV_X1 U8848 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9425) );
  NOR2_X1 U8849 ( .A1(n7032), .A2(n9425), .ZN(P2_U3240) );
  INV_X1 U8850 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n7020) );
  NOR2_X1 U8851 ( .A1(n7032), .A2(n7020), .ZN(P2_U3255) );
  INV_X1 U8852 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n7021) );
  NOR2_X1 U8853 ( .A1(n7032), .A2(n7021), .ZN(P2_U3254) );
  INV_X1 U8854 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7022) );
  NOR2_X1 U8855 ( .A1(n7032), .A2(n7022), .ZN(P2_U3253) );
  INV_X1 U8856 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7023) );
  NOR2_X1 U8857 ( .A1(n7032), .A2(n7023), .ZN(P2_U3252) );
  INV_X1 U8858 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n7024) );
  NOR2_X1 U8859 ( .A1(n7032), .A2(n7024), .ZN(P2_U3256) );
  INV_X1 U8860 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n7025) );
  NOR2_X1 U8861 ( .A1(n7032), .A2(n7025), .ZN(P2_U3238) );
  INV_X1 U8862 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n7026) );
  NOR2_X1 U8863 ( .A1(n7032), .A2(n7026), .ZN(P2_U3246) );
  INV_X1 U8864 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n7027) );
  NOR2_X1 U8865 ( .A1(n7032), .A2(n7027), .ZN(P2_U3245) );
  INV_X1 U8866 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9172) );
  NOR2_X1 U8867 ( .A1(n7032), .A2(n9172), .ZN(P2_U3241) );
  INV_X1 U8868 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n7028) );
  NOR2_X1 U8869 ( .A1(n7032), .A2(n7028), .ZN(P2_U3248) );
  INV_X1 U8870 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U8871 ( .A1(n7032), .A2(n7029), .ZN(P2_U3236) );
  INV_X1 U8872 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U8873 ( .A1(n7032), .A2(n7030), .ZN(P2_U3244) );
  INV_X1 U8874 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n7031) );
  NOR2_X1 U8875 ( .A1(n7032), .A2(n7031), .ZN(P2_U3234) );
  XNOR2_X1 U8876 ( .A(n7034), .B(n7033), .ZN(n7035) );
  XOR2_X1 U8877 ( .A(n7036), .B(n7035), .Z(n7045) );
  OR2_X1 U8878 ( .A1(n4549), .A2(P1_U3086), .ZN(n7649) );
  INV_X1 U8879 ( .A(n7649), .ZN(n7039) );
  AOI211_X1 U8880 ( .C1(n7039), .C2(n7038), .A(n10458), .B(n7037), .ZN(n7298)
         );
  NAND2_X1 U8881 ( .A1(n5891), .A2(n9666), .ZN(n7041) );
  NAND2_X1 U8882 ( .A1(n9986), .A2(n9667), .ZN(n7040) );
  AND2_X1 U8883 ( .A1(n7041), .A2(n7040), .ZN(n7492) );
  OAI22_X1 U8884 ( .A1(n7298), .A2(n7042), .B1(n7492), .B2(n10492), .ZN(n7043)
         );
  AOI21_X1 U8885 ( .B1(n5897), .B2(n10502), .A(n7043), .ZN(n7044) );
  OAI21_X1 U8886 ( .B1(n7045), .B2(n10535), .A(n7044), .ZN(P1_U3222) );
  NAND2_X1 U8887 ( .A1(n7345), .A2(n7046), .ZN(n7047) );
  NAND2_X1 U8888 ( .A1(n7048), .A2(n7047), .ZN(n7052) );
  NAND2_X1 U8889 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  INV_X1 U8890 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8891 ( .A1(n10683), .A2(n7053), .ZN(n7054) );
  OAI21_X1 U8892 ( .B1(n10683), .B2(n7055), .A(n7054), .ZN(P2_U3390) );
  XNOR2_X1 U8893 ( .A(n7056), .B(n8274), .ZN(n7365) );
  OAI21_X1 U8894 ( .B1(n8274), .B2(n7058), .A(n7057), .ZN(n7060) );
  OAI22_X1 U8895 ( .A1(n6304), .A2(n8953), .B1(n8675), .B2(n8993), .ZN(n7059)
         );
  AOI21_X1 U8896 ( .B1(n7060), .B2(n9017), .A(n7059), .ZN(n7061) );
  OAI21_X1 U8897 ( .B1(n7365), .B2(n7653), .A(n7061), .ZN(n7367) );
  OAI22_X1 U8898 ( .A1(n7365), .A2(n7731), .B1(n7366), .B2(n9454), .ZN(n7062)
         );
  NOR2_X1 U8899 ( .A1(n7367), .A2(n7062), .ZN(n10669) );
  INV_X1 U8900 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7063) );
  OR2_X1 U8901 ( .A1(n9456), .A2(n7063), .ZN(n7064) );
  OAI21_X1 U8902 ( .B1(n10669), .B2(n4671), .A(n7064), .ZN(P2_U3461) );
  AND2_X1 U8903 ( .A1(n8287), .A2(n8279), .ZN(n8276) );
  XNOR2_X1 U8904 ( .A(n7065), .B(n8276), .ZN(n7066) );
  OAI222_X1 U8905 ( .A1(n8993), .A2(n6304), .B1(n8953), .B2(n7324), .C1(n8990), 
        .C2(n7066), .ZN(n7894) );
  INV_X1 U8906 ( .A(n8276), .ZN(n8191) );
  XNOR2_X1 U8907 ( .A(n7067), .B(n8191), .ZN(n7898) );
  INV_X1 U8908 ( .A(n9449), .ZN(n9448) );
  INV_X1 U8909 ( .A(n7895), .ZN(n7170) );
  OAI22_X1 U8910 ( .A1(n7898), .A2(n9448), .B1(n7170), .B2(n9454), .ZN(n7068)
         );
  NOR2_X1 U8911 ( .A1(n7894), .A2(n7068), .ZN(n10672) );
  OR2_X1 U8912 ( .A1(n9456), .A2(n7069), .ZN(n7070) );
  OAI21_X1 U8913 ( .B1(n10672), .B2(n4671), .A(n7070), .ZN(P2_U3463) );
  OAI21_X1 U8914 ( .B1(n7072), .B2(n7075), .A(n7071), .ZN(n7078) );
  INV_X1 U8915 ( .A(n8677), .ZN(n7101) );
  INV_X1 U8916 ( .A(n4669), .ZN(n8269) );
  OAI22_X1 U8917 ( .A1(n7101), .A2(n8993), .B1(n8269), .B2(n8953), .ZN(n7077)
         );
  INV_X1 U8918 ( .A(n7073), .ZN(n7074) );
  AOI21_X1 U8919 ( .B1(n8261), .B2(n7075), .A(n7074), .ZN(n7381) );
  NOR2_X1 U8920 ( .A1(n7381), .A2(n7653), .ZN(n7076) );
  AOI211_X1 U8921 ( .C1(n9017), .C2(n7078), .A(n7077), .B(n7076), .ZN(n7374)
         );
  INV_X1 U8922 ( .A(n7374), .ZN(n7081) );
  OAI22_X1 U8923 ( .A1(n7381), .A2(n7731), .B1(n7079), .B2(n9454), .ZN(n7080)
         );
  NOR2_X1 U8924 ( .A1(n7081), .A2(n7080), .ZN(n10667) );
  OR2_X1 U8925 ( .A1(n9456), .A2(n6269), .ZN(n7082) );
  OAI21_X1 U8926 ( .B1(n10667), .B2(n4671), .A(n7082), .ZN(P2_U3460) );
  NAND2_X1 U8927 ( .A1(n7083), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8413) );
  INV_X1 U8928 ( .A(n7085), .ZN(n7087) );
  OAI22_X1 U8929 ( .A1(n8648), .A2(n7697), .B1(n8269), .B2(n8641), .ZN(n7086)
         );
  AOI211_X1 U8930 ( .C1(n8639), .C2(n8672), .A(n7087), .B(n7086), .ZN(n7096)
         );
  NAND2_X1 U8931 ( .A1(n7088), .A2(n8269), .ZN(n7089) );
  XNOR2_X1 U8932 ( .A(n7159), .B(n8673), .ZN(n7092) );
  AOI21_X1 U8933 ( .B1(n7091), .B2(n7092), .A(n8632), .ZN(n7094) );
  INV_X1 U8934 ( .A(n7092), .ZN(n7093) );
  NAND2_X1 U8935 ( .A1(n7094), .A2(n7161), .ZN(n7095) );
  OAI211_X1 U8936 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8524), .A(n7096), .B(
        n7095), .ZN(P2_U3158) );
  INV_X1 U8937 ( .A(n7097), .ZN(n7098) );
  AOI21_X1 U8938 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n7106) );
  OAI22_X1 U8939 ( .A1(n8627), .A2(n8269), .B1(n7101), .B2(n8641), .ZN(n7104)
         );
  NOR2_X1 U8940 ( .A1(n7102), .A2(n7376), .ZN(n7103) );
  AOI211_X1 U8941 ( .C1(n7378), .C2(n8629), .A(n7104), .B(n7103), .ZN(n7105)
         );
  OAI21_X1 U8942 ( .B1(n8632), .B2(n7106), .A(n7105), .ZN(P2_U3162) );
  NOR2_X1 U8943 ( .A1(n7252), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7107) );
  AOI21_X1 U8944 ( .B1(n7252), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7107), .ZN(
        n7113) );
  OAI21_X1 U8945 ( .B1(n7109), .B2(n7779), .A(n7108), .ZN(n10020) );
  INV_X1 U8946 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7110) );
  MUX2_X1 U8947 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7110), .S(n10017), .Z(n10019) );
  NAND2_X1 U8948 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  INV_X1 U8949 ( .A(n10018), .ZN(n7111) );
  NAND2_X1 U8950 ( .A1(n7112), .A2(n7113), .ZN(n7251) );
  OAI21_X1 U8951 ( .B1(n7113), .B2(n7112), .A(n7251), .ZN(n7126) );
  AOI21_X1 U8952 ( .B1(n7115), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7114), .ZN(
        n10013) );
  INV_X1 U8953 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7116) );
  MUX2_X1 U8954 ( .A(n7116), .B(P1_REG1_REG_8__SCAN_IN), .S(n10017), .Z(n10012) );
  NOR2_X1 U8955 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  MUX2_X1 U8956 ( .A(n7117), .B(P1_REG1_REG_9__SCAN_IN), .S(n7124), .Z(n7118)
         );
  NAND2_X1 U8957 ( .A1(n7119), .A2(n7118), .ZN(n7248) );
  OAI21_X1 U8958 ( .B1(n7119), .B2(n7118), .A(n7248), .ZN(n7120) );
  NAND2_X1 U8959 ( .A1(n7120), .A2(n10087), .ZN(n7123) );
  NOR2_X1 U8960 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7121), .ZN(n7741) );
  AOI21_X1 U8961 ( .B1(n10055), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7741), .ZN(
        n7122) );
  OAI211_X1 U8962 ( .C1(n10089), .C2(n7124), .A(n7123), .B(n7122), .ZN(n7125)
         );
  AOI21_X1 U8963 ( .B1(n10093), .B2(n7126), .A(n7125), .ZN(n7127) );
  INV_X1 U8964 ( .A(n7127), .ZN(P1_U3252) );
  INV_X1 U8965 ( .A(n7703), .ZN(n7133) );
  OAI21_X1 U8966 ( .B1(n7130), .B2(n7129), .A(n7128), .ZN(n7131) );
  INV_X1 U8967 ( .A(n8993), .ZN(n9012) );
  AOI222_X1 U8968 ( .A1(n9017), .A2(n7131), .B1(n4669), .B2(n9012), .C1(n8672), 
        .C2(n9014), .ZN(n7699) );
  OAI21_X1 U8969 ( .B1(n7697), .B2(n9454), .A(n7699), .ZN(n7132) );
  AOI21_X1 U8970 ( .B1(n7133), .B2(n9449), .A(n7132), .ZN(n10670) );
  OR2_X1 U8971 ( .A1(n9456), .A2(n6291), .ZN(n7134) );
  OAI21_X1 U8972 ( .B1(n10670), .B2(n4671), .A(n7134), .ZN(P2_U3462) );
  INV_X1 U8973 ( .A(n7137), .ZN(n7138) );
  AOI21_X1 U8974 ( .B1(n7135), .B2(n7136), .A(n7138), .ZN(n7142) );
  AOI22_X1 U8975 ( .A1(n9667), .A2(n9984), .B1(n9987), .B2(n9666), .ZN(n7183)
         );
  OAI22_X1 U8976 ( .A1(n7298), .A2(n7502), .B1(n7183), .B2(n10492), .ZN(n7139)
         );
  AOI21_X1 U8977 ( .B1(n7140), .B2(n10502), .A(n7139), .ZN(n7141) );
  OAI21_X1 U8978 ( .B1(n7142), .B2(n10535), .A(n7141), .ZN(P1_U3237) );
  INV_X1 U8979 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U8980 ( .A1(n7143), .A2(n5049), .ZN(n7219) );
  AOI21_X1 U8981 ( .B1(n7418), .B2(n7144), .A(n7216), .ZN(n7158) );
  INV_X1 U8982 ( .A(n7145), .ZN(n7147) );
  AOI21_X1 U8983 ( .B1(n7148), .B2(n7147), .A(n7146), .ZN(n7223) );
  MUX2_X1 U8984 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8798), .Z(n7221) );
  XOR2_X1 U8985 ( .A(n7151), .B(n7221), .Z(n7222) );
  XNOR2_X1 U8986 ( .A(n7223), .B(n7222), .ZN(n7149) );
  NAND2_X1 U8987 ( .A1(n7149), .A2(n10652), .ZN(n7157) );
  OAI21_X1 U8988 ( .B1(n7152), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7231), .ZN(
        n7155) );
  INV_X1 U8989 ( .A(n8841), .ZN(n10664) );
  NAND2_X1 U8990 ( .A1(n8839), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7153) );
  NAND2_X1 U8991 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7430) );
  OAI211_X1 U8992 ( .C1(n8837), .C2(n5049), .A(n7153), .B(n7430), .ZN(n7154)
         );
  AOI21_X1 U8993 ( .B1(n7155), .B2(n10664), .A(n7154), .ZN(n7156) );
  OAI211_X1 U8994 ( .C1(n7158), .C2(n8806), .A(n7157), .B(n7156), .ZN(P2_U3189) );
  NAND2_X1 U8995 ( .A1(n7159), .A2(n8673), .ZN(n7160) );
  XNOR2_X1 U8996 ( .A(n7162), .B(n7895), .ZN(n7163) );
  NAND2_X1 U8997 ( .A1(n7163), .A2(n7282), .ZN(n7274) );
  INV_X1 U8998 ( .A(n7163), .ZN(n7164) );
  NAND2_X1 U8999 ( .A1(n7164), .A2(n8672), .ZN(n7165) );
  AND2_X1 U9000 ( .A1(n7274), .A2(n7165), .ZN(n7166) );
  OAI21_X1 U9001 ( .B1(n7167), .B2(n7166), .A(n7275), .ZN(n7168) );
  NAND2_X1 U9002 ( .A1(n7168), .A2(n8635), .ZN(n7174) );
  INV_X1 U9003 ( .A(n7169), .ZN(n7172) );
  OAI22_X1 U9004 ( .A1(n8648), .A2(n7170), .B1(n6304), .B2(n8641), .ZN(n7171)
         );
  AOI211_X1 U9005 ( .C1(n8639), .C2(n8671), .A(n7172), .B(n7171), .ZN(n7173)
         );
  OAI211_X1 U9006 ( .C1(n7897), .C2(n8524), .A(n7174), .B(n7173), .ZN(P2_U3170) );
  INV_X1 U9007 ( .A(n7175), .ZN(n7178) );
  INV_X1 U9008 ( .A(n8057), .ZN(n10032) );
  OAI222_X1 U9009 ( .A1(n10470), .A2(n7176), .B1(n10472), .B2(n7178), .C1(
        n10032), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI222_X1 U9010 ( .A1(P2_U3151), .A2(n4659), .B1(n9524), .B2(n7178), .C1(
        n7177), .C2(n8484), .ZN(P2_U3280) );
  INV_X1 U9011 ( .A(n7179), .ZN(n7182) );
  INV_X1 U9012 ( .A(n8054), .ZN(n7867) );
  OAI222_X1 U9013 ( .A1(n10470), .A2(n7180), .B1(n10472), .B2(n7182), .C1(
        P1_U3086), .C2(n7867), .ZN(P1_U3341) );
  OAI222_X1 U9014 ( .A1(n8732), .A2(P2_U3151), .B1(n9524), .B2(n7182), .C1(
        n7181), .C2(n8484), .ZN(P2_U3281) );
  XNOR2_X1 U9015 ( .A(n9701), .B(n7188), .ZN(n7184) );
  OAI21_X1 U9016 ( .B1(n7184), .B2(n10302), .A(n7183), .ZN(n7499) );
  INV_X1 U9017 ( .A(n7200), .ZN(n7187) );
  AOI21_X1 U9018 ( .B1(n5408), .B2(n7185), .A(n7503), .ZN(n7186) );
  NOR3_X1 U9019 ( .A1(n7187), .A2(n7186), .A3(n10308), .ZN(n7505) );
  NOR2_X1 U9020 ( .A1(n7499), .A2(n7505), .ZN(n7449) );
  INV_X1 U9021 ( .A(n10381), .ZN(n10391) );
  OR2_X1 U9022 ( .A1(n7189), .A2(n7188), .ZN(n7190) );
  NAND2_X1 U9023 ( .A1(n7191), .A2(n7190), .ZN(n7498) );
  INV_X1 U9024 ( .A(n10392), .ZN(n10356) );
  OAI22_X1 U9025 ( .A1(n10356), .A2(n7503), .B1(n10643), .B2(n7192), .ZN(n7193) );
  AOI21_X1 U9026 ( .B1(n10391), .B2(n7498), .A(n7193), .ZN(n7194) );
  OAI21_X1 U9027 ( .B1(n7449), .B2(n10641), .A(n7194), .ZN(P1_U3524) );
  OAI21_X1 U9028 ( .B1(n7196), .B2(n9684), .A(n7195), .ZN(n7199) );
  NAND2_X1 U9029 ( .A1(n9986), .A2(n9666), .ZN(n7198) );
  NAND2_X1 U9030 ( .A1(n9983), .A2(n9667), .ZN(n7197) );
  NAND2_X1 U9031 ( .A1(n7198), .A2(n7197), .ZN(n9550) );
  AOI21_X1 U9032 ( .B1(n7199), .B2(n10285), .A(n9550), .ZN(n7438) );
  AOI21_X1 U9033 ( .B1(n7200), .B2(n4561), .A(n10308), .ZN(n7201) );
  NAND2_X1 U9034 ( .A1(n7201), .A2(n7290), .ZN(n7440) );
  AND2_X1 U9035 ( .A1(n7438), .A2(n7440), .ZN(n7454) );
  OAI21_X1 U9036 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7452) );
  OAI22_X1 U9037 ( .A1(n10356), .A2(n7450), .B1(n10643), .B2(n6710), .ZN(n7205) );
  AOI21_X1 U9038 ( .B1(n7452), .B2(n10391), .A(n7205), .ZN(n7206) );
  OAI21_X1 U9039 ( .B1(n7454), .B2(n10641), .A(n7206), .ZN(P1_U3525) );
  AND2_X1 U9040 ( .A1(n8285), .A2(n8282), .ZN(n8195) );
  XNOR2_X1 U9041 ( .A(n7207), .B(n8195), .ZN(n7208) );
  OAI222_X1 U9042 ( .A1(n8953), .A2(n8247), .B1(n8993), .B2(n7324), .C1(n8990), 
        .C2(n7208), .ZN(n7655) );
  NAND2_X1 U9043 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  XOR2_X1 U9044 ( .A(n8195), .B(n7211), .Z(n7663) );
  INV_X1 U9045 ( .A(n7660), .ZN(n7329) );
  OAI22_X1 U9046 ( .A1(n7663), .A2(n9448), .B1(n7329), .B2(n9454), .ZN(n7212)
         );
  NOR2_X1 U9047 ( .A1(n7655), .A2(n7212), .ZN(n10675) );
  INV_X1 U9048 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7213) );
  OR2_X1 U9049 ( .A1(n9456), .A2(n7213), .ZN(n7214) );
  OAI21_X1 U9050 ( .B1(n10675), .B2(n4671), .A(n7214), .ZN(P2_U3465) );
  INV_X1 U9051 ( .A(n7219), .ZN(n7215) );
  XNOR2_X1 U9052 ( .A(n7228), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7217) );
  NOR3_X1 U9053 ( .A1(n7216), .A2(n7215), .A3(n7217), .ZN(n7220) );
  INV_X1 U9054 ( .A(n7217), .ZN(n7218) );
  NOR2_X1 U9055 ( .A1(n7220), .A2(n7471), .ZN(n7238) );
  OAI22_X1 U9056 ( .A1(n7223), .A2(n7222), .B1(n7221), .B2(n5049), .ZN(n7225)
         );
  MUX2_X1 U9057 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8798), .Z(n7463) );
  XNOR2_X1 U9058 ( .A(n7463), .B(n7228), .ZN(n7224) );
  NAND2_X1 U9059 ( .A1(n7225), .A2(n7224), .ZN(n7464) );
  OAI21_X1 U9060 ( .B1(n7225), .B2(n7224), .A(n7464), .ZN(n7226) );
  NAND2_X1 U9061 ( .A1(n7226), .A2(n10652), .ZN(n7237) );
  NAND2_X1 U9062 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7556) );
  OAI21_X1 U9063 ( .B1(n8837), .B2(n7472), .A(n7556), .ZN(n7235) );
  INV_X1 U9064 ( .A(n7227), .ZN(n7229) );
  MUX2_X1 U9065 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7666), .S(n7228), .Z(n7230)
         );
  INV_X1 U9066 ( .A(n7461), .ZN(n7233) );
  NAND3_X1 U9067 ( .A1(n7231), .A2(n7230), .A3(n7229), .ZN(n7232) );
  AOI21_X1 U9068 ( .B1(n7233), .B2(n7232), .A(n8841), .ZN(n7234) );
  AOI211_X1 U9069 ( .C1(n8839), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7235), .B(
        n7234), .ZN(n7236) );
  OAI211_X1 U9070 ( .C1(n7238), .C2(n8806), .A(n7237), .B(n7236), .ZN(P2_U3190) );
  INV_X1 U9071 ( .A(n7239), .ZN(n7241) );
  AOI21_X1 U9072 ( .B1(n7241), .B2(n9811), .A(n7240), .ZN(n7246) );
  NOR2_X1 U9073 ( .A1(n10275), .A2(n10308), .ZN(n10110) );
  OAI21_X1 U9074 ( .B1(n10278), .B2(n10110), .A(n7488), .ZN(n7245) );
  OAI22_X1 U9075 ( .A1(n10241), .A2(n7242), .B1(n7297), .B2(n10270), .ZN(n7243) );
  INV_X1 U9076 ( .A(n7243), .ZN(n7244) );
  OAI211_X1 U9077 ( .C1(n10563), .C2(n7246), .A(n7245), .B(n7244), .ZN(
        P1_U3293) );
  INV_X1 U9078 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7247) );
  MUX2_X1 U9079 ( .A(n7247), .B(P1_REG1_REG_10__SCAN_IN), .S(n7356), .Z(n7250)
         );
  OAI21_X1 U9080 ( .B1(n7252), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7248), .ZN(
        n7249) );
  NOR2_X1 U9081 ( .A1(n7249), .A2(n7250), .ZN(n7351) );
  AOI211_X1 U9082 ( .C1(n7250), .C2(n7249), .A(n10090), .B(n7351), .ZN(n7259)
         );
  OAI21_X1 U9083 ( .B1(n7252), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7251), .ZN(
        n7255) );
  INV_X1 U9084 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7253) );
  MUX2_X1 U9085 ( .A(n7253), .B(P1_REG2_REG_10__SCAN_IN), .S(n7356), .Z(n7254)
         );
  NOR2_X1 U9086 ( .A1(n7254), .A2(n7255), .ZN(n7355) );
  AOI211_X1 U9087 ( .C1(n7255), .C2(n7254), .A(n7355), .B(n10037), .ZN(n7258)
         );
  INV_X1 U9088 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U9089 ( .A1(n10072), .A2(n7356), .ZN(n7256) );
  NAND2_X1 U9090 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10476) );
  OAI211_X1 U9091 ( .C1(n8144), .C2(n10099), .A(n7256), .B(n10476), .ZN(n7257)
         );
  OR3_X1 U9092 ( .A1(n7259), .A2(n7258), .A3(n7257), .ZN(P1_U3253) );
  NAND2_X1 U9093 ( .A1(n7262), .A2(n10449), .ZN(n7263) );
  OAI21_X1 U9094 ( .B1(n10449), .B2(n5413), .A(n7263), .ZN(P1_U3453) );
  XNOR2_X1 U9095 ( .A(n7264), .B(n7266), .ZN(n7388) );
  NOR2_X1 U9096 ( .A1(n7388), .A2(n7731), .ZN(n7270) );
  XNOR2_X1 U9097 ( .A(n7265), .B(n7266), .ZN(n7268) );
  OAI22_X1 U9098 ( .A1(n7431), .A2(n8953), .B1(n7282), .B2(n8993), .ZN(n7267)
         );
  AOI21_X1 U9099 ( .B1(n7268), .B2(n9017), .A(n7267), .ZN(n7269) );
  OAI21_X1 U9100 ( .B1(n7653), .B2(n7388), .A(n7269), .ZN(n7382) );
  AOI211_X1 U9101 ( .C1(n9443), .C2(n7385), .A(n7270), .B(n7382), .ZN(n10673)
         );
  OR2_X1 U9102 ( .A1(n10673), .A2(n4671), .ZN(n7271) );
  OAI21_X1 U9103 ( .B1(n9456), .B2(n8687), .A(n7271), .ZN(P2_U3464) );
  INV_X1 U9104 ( .A(n7275), .ZN(n7273) );
  INV_X1 U9105 ( .A(n7274), .ZN(n7272) );
  INV_X4 U9106 ( .A(n8517), .ZN(n8546) );
  XNOR2_X1 U9107 ( .A(n8546), .B(n7385), .ZN(n7316) );
  XNOR2_X1 U9108 ( .A(n7316), .B(n8671), .ZN(n7276) );
  NOR3_X1 U9109 ( .A1(n7273), .A2(n7272), .A3(n7276), .ZN(n7279) );
  NAND2_X1 U9110 ( .A1(n7277), .A2(n7276), .ZN(n7318) );
  INV_X1 U9111 ( .A(n7318), .ZN(n7278) );
  OAI21_X1 U9112 ( .B1(n7279), .B2(n7278), .A(n8635), .ZN(n7285) );
  NAND2_X1 U9113 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8682) );
  INV_X1 U9114 ( .A(n8682), .ZN(n7280) );
  AOI21_X1 U9115 ( .B1(n8639), .B2(n8670), .A(n7280), .ZN(n7281) );
  OAI21_X1 U9116 ( .B1(n7282), .B2(n8641), .A(n7281), .ZN(n7283) );
  AOI21_X1 U9117 ( .B1(n7385), .B2(n8629), .A(n7283), .ZN(n7284) );
  OAI211_X1 U9118 ( .C1(n7383), .C2(n8524), .A(n7285), .B(n7284), .ZN(P2_U3167) );
  XNOR2_X1 U9119 ( .A(n7286), .B(n7292), .ZN(n7289) );
  NAND2_X1 U9120 ( .A1(n9984), .A2(n9666), .ZN(n7288) );
  NAND2_X1 U9121 ( .A1(n9982), .A2(n9667), .ZN(n7287) );
  AND2_X1 U9122 ( .A1(n7288), .A2(n7287), .ZN(n7311) );
  OAI21_X1 U9123 ( .B1(n7289), .B2(n10302), .A(n7311), .ZN(n7516) );
  AOI211_X1 U9124 ( .C1(n7313), .C2(n7290), .A(n10308), .B(n4580), .ZN(n7515)
         );
  NOR2_X1 U9125 ( .A1(n7516), .A2(n7515), .ZN(n7446) );
  OAI21_X1 U9126 ( .B1(n7293), .B2(n7292), .A(n7291), .ZN(n7509) );
  OAI22_X1 U9127 ( .A1(n10356), .A2(n7513), .B1(n10643), .B2(n9397), .ZN(n7294) );
  AOI21_X1 U9128 ( .B1(n7509), .B2(n10391), .A(n7294), .ZN(n7295) );
  OAI21_X1 U9129 ( .B1(n7446), .B2(n10641), .A(n7295), .ZN(P1_U3526) );
  OAI22_X1 U9130 ( .A1(n7298), .A2(n7297), .B1(n10492), .B2(n7296), .ZN(n7299)
         );
  AOI21_X1 U9131 ( .B1(n7488), .B2(n10515), .A(n7299), .ZN(n7300) );
  OAI21_X1 U9132 ( .B1(n10535), .B2(n7301), .A(n7300), .ZN(P1_U3232) );
  INV_X1 U9133 ( .A(n7302), .ZN(n7304) );
  OAI222_X1 U9134 ( .A1(n8772), .A2(P2_U3151), .B1(n9524), .B2(n7304), .C1(
        n7303), .C2(n8484), .ZN(P2_U3279) );
  INV_X1 U9135 ( .A(n10049), .ZN(n10045) );
  OAI222_X1 U9136 ( .A1(n10470), .A2(n7305), .B1(n10472), .B2(n7304), .C1(
        P1_U3086), .C2(n10045), .ZN(P1_U3339) );
  AOI21_X1 U9137 ( .B1(n7307), .B2(n7306), .A(n10535), .ZN(n7309) );
  NAND2_X1 U9138 ( .A1(n7309), .A2(n7308), .ZN(n7315) );
  OAI21_X1 U9139 ( .B1(n10492), .B2(n7311), .A(n7310), .ZN(n7312) );
  AOI21_X1 U9140 ( .B1(n7313), .B2(n10515), .A(n7312), .ZN(n7314) );
  OAI211_X1 U9141 ( .C1(n10547), .C2(n7510), .A(n7315), .B(n7314), .ZN(
        P1_U3230) );
  NAND2_X1 U9142 ( .A1(n7316), .A2(n7324), .ZN(n7317) );
  XNOR2_X1 U9143 ( .A(n8546), .B(n7660), .ZN(n7419) );
  XNOR2_X1 U9144 ( .A(n7419), .B(n8670), .ZN(n7319) );
  OAI211_X1 U9145 ( .C1(n7320), .C2(n7319), .A(n7422), .B(n8635), .ZN(n7328)
         );
  INV_X1 U9146 ( .A(n7658), .ZN(n7326) );
  INV_X1 U9147 ( .A(n7321), .ZN(n7322) );
  AOI21_X1 U9148 ( .B1(n8639), .B2(n8669), .A(n7322), .ZN(n7323) );
  OAI21_X1 U9149 ( .B1(n7324), .B2(n8641), .A(n7323), .ZN(n7325) );
  AOI21_X1 U9150 ( .B1(n8645), .B2(n7326), .A(n7325), .ZN(n7327) );
  OAI211_X1 U9151 ( .C1(n7329), .C2(n8648), .A(n7328), .B(n7327), .ZN(P2_U3179) );
  INV_X1 U9152 ( .A(n8797), .ZN(n8783) );
  INV_X1 U9153 ( .A(n7330), .ZN(n7332) );
  OAI222_X1 U9154 ( .A1(P2_U3151), .A2(n8783), .B1(n9524), .B2(n7332), .C1(
        n7331), .C2(n8484), .ZN(P2_U3278) );
  INV_X1 U9155 ( .A(n10064), .ZN(n10057) );
  OAI222_X1 U9156 ( .A1(n10470), .A2(n7333), .B1(P1_U3086), .B2(n10057), .C1(
        n7332), .C2(n10472), .ZN(P1_U3338) );
  INV_X1 U9157 ( .A(n7334), .ZN(n7337) );
  AOI22_X1 U9158 ( .A1(n10075), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10464), .ZN(n7335) );
  OAI21_X1 U9159 ( .B1(n7337), .B2(n10472), .A(n7335), .ZN(P1_U3337) );
  AOI22_X1 U9160 ( .A1(n8833), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9522), .ZN(n7336) );
  OAI21_X1 U9161 ( .B1(n7337), .B2(n9524), .A(n7336), .ZN(P2_U3277) );
  INV_X1 U9162 ( .A(n7338), .ZN(n7342) );
  NOR2_X1 U9163 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  NOR2_X2 U9164 ( .A1(n7343), .A2(n8905), .ZN(n9023) );
  AOI22_X1 U9165 ( .A1(n9023), .A2(n7344), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8999), .ZN(n7350) );
  INV_X1 U9166 ( .A(n7345), .ZN(n7346) );
  NOR3_X1 U9167 ( .A1(n7346), .A2(n8188), .A3(n9443), .ZN(n7347) );
  OAI21_X1 U9168 ( .B1(n7348), .B2(n7347), .A(n9020), .ZN(n7349) );
  OAI211_X1 U9169 ( .C1(n6282), .C2(n9020), .A(n7350), .B(n7349), .ZN(P2_U3233) );
  INV_X1 U9170 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7352) );
  MUX2_X1 U9171 ( .A(n7352), .B(P1_REG1_REG_11__SCAN_IN), .S(n7395), .Z(n7353)
         );
  NOR2_X1 U9172 ( .A1(n7354), .A2(n7353), .ZN(n7389) );
  AOI211_X1 U9173 ( .C1(n7354), .C2(n7353), .A(n10090), .B(n7389), .ZN(n7363)
         );
  AOI22_X1 U9174 ( .A1(n7395), .A2(n7926), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7357), .ZN(n7358) );
  NOR2_X1 U9175 ( .A1(n7359), .A2(n7358), .ZN(n7394) );
  AOI211_X1 U9176 ( .C1(n7359), .C2(n7358), .A(n7394), .B(n10037), .ZN(n7362)
         );
  INV_X1 U9177 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U9178 ( .A1(n10072), .A2(n7395), .ZN(n7360) );
  NAND2_X1 U9179 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10506) );
  OAI211_X1 U9180 ( .C1(n8123), .C2(n10099), .A(n7360), .B(n10506), .ZN(n7361)
         );
  OR3_X1 U9181 ( .A1(n7363), .A2(n7362), .A3(n7361), .ZN(P1_U3254) );
  OR2_X1 U9182 ( .A1(n6622), .A2(n7364), .ZN(n7652) );
  INV_X1 U9183 ( .A(n7652), .ZN(n7373) );
  INV_X1 U9184 ( .A(n7365), .ZN(n7369) );
  OAI22_X1 U9185 ( .A1(n9018), .A2(n6939), .B1(n7366), .B2(n8905), .ZN(n7368)
         );
  AOI211_X1 U9186 ( .C1(n7373), .C2(n7369), .A(n7368), .B(n7367), .ZN(n7370)
         );
  MUX2_X1 U9187 ( .A(n7371), .B(n7370), .S(n9020), .Z(n7372) );
  INV_X1 U9188 ( .A(n7372), .ZN(P2_U3231) );
  NAND2_X1 U9189 ( .A1(n9020), .A2(n7373), .ZN(n7578) );
  MUX2_X1 U9190 ( .A(n7375), .B(n7374), .S(n9020), .Z(n7380) );
  NOR2_X1 U9191 ( .A1(n9018), .A2(n7376), .ZN(n7377) );
  AOI21_X1 U9192 ( .B1(n9023), .B2(n7378), .A(n7377), .ZN(n7379) );
  OAI211_X1 U9193 ( .C1(n7381), .C2(n7578), .A(n7380), .B(n7379), .ZN(P2_U3232) );
  NAND2_X1 U9194 ( .A1(n7382), .A2(n9020), .ZN(n7387) );
  OAI22_X1 U9195 ( .A1(n9020), .A2(n6333), .B1(n7383), .B2(n9018), .ZN(n7384)
         );
  AOI21_X1 U9196 ( .B1(n9023), .B2(n7385), .A(n7384), .ZN(n7386) );
  OAI211_X1 U9197 ( .C1(n7388), .C2(n7578), .A(n7387), .B(n7386), .ZN(P2_U3228) );
  INV_X1 U9198 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7390) );
  AOI22_X1 U9199 ( .A1(n7709), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7390), .B2(
        n7401), .ZN(n7391) );
  NAND2_X1 U9200 ( .A1(n7392), .A2(n7391), .ZN(n7708) );
  OAI21_X1 U9201 ( .B1(n7392), .B2(n7391), .A(n7708), .ZN(n7403) );
  NOR2_X1 U9202 ( .A1(n7709), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7393) );
  AOI21_X1 U9203 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7709), .A(n7393), .ZN(
        n7397) );
  AOI21_X1 U9204 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7395), .A(n7394), .ZN(
        n7396) );
  NAND2_X1 U9205 ( .A1(n7397), .A2(n7396), .ZN(n7704) );
  OAI21_X1 U9206 ( .B1(n7397), .B2(n7396), .A(n7704), .ZN(n7398) );
  NAND2_X1 U9207 ( .A1(n7398), .A2(n10093), .ZN(n7400) );
  AND2_X1 U9208 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10489) );
  AOI21_X1 U9209 ( .B1(n10055), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10489), .ZN(
        n7399) );
  OAI211_X1 U9210 ( .C1(n10089), .C2(n7401), .A(n7400), .B(n7399), .ZN(n7402)
         );
  AOI21_X1 U9211 ( .B1(n10087), .B2(n7403), .A(n7402), .ZN(n7404) );
  INV_X1 U9212 ( .A(n7404), .ZN(P1_U3255) );
  XNOR2_X1 U9213 ( .A(n7405), .B(n6364), .ZN(n7411) );
  INV_X1 U9214 ( .A(n7411), .ZN(n7554) );
  NOR2_X1 U9215 ( .A1(n7554), .A2(n7731), .ZN(n7416) );
  NAND2_X1 U9216 ( .A1(n7407), .A2(n8298), .ZN(n7408) );
  NAND2_X1 U9217 ( .A1(n7406), .A2(n7408), .ZN(n7409) );
  NAND2_X1 U9218 ( .A1(n7409), .A2(n9017), .ZN(n7414) );
  AOI22_X1 U9219 ( .A1(n9014), .A2(n8668), .B1(n8670), .B2(n9012), .ZN(n7413)
         );
  INV_X1 U9220 ( .A(n7653), .ZN(n7410) );
  NAND2_X1 U9221 ( .A1(n7411), .A2(n7410), .ZN(n7412) );
  AND3_X1 U9222 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(n7549) );
  INV_X1 U9223 ( .A(n7549), .ZN(n7415) );
  AOI211_X1 U9224 ( .C1(n9443), .C2(n8248), .A(n7416), .B(n7415), .ZN(n10677)
         );
  OR2_X1 U9225 ( .A1(n10677), .A2(n4671), .ZN(n7417) );
  OAI21_X1 U9226 ( .B1(n9456), .B2(n7418), .A(n7417), .ZN(P2_U3466) );
  INV_X1 U9227 ( .A(n7419), .ZN(n7420) );
  NAND2_X1 U9228 ( .A1(n7420), .A2(n8670), .ZN(n7421) );
  XNOR2_X1 U9229 ( .A(n8248), .B(n8546), .ZN(n7423) );
  NAND2_X1 U9230 ( .A1(n7423), .A2(n8247), .ZN(n7563) );
  INV_X1 U9231 ( .A(n7423), .ZN(n7424) );
  NAND2_X1 U9232 ( .A1(n7424), .A2(n8669), .ZN(n7425) );
  NAND2_X1 U9233 ( .A1(n7563), .A2(n7425), .ZN(n7428) );
  INV_X1 U9234 ( .A(n7428), .ZN(n7426) );
  INV_X1 U9235 ( .A(n7560), .ZN(n7427) );
  AOI21_X1 U9236 ( .B1(n7429), .B2(n7428), .A(n7427), .ZN(n7437) );
  INV_X1 U9237 ( .A(n7430), .ZN(n7433) );
  NOR2_X1 U9238 ( .A1(n8641), .A2(n7431), .ZN(n7432) );
  AOI211_X1 U9239 ( .C1(n8639), .C2(n8668), .A(n7433), .B(n7432), .ZN(n7434)
         );
  OAI21_X1 U9240 ( .B1(n8524), .B2(n7550), .A(n7434), .ZN(n7435) );
  AOI21_X1 U9241 ( .B1(n8248), .B2(n8629), .A(n7435), .ZN(n7436) );
  OAI21_X1 U9242 ( .B1(n7437), .B2(n8632), .A(n7436), .ZN(P2_U3153) );
  MUX2_X1 U9243 ( .A(n6706), .B(n7438), .S(n5878), .Z(n7443) );
  AOI22_X1 U9244 ( .A1(n10278), .A2(n4561), .B1(n5460), .B2(n10551), .ZN(n7439) );
  OAI21_X1 U9245 ( .B1(n10275), .B2(n7440), .A(n7439), .ZN(n7441) );
  AOI21_X1 U9246 ( .B1(n7452), .B2(n10560), .A(n7441), .ZN(n7442) );
  NAND2_X1 U9247 ( .A1(n7443), .A2(n7442), .ZN(P1_U3290) );
  INV_X1 U9248 ( .A(n10447), .ZN(n10451) );
  OAI22_X1 U9249 ( .A1(n10425), .A2(n7513), .B1(n10449), .B2(n5463), .ZN(n7444) );
  AOI21_X1 U9250 ( .B1(n7509), .B2(n10451), .A(n7444), .ZN(n7445) );
  OAI21_X1 U9251 ( .B1(n7446), .B2(n10634), .A(n7445), .ZN(P1_U3465) );
  OAI22_X1 U9252 ( .A1(n10425), .A2(n7503), .B1(n10449), .B2(n5426), .ZN(n7447) );
  AOI21_X1 U9253 ( .B1(n10451), .B2(n7498), .A(n7447), .ZN(n7448) );
  OAI21_X1 U9254 ( .B1(n7449), .B2(n10634), .A(n7448), .ZN(P1_U3459) );
  OAI22_X1 U9255 ( .A1(n10425), .A2(n7450), .B1(n10449), .B2(n5443), .ZN(n7451) );
  AOI21_X1 U9256 ( .B1(n7452), .B2(n10451), .A(n7451), .ZN(n7453) );
  OAI21_X1 U9257 ( .B1(n7454), .B2(n10634), .A(n7453), .ZN(P1_U3462) );
  INV_X1 U9258 ( .A(n8243), .ZN(n8245) );
  NAND2_X1 U9259 ( .A1(n8245), .A2(n8250), .ZN(n8197) );
  XOR2_X1 U9260 ( .A(n7455), .B(n8197), .Z(n7456) );
  OAI222_X1 U9261 ( .A1(n8993), .A2(n8247), .B1(n8953), .B2(n7885), .C1(n8990), 
        .C2(n7456), .ZN(n7664) );
  XOR2_X1 U9262 ( .A(n8197), .B(n7457), .Z(n7672) );
  OAI22_X1 U9263 ( .A1(n7672), .A2(n9448), .B1(n7458), .B2(n9454), .ZN(n7459)
         );
  NOR2_X1 U9264 ( .A1(n7664), .A2(n7459), .ZN(n10678) );
  OR2_X1 U9265 ( .A1(n9456), .A2(n4748), .ZN(n7460) );
  OAI21_X1 U9266 ( .B1(n10678), .B2(n4671), .A(n7460), .ZN(P2_U3467) );
  XNOR2_X1 U9267 ( .A(n7612), .B(n7613), .ZN(n7462) );
  AOI21_X1 U9268 ( .B1(n7462), .B2(n6390), .A(n7614), .ZN(n7478) );
  MUX2_X1 U9269 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8798), .Z(n7621) );
  XNOR2_X1 U9270 ( .A(n7621), .B(n7613), .ZN(n7467) );
  OR2_X1 U9271 ( .A1(n7463), .A2(n7472), .ZN(n7465) );
  NAND2_X1 U9272 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NAND2_X1 U9273 ( .A1(n7467), .A2(n7466), .ZN(n7622) );
  OAI21_X1 U9274 ( .B1(n7467), .B2(n7466), .A(n7622), .ZN(n7468) );
  NAND2_X1 U9275 ( .A1(n10652), .A2(n7468), .ZN(n7470) );
  AND2_X1 U9276 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7641) );
  INV_X1 U9277 ( .A(n7641), .ZN(n7469) );
  OAI211_X1 U9278 ( .C1(n8837), .C2(n7620), .A(n7470), .B(n7469), .ZN(n7476)
         );
  NOR2_X1 U9279 ( .A1(n6387), .A2(n7473), .ZN(n7606) );
  AOI21_X1 U9280 ( .B1(n6387), .B2(n7473), .A(n7606), .ZN(n7474) );
  NOR2_X1 U9281 ( .A1(n7474), .A2(n8806), .ZN(n7475) );
  AOI211_X1 U9282 ( .C1(n8839), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7476), .B(
        n7475), .ZN(n7477) );
  OAI21_X1 U9283 ( .B1(n7478), .B2(n8841), .A(n7477), .ZN(P2_U3191) );
  XNOR2_X1 U9284 ( .A(n7479), .B(n8198), .ZN(n7524) );
  XNOR2_X1 U9285 ( .A(n7480), .B(n8198), .ZN(n7481) );
  NAND2_X1 U9286 ( .A1(n7481), .A2(n9017), .ZN(n7483) );
  AOI22_X1 U9287 ( .A1(n9014), .A2(n8666), .B1(n8668), .B2(n9012), .ZN(n7482)
         );
  OAI211_X1 U9288 ( .C1(n7653), .C2(n7524), .A(n7483), .B(n7482), .ZN(n7520)
         );
  INV_X1 U9289 ( .A(n7637), .ZN(n7647) );
  OAI22_X1 U9290 ( .A1(n7524), .A2(n7731), .B1(n7647), .B2(n9454), .ZN(n7484)
         );
  NOR2_X1 U9291 ( .A1(n7520), .A2(n7484), .ZN(n10679) );
  NAND2_X1 U9292 ( .A1(n4671), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7485) );
  OAI21_X1 U9293 ( .B1(n10679), .B2(n4671), .A(n7485), .ZN(P2_U3468) );
  OAI21_X1 U9294 ( .B1(n5833), .B2(n7487), .A(n7486), .ZN(n10600) );
  INV_X1 U9295 ( .A(n10600), .ZN(n10597) );
  XNOR2_X1 U9296 ( .A(n5897), .B(n7488), .ZN(n7489) );
  NOR2_X1 U9297 ( .A1(n7489), .A2(n10308), .ZN(n10595) );
  XNOR2_X1 U9298 ( .A(n9812), .B(n7490), .ZN(n7491) );
  NAND2_X1 U9299 ( .A1(n7491), .A2(n10285), .ZN(n7493) );
  NAND2_X1 U9300 ( .A1(n7493), .A2(n7492), .ZN(n10599) );
  AOI21_X1 U9301 ( .B1(n10595), .B2(n9938), .A(n10599), .ZN(n7495) );
  MUX2_X1 U9302 ( .A(n7495), .B(n7494), .S(n10553), .Z(n7497) );
  AOI22_X1 U9303 ( .A1(n10278), .A2(n5897), .B1(n10551), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7496) );
  OAI211_X1 U9304 ( .C1(n10259), .C2(n10597), .A(n7497), .B(n7496), .ZN(
        P1_U3292) );
  INV_X1 U9305 ( .A(n7498), .ZN(n7508) );
  INV_X1 U9306 ( .A(n7499), .ZN(n7500) );
  MUX2_X1 U9307 ( .A(n7501), .B(n7500), .S(n5878), .Z(n7507) );
  OAI22_X1 U9308 ( .A1(n10556), .A2(n7503), .B1(n10270), .B2(n7502), .ZN(n7504) );
  AOI21_X1 U9309 ( .B1(n10548), .B2(n7505), .A(n7504), .ZN(n7506) );
  OAI211_X1 U9310 ( .C1(n10259), .C2(n7508), .A(n7507), .B(n7506), .ZN(
        P1_U3291) );
  INV_X1 U9311 ( .A(n7509), .ZN(n7519) );
  INV_X1 U9312 ( .A(n7510), .ZN(n7511) );
  AOI22_X1 U9313 ( .A1(n10553), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7511), .B2(
        n10551), .ZN(n7512) );
  OAI21_X1 U9314 ( .B1(n10556), .B2(n7513), .A(n7512), .ZN(n7514) );
  AOI21_X1 U9315 ( .B1(n7515), .B2(n10548), .A(n7514), .ZN(n7518) );
  NAND2_X1 U9316 ( .A1(n7516), .A2(n5878), .ZN(n7517) );
  OAI211_X1 U9317 ( .C1(n7519), .C2(n10259), .A(n7518), .B(n7517), .ZN(
        P1_U3289) );
  NAND2_X1 U9318 ( .A1(n7520), .A2(n9020), .ZN(n7523) );
  OAI22_X1 U9319 ( .A1(n9020), .A2(n6390), .B1(n7640), .B2(n9018), .ZN(n7521)
         );
  AOI21_X1 U9320 ( .B1(n9023), .B2(n7637), .A(n7521), .ZN(n7522) );
  OAI211_X1 U9321 ( .C1(n7524), .C2(n7578), .A(n7523), .B(n7522), .ZN(P2_U3224) );
  OAI21_X1 U9322 ( .B1(n7526), .B2(n9815), .A(n7525), .ZN(n10605) );
  OAI211_X1 U9323 ( .C1(n4580), .C2(n10602), .A(n7594), .B(n10319), .ZN(n10601) );
  INV_X1 U9324 ( .A(n7586), .ZN(n7527) );
  AOI22_X1 U9325 ( .A1(n10278), .A2(n9690), .B1(n10551), .B2(n7527), .ZN(n7528) );
  OAI21_X1 U9326 ( .B1(n10601), .B2(n10275), .A(n7528), .ZN(n7535) );
  XNOR2_X1 U9327 ( .A(n7529), .B(n9815), .ZN(n7533) );
  NAND2_X1 U9328 ( .A1(n9981), .A2(n9667), .ZN(n7531) );
  NAND2_X1 U9329 ( .A1(n9983), .A2(n9666), .ZN(n7530) );
  NAND2_X1 U9330 ( .A1(n7531), .A2(n7530), .ZN(n7583) );
  INV_X1 U9331 ( .A(n7583), .ZN(n7532) );
  OAI21_X1 U9332 ( .B1(n7533), .B2(n10302), .A(n7532), .ZN(n10603) );
  MUX2_X1 U9333 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10603), .S(n5878), .Z(n7534)
         );
  AOI211_X1 U9334 ( .C1(n10560), .C2(n10605), .A(n7535), .B(n7534), .ZN(n7536)
         );
  INV_X1 U9335 ( .A(n7536), .ZN(P1_U3288) );
  OAI21_X1 U9336 ( .B1(n7539), .B2(n7538), .A(n7537), .ZN(n7546) );
  NAND2_X1 U9337 ( .A1(n9979), .A2(n9667), .ZN(n7541) );
  NAND2_X1 U9338 ( .A1(n9981), .A2(n9666), .ZN(n7540) );
  NAND2_X1 U9339 ( .A1(n7541), .A2(n7540), .ZN(n7774) );
  AOI21_X1 U9340 ( .B1(n10541), .B2(n7774), .A(n7542), .ZN(n7544) );
  NAND2_X1 U9341 ( .A1(n10515), .A2(n10607), .ZN(n7543) );
  OAI211_X1 U9342 ( .C1(n10547), .C2(n7783), .A(n7544), .B(n7543), .ZN(n7545)
         );
  AOI21_X1 U9343 ( .B1(n7546), .B2(n10527), .A(n7545), .ZN(n7547) );
  INV_X1 U9344 ( .A(n7547), .ZN(P1_U3213) );
  INV_X1 U9345 ( .A(n7548), .ZN(n7648) );
  OAI222_X1 U9346 ( .A1(n10470), .A2(n9174), .B1(n10472), .B2(n7648), .C1(
        P1_U3086), .C2(n9938), .ZN(P1_U3336) );
  MUX2_X1 U9347 ( .A(n7549), .B(n4753), .S(n9000), .Z(n7553) );
  INV_X1 U9348 ( .A(n7550), .ZN(n7551) );
  AOI22_X1 U9349 ( .A1(n9023), .A2(n8248), .B1(n8999), .B2(n7551), .ZN(n7552)
         );
  OAI211_X1 U9350 ( .C1(n7554), .C2(n7578), .A(n7553), .B(n7552), .ZN(P2_U3226) );
  NAND2_X1 U9351 ( .A1(n8676), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7555) );
  OAI21_X1 U9352 ( .B1(n8186), .B2(n8676), .A(n7555), .ZN(P2_U3521) );
  INV_X1 U9353 ( .A(n7556), .ZN(n7558) );
  NOR2_X1 U9354 ( .A1(n8641), .A2(n8247), .ZN(n7557) );
  AOI211_X1 U9355 ( .C1(n8639), .C2(n8667), .A(n7558), .B(n7557), .ZN(n7559)
         );
  OAI21_X1 U9356 ( .B1(n8524), .B2(n7667), .A(n7559), .ZN(n7567) );
  NAND2_X1 U9357 ( .A1(n7560), .A2(n7563), .ZN(n7561) );
  XNOR2_X1 U9358 ( .A(n7669), .B(n8546), .ZN(n7634) );
  XNOR2_X1 U9359 ( .A(n7634), .B(n8668), .ZN(n7562) );
  NAND2_X1 U9360 ( .A1(n7561), .A2(n7562), .ZN(n7636) );
  INV_X1 U9361 ( .A(n7562), .ZN(n7564) );
  NAND3_X1 U9362 ( .A1(n7560), .A2(n7564), .A3(n7563), .ZN(n7565) );
  AOI21_X1 U9363 ( .B1(n7636), .B2(n7565), .A(n8632), .ZN(n7566) );
  AOI211_X1 U9364 ( .C1(n7669), .C2(n8629), .A(n7567), .B(n7566), .ZN(n7568)
         );
  INV_X1 U9365 ( .A(n7568), .ZN(P2_U3161) );
  NAND2_X1 U9366 ( .A1(n8304), .A2(n8252), .ZN(n8200) );
  INV_X1 U9367 ( .A(n8200), .ZN(n7569) );
  XNOR2_X1 U9368 ( .A(n7570), .B(n7569), .ZN(n7732) );
  XNOR2_X1 U9369 ( .A(n7571), .B(n8200), .ZN(n7572) );
  NAND2_X1 U9370 ( .A1(n7572), .A2(n9017), .ZN(n7574) );
  AOI22_X1 U9371 ( .A1(n9014), .A2(n8665), .B1(n8667), .B2(n9012), .ZN(n7573)
         );
  OAI211_X1 U9372 ( .C1(n7732), .C2(n7653), .A(n7574), .B(n7573), .ZN(n7733)
         );
  NAND2_X1 U9373 ( .A1(n7733), .A2(n9020), .ZN(n7577) );
  OAI22_X1 U9374 ( .A1(n9020), .A2(n7615), .B1(n7889), .B2(n9018), .ZN(n7575)
         );
  AOI21_X1 U9375 ( .B1(n9023), .B2(n7891), .A(n7575), .ZN(n7576) );
  OAI211_X1 U9376 ( .C1(n7732), .C2(n7578), .A(n7577), .B(n7576), .ZN(P2_U3223) );
  NOR2_X1 U9377 ( .A1(n7580), .A2(n7579), .ZN(n10531) );
  AOI21_X1 U9378 ( .B1(n7580), .B2(n7579), .A(n10531), .ZN(n7581) );
  NAND2_X1 U9379 ( .A1(n7581), .A2(n7582), .ZN(n10534) );
  OAI21_X1 U9380 ( .B1(n7582), .B2(n7581), .A(n10534), .ZN(n7589) );
  NOR2_X1 U9381 ( .A1(n10543), .A2(n10602), .ZN(n7588) );
  NAND2_X1 U9382 ( .A1(n10541), .A2(n7583), .ZN(n7585) );
  OAI211_X1 U9383 ( .C1(n10547), .C2(n7586), .A(n7585), .B(n7584), .ZN(n7587)
         );
  AOI211_X1 U9384 ( .C1(n7589), .C2(n10527), .A(n7588), .B(n7587), .ZN(n7590)
         );
  INV_X1 U9385 ( .A(n7590), .ZN(P1_U3227) );
  OAI21_X1 U9386 ( .B1(n7592), .B2(n7595), .A(n7591), .ZN(n10559) );
  INV_X1 U9387 ( .A(n7780), .ZN(n7593) );
  AOI211_X1 U9388 ( .C1(n9698), .C2(n7594), .A(n10308), .B(n7593), .ZN(n10549)
         );
  XNOR2_X1 U9389 ( .A(n7749), .B(n7595), .ZN(n7598) );
  NAND2_X1 U9390 ( .A1(n9982), .A2(n9666), .ZN(n7597) );
  NAND2_X1 U9391 ( .A1(n9980), .A2(n9667), .ZN(n7596) );
  NAND2_X1 U9392 ( .A1(n7597), .A2(n7596), .ZN(n10540) );
  AOI21_X1 U9393 ( .B1(n7598), .B2(n10285), .A(n10540), .ZN(n10562) );
  INV_X1 U9394 ( .A(n10562), .ZN(n7599) );
  AOI211_X1 U9395 ( .C1(n10622), .C2(n10559), .A(n10549), .B(n7599), .ZN(n7604) );
  INV_X1 U9396 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7600) );
  OAI22_X1 U9397 ( .A1(n10425), .A2(n10557), .B1(n10449), .B2(n7600), .ZN(
        n7601) );
  INV_X1 U9398 ( .A(n7601), .ZN(n7602) );
  OAI21_X1 U9399 ( .B1(n7604), .B2(n10634), .A(n7602), .ZN(P1_U3471) );
  AOI22_X1 U9400 ( .A1(n10392), .A2(n9698), .B1(n10641), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7603) );
  OAI21_X1 U9401 ( .B1(n7604), .B2(n10641), .A(n7603), .ZN(P1_U3528) );
  OR2_X1 U9402 ( .A1(n7627), .A2(n7607), .ZN(n7676) );
  NAND2_X1 U9403 ( .A1(n7627), .A2(n7607), .ZN(n7608) );
  NAND2_X1 U9404 ( .A1(n7676), .A2(n7608), .ZN(n7609) );
  NAND2_X1 U9405 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  AOI21_X1 U9406 ( .B1(n7677), .B2(n7611), .A(n8806), .ZN(n7632) );
  OR2_X1 U9407 ( .A1(n7627), .A2(n7615), .ZN(n7673) );
  NAND2_X1 U9408 ( .A1(n7627), .A2(n7615), .ZN(n7616) );
  NAND2_X1 U9409 ( .A1(n7673), .A2(n7616), .ZN(n7617) );
  NAND2_X1 U9410 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  AOI21_X1 U9411 ( .B1(n7674), .B2(n7619), .A(n8841), .ZN(n7631) );
  INV_X1 U9412 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8143) );
  MUX2_X1 U9413 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8798), .Z(n7681) );
  XNOR2_X1 U9414 ( .A(n7681), .B(n7627), .ZN(n7625) );
  OR2_X1 U9415 ( .A1(n7621), .A2(n7620), .ZN(n7623) );
  NAND2_X1 U9416 ( .A1(n7623), .A2(n7622), .ZN(n7624) );
  NAND2_X1 U9417 ( .A1(n7625), .A2(n7624), .ZN(n7682) );
  OAI21_X1 U9418 ( .B1(n7625), .B2(n7624), .A(n7682), .ZN(n7626) );
  INV_X1 U9419 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9165) );
  NOR2_X1 U9420 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9165), .ZN(n7887) );
  AOI21_X1 U9421 ( .B1(n10652), .B2(n7626), .A(n7887), .ZN(n7629) );
  NAND2_X1 U9422 ( .A1(n10650), .A2(n7627), .ZN(n7628) );
  OAI211_X1 U9423 ( .C1(n8143), .C2(n10657), .A(n7629), .B(n7628), .ZN(n7630)
         );
  OR3_X1 U9424 ( .A1(n7632), .A2(n7631), .A3(n7630), .ZN(P2_U3192) );
  NAND2_X1 U9425 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  XNOR2_X1 U9426 ( .A(n7637), .B(n8546), .ZN(n7879) );
  XNOR2_X1 U9427 ( .A(n7879), .B(n8667), .ZN(n7638) );
  OAI211_X1 U9428 ( .C1(n7639), .C2(n7638), .A(n7882), .B(n8635), .ZN(n7646)
         );
  INV_X1 U9429 ( .A(n7640), .ZN(n7644) );
  AOI21_X1 U9430 ( .B1(n8624), .B2(n8668), .A(n7641), .ZN(n7642) );
  OAI21_X1 U9431 ( .B1(n7960), .B2(n8627), .A(n7642), .ZN(n7643) );
  AOI21_X1 U9432 ( .B1(n8645), .B2(n7644), .A(n7643), .ZN(n7645) );
  OAI211_X1 U9433 ( .C1(n7647), .C2(n8648), .A(n7646), .B(n7645), .ZN(P2_U3171) );
  OAI222_X1 U9434 ( .A1(P2_U3151), .A2(n6622), .B1(n9524), .B2(n7648), .C1(
        n9185), .C2(n8484), .ZN(P2_U3276) );
  NAND2_X1 U9435 ( .A1(n7694), .A2(n7936), .ZN(n7650) );
  OAI211_X1 U9436 ( .C1(n10470), .C2(n7651), .A(n7650), .B(n7649), .ZN(
        P1_U3335) );
  AND2_X1 U9437 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  INV_X1 U9438 ( .A(n7655), .ZN(n7656) );
  MUX2_X1 U9439 ( .A(n7657), .B(n7656), .S(n9020), .Z(n7662) );
  NOR2_X1 U9440 ( .A1(n9018), .A2(n7658), .ZN(n7659) );
  AOI21_X1 U9441 ( .B1(n9023), .B2(n7660), .A(n7659), .ZN(n7661) );
  OAI211_X1 U9442 ( .C1(n9026), .C2(n7663), .A(n7662), .B(n7661), .ZN(P2_U3227) );
  INV_X1 U9443 ( .A(n7664), .ZN(n7665) );
  MUX2_X1 U9444 ( .A(n7666), .B(n7665), .S(n9020), .Z(n7671) );
  INV_X1 U9445 ( .A(n7667), .ZN(n7668) );
  AOI22_X1 U9446 ( .A1(n9023), .A2(n7669), .B1(n8999), .B2(n7668), .ZN(n7670)
         );
  OAI211_X1 U9447 ( .C1(n7672), .C2(n9026), .A(n7671), .B(n7670), .ZN(P2_U3225) );
  AOI21_X1 U9448 ( .B1(n7675), .B2(n6415), .A(n7809), .ZN(n7693) );
  NOR2_X1 U9449 ( .A1(n6414), .A2(n7678), .ZN(n7826) );
  AOI21_X1 U9450 ( .B1(n6414), .B2(n7678), .A(n7826), .ZN(n7679) );
  NOR2_X1 U9451 ( .A1(n7679), .A2(n8806), .ZN(n7691) );
  INV_X1 U9452 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7689) );
  MUX2_X1 U9453 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8798), .Z(n7814) );
  XNOR2_X1 U9454 ( .A(n7814), .B(n7825), .ZN(n7685) );
  OR2_X1 U9455 ( .A1(n7681), .A2(n7680), .ZN(n7683) );
  NAND2_X1 U9456 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U9457 ( .A1(n7685), .A2(n7684), .ZN(n7816) );
  OAI21_X1 U9458 ( .B1(n7685), .B2(n7684), .A(n7816), .ZN(n7686) );
  AND2_X1 U9459 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7963) );
  AOI21_X1 U9460 ( .B1(n10652), .B2(n7686), .A(n7963), .ZN(n7688) );
  NAND2_X1 U9461 ( .A1(n10650), .A2(n7825), .ZN(n7687) );
  OAI211_X1 U9462 ( .C1(n7689), .C2(n10657), .A(n7688), .B(n7687), .ZN(n7690)
         );
  NOR2_X1 U9463 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  OAI21_X1 U9464 ( .B1(n7693), .B2(n8841), .A(n7692), .ZN(P2_U3193) );
  INV_X1 U9465 ( .A(n7694), .ZN(n7696) );
  OAI222_X1 U9466 ( .A1(n8406), .A2(P2_U3151), .B1(n9524), .B2(n7696), .C1(
        n7695), .C2(n8484), .ZN(P2_U3275) );
  NAND2_X1 U9467 ( .A1(n9023), .A2(n6303), .ZN(n7698) );
  OAI21_X1 U9468 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n9018), .A(n7698), .ZN(
        n7701) );
  NOR2_X1 U9469 ( .A1(n7699), .A2(n9022), .ZN(n7700) );
  AOI211_X1 U9470 ( .C1(n9000), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7701), .B(
        n7700), .ZN(n7702) );
  OAI21_X1 U9471 ( .B1(n9026), .B2(n7703), .A(n7702), .ZN(P2_U3230) );
  OAI21_X1 U9472 ( .B1(n7709), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7704), .ZN(
        n7707) );
  AOI22_X1 U9473 ( .A1(n7871), .A2(n8451), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7705), .ZN(n7706) );
  NOR2_X1 U9474 ( .A1(n7706), .A2(n7707), .ZN(n7866) );
  AOI211_X1 U9475 ( .C1(n7707), .C2(n7706), .A(n7866), .B(n10037), .ZN(n7717)
         );
  OAI21_X1 U9476 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7709), .A(n7708), .ZN(
        n7712) );
  INV_X1 U9477 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8464) );
  NOR2_X1 U9478 ( .A1(n7871), .A2(n8464), .ZN(n7710) );
  AOI21_X1 U9479 ( .B1(n8464), .B2(n7871), .A(n7710), .ZN(n7711) );
  NOR2_X1 U9480 ( .A1(n7711), .A2(n7712), .ZN(n7870) );
  AOI211_X1 U9481 ( .C1(n7712), .C2(n7711), .A(n7870), .B(n10090), .ZN(n7716)
         );
  INV_X1 U9482 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U9483 ( .A1(n10072), .A2(n7871), .ZN(n7714) );
  NAND2_X1 U9484 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7713) );
  OAI211_X1 U9485 ( .C1(n9288), .C2(n10099), .A(n7714), .B(n7713), .ZN(n7715)
         );
  OR3_X1 U9486 ( .A1(n7717), .A2(n7716), .A3(n7715), .ZN(P1_U3256) );
  XNOR2_X1 U9487 ( .A(n7726), .B(n8665), .ZN(n8201) );
  NAND2_X1 U9488 ( .A1(n7718), .A2(n8252), .ZN(n7719) );
  XOR2_X1 U9489 ( .A(n8201), .B(n7719), .Z(n7727) );
  XNOR2_X1 U9490 ( .A(n4658), .B(n8201), .ZN(n7721) );
  OAI222_X1 U9491 ( .A1(n8953), .A2(n7965), .B1(n8993), .B2(n7960), .C1(n7721), 
        .C2(n8990), .ZN(n7729) );
  NAND2_X1 U9492 ( .A1(n7729), .A2(n9020), .ZN(n7725) );
  INV_X1 U9493 ( .A(n7967), .ZN(n7722) );
  OAI22_X1 U9494 ( .A1(n9020), .A2(n6415), .B1(n7722), .B2(n9018), .ZN(n7723)
         );
  AOI21_X1 U9495 ( .B1(n9023), .B2(n7726), .A(n7723), .ZN(n7724) );
  OAI211_X1 U9496 ( .C1(n7727), .C2(n9026), .A(n7725), .B(n7724), .ZN(P2_U3222) );
  OAI22_X1 U9497 ( .A1(n7727), .A2(n9448), .B1(n5010), .B2(n9454), .ZN(n7728)
         );
  NOR2_X1 U9498 ( .A1(n7729), .A2(n7728), .ZN(n10684) );
  NAND2_X1 U9499 ( .A1(n4671), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7730) );
  OAI21_X1 U9500 ( .B1(n10684), .B2(n4671), .A(n7730), .ZN(P2_U3470) );
  NOR2_X1 U9501 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  AOI211_X1 U9502 ( .C1(n9443), .C2(n7891), .A(n7734), .B(n7733), .ZN(n10681)
         );
  OR2_X1 U9503 ( .A1(n10681), .A2(n4671), .ZN(n7735) );
  OAI21_X1 U9504 ( .B1(n9456), .B2(n7607), .A(n7735), .ZN(P2_U3469) );
  NAND2_X1 U9505 ( .A1(n7736), .A2(n10527), .ZN(n7747) );
  AOI21_X1 U9506 ( .B1(n7737), .B2(n7739), .A(n7738), .ZN(n7746) );
  NAND2_X1 U9507 ( .A1(n9977), .A2(n9667), .ZN(n7758) );
  NAND2_X1 U9508 ( .A1(n9979), .A2(n9666), .ZN(n7753) );
  NAND2_X1 U9509 ( .A1(n7758), .A2(n7753), .ZN(n7740) );
  NAND2_X1 U9510 ( .A1(n10541), .A2(n7740), .ZN(n7743) );
  INV_X1 U9511 ( .A(n7741), .ZN(n7742) );
  OAI211_X1 U9512 ( .C1(n10547), .C2(n7760), .A(n7743), .B(n7742), .ZN(n7744)
         );
  AOI21_X1 U9513 ( .B1(n4559), .B2(n10515), .A(n7744), .ZN(n7745) );
  OAI21_X1 U9514 ( .B1(n7747), .B2(n7746), .A(n7745), .ZN(P1_U3231) );
  INV_X1 U9515 ( .A(n9706), .ZN(n7748) );
  OR2_X1 U9516 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  NAND2_X1 U9517 ( .A1(n7750), .A2(n9882), .ZN(n7773) );
  AND2_X1 U9518 ( .A1(n7773), .A2(n9711), .ZN(n7772) );
  INV_X1 U9519 ( .A(n7751), .ZN(n9715) );
  OAI21_X1 U9520 ( .B1(n7772), .B2(n9715), .A(n9714), .ZN(n7752) );
  XOR2_X1 U9521 ( .A(n7756), .B(n7752), .Z(n7754) );
  OAI21_X1 U9522 ( .B1(n7754), .B2(n10302), .A(n7753), .ZN(n10619) );
  INV_X1 U9523 ( .A(n10619), .ZN(n7767) );
  OAI21_X1 U9524 ( .B1(n7757), .B2(n7756), .A(n7755), .ZN(n10621) );
  OAI211_X1 U9525 ( .C1(n10618), .C2(n7857), .A(n7801), .B(n10319), .ZN(n7759)
         );
  AND2_X1 U9526 ( .A1(n7759), .A2(n7758), .ZN(n10616) );
  INV_X1 U9527 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7761) );
  OAI22_X1 U9528 ( .A1(n5878), .A2(n7761), .B1(n7760), .B2(n10270), .ZN(n7762)
         );
  AOI21_X1 U9529 ( .B1(n10278), .B2(n4559), .A(n7762), .ZN(n7764) );
  OAI21_X1 U9530 ( .B1(n10616), .B2(n10275), .A(n7764), .ZN(n7765) );
  AOI21_X1 U9531 ( .B1(n10621), .B2(n10560), .A(n7765), .ZN(n7766) );
  OAI21_X1 U9532 ( .B1(n10563), .B2(n7767), .A(n7766), .ZN(P1_U3284) );
  OR2_X1 U9533 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  NAND2_X1 U9534 ( .A1(n7771), .A2(n7770), .ZN(n10612) );
  INV_X1 U9535 ( .A(n10612), .ZN(n7788) );
  INV_X1 U9536 ( .A(n7772), .ZN(n7851) );
  OAI21_X1 U9537 ( .B1(n9711), .B2(n7773), .A(n7851), .ZN(n7775) );
  AOI21_X1 U9538 ( .B1(n7775), .B2(n10285), .A(n7774), .ZN(n7778) );
  INV_X1 U9539 ( .A(n7776), .ZN(n10633) );
  NAND2_X1 U9540 ( .A1(n10612), .A2(n10633), .ZN(n7777) );
  AND2_X1 U9541 ( .A1(n7778), .A2(n7777), .ZN(n10614) );
  MUX2_X1 U9542 ( .A(n10614), .B(n7779), .S(n10553), .Z(n7787) );
  NAND2_X1 U9543 ( .A1(n7780), .A2(n10607), .ZN(n7781) );
  NAND2_X1 U9544 ( .A1(n7781), .A2(n10319), .ZN(n7782) );
  NOR2_X1 U9545 ( .A1(n7856), .A2(n7782), .ZN(n10609) );
  INV_X1 U9546 ( .A(n10607), .ZN(n7784) );
  OAI22_X1 U9547 ( .A1(n10556), .A2(n7784), .B1(n7783), .B2(n10270), .ZN(n7785) );
  AOI21_X1 U9548 ( .B1(n10609), .B2(n10548), .A(n7785), .ZN(n7786) );
  OAI211_X1 U9549 ( .C1(n7788), .C2(n7862), .A(n7787), .B(n7786), .ZN(P1_U3286) );
  INV_X1 U9550 ( .A(n7789), .ZN(n7791) );
  OAI222_X1 U9551 ( .A1(n8262), .A2(P2_U3151), .B1(n9524), .B2(n7791), .C1(
        n9264), .C2(n8484), .ZN(P2_U3274) );
  OAI222_X1 U9552 ( .A1(P1_U3086), .A2(n9807), .B1(n10472), .B2(n7791), .C1(
        n7790), .C2(n10470), .ZN(P1_U3334) );
  NAND3_X1 U9553 ( .A1(n7792), .A2(n9887), .A3(n7798), .ZN(n7793) );
  AOI21_X1 U9554 ( .B1(n7916), .B2(n7793), .A(n10302), .ZN(n7796) );
  NAND2_X1 U9555 ( .A1(n9978), .A2(n9666), .ZN(n7795) );
  NAND2_X1 U9556 ( .A1(n9976), .A2(n9667), .ZN(n7794) );
  NAND2_X1 U9557 ( .A1(n7795), .A2(n7794), .ZN(n10478) );
  INV_X1 U9558 ( .A(n7837), .ZN(n7807) );
  OAI21_X1 U9559 ( .B1(n7799), .B2(n7798), .A(n7797), .ZN(n7839) );
  NAND2_X1 U9560 ( .A1(n7839), .A2(n10560), .ZN(n7806) );
  AOI211_X1 U9561 ( .C1(n10486), .C2(n7801), .A(n10308), .B(n7800), .ZN(n7838)
         );
  INV_X1 U9562 ( .A(n10486), .ZN(n7802) );
  NOR2_X1 U9563 ( .A1(n7802), .A2(n10556), .ZN(n7804) );
  OAI22_X1 U9564 ( .A1(n10241), .A2(n7253), .B1(n10488), .B2(n10270), .ZN(
        n7803) );
  AOI211_X1 U9565 ( .C1(n7838), .C2(n10548), .A(n7804), .B(n7803), .ZN(n7805)
         );
  OAI211_X1 U9566 ( .C1(n10563), .C2(n7807), .A(n7806), .B(n7805), .ZN(
        P1_U3283) );
  NOR2_X1 U9567 ( .A1(n7825), .A2(n7808), .ZN(n7810) );
  XNOR2_X1 U9568 ( .A(n7829), .B(n7811), .ZN(n7812) );
  NOR2_X1 U9569 ( .A1(n7813), .A2(n7812), .ZN(n7985) );
  AOI21_X1 U9570 ( .B1(n7813), .B2(n7812), .A(n7985), .ZN(n7836) );
  MUX2_X1 U9571 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8798), .Z(n7989) );
  XNOR2_X1 U9572 ( .A(n7829), .B(n7989), .ZN(n7819) );
  INV_X1 U9573 ( .A(n7814), .ZN(n7815) );
  NAND2_X1 U9574 ( .A1(n7825), .A2(n7815), .ZN(n7817) );
  NAND2_X1 U9575 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  NAND2_X1 U9576 ( .A1(n7819), .A2(n7818), .ZN(n7990) );
  OAI21_X1 U9577 ( .B1(n7819), .B2(n7818), .A(n7990), .ZN(n7820) );
  NAND2_X1 U9578 ( .A1(n10652), .A2(n7820), .ZN(n7823) );
  NOR2_X1 U9579 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7821), .ZN(n8025) );
  INV_X1 U9580 ( .A(n8025), .ZN(n7822) );
  OAI211_X1 U9581 ( .C1(n8837), .C2(n7988), .A(n7823), .B(n7822), .ZN(n7834)
         );
  NOR2_X1 U9582 ( .A1(n7825), .A2(n7824), .ZN(n7827) );
  AOI22_X1 U9583 ( .A1(n7829), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n7828), .B2(
        n7988), .ZN(n7830) );
  AOI21_X1 U9584 ( .B1(n7831), .B2(n7830), .A(n7983), .ZN(n7832) );
  NOR2_X1 U9585 ( .A1(n7832), .A2(n8806), .ZN(n7833) );
  AOI211_X1 U9586 ( .C1(n8839), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7834), .B(
        n7833), .ZN(n7835) );
  OAI21_X1 U9587 ( .B1(n7836), .B2(n8841), .A(n7835), .ZN(P2_U3194) );
  AOI211_X1 U9588 ( .C1(n7839), .C2(n10622), .A(n7838), .B(n7837), .ZN(n7843)
         );
  AOI22_X1 U9589 ( .A1(n10486), .A2(n10392), .B1(n10641), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7840) );
  OAI21_X1 U9590 ( .B1(n7843), .B2(n10641), .A(n7840), .ZN(P1_U3532) );
  NOR2_X1 U9591 ( .A1(n10449), .A2(n5546), .ZN(n7841) );
  AOI21_X1 U9592 ( .B1(n10486), .B2(n10453), .A(n7841), .ZN(n7842) );
  OAI21_X1 U9593 ( .B1(n7843), .B2(n10634), .A(n7842), .ZN(P1_U3483) );
  OAI21_X1 U9594 ( .B1(n7845), .B2(n7852), .A(n7844), .ZN(n7861) );
  OAI22_X1 U9595 ( .A1(n7849), .A2(n7848), .B1(n7847), .B2(n7846), .ZN(n10523)
         );
  NAND2_X1 U9596 ( .A1(n7851), .A2(n7850), .ZN(n7853) );
  XNOR2_X1 U9597 ( .A(n7853), .B(n7852), .ZN(n7854) );
  NOR2_X1 U9598 ( .A1(n7854), .A2(n10302), .ZN(n7855) );
  AOI211_X1 U9599 ( .C1(n10633), .C2(n7861), .A(n10523), .B(n7855), .ZN(n7953)
         );
  INV_X1 U9600 ( .A(n7856), .ZN(n7858) );
  AOI21_X1 U9601 ( .B1(n7950), .B2(n7858), .A(n7857), .ZN(n7951) );
  INV_X1 U9602 ( .A(n10530), .ZN(n7859) );
  AOI22_X1 U9603 ( .A1(n10553), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7859), .B2(
        n10551), .ZN(n7860) );
  OAI21_X1 U9604 ( .B1(n10556), .B2(n10525), .A(n7860), .ZN(n7864) );
  INV_X1 U9605 ( .A(n7861), .ZN(n7954) );
  NOR2_X1 U9606 ( .A1(n7954), .A2(n7862), .ZN(n7863) );
  AOI211_X1 U9607 ( .C1(n7951), .C2(n10110), .A(n7864), .B(n7863), .ZN(n7865)
         );
  OAI21_X1 U9608 ( .B1(n10563), .B2(n7953), .A(n7865), .ZN(P1_U3285) );
  AOI22_X1 U9609 ( .A1(n8054), .A2(n8068), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7867), .ZN(n7868) );
  NOR2_X1 U9610 ( .A1(n7869), .A2(n7868), .ZN(n8050) );
  AOI211_X1 U9611 ( .C1(n7869), .C2(n7868), .A(n8050), .B(n10037), .ZN(n7878)
         );
  XNOR2_X1 U9612 ( .A(n8054), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7872) );
  NOR2_X1 U9613 ( .A1(n7873), .A2(n7872), .ZN(n8053) );
  AOI211_X1 U9614 ( .C1(n7873), .C2(n7872), .A(n8053), .B(n10090), .ZN(n7877)
         );
  INV_X1 U9615 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U9616 ( .A1(n10072), .A2(n8054), .ZN(n7875) );
  NAND2_X1 U9617 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n7874) );
  OAI211_X1 U9618 ( .C1(n9292), .C2(n10099), .A(n7875), .B(n7874), .ZN(n7876)
         );
  OR3_X1 U9619 ( .A1(n7878), .A2(n7877), .A3(n7876), .ZN(P1_U3257) );
  XOR2_X1 U9620 ( .A(n8546), .B(n7891), .Z(n7884) );
  INV_X1 U9621 ( .A(n7879), .ZN(n7880) );
  NAND2_X1 U9622 ( .A1(n7880), .A2(n8667), .ZN(n7881) );
  AOI21_X1 U9623 ( .B1(n7884), .B2(n7883), .A(n7959), .ZN(n7893) );
  NOR2_X1 U9624 ( .A1(n8641), .A2(n7885), .ZN(n7886) );
  AOI211_X1 U9625 ( .C1(n8639), .C2(n8665), .A(n7887), .B(n7886), .ZN(n7888)
         );
  OAI21_X1 U9626 ( .B1(n8524), .B2(n7889), .A(n7888), .ZN(n7890) );
  AOI21_X1 U9627 ( .B1(n7891), .B2(n8629), .A(n7890), .ZN(n7892) );
  OAI21_X1 U9628 ( .B1(n7893), .B2(n8632), .A(n7892), .ZN(P2_U3157) );
  INV_X1 U9629 ( .A(n7894), .ZN(n7902) );
  NAND2_X1 U9630 ( .A1(n9023), .A2(n7895), .ZN(n7896) );
  OAI21_X1 U9631 ( .B1(n7897), .B2(n9018), .A(n7896), .ZN(n7900) );
  NOR2_X1 U9632 ( .A1(n9026), .A2(n7898), .ZN(n7899) );
  AOI211_X1 U9633 ( .C1(n9022), .C2(P2_REG2_REG_4__SCAN_IN), .A(n7900), .B(
        n7899), .ZN(n7901) );
  OAI21_X1 U9634 ( .B1(n9022), .B2(n7902), .A(n7901), .ZN(P2_U3229) );
  XOR2_X1 U9635 ( .A(n8314), .B(n7903), .Z(n7904) );
  OAI222_X1 U9636 ( .A1(n8993), .A2(n8028), .B1(n8953), .B2(n8113), .C1(n7904), 
        .C2(n8990), .ZN(n7911) );
  INV_X1 U9637 ( .A(n7911), .ZN(n7910) );
  XOR2_X1 U9638 ( .A(n7905), .B(n8314), .Z(n7912) );
  INV_X1 U9639 ( .A(n8030), .ZN(n7907) );
  AOI22_X1 U9640 ( .A1(n9000), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8999), .B2(
        n8024), .ZN(n7906) );
  OAI21_X1 U9641 ( .B1(n7907), .B2(n9002), .A(n7906), .ZN(n7908) );
  AOI21_X1 U9642 ( .B1(n7912), .B2(n9004), .A(n7908), .ZN(n7909) );
  OAI21_X1 U9643 ( .B1(n7910), .B2(n9022), .A(n7909), .ZN(P2_U3221) );
  AOI21_X1 U9644 ( .B1(n9449), .B2(n7912), .A(n7911), .ZN(n7915) );
  AOI22_X1 U9645 ( .A1(n8030), .A2(n9028), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n4671), .ZN(n7913) );
  OAI21_X1 U9646 ( .B1(n7915), .B2(n4671), .A(n7913), .ZN(P2_U3471) );
  NOR2_X1 U9647 ( .A1(n10685), .A2(n9454), .ZN(n9467) );
  AOI22_X1 U9648 ( .A1(n8030), .A2(n9467), .B1(P2_REG0_REG_12__SCAN_IN), .B2(
        n10685), .ZN(n7914) );
  OAI21_X1 U9649 ( .B1(n7915), .B2(n10685), .A(n7914), .ZN(P2_U3426) );
  INV_X1 U9650 ( .A(n7923), .ZN(n9819) );
  AOI21_X1 U9651 ( .B1(n7916), .B2(n9736), .A(n9819), .ZN(n7917) );
  NOR2_X1 U9652 ( .A1(n7917), .A2(n10302), .ZN(n7921) );
  NAND2_X1 U9653 ( .A1(n9975), .A2(n9667), .ZN(n7919) );
  NAND2_X1 U9654 ( .A1(n9977), .A2(n9666), .ZN(n7918) );
  NAND2_X1 U9655 ( .A1(n7919), .A2(n7918), .ZN(n10508) );
  AOI21_X1 U9656 ( .B1(n7921), .B2(n7920), .A(n10508), .ZN(n10628) );
  OAI21_X1 U9657 ( .B1(n7924), .B2(n7923), .A(n7922), .ZN(n10632) );
  NAND2_X1 U9658 ( .A1(n10632), .A2(n10560), .ZN(n7930) );
  INV_X1 U9659 ( .A(n7976), .ZN(n7925) );
  AOI211_X1 U9660 ( .C1(n10625), .C2(n4841), .A(n10308), .B(n7925), .ZN(n10624) );
  NOR2_X1 U9661 ( .A1(n5828), .A2(n10556), .ZN(n7928) );
  OAI22_X1 U9662 ( .A1(n5878), .A2(n7926), .B1(n10517), .B2(n10270), .ZN(n7927) );
  AOI211_X1 U9663 ( .C1(n10624), .C2(n10548), .A(n7928), .B(n7927), .ZN(n7929)
         );
  OAI211_X1 U9664 ( .C1(n10563), .C2(n10628), .A(n7930), .B(n7929), .ZN(
        P1_U3282) );
  INV_X1 U9665 ( .A(n7931), .ZN(n7934) );
  OAI222_X1 U9666 ( .A1(P2_U3151), .A2(n7932), .B1(n9524), .B2(n7934), .C1(
        n9186), .C2(n8484), .ZN(P2_U3273) );
  OAI222_X1 U9667 ( .A1(n10470), .A2(n7935), .B1(n10472), .B2(n7934), .C1(
        P1_U3086), .C2(n7933), .ZN(P1_U3333) );
  NAND2_X1 U9668 ( .A1(n7940), .A2(n7936), .ZN(n7938) );
  OR2_X1 U9669 ( .A1(n7937), .A2(P1_U3086), .ZN(n9940) );
  OAI211_X1 U9670 ( .C1(n7939), .C2(n10470), .A(n7938), .B(n9940), .ZN(
        P1_U3332) );
  NAND2_X1 U9671 ( .A1(n7940), .A2(n8119), .ZN(n7941) );
  OAI211_X1 U9672 ( .C1(n7942), .C2(n8484), .A(n7941), .B(n8413), .ZN(P2_U3272) );
  INV_X1 U9673 ( .A(n8905), .ZN(n8898) );
  XNOR2_X1 U9674 ( .A(n7943), .B(n8205), .ZN(n7944) );
  OAI222_X1 U9675 ( .A1(n8993), .A2(n7965), .B1(n8953), .B2(n8642), .C1(n7944), 
        .C2(n8990), .ZN(n8008) );
  AOI21_X1 U9676 ( .B1(n8898), .B2(n8318), .A(n8008), .ZN(n7949) );
  AOI22_X1 U9677 ( .A1(n9000), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8999), .B2(
        n8093), .ZN(n7948) );
  XNOR2_X1 U9678 ( .A(n7946), .B(n7945), .ZN(n8009) );
  NAND2_X1 U9679 ( .A1(n8009), .A2(n9004), .ZN(n7947) );
  OAI211_X1 U9680 ( .C1(n7949), .C2(n9022), .A(n7948), .B(n7947), .ZN(P2_U3220) );
  AOI22_X1 U9681 ( .A1(n7951), .A2(n10319), .B1(n10626), .B2(n7950), .ZN(n7952) );
  OAI211_X1 U9682 ( .C1(n7954), .C2(n10629), .A(n7953), .B(n7952), .ZN(n7956)
         );
  NAND2_X1 U9683 ( .A1(n7956), .A2(n10643), .ZN(n7955) );
  OAI21_X1 U9684 ( .B1(n10643), .B2(n7116), .A(n7955), .ZN(P1_U3530) );
  NAND2_X1 U9685 ( .A1(n7956), .A2(n10449), .ZN(n7957) );
  OAI21_X1 U9686 ( .B1(n10449), .B2(n5510), .A(n7957), .ZN(P1_U3477) );
  INV_X1 U9687 ( .A(n7958), .ZN(n7961) );
  XNOR2_X1 U9688 ( .A(n8201), .B(n8546), .ZN(n8023) );
  OAI211_X1 U9689 ( .C1(n7962), .C2(n8023), .A(n8022), .B(n8635), .ZN(n7969)
         );
  AOI21_X1 U9690 ( .B1(n8624), .B2(n8666), .A(n7963), .ZN(n7964) );
  OAI21_X1 U9691 ( .B1(n7965), .B2(n8627), .A(n7964), .ZN(n7966) );
  AOI21_X1 U9692 ( .B1(n8645), .B2(n7967), .A(n7966), .ZN(n7968) );
  OAI211_X1 U9693 ( .C1(n5010), .C2(n8648), .A(n7969), .B(n7968), .ZN(P2_U3176) );
  OAI211_X1 U9694 ( .C1(n9821), .C2(n7970), .A(n8441), .B(n10285), .ZN(n7973)
         );
  NAND2_X1 U9695 ( .A1(n9974), .A2(n9667), .ZN(n7972) );
  NAND2_X1 U9696 ( .A1(n9976), .A2(n9666), .ZN(n7971) );
  AND2_X1 U9697 ( .A1(n7972), .A2(n7971), .ZN(n10491) );
  NAND2_X1 U9698 ( .A1(n7973), .A2(n10491), .ZN(n8014) );
  INV_X1 U9699 ( .A(n8014), .ZN(n7982) );
  NAND2_X1 U9700 ( .A1(n7975), .A2(n7974), .ZN(n8447) );
  OAI21_X1 U9701 ( .B1(n7975), .B2(n7974), .A(n8447), .ZN(n8016) );
  NAND2_X1 U9702 ( .A1(n8016), .A2(n10560), .ZN(n7981) );
  AOI211_X1 U9703 ( .C1(n10503), .C2(n7976), .A(n10308), .B(n8453), .ZN(n8015)
         );
  NOR2_X1 U9704 ( .A1(n4837), .A2(n10556), .ZN(n7979) );
  OAI22_X1 U9705 ( .A1(n5878), .A2(n7977), .B1(n10505), .B2(n10270), .ZN(n7978) );
  AOI211_X1 U9706 ( .C1(n8015), .C2(n10548), .A(n7979), .B(n7978), .ZN(n7980)
         );
  OAI211_X1 U9707 ( .C1(n10553), .C2(n7982), .A(n7981), .B(n7980), .ZN(
        P1_U3281) );
  AOI21_X1 U9708 ( .B1(n8010), .B2(n7984), .A(n8714), .ZN(n8000) );
  AOI21_X1 U9709 ( .B1(n7987), .B2(n7986), .A(n8698), .ZN(n7997) );
  MUX2_X1 U9710 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8798), .Z(n8703) );
  XNOR2_X1 U9711 ( .A(n8713), .B(n8703), .ZN(n7993) );
  OR2_X1 U9712 ( .A1(n7989), .A2(n7988), .ZN(n7991) );
  NAND2_X1 U9713 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  NAND2_X1 U9714 ( .A1(n7993), .A2(n7992), .ZN(n8705) );
  OAI21_X1 U9715 ( .B1(n7993), .B2(n7992), .A(n8705), .ZN(n7994) );
  AOI22_X1 U9716 ( .A1(n10650), .A2(n8713), .B1(n10652), .B2(n7994), .ZN(n7996) );
  AND2_X1 U9717 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8090) );
  INV_X1 U9718 ( .A(n8090), .ZN(n7995) );
  OAI211_X1 U9719 ( .C1(n7997), .C2(n8841), .A(n7996), .B(n7995), .ZN(n7998)
         );
  AOI21_X1 U9720 ( .B1(n8839), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7998), .ZN(
        n7999) );
  OAI21_X1 U9721 ( .B1(n8000), .B2(n8806), .A(n7999), .ZN(P2_U3195) );
  XOR2_X1 U9722 ( .A(n8326), .B(n8001), .Z(n8002) );
  AOI222_X1 U9723 ( .A1(n9017), .A2(n8002), .B1(n8662), .B2(n9012), .C1(n8661), 
        .C2(n9014), .ZN(n9453) );
  INV_X1 U9724 ( .A(n8644), .ZN(n8003) );
  OAI22_X1 U9725 ( .A1(n9020), .A2(n9270), .B1(n8003), .B2(n9018), .ZN(n8004)
         );
  AOI21_X1 U9726 ( .B1(n8634), .B2(n9023), .A(n8004), .ZN(n8007) );
  INV_X1 U9727 ( .A(n8326), .ZN(n8005) );
  NAND2_X1 U9728 ( .A1(n4646), .A2(n8005), .ZN(n9451) );
  NAND3_X1 U9729 ( .A1(n9451), .A2(n9004), .A3(n9450), .ZN(n8006) );
  OAI211_X1 U9730 ( .C1(n9453), .C2(n9000), .A(n8007), .B(n8006), .ZN(P2_U3218) );
  INV_X1 U9731 ( .A(n8318), .ZN(n8096) );
  AOI21_X1 U9732 ( .B1(n8009), .B2(n9449), .A(n8008), .ZN(n8012) );
  MUX2_X1 U9733 ( .A(n8010), .B(n8012), .S(n9456), .Z(n8011) );
  OAI21_X1 U9734 ( .B1(n8096), .B2(n9442), .A(n8011), .ZN(P2_U3472) );
  MUX2_X1 U9735 ( .A(n9402), .B(n8012), .S(n10683), .Z(n8013) );
  OAI21_X1 U9736 ( .B1(n8096), .B2(n9514), .A(n8013), .ZN(P2_U3429) );
  AOI211_X1 U9737 ( .C1(n8016), .C2(n10622), .A(n8015), .B(n8014), .ZN(n8021)
         );
  INV_X1 U9738 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8017) );
  NOR2_X1 U9739 ( .A1(n10449), .A2(n8017), .ZN(n8018) );
  AOI21_X1 U9740 ( .B1(n10503), .B2(n10453), .A(n8018), .ZN(n8019) );
  OAI21_X1 U9741 ( .B1(n8021), .B2(n10634), .A(n8019), .ZN(P1_U3489) );
  AOI22_X1 U9742 ( .A1(n10503), .A2(n10392), .B1(n10641), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n8020) );
  OAI21_X1 U9743 ( .B1(n8021), .B2(n10641), .A(n8020), .ZN(P1_U3534) );
  XNOR2_X1 U9744 ( .A(n8030), .B(n8546), .ZN(n8084) );
  XNOR2_X1 U9745 ( .A(n8084), .B(n8664), .ZN(n8082) );
  XNOR2_X1 U9746 ( .A(n8083), .B(n8082), .ZN(n8032) );
  NAND2_X1 U9747 ( .A1(n8645), .A2(n8024), .ZN(n8027) );
  AOI21_X1 U9748 ( .B1(n8639), .B2(n8663), .A(n8025), .ZN(n8026) );
  OAI211_X1 U9749 ( .C1(n8028), .C2(n8641), .A(n8027), .B(n8026), .ZN(n8029)
         );
  AOI21_X1 U9750 ( .B1(n8030), .B2(n8629), .A(n8029), .ZN(n8031) );
  OAI21_X1 U9751 ( .B1(n8032), .B2(n8632), .A(n8031), .ZN(P2_U3164) );
  INV_X1 U9752 ( .A(n8033), .ZN(n8470) );
  OAI222_X1 U9753 ( .A1(n8035), .A2(P1_U3086), .B1(n10472), .B2(n8470), .C1(
        n8034), .C2(n10470), .ZN(P1_U3331) );
  NOR2_X1 U9754 ( .A1(n8118), .A2(n8905), .ZN(n8038) );
  AND2_X1 U9755 ( .A1(n8323), .A2(n8324), .ZN(n8320) );
  XNOR2_X1 U9756 ( .A(n8036), .B(n8320), .ZN(n8037) );
  OAI222_X1 U9757 ( .A1(n8993), .A2(n8113), .B1(n8953), .B2(n8575), .C1(n8990), 
        .C2(n8037), .ZN(n8042) );
  AOI211_X1 U9758 ( .C1(n8999), .C2(n8115), .A(n8038), .B(n8042), .ZN(n8041)
         );
  INV_X1 U9759 ( .A(n8320), .ZN(n8204) );
  XNOR2_X1 U9760 ( .A(n8039), .B(n8204), .ZN(n8043) );
  AOI22_X1 U9761 ( .A1(n8043), .A2(n9004), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9022), .ZN(n8040) );
  OAI21_X1 U9762 ( .B1(n8041), .B2(n9022), .A(n8040), .ZN(P2_U3219) );
  AOI21_X1 U9763 ( .B1(n9449), .B2(n8043), .A(n8042), .ZN(n8045) );
  MUX2_X1 U9764 ( .A(n8701), .B(n8045), .S(n9456), .Z(n8044) );
  OAI21_X1 U9765 ( .B1(n8118), .B2(n9442), .A(n8044), .ZN(P2_U3473) );
  MUX2_X1 U9766 ( .A(n8046), .B(n8045), .S(n10683), .Z(n8047) );
  OAI21_X1 U9767 ( .B1(n8118), .B2(n9514), .A(n8047), .ZN(P2_U3432) );
  INV_X1 U9768 ( .A(n8048), .ZN(n8416) );
  OAI222_X1 U9769 ( .A1(n5792), .A2(P1_U3086), .B1(n10472), .B2(n8416), .C1(
        n8049), .C2(n10470), .ZN(P1_U3330) );
  XOR2_X1 U9770 ( .A(n10033), .B(n8057), .Z(n8052) );
  INV_X1 U9771 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8051) );
  NOR2_X1 U9772 ( .A1(n8051), .A2(n8052), .ZN(n10034) );
  AOI211_X1 U9773 ( .C1(n8052), .C2(n8051), .A(n10034), .B(n10037), .ZN(n8062)
         );
  XNOR2_X1 U9774 ( .A(n10032), .B(n10024), .ZN(n8056) );
  NOR2_X1 U9775 ( .A1(n8055), .A2(n8056), .ZN(n10025) );
  AOI211_X1 U9776 ( .C1(n8056), .C2(n8055), .A(n10025), .B(n10090), .ZN(n8061)
         );
  INV_X1 U9777 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U9778 ( .A1(n10072), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U9779 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n8058) );
  OAI211_X1 U9780 ( .C1(n9255), .C2(n10099), .A(n8059), .B(n8058), .ZN(n8060)
         );
  OR3_X1 U9781 ( .A1(n8062), .A2(n8061), .A3(n8060), .ZN(P1_U3258) );
  AOI21_X1 U9782 ( .B1(n8063), .B2(n9743), .A(n10302), .ZN(n8066) );
  NAND2_X1 U9783 ( .A1(n9972), .A2(n9667), .ZN(n8065) );
  NAND2_X1 U9784 ( .A1(n9974), .A2(n9666), .ZN(n8064) );
  NAND2_X1 U9785 ( .A1(n8065), .A2(n8064), .ZN(n9530) );
  AOI21_X1 U9786 ( .B1(n8066), .B2(n10299), .A(n9530), .ZN(n8075) );
  XNOR2_X1 U9787 ( .A(n8067), .B(n9743), .ZN(n8078) );
  NAND2_X1 U9788 ( .A1(n8078), .A2(n10560), .ZN(n8073) );
  OAI22_X1 U9789 ( .A1(n5878), .A2(n8068), .B1(n9532), .B2(n10270), .ZN(n8071)
         );
  INV_X1 U9790 ( .A(n8452), .ZN(n8069) );
  OAI211_X1 U9791 ( .C1(n8069), .C2(n8076), .A(n10319), .B(n10309), .ZN(n8074)
         );
  NOR2_X1 U9792 ( .A1(n8074), .A2(n10275), .ZN(n8070) );
  AOI211_X1 U9793 ( .C1(n10278), .C2(n9534), .A(n8071), .B(n8070), .ZN(n8072)
         );
  OAI211_X1 U9794 ( .C1(n10563), .C2(n8075), .A(n8073), .B(n8072), .ZN(
        P1_U3279) );
  OAI211_X1 U9795 ( .C1(n8076), .C2(n10617), .A(n8075), .B(n8074), .ZN(n8077)
         );
  AOI21_X1 U9796 ( .B1(n8078), .B2(n10622), .A(n8077), .ZN(n8081) );
  NAND2_X1 U9797 ( .A1(n10634), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8079) );
  OAI21_X1 U9798 ( .B1(n8081), .B2(n10634), .A(n8079), .ZN(P1_U3495) );
  NAND2_X1 U9799 ( .A1(n10641), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8080) );
  OAI21_X1 U9800 ( .B1(n8081), .B2(n10641), .A(n8080), .ZN(P1_U3536) );
  INV_X1 U9801 ( .A(n8084), .ZN(n8085) );
  XNOR2_X1 U9802 ( .A(n8318), .B(n8517), .ZN(n8086) );
  NOR2_X1 U9803 ( .A1(n8086), .A2(n8663), .ZN(n8106) );
  AOI21_X1 U9804 ( .B1(n8086), .B2(n8663), .A(n8106), .ZN(n8087) );
  OAI21_X1 U9805 ( .B1(n8088), .B2(n8087), .A(n8110), .ZN(n8089) );
  NAND2_X1 U9806 ( .A1(n8089), .A2(n8635), .ZN(n8095) );
  AOI21_X1 U9807 ( .B1(n8624), .B2(n8664), .A(n8090), .ZN(n8091) );
  OAI21_X1 U9808 ( .B1(n8642), .B2(n8627), .A(n8091), .ZN(n8092) );
  AOI21_X1 U9809 ( .B1(n8645), .B2(n8093), .A(n8092), .ZN(n8094) );
  OAI211_X1 U9810 ( .C1(n8096), .C2(n8648), .A(n8095), .B(n8094), .ZN(P2_U3174) );
  INV_X1 U9811 ( .A(n8097), .ZN(n8101) );
  OAI222_X1 U9812 ( .A1(n8099), .A2(P1_U3086), .B1(n10472), .B2(n8101), .C1(
        n8098), .C2(n10470), .ZN(P1_U3329) );
  OAI222_X1 U9813 ( .A1(n8102), .A2(P2_U3151), .B1(n9524), .B2(n8101), .C1(
        n8100), .C2(n8484), .ZN(P2_U3269) );
  INV_X1 U9814 ( .A(n8103), .ZN(n8157) );
  AOI21_X1 U9815 ( .B1(n9522), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8104), .ZN(
        n8105) );
  OAI21_X1 U9816 ( .B1(n8157), .B2(n9524), .A(n8105), .ZN(P2_U3268) );
  INV_X1 U9817 ( .A(n8106), .ZN(n8108) );
  XNOR2_X1 U9818 ( .A(n8107), .B(n8517), .ZN(n8493) );
  XNOR2_X1 U9819 ( .A(n8493), .B(n8662), .ZN(n8109) );
  AND3_X1 U9820 ( .A1(n8110), .A2(n8109), .A3(n8108), .ZN(n8111) );
  OAI21_X1 U9821 ( .B1(n8494), .B2(n8111), .A(n8635), .ZN(n8117) );
  NAND2_X1 U9822 ( .A1(n8639), .A2(n9013), .ZN(n8112) );
  NAND2_X1 U9823 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U9824 ( .C1(n8113), .C2(n8641), .A(n8112), .B(n8710), .ZN(n8114)
         );
  AOI21_X1 U9825 ( .B1(n8645), .B2(n8115), .A(n8114), .ZN(n8116) );
  OAI211_X1 U9826 ( .C1(n8118), .C2(n8648), .A(n8117), .B(n8116), .ZN(P2_U3155) );
  NAND2_X1 U9827 ( .A1(n8159), .A2(n8119), .ZN(n8121) );
  OAI211_X1 U9828 ( .C1(n8484), .C2(n8122), .A(n8121), .B(n8120), .ZN(P2_U3267) );
  INV_X1 U9829 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U9830 ( .A1(n10710), .A2(n10711), .ZN(n10709) );
  NAND2_X1 U9831 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n8147) );
  XNOR2_X1 U9832 ( .A(n8123), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n10715) );
  NOR2_X1 U9833 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10716) );
  AOI22_X1 U9834 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9412), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n8129), .ZN(n10738) );
  NAND2_X1 U9835 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8127) );
  INV_X1 U9836 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9999) );
  XNOR2_X1 U9837 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n9999), .ZN(n10736) );
  NAND2_X1 U9838 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8125) );
  XOR2_X1 U9839 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10734) );
  AOI21_X1 U9840 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10686) );
  NAND3_X1 U9841 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10688) );
  OAI21_X1 U9842 ( .B1(n10686), .B2(n10690), .A(n10688), .ZN(n10733) );
  NAND2_X1 U9843 ( .A1(n10734), .A2(n10733), .ZN(n8124) );
  NAND2_X1 U9844 ( .A1(n8125), .A2(n8124), .ZN(n10735) );
  NAND2_X1 U9845 ( .A1(n10736), .A2(n10735), .ZN(n8126) );
  NAND2_X1 U9846 ( .A1(n8127), .A2(n8126), .ZN(n10737) );
  NOR2_X1 U9847 ( .A1(n10738), .A2(n10737), .ZN(n8128) );
  AOI21_X1 U9848 ( .B1(n8129), .B2(n9412), .A(n8128), .ZN(n8130) );
  NOR2_X1 U9849 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8130), .ZN(n10722) );
  AND2_X1 U9850 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8130), .ZN(n10721) );
  NOR2_X1 U9851 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10721), .ZN(n8131) );
  NOR2_X1 U9852 ( .A1(n10722), .A2(n8131), .ZN(n8133) );
  NAND2_X1 U9853 ( .A1(n8133), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8135) );
  XNOR2_X1 U9854 ( .A(n8133), .B(n8132), .ZN(n10720) );
  NAND2_X1 U9855 ( .A1(n10720), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U9856 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  AND2_X1 U9857 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8136), .ZN(n8137) );
  XNOR2_X1 U9858 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8136), .ZN(n10728) );
  NOR2_X1 U9859 ( .A1(n10729), .A2(n10728), .ZN(n10727) );
  NOR2_X1 U9860 ( .A1(n8138), .A2(n10015), .ZN(n8139) );
  INV_X1 U9861 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10732) );
  XOR2_X1 U9862 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8138), .Z(n10731) );
  NOR2_X1 U9863 ( .A1(n10732), .A2(n10731), .ZN(n10730) );
  INV_X1 U9864 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n8140) );
  NOR2_X1 U9865 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  INV_X1 U9866 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10726) );
  XOR2_X1 U9867 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8141), .Z(n10725) );
  NOR2_X1 U9868 ( .A1(n10726), .A2(n10725), .ZN(n10724) );
  NOR2_X1 U9869 ( .A1(n8142), .A2(n10724), .ZN(n10719) );
  NOR2_X1 U9870 ( .A1(n8144), .A2(n8143), .ZN(n10717) );
  INV_X1 U9871 ( .A(n10717), .ZN(n8145) );
  OAI21_X1 U9872 ( .B1(n10716), .B2(n10719), .A(n8145), .ZN(n10714) );
  NAND2_X1 U9873 ( .A1(n10715), .A2(n10714), .ZN(n8146) );
  NAND2_X1 U9874 ( .A1(n8147), .A2(n8146), .ZN(n10712) );
  AOI22_X1 U9875 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .B1(n10709), .B2(n10712), .ZN(n10708) );
  INV_X1 U9876 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8148) );
  AOI22_X1 U9877 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8148), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(n9288), .ZN(n10707) );
  NOR2_X1 U9878 ( .A1(n10708), .A2(n10707), .ZN(n10706) );
  AOI21_X1 U9879 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10706), .ZN(n10705) );
  INV_X1 U9880 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8149) );
  AOI22_X1 U9881 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n8149), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(n9292), .ZN(n10704) );
  NOR2_X1 U9882 ( .A1(n10705), .A2(n10704), .ZN(n10703) );
  AOI21_X1 U9883 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10703), .ZN(n10702) );
  INV_X1 U9884 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8735) );
  AOI22_X1 U9885 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n8735), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n9255), .ZN(n10701) );
  NOR2_X1 U9886 ( .A1(n10702), .A2(n10701), .ZN(n10700) );
  AOI21_X1 U9887 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10700), .ZN(n10699) );
  NAND2_X1 U9888 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8150) );
  OAI21_X1 U9889 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n8150), .ZN(n10698) );
  NOR2_X1 U9890 ( .A1(n10699), .A2(n10698), .ZN(n10697) );
  AOI21_X1 U9891 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10697), .ZN(n10696) );
  INV_X1 U9892 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8151) );
  INV_X1 U9893 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9160) );
  AOI22_X1 U9894 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8151), .B1(
        P2_ADDR_REG_17__SCAN_IN), .B2(n9160), .ZN(n10695) );
  NOR2_X1 U9895 ( .A1(n10696), .A2(n10695), .ZN(n10694) );
  AOI21_X1 U9896 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10694), .ZN(n8152) );
  INV_X1 U9897 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U9898 ( .A1(n8152), .A2(n10063), .ZN(n8153) );
  INV_X1 U9899 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10693) );
  XOR2_X1 U9900 ( .A(n8152), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n10692) );
  NOR2_X1 U9901 ( .A1(n10693), .A2(n10692), .ZN(n10691) );
  NOR2_X1 U9902 ( .A1(n8153), .A2(n10691), .ZN(n8156) );
  XNOR2_X1 U9903 ( .A(n8154), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8155) );
  XNOR2_X1 U9904 ( .A(n8156), .B(n8155), .ZN(ADD_1068_U4) );
  OAI222_X1 U9905 ( .A1(n10470), .A2(n8158), .B1(P1_U3086), .B2(n4558), .C1(
        n10472), .C2(n8157), .ZN(P1_U3328) );
  INV_X1 U9906 ( .A(n8159), .ZN(n8160) );
  OAI222_X1 U9907 ( .A1(n10470), .A2(n8161), .B1(P1_U3086), .B2(n5871), .C1(
        n10472), .C2(n8160), .ZN(P1_U3327) );
  INV_X1 U9908 ( .A(n8162), .ZN(n8164) );
  NAND2_X1 U9909 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  MUX2_X1 U9910 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8171), .Z(n8167) );
  XNOR2_X1 U9911 ( .A(n8167), .B(SI_30_), .ZN(n8182) );
  OAI22_X1 U9912 ( .A1(n8183), .A2(n8182), .B1(SI_30_), .B2(n8167), .ZN(n8170)
         );
  INV_X1 U9913 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9674) );
  MUX2_X1 U9914 ( .A(n9674), .B(n6765), .S(n8171), .Z(n8168) );
  XNOR2_X1 U9915 ( .A(n8168), .B(SI_31_), .ZN(n8169) );
  XNOR2_X1 U9916 ( .A(n8170), .B(n8169), .ZN(n9673) );
  MUX2_X1 U9917 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9673), .S(n8171), .Z(n8173) );
  INV_X1 U9918 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U9919 ( .A1(n8174), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8177) );
  INV_X1 U9920 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8175) );
  OR2_X1 U9921 ( .A1(n6270), .A2(n8175), .ZN(n8176) );
  OAI211_X1 U9922 ( .C1(n8178), .C2(n6569), .A(n8177), .B(n8176), .ZN(n8179)
         );
  INV_X1 U9923 ( .A(n8179), .ZN(n8180) );
  AND2_X1 U9924 ( .A1(n8226), .A2(n8849), .ZN(n8401) );
  INV_X1 U9925 ( .A(n8401), .ZN(n8220) );
  NAND2_X1 U9926 ( .A1(n9789), .A2(n4541), .ZN(n8185) );
  INV_X1 U9927 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8417) );
  OR2_X1 U9928 ( .A1(n6276), .A2(n8417), .ZN(n8184) );
  NAND2_X1 U9929 ( .A1(n8185), .A2(n8184), .ZN(n9029) );
  OR2_X1 U9930 ( .A1(n9029), .A2(n8186), .ZN(n8399) );
  NAND2_X1 U9931 ( .A1(n9029), .A2(n8186), .ZN(n8232) );
  NAND2_X1 U9932 ( .A1(n8378), .A2(n8379), .ZN(n8888) );
  INV_X1 U9933 ( .A(n8888), .ZN(n8884) );
  INV_X1 U9934 ( .A(n8988), .ZN(n8997) );
  INV_X1 U9935 ( .A(n8980), .ZN(n8210) );
  NAND4_X1 U9936 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n8192)
         );
  NOR2_X1 U9937 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  NAND4_X1 U9938 ( .A1(n8298), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n8196)
         );
  OR3_X1 U9939 ( .A1(n8198), .A2(n8197), .A3(n8196), .ZN(n8199) );
  NOR2_X1 U9940 ( .A1(n8200), .A2(n8199), .ZN(n8202) );
  NAND3_X1 U9941 ( .A1(n8314), .A2(n8202), .A3(n8201), .ZN(n8203) );
  NOR2_X1 U9942 ( .A1(n8204), .A2(n8203), .ZN(n8206) );
  NAND3_X1 U9943 ( .A1(n8326), .A2(n8206), .A3(n8205), .ZN(n8207) );
  NOR2_X1 U9944 ( .A1(n8208), .A2(n8207), .ZN(n8209) );
  NAND4_X1 U9945 ( .A1(n8963), .A2(n8997), .A3(n8210), .A4(n8209), .ZN(n8211)
         );
  NOR2_X1 U9946 ( .A1(n8955), .A2(n8211), .ZN(n8212) );
  NAND4_X1 U9947 ( .A1(n8920), .A2(n8931), .A3(n8940), .A4(n8212), .ZN(n8214)
         );
  NAND2_X1 U9948 ( .A1(n8363), .A2(n8213), .ZN(n8914) );
  NOR2_X1 U9949 ( .A1(n8214), .A2(n8914), .ZN(n8215) );
  NAND4_X1 U9950 ( .A1(n8877), .A2(n8884), .A3(n8900), .A4(n8215), .ZN(n8216)
         );
  NOR2_X1 U9951 ( .A1(n8868), .A2(n8216), .ZN(n8217) );
  AND4_X1 U9952 ( .A1(n8399), .A2(n8232), .A3(n8223), .A4(n8217), .ZN(n8219)
         );
  INV_X1 U9953 ( .A(n8849), .ZN(n8649) );
  AND2_X1 U9954 ( .A1(n9459), .A2(n8649), .ZN(n8404) );
  INV_X1 U9955 ( .A(n8404), .ZN(n8218) );
  NAND3_X1 U9956 ( .A1(n8220), .A2(n8219), .A3(n8218), .ZN(n8231) );
  AND2_X1 U9957 ( .A1(n8232), .A2(n8221), .ZN(n8388) );
  INV_X1 U9958 ( .A(n8388), .ZN(n8222) );
  AOI21_X1 U9959 ( .B1(n8224), .B2(n8223), .A(n8222), .ZN(n8225) );
  NOR2_X1 U9960 ( .A1(n8225), .A2(n8401), .ZN(n8228) );
  INV_X1 U9961 ( .A(n9029), .ZN(n9462) );
  AOI21_X1 U9962 ( .B1(n8849), .B2(n9462), .A(n8226), .ZN(n8227) );
  OAI22_X1 U9963 ( .A1(n8228), .A2(n8227), .B1(n9459), .B2(n8399), .ZN(n8230)
         );
  INV_X1 U9964 ( .A(n8232), .ZN(n8398) );
  MUX2_X1 U9965 ( .A(n8652), .B(n8518), .S(n8402), .Z(n8382) );
  NAND2_X1 U9966 ( .A1(n8911), .A2(n8233), .ZN(n8236) );
  NAND2_X1 U9967 ( .A1(n8362), .A2(n8234), .ZN(n8235) );
  MUX2_X1 U9968 ( .A(n8236), .B(n8235), .S(n8392), .Z(n8237) );
  INV_X1 U9969 ( .A(n8237), .ZN(n8361) );
  NAND2_X1 U9970 ( .A1(n8357), .A2(n8346), .ZN(n8238) );
  NAND3_X1 U9971 ( .A1(n8238), .A2(n8402), .A3(n8349), .ZN(n8239) );
  NAND2_X1 U9972 ( .A1(n8239), .A2(n8952), .ZN(n8240) );
  NAND2_X1 U9973 ( .A1(n9501), .A2(n8240), .ZN(n8356) );
  NOR2_X1 U9974 ( .A1(n8658), .A2(n8392), .ZN(n8347) );
  NAND2_X1 U9975 ( .A1(n8560), .A2(n8347), .ZN(n8345) );
  NAND2_X1 U9976 ( .A1(n8346), .A2(n8337), .ZN(n8242) );
  AOI21_X1 U9977 ( .B1(n8392), .B2(n8242), .A(n8241), .ZN(n8344) );
  AND2_X1 U9978 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  OAI211_X1 U9979 ( .C1(n8257), .C2(n8246), .A(n8304), .B(n4588), .ZN(n8255)
         );
  NAND2_X1 U9980 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  AND2_X1 U9981 ( .A1(n8250), .A2(n8249), .ZN(n8253) );
  OAI211_X1 U9982 ( .C1(n8257), .C2(n8253), .A(n8252), .B(n8251), .ZN(n8254)
         );
  MUX2_X1 U9983 ( .A(n8255), .B(n8254), .S(n8392), .Z(n8256) );
  INV_X1 U9984 ( .A(n8256), .ZN(n8301) );
  INV_X1 U9985 ( .A(n8257), .ZN(n8299) );
  NAND2_X1 U9986 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U9987 ( .A1(n8260), .A2(n8263), .ZN(n8265) );
  NAND3_X1 U9988 ( .A1(n8263), .A2(n8262), .A3(n8261), .ZN(n8264) );
  NAND2_X1 U9989 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  MUX2_X1 U9990 ( .A(n8266), .B(n8265), .S(n8392), .Z(n8275) );
  NAND2_X1 U9991 ( .A1(n8286), .A2(n8267), .ZN(n8271) );
  OAI21_X1 U9992 ( .B1(n8269), .B2(n8268), .A(n8278), .ZN(n8270) );
  MUX2_X1 U9993 ( .A(n8271), .B(n8270), .S(n8392), .Z(n8272) );
  INV_X1 U9994 ( .A(n8272), .ZN(n8273) );
  OAI21_X1 U9995 ( .B1(n8275), .B2(n8274), .A(n8273), .ZN(n8277) );
  NAND2_X1 U9996 ( .A1(n8277), .A2(n8276), .ZN(n8292) );
  INV_X1 U9997 ( .A(n8278), .ZN(n8280) );
  OAI211_X1 U9998 ( .C1(n8292), .C2(n8280), .A(n8294), .B(n8279), .ZN(n8284)
         );
  NAND2_X1 U9999 ( .A1(n8285), .A2(n8281), .ZN(n8289) );
  NAND2_X1 U10000 ( .A1(n8289), .A2(n8282), .ZN(n8283) );
  NAND2_X1 U10001 ( .A1(n8284), .A2(n8283), .ZN(n8296) );
  INV_X1 U10002 ( .A(n8286), .ZN(n8291) );
  INV_X1 U10003 ( .A(n8287), .ZN(n8288) );
  NOR2_X1 U10004 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  OAI21_X1 U10005 ( .B1(n8292), .B2(n8291), .A(n8290), .ZN(n8293) );
  OAI21_X1 U10006 ( .B1(n8294), .B2(n5063), .A(n8293), .ZN(n8295) );
  MUX2_X1 U10007 ( .A(n8296), .B(n8295), .S(n8392), .Z(n8297) );
  NAND3_X1 U10008 ( .A1(n8299), .A2(n8298), .A3(n8297), .ZN(n8300) );
  NAND2_X1 U10009 ( .A1(n8301), .A2(n8300), .ZN(n8305) );
  INV_X1 U10010 ( .A(n8308), .ZN(n8302) );
  AOI21_X1 U10011 ( .B1(n8305), .B2(n8303), .A(n8302), .ZN(n8310) );
  NAND2_X1 U10012 ( .A1(n8305), .A2(n8304), .ZN(n8307) );
  NAND2_X1 U10013 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  MUX2_X1 U10014 ( .A(n8312), .B(n8311), .S(n8392), .Z(n8313) );
  MUX2_X1 U10015 ( .A(n8663), .B(n8318), .S(n8392), .Z(n8315) );
  AOI21_X1 U10016 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(n8322) );
  AND3_X1 U10017 ( .A1(n8319), .A2(n8663), .A3(n8318), .ZN(n8321) );
  OAI21_X1 U10018 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8327) );
  MUX2_X1 U10019 ( .A(n8324), .B(n8323), .S(n8392), .Z(n8325) );
  MUX2_X1 U10020 ( .A(n8329), .B(n8328), .S(n8392), .Z(n8330) );
  INV_X1 U10021 ( .A(n8331), .ZN(n8334) );
  INV_X1 U10022 ( .A(n8332), .ZN(n8333) );
  MUX2_X1 U10023 ( .A(n8334), .B(n8333), .S(n8392), .Z(n8335) );
  NOR2_X1 U10024 ( .A1(n8988), .A2(n8335), .ZN(n8339) );
  AOI21_X1 U10025 ( .B1(n8337), .B2(n8336), .A(n8392), .ZN(n8338) );
  AND2_X1 U10026 ( .A1(n8341), .A2(n8340), .ZN(n8342) );
  OR2_X1 U10027 ( .A1(n8349), .A2(n8392), .ZN(n8352) );
  NAND4_X1 U10028 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8352), .ZN(n8355)
         );
  NAND3_X1 U10029 ( .A1(n8357), .A2(n8402), .A3(n8346), .ZN(n8353) );
  INV_X1 U10030 ( .A(n8347), .ZN(n8351) );
  NAND3_X1 U10031 ( .A1(n8349), .A2(n8392), .A3(n8348), .ZN(n8350) );
  NAND4_X1 U10032 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n8354)
         );
  NAND2_X1 U10033 ( .A1(n8358), .A2(n8357), .ZN(n8359) );
  AND2_X1 U10034 ( .A1(n8363), .A2(n8362), .ZN(n8365) );
  AOI21_X1 U10035 ( .B1(n8368), .B2(n8365), .A(n8364), .ZN(n8370) );
  AOI21_X1 U10036 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8369) );
  MUX2_X1 U10037 ( .A(n8370), .B(n8369), .S(n8392), .Z(n8371) );
  NAND2_X1 U10038 ( .A1(n8371), .A2(n8900), .ZN(n8377) );
  INV_X1 U10039 ( .A(n8372), .ZN(n8373) );
  MUX2_X1 U10040 ( .A(n8374), .B(n8373), .S(n8402), .Z(n8375) );
  NOR2_X1 U10041 ( .A1(n8888), .A2(n8375), .ZN(n8376) );
  NAND2_X1 U10042 ( .A1(n8377), .A2(n8376), .ZN(n8381) );
  MUX2_X1 U10043 ( .A(n8379), .B(n8378), .S(n8392), .Z(n8380) );
  INV_X1 U10044 ( .A(n8387), .ZN(n8397) );
  MUX2_X1 U10045 ( .A(n8876), .B(n9474), .S(n8402), .Z(n8384) );
  INV_X1 U10046 ( .A(n8384), .ZN(n8396) );
  OR2_X1 U10047 ( .A1(n8385), .A2(n8384), .ZN(n8386) );
  OAI21_X1 U10048 ( .B1(n8391), .B2(n8651), .A(n8388), .ZN(n8394) );
  AND2_X1 U10049 ( .A1(n8399), .A2(n8389), .ZN(n8390) );
  OAI21_X1 U10050 ( .B1(n8391), .B2(n8552), .A(n8390), .ZN(n8393) );
  AOI211_X1 U10051 ( .C1(n8402), .C2(n8399), .A(n8398), .B(n8403), .ZN(n8400)
         );
  NAND3_X1 U10052 ( .A1(n8409), .A2(n8408), .A3(n8798), .ZN(n8410) );
  OAI211_X1 U10053 ( .C1(n8411), .C2(n8413), .A(n8410), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8412) );
  OAI21_X1 U10054 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(P2_U3296) );
  OAI222_X1 U10055 ( .A1(n6641), .A2(P2_U3151), .B1(n9524), .B2(n8416), .C1(
        n8415), .C2(n8484), .ZN(P2_U3270) );
  INV_X1 U10056 ( .A(n9789), .ZN(n10468) );
  OAI222_X1 U10057 ( .A1(n6191), .A2(P2_U3151), .B1(n9524), .B2(n10468), .C1(
        n8417), .C2(n8484), .ZN(P2_U3265) );
  XNOR2_X1 U10058 ( .A(n8418), .B(n8423), .ZN(n8440) );
  INV_X1 U10059 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8427) );
  INV_X1 U10060 ( .A(n10137), .ZN(n8420) );
  INV_X1 U10061 ( .A(n10121), .ZN(n8419) );
  AOI211_X1 U10062 ( .C1(n8479), .C2(n8420), .A(n10308), .B(n8419), .ZN(n8432)
         );
  OAI21_X1 U10063 ( .B1(n8423), .B2(n8422), .A(n8421), .ZN(n8424) );
  NAND2_X1 U10064 ( .A1(n8424), .A2(n10285), .ZN(n8426) );
  AND2_X1 U10065 ( .A1(n9961), .A2(n9666), .ZN(n8425) );
  AOI21_X1 U10066 ( .B1(n9959), .B2(n9667), .A(n8425), .ZN(n8477) );
  NAND2_X1 U10067 ( .A1(n8426), .A2(n8477), .ZN(n8438) );
  AOI211_X1 U10068 ( .C1(n10626), .C2(n8479), .A(n8432), .B(n8438), .ZN(n8429)
         );
  MUX2_X1 U10069 ( .A(n8427), .B(n8429), .S(n10449), .Z(n8428) );
  OAI21_X1 U10070 ( .B1(n8440), .B2(n10447), .A(n8428), .ZN(P1_U3517) );
  INV_X1 U10071 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8430) );
  MUX2_X1 U10072 ( .A(n8430), .B(n8429), .S(n10643), .Z(n8431) );
  OAI21_X1 U10073 ( .B1(n8440), .B2(n10381), .A(n8431), .ZN(P1_U3549) );
  NAND2_X1 U10074 ( .A1(n8432), .A2(n10548), .ZN(n8435) );
  INV_X1 U10075 ( .A(n8433), .ZN(n8475) );
  AOI22_X1 U10076 ( .A1(n8475), .A2(n10551), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10563), .ZN(n8434) );
  OAI211_X1 U10077 ( .C1(n8436), .C2(n10556), .A(n8435), .B(n8434), .ZN(n8437)
         );
  AOI21_X1 U10078 ( .B1(n10241), .B2(n8438), .A(n8437), .ZN(n8439) );
  OAI21_X1 U10079 ( .B1(n8440), .B2(n10259), .A(n8439), .ZN(P1_U3266) );
  NAND2_X1 U10080 ( .A1(n8441), .A2(n9739), .ZN(n8442) );
  XNOR2_X1 U10081 ( .A(n8442), .B(n9823), .ZN(n8446) );
  NAND2_X1 U10082 ( .A1(n9973), .A2(n9667), .ZN(n8444) );
  NAND2_X1 U10083 ( .A1(n9975), .A2(n9666), .ZN(n8443) );
  AND2_X1 U10084 ( .A1(n8444), .A2(n8443), .ZN(n9624) );
  INV_X1 U10085 ( .A(n9624), .ZN(n8445) );
  AOI21_X1 U10086 ( .B1(n8446), .B2(n10285), .A(n8445), .ZN(n8461) );
  NAND2_X1 U10087 ( .A1(n8448), .A2(n8447), .ZN(n8450) );
  OAI21_X1 U10088 ( .B1(n8450), .B2(n9823), .A(n8449), .ZN(n8459) );
  NAND2_X1 U10089 ( .A1(n8459), .A2(n10560), .ZN(n8458) );
  OAI22_X1 U10090 ( .A1(n5878), .A2(n8451), .B1(n9622), .B2(n10270), .ZN(n8455) );
  OAI211_X1 U10091 ( .C1(n8453), .C2(n9629), .A(n8452), .B(n10319), .ZN(n8460)
         );
  NOR2_X1 U10092 ( .A1(n8460), .A2(n10275), .ZN(n8454) );
  AOI211_X1 U10093 ( .C1(n10278), .C2(n8456), .A(n8455), .B(n8454), .ZN(n8457)
         );
  OAI211_X1 U10094 ( .C1(n10563), .C2(n8461), .A(n8458), .B(n8457), .ZN(
        P1_U3280) );
  INV_X1 U10095 ( .A(n8459), .ZN(n8468) );
  NAND2_X1 U10096 ( .A1(n8461), .A2(n8460), .ZN(n8466) );
  INV_X1 U10097 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9408) );
  OAI22_X1 U10098 ( .A1(n9629), .A2(n10425), .B1(n10449), .B2(n9408), .ZN(
        n8462) );
  AOI21_X1 U10099 ( .B1(n8466), .B2(n10449), .A(n8462), .ZN(n8463) );
  OAI21_X1 U10100 ( .B1(n8468), .B2(n10447), .A(n8463), .ZN(P1_U3492) );
  OAI22_X1 U10101 ( .A1(n9629), .A2(n10356), .B1(n10643), .B2(n8464), .ZN(
        n8465) );
  AOI21_X1 U10102 ( .B1(n8466), .B2(n10643), .A(n8465), .ZN(n8467) );
  OAI21_X1 U10103 ( .B1(n8468), .B2(n10381), .A(n8467), .ZN(P1_U3535) );
  OAI222_X1 U10104 ( .A1(n6645), .A2(P2_U3151), .B1(n9524), .B2(n8470), .C1(
        n8469), .C2(n8484), .ZN(P2_U3271) );
  NAND2_X1 U10105 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  AND2_X1 U10106 ( .A1(n8474), .A2(n8473), .ZN(n8481) );
  AOI22_X1 U10107 ( .A1(n8475), .A2(n9638), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8476) );
  OAI21_X1 U10108 ( .B1(n8477), .B2(n10492), .A(n8476), .ZN(n8478) );
  AOI21_X1 U10109 ( .B1(n8479), .B2(n10502), .A(n8478), .ZN(n8480) );
  OAI21_X1 U10110 ( .B1(n8481), .B2(n10535), .A(n8480), .ZN(P1_U3214) );
  OAI222_X1 U10111 ( .A1(n8484), .A2(n8483), .B1(P2_U3151), .B2(n8482), .C1(
        n10471), .C2(n9524), .ZN(P2_U3266) );
  MUX2_X1 U10112 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n8488), .S(n10449), .Z(
        n8487) );
  OAI21_X1 U10113 ( .B1(n8491), .B2(n10381), .A(n8490), .ZN(P1_U3551) );
  XNOR2_X1 U10114 ( .A(n8630), .B(n8546), .ZN(n8516) );
  XNOR2_X1 U10115 ( .A(n8492), .B(n8546), .ZN(n8504) );
  INV_X1 U10116 ( .A(n8493), .ZN(n8495) );
  XNOR2_X1 U10117 ( .A(n8634), .B(n8546), .ZN(n8497) );
  XNOR2_X1 U10118 ( .A(n8497), .B(n9013), .ZN(n8637) );
  XNOR2_X1 U10119 ( .A(n9444), .B(n8517), .ZN(n8496) );
  NOR2_X1 U10120 ( .A1(n8496), .A2(n8661), .ZN(n8499) );
  AOI21_X1 U10121 ( .B1(n8496), .B2(n8661), .A(n8499), .ZN(n8570) );
  INV_X1 U10122 ( .A(n8497), .ZN(n8498) );
  NAND2_X1 U10123 ( .A1(n8498), .A2(n9013), .ZN(n8571) );
  INV_X1 U10124 ( .A(n8499), .ZN(n8582) );
  XNOR2_X1 U10125 ( .A(n8580), .B(n8546), .ZN(n8500) );
  NAND2_X1 U10126 ( .A1(n8500), .A2(n8975), .ZN(n8503) );
  INV_X1 U10127 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U10128 ( .A1(n8501), .A2(n9015), .ZN(n8502) );
  NAND2_X1 U10129 ( .A1(n8503), .A2(n8502), .ZN(n8581) );
  INV_X1 U10130 ( .A(n8503), .ZN(n8614) );
  XNOR2_X1 U10131 ( .A(n8504), .B(n8660), .ZN(n8613) );
  XNOR2_X1 U10132 ( .A(n8967), .B(n8517), .ZN(n8536) );
  INV_X1 U10133 ( .A(n8536), .ZN(n8505) );
  XNOR2_X1 U10134 ( .A(n9062), .B(n8546), .ZN(n8506) );
  XNOR2_X1 U10135 ( .A(n8506), .B(n8964), .ZN(n8598) );
  INV_X1 U10136 ( .A(n8506), .ZN(n8507) );
  XNOR2_X1 U10137 ( .A(n8560), .B(n8546), .ZN(n8508) );
  XNOR2_X1 U10138 ( .A(n8508), .B(n8658), .ZN(n8556) );
  XNOR2_X1 U10139 ( .A(n8604), .B(n8546), .ZN(n8509) );
  XNOR2_X1 U10140 ( .A(n8509), .B(n8657), .ZN(n8606) );
  XNOR2_X1 U10141 ( .A(n8533), .B(n8517), .ZN(n8512) );
  OAI22_X2 U10142 ( .A1(n8529), .A2(n8656), .B1(n8512), .B2(n8511), .ZN(n8589)
         );
  XNOR2_X1 U10143 ( .A(n8594), .B(n8546), .ZN(n8513) );
  XNOR2_X1 U10144 ( .A(n8513), .B(n8655), .ZN(n8590) );
  XNOR2_X1 U10145 ( .A(n9043), .B(n8546), .ZN(n8514) );
  XOR2_X1 U10146 ( .A(n8654), .B(n8514), .Z(n8564) );
  INV_X1 U10147 ( .A(n8514), .ZN(n8515) );
  XNOR2_X1 U10148 ( .A(n8516), .B(n8653), .ZN(n8623) );
  XNOR2_X1 U10149 ( .A(n8518), .B(n8517), .ZN(n8519) );
  NAND2_X1 U10150 ( .A1(n8519), .A2(n8652), .ZN(n8544) );
  OAI21_X1 U10151 ( .B1(n8519), .B2(n8652), .A(n8544), .ZN(n8520) );
  AOI21_X1 U10152 ( .B1(n8521), .B2(n8520), .A(n8632), .ZN(n8522) );
  NAND2_X1 U10153 ( .A1(n8522), .A2(n8545), .ZN(n8528) );
  INV_X1 U10154 ( .A(n8879), .ZN(n8525) );
  AOI22_X1 U10155 ( .A1(n8653), .A2(n8624), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8523) );
  OAI21_X1 U10156 ( .B1(n8525), .B2(n8524), .A(n8523), .ZN(n8526) );
  AOI21_X1 U10157 ( .B1(n8651), .B2(n8639), .A(n8526), .ZN(n8527) );
  OAI211_X1 U10158 ( .C1(n9477), .C2(n8648), .A(n8528), .B(n8527), .ZN(
        P2_U3154) );
  XNOR2_X1 U10159 ( .A(n8529), .B(n8929), .ZN(n8535) );
  AOI22_X1 U10160 ( .A1(n8657), .A2(n8624), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8531) );
  NAND2_X1 U10161 ( .A1(n8645), .A2(n8922), .ZN(n8530) );
  OAI211_X1 U10162 ( .C1(n8919), .C2(n8627), .A(n8531), .B(n8530), .ZN(n8532)
         );
  AOI21_X1 U10163 ( .B1(n8533), .B2(n8629), .A(n8532), .ZN(n8534) );
  OAI21_X1 U10164 ( .B1(n8535), .B2(n8632), .A(n8534), .ZN(P2_U3156) );
  XNOR2_X1 U10165 ( .A(n8536), .B(n8977), .ZN(n8537) );
  XNOR2_X1 U10166 ( .A(n8538), .B(n8537), .ZN(n8543) );
  NAND2_X1 U10167 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U10168 ( .A1(n8624), .A2(n8660), .ZN(n8539) );
  OAI211_X1 U10169 ( .C1(n8627), .C2(n8964), .A(n8836), .B(n8539), .ZN(n8540)
         );
  AOI21_X1 U10170 ( .B1(n8645), .B2(n8968), .A(n8540), .ZN(n8542) );
  NAND2_X1 U10171 ( .A1(n8967), .A2(n8629), .ZN(n8541) );
  OAI211_X1 U10172 ( .C1(n8543), .C2(n8632), .A(n8542), .B(n8541), .ZN(
        P2_U3159) );
  XOR2_X1 U10173 ( .A(n8546), .B(n8868), .Z(n8547) );
  XNOR2_X1 U10174 ( .A(n8548), .B(n8547), .ZN(n8554) );
  NAND2_X1 U10175 ( .A1(n8650), .A2(n8639), .ZN(n8550) );
  AOI22_X1 U10176 ( .A1(n8870), .A2(n8645), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8549) );
  OAI211_X1 U10177 ( .C1(n8887), .C2(n8641), .A(n8550), .B(n8549), .ZN(n8551)
         );
  AOI21_X1 U10178 ( .B1(n8552), .B2(n8629), .A(n8551), .ZN(n8553) );
  OAI21_X1 U10179 ( .B1(n8554), .B2(n8632), .A(n8553), .ZN(P2_U3160) );
  XOR2_X1 U10180 ( .A(n8556), .B(n8555), .Z(n8562) );
  NAND2_X1 U10181 ( .A1(n8645), .A2(n8942), .ZN(n8558) );
  AOI22_X1 U10182 ( .A1(n8657), .A2(n8639), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8557) );
  OAI211_X1 U10183 ( .C1(n8964), .C2(n8641), .A(n8558), .B(n8557), .ZN(n8559)
         );
  AOI21_X1 U10184 ( .B1(n8560), .B2(n8629), .A(n8559), .ZN(n8561) );
  OAI21_X1 U10185 ( .B1(n8562), .B2(n8632), .A(n8561), .ZN(P2_U3163) );
  XOR2_X1 U10186 ( .A(n8564), .B(n8563), .Z(n8569) );
  AOI22_X1 U10187 ( .A1(n8655), .A2(n8624), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8566) );
  NAND2_X1 U10188 ( .A1(n8899), .A2(n8645), .ZN(n8565) );
  OAI211_X1 U10189 ( .C1(n8897), .C2(n8627), .A(n8566), .B(n8565), .ZN(n8567)
         );
  AOI21_X1 U10190 ( .B1(n9043), .B2(n8629), .A(n8567), .ZN(n8568) );
  OAI21_X1 U10191 ( .B1(n8569), .B2(n8632), .A(n8568), .ZN(P2_U3165) );
  INV_X1 U10192 ( .A(n9444), .ZN(n8579) );
  INV_X1 U10193 ( .A(n8583), .ZN(n8573) );
  AOI21_X1 U10194 ( .B1(n8636), .B2(n8571), .A(n8570), .ZN(n8572) );
  OAI21_X1 U10195 ( .B1(n8573), .B2(n8572), .A(n8635), .ZN(n8578) );
  NAND2_X1 U10196 ( .A1(n8639), .A2(n9015), .ZN(n8574) );
  NAND2_X1 U10197 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8760) );
  OAI211_X1 U10198 ( .C1(n8575), .C2(n8641), .A(n8574), .B(n8760), .ZN(n8576)
         );
  AOI21_X1 U10199 ( .B1(n8645), .B2(n9009), .A(n8576), .ZN(n8577) );
  OAI211_X1 U10200 ( .C1(n8579), .C2(n8648), .A(n8578), .B(n8577), .ZN(
        P2_U3166) );
  AND3_X1 U10201 ( .A1(n8583), .A2(n8582), .A3(n8581), .ZN(n8584) );
  OAI21_X1 U10202 ( .B1(n8615), .B2(n8584), .A(n8635), .ZN(n8588) );
  NAND2_X1 U10203 ( .A1(n8639), .A2(n8660), .ZN(n8585) );
  NAND2_X1 U10204 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8779) );
  OAI211_X1 U10205 ( .C1(n8992), .C2(n8641), .A(n8585), .B(n8779), .ZN(n8586)
         );
  AOI21_X1 U10206 ( .B1(n8645), .B2(n8998), .A(n8586), .ZN(n8587) );
  OAI211_X1 U10207 ( .C1(n9515), .C2(n8648), .A(n8588), .B(n8587), .ZN(
        P2_U3168) );
  XOR2_X1 U10208 ( .A(n8590), .B(n8589), .Z(n8596) );
  AOI22_X1 U10209 ( .A1(n8656), .A2(n8624), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8592) );
  NAND2_X1 U10210 ( .A1(n8645), .A2(n8910), .ZN(n8591) );
  OAI211_X1 U10211 ( .C1(n8908), .C2(n8627), .A(n8592), .B(n8591), .ZN(n8593)
         );
  AOI21_X1 U10212 ( .B1(n8594), .B2(n8629), .A(n8593), .ZN(n8595) );
  OAI21_X1 U10213 ( .B1(n8596), .B2(n8632), .A(n8595), .ZN(P2_U3169) );
  XOR2_X1 U10214 ( .A(n8598), .B(n8597), .Z(n8603) );
  NAND2_X1 U10215 ( .A1(n8645), .A2(n8954), .ZN(n8600) );
  AOI22_X1 U10216 ( .A1(n8658), .A2(n8639), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8599) );
  OAI211_X1 U10217 ( .C1(n8951), .C2(n8641), .A(n8600), .B(n8599), .ZN(n8601)
         );
  AOI21_X1 U10218 ( .B1(n9062), .B2(n8629), .A(n8601), .ZN(n8602) );
  OAI21_X1 U10219 ( .B1(n8603), .B2(n8632), .A(n8602), .ZN(P2_U3173) );
  OAI211_X1 U10220 ( .C1(n8607), .C2(n8606), .A(n8605), .B(n8635), .ZN(n8611)
         );
  AOI22_X1 U10221 ( .A1(n8658), .A2(n8624), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8608) );
  OAI21_X1 U10222 ( .B1(n8929), .B2(n8627), .A(n8608), .ZN(n8609) );
  AOI21_X1 U10223 ( .B1(n8932), .B2(n8645), .A(n8609), .ZN(n8610) );
  OAI211_X1 U10224 ( .C1(n9497), .C2(n8648), .A(n8611), .B(n8610), .ZN(
        P2_U3175) );
  INV_X1 U10225 ( .A(n8612), .ZN(n8617) );
  NOR3_X1 U10226 ( .A1(n8615), .A2(n8614), .A3(n8613), .ZN(n8616) );
  OAI21_X1 U10227 ( .B1(n8617), .B2(n8616), .A(n8635), .ZN(n8621) );
  NAND2_X1 U10228 ( .A1(n8639), .A2(n8977), .ZN(n8618) );
  NAND2_X1 U10229 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8819) );
  OAI211_X1 U10230 ( .C1(n8975), .C2(n8641), .A(n8618), .B(n8819), .ZN(n8619)
         );
  AOI21_X1 U10231 ( .B1(n8645), .B2(n8983), .A(n8619), .ZN(n8620) );
  OAI211_X1 U10232 ( .C1(n9071), .C2(n8648), .A(n8621), .B(n8620), .ZN(
        P2_U3178) );
  XOR2_X1 U10233 ( .A(n8623), .B(n8622), .Z(n8633) );
  AOI22_X1 U10234 ( .A1(n8654), .A2(n8624), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8626) );
  NAND2_X1 U10235 ( .A1(n8890), .A2(n8645), .ZN(n8625) );
  OAI211_X1 U10236 ( .C1(n8887), .C2(n8627), .A(n8626), .B(n8625), .ZN(n8628)
         );
  AOI21_X1 U10237 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8631) );
  OAI21_X1 U10238 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(P2_U3180) );
  INV_X1 U10239 ( .A(n8634), .ZN(n9455) );
  OAI211_X1 U10240 ( .C1(n8638), .C2(n8637), .A(n8636), .B(n8635), .ZN(n8647)
         );
  NAND2_X1 U10241 ( .A1(n8639), .A2(n8661), .ZN(n8640) );
  NAND2_X1 U10242 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8736) );
  OAI211_X1 U10243 ( .C1(n8642), .C2(n8641), .A(n8640), .B(n8736), .ZN(n8643)
         );
  AOI21_X1 U10244 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8646) );
  OAI211_X1 U10245 ( .C1(n9455), .C2(n8648), .A(n8647), .B(n8646), .ZN(
        P2_U3181) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8649), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10247 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8650), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10248 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8651), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10249 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8652), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10250 ( .A(n8653), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8676), .Z(
        P2_U3517) );
  MUX2_X1 U10251 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8654), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10252 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8655), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10253 ( .A(n8656), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8676), .Z(
        P2_U3514) );
  MUX2_X1 U10254 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8657), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10255 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8658), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10256 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8659), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10257 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8977), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10258 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8660), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10259 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9015), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10260 ( .A(n8661), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8676), .Z(
        P2_U3507) );
  MUX2_X1 U10261 ( .A(n9013), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8676), .Z(
        P2_U3506) );
  MUX2_X1 U10262 ( .A(n8662), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8676), .Z(
        P2_U3505) );
  MUX2_X1 U10263 ( .A(n8663), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8676), .Z(
        P2_U3504) );
  MUX2_X1 U10264 ( .A(n8664), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8676), .Z(
        P2_U3503) );
  MUX2_X1 U10265 ( .A(n8665), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8676), .Z(
        P2_U3502) );
  MUX2_X1 U10266 ( .A(n8666), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8676), .Z(
        P2_U3501) );
  MUX2_X1 U10267 ( .A(n8667), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8676), .Z(
        P2_U3500) );
  MUX2_X1 U10268 ( .A(n8668), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8676), .Z(
        P2_U3499) );
  MUX2_X1 U10269 ( .A(n8669), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8676), .Z(
        P2_U3498) );
  MUX2_X1 U10270 ( .A(n8670), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8676), .Z(
        P2_U3497) );
  MUX2_X1 U10271 ( .A(n8671), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8676), .Z(
        P2_U3496) );
  MUX2_X1 U10272 ( .A(n8672), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8676), .Z(
        P2_U3495) );
  MUX2_X1 U10273 ( .A(n8673), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8676), .Z(
        P2_U3494) );
  MUX2_X1 U10274 ( .A(n4669), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8676), .Z(
        P2_U3493) );
  MUX2_X1 U10275 ( .A(n6280), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8676), .Z(
        P2_U3492) );
  MUX2_X1 U10276 ( .A(n8677), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8676), .Z(
        P2_U3491) );
  OAI211_X1 U10277 ( .C1(n8680), .C2(n8679), .A(n8678), .B(n10652), .ZN(n8696)
         );
  INV_X1 U10278 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n8681) );
  OR2_X1 U10279 ( .A1(n10657), .A2(n8681), .ZN(n8683) );
  OAI211_X1 U10280 ( .C1(n8837), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8685)
         );
  INV_X1 U10281 ( .A(n8685), .ZN(n8695) );
  NAND2_X1 U10282 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U10283 ( .A1(n4745), .A2(n8689), .ZN(n8693) );
  OAI21_X1 U10284 ( .B1(n8691), .B2(P2_REG2_REG_5__SCAN_IN), .A(n8690), .ZN(
        n8692) );
  AOI22_X1 U10285 ( .A1(n10648), .A2(n8693), .B1(n10664), .B2(n8692), .ZN(
        n8694) );
  NAND3_X1 U10286 ( .A1(n8696), .A2(n8695), .A3(n8694), .ZN(P2_U3187) );
  NOR2_X1 U10287 ( .A1(n8713), .A2(n8697), .ZN(n8699) );
  MUX2_X1 U10288 ( .A(n8702), .B(P2_REG2_REG_14__SCAN_IN), .S(n8732), .Z(n8700) );
  AOI21_X1 U10289 ( .B1(n4639), .B2(n8700), .A(n8731), .ZN(n8722) );
  MUX2_X1 U10290 ( .A(n8702), .B(n8701), .S(n8798), .Z(n8725) );
  XNOR2_X1 U10291 ( .A(n8732), .B(n8725), .ZN(n8708) );
  INV_X1 U10292 ( .A(n8703), .ZN(n8704) );
  NAND2_X1 U10293 ( .A1(n8713), .A2(n8704), .ZN(n8706) );
  NAND2_X1 U10294 ( .A1(n8706), .A2(n8705), .ZN(n8707) );
  NAND2_X1 U10295 ( .A1(n8708), .A2(n8707), .ZN(n8727) );
  OAI21_X1 U10296 ( .B1(n8708), .B2(n8707), .A(n8727), .ZN(n8709) );
  NAND2_X1 U10297 ( .A1(n10652), .A2(n8709), .ZN(n8711) );
  OAI211_X1 U10298 ( .C1(n8837), .C2(n8732), .A(n8711), .B(n8710), .ZN(n8720)
         );
  NOR2_X1 U10299 ( .A1(n8713), .A2(n8712), .ZN(n8715) );
  NAND2_X1 U10300 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8732), .ZN(n8716) );
  OAI21_X1 U10301 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8732), .A(n8716), .ZN(
        n8717) );
  AOI21_X1 U10302 ( .B1(n4643), .B2(n8717), .A(n8723), .ZN(n8718) );
  NOR2_X1 U10303 ( .A1(n8718), .A2(n8806), .ZN(n8719) );
  AOI211_X1 U10304 ( .C1(n8839), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8720), .B(
        n8719), .ZN(n8721) );
  OAI21_X1 U10305 ( .B1(n8722), .B2(n8841), .A(n8721), .ZN(P2_U3196) );
  INV_X1 U10306 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9400) );
  AOI21_X1 U10307 ( .B1(n9400), .B2(n8724), .A(n8749), .ZN(n8742) );
  MUX2_X1 U10308 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8798), .Z(n8754) );
  XNOR2_X1 U10309 ( .A(n8748), .B(n8754), .ZN(n8730) );
  INV_X1 U10310 ( .A(n8732), .ZN(n8726) );
  NAND2_X1 U10311 ( .A1(n8726), .A2(n8725), .ZN(n8728) );
  NAND2_X1 U10312 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND2_X1 U10313 ( .A1(n8730), .A2(n8729), .ZN(n8755) );
  OAI21_X1 U10314 ( .B1(n8730), .B2(n8729), .A(n8755), .ZN(n8740) );
  AOI21_X1 U10315 ( .B1(n8733), .B2(n9270), .A(n8744), .ZN(n8734) );
  NOR2_X1 U10316 ( .A1(n8734), .A2(n8841), .ZN(n8739) );
  OR2_X1 U10317 ( .A1(n10657), .A2(n8735), .ZN(n8737) );
  OAI211_X1 U10318 ( .C1(n8837), .C2(n4659), .A(n8737), .B(n8736), .ZN(n8738)
         );
  AOI211_X1 U10319 ( .C1(n10652), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  OAI21_X1 U10320 ( .B1(n8742), .B2(n8806), .A(n8741), .ZN(P2_U3197) );
  NAND2_X1 U10321 ( .A1(n8772), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8767) );
  OAI21_X1 U10322 ( .B1(n8772), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8767), .ZN(
        n8746) );
  AOI21_X1 U10323 ( .B1(n4642), .B2(n8746), .A(n8769), .ZN(n8766) );
  NAND2_X1 U10324 ( .A1(n8772), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8781) );
  OAI21_X1 U10325 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8772), .A(n8781), .ZN(
        n8750) );
  NAND2_X1 U10326 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  AOI21_X1 U10327 ( .B1(n8782), .B2(n8752), .A(n8806), .ZN(n8764) );
  INV_X1 U10328 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8753) );
  NOR2_X1 U10329 ( .A1(n10657), .A2(n8753), .ZN(n8763) );
  MUX2_X1 U10330 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8798), .Z(n8773) );
  XOR2_X1 U10331 ( .A(n8773), .B(n8772), .Z(n8758) );
  OR2_X1 U10332 ( .A1(n8754), .A2(n4659), .ZN(n8756) );
  NAND2_X1 U10333 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U10334 ( .A1(n8758), .A2(n8757), .ZN(n8774) );
  OAI21_X1 U10335 ( .B1(n8758), .B2(n8757), .A(n8774), .ZN(n8759) );
  NAND2_X1 U10336 ( .A1(n8759), .A2(n10652), .ZN(n8761) );
  OAI211_X1 U10337 ( .C1(n8837), .C2(n8772), .A(n8761), .B(n8760), .ZN(n8762)
         );
  NOR3_X1 U10338 ( .A1(n8764), .A2(n8763), .A3(n8762), .ZN(n8765) );
  OAI21_X1 U10339 ( .B1(n8766), .B2(n8841), .A(n8765), .ZN(P2_U3198) );
  INV_X1 U10340 ( .A(n8767), .ZN(n8768) );
  NOR2_X1 U10341 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  AOI21_X1 U10342 ( .B1(n6495), .B2(n8771), .A(n8791), .ZN(n8790) );
  MUX2_X1 U10343 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8798), .Z(n8793) );
  XNOR2_X1 U10344 ( .A(n8797), .B(n8793), .ZN(n8777) );
  OR2_X1 U10345 ( .A1(n8773), .A2(n8772), .ZN(n8775) );
  NAND2_X1 U10346 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  NAND2_X1 U10347 ( .A1(n8777), .A2(n8776), .ZN(n8794) );
  OAI21_X1 U10348 ( .B1(n8777), .B2(n8776), .A(n8794), .ZN(n8778) );
  NAND2_X1 U10349 ( .A1(n10652), .A2(n8778), .ZN(n8780) );
  OAI211_X1 U10350 ( .C1(n8837), .C2(n8783), .A(n8780), .B(n8779), .ZN(n8788)
         );
  NAND2_X1 U10351 ( .A1(n8782), .A2(n8781), .ZN(n8784) );
  AOI21_X1 U10352 ( .B1(n8785), .B2(n9440), .A(n8804), .ZN(n8786) );
  NOR2_X1 U10353 ( .A1(n8786), .A2(n8806), .ZN(n8787) );
  AOI211_X1 U10354 ( .C1(n8839), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8788), .B(
        n8787), .ZN(n8789) );
  OAI21_X1 U10355 ( .B1(n8790), .B2(n8841), .A(n8789), .ZN(P2_U3199) );
  OR2_X1 U10356 ( .A1(n8841), .A2(n8817), .ZN(n8811) );
  INV_X1 U10357 ( .A(n8793), .ZN(n8796) );
  INV_X1 U10358 ( .A(n8794), .ZN(n8795) );
  AOI21_X1 U10359 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8799) );
  MUX2_X1 U10360 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8798), .Z(n8800) );
  AND2_X1 U10361 ( .A1(n8799), .A2(n8800), .ZN(n8824) );
  INV_X1 U10362 ( .A(n8799), .ZN(n8802) );
  INV_X1 U10363 ( .A(n8800), .ZN(n8801) );
  NAND2_X1 U10364 ( .A1(n8802), .A2(n8801), .ZN(n8823) );
  INV_X1 U10365 ( .A(n8823), .ZN(n8803) );
  NOR2_X1 U10366 ( .A1(n8824), .A2(n8803), .ZN(n8809) );
  AOI21_X1 U10367 ( .B1(n8809), .B2(P2_U3893), .A(n10650), .ZN(n8807) );
  INV_X1 U10368 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8814) );
  INV_X1 U10369 ( .A(n8809), .ZN(n8810) );
  NAND2_X1 U10370 ( .A1(n10652), .A2(n8810), .ZN(n8812) );
  INV_X1 U10371 ( .A(n8833), .ZN(n8828) );
  MUX2_X1 U10372 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8814), .S(n8833), .Z(n8816) );
  MUX2_X1 U10373 ( .A(n8832), .B(P2_REG2_REG_18__SCAN_IN), .S(n8833), .Z(n8818) );
  NAND2_X1 U10374 ( .A1(n8818), .A2(n8817), .ZN(n8831) );
  OAI21_X1 U10375 ( .B1(n8831), .B2(n8841), .A(n8819), .ZN(n8820) );
  AOI21_X1 U10376 ( .B1(n10648), .B2(n8827), .A(n8820), .ZN(n8821) );
  XNOR2_X1 U10377 ( .A(n6622), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8829) );
  XNOR2_X1 U10378 ( .A(n6622), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8834) );
  MUX2_X1 U10379 ( .A(n8829), .B(n8834), .S(n8822), .Z(n8826) );
  OAI21_X1 U10380 ( .B1(n8824), .B2(n8828), .A(n8823), .ZN(n8825) );
  XNOR2_X1 U10381 ( .A(n8826), .B(n8825), .ZN(n8847) );
  XNOR2_X1 U10382 ( .A(n8830), .B(n8829), .ZN(n8844) );
  OAI21_X1 U10383 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8835) );
  XNOR2_X1 U10384 ( .A(n8835), .B(n8834), .ZN(n8842) );
  OAI21_X1 U10385 ( .B1(n8837), .B2(n6622), .A(n8836), .ZN(n8838) );
  AOI21_X1 U10386 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n8839), .A(n8838), .ZN(
        n8840) );
  OAI21_X1 U10387 ( .B1(n8842), .B2(n8841), .A(n8840), .ZN(n8843) );
  AOI21_X1 U10388 ( .B1(n8844), .B2(n10648), .A(n8843), .ZN(n8845) );
  OAI21_X1 U10389 ( .B1(n8847), .B2(n8846), .A(n8845), .ZN(P2_U3201) );
  NAND2_X1 U10390 ( .A1(n8850), .A2(n8999), .ZN(n8855) );
  OAI21_X1 U10391 ( .B1(n9000), .B2(n9457), .A(n8855), .ZN(n8852) );
  AOI21_X1 U10392 ( .B1(n9022), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8852), .ZN(
        n8851) );
  OAI21_X1 U10393 ( .B1(n9459), .B2(n9002), .A(n8851), .ZN(P2_U3202) );
  AOI21_X1 U10394 ( .B1(n9022), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8852), .ZN(
        n8853) );
  OAI21_X1 U10395 ( .B1(n9462), .B2(n9002), .A(n8853), .ZN(P2_U3203) );
  INV_X1 U10396 ( .A(n8854), .ZN(n8861) );
  NAND2_X1 U10397 ( .A1(n9468), .A2(n9023), .ZN(n8856) );
  OAI211_X1 U10398 ( .C1(n9020), .C2(n8857), .A(n8856), .B(n8855), .ZN(n8858)
         );
  AOI21_X1 U10399 ( .B1(n8859), .B2(n9004), .A(n8858), .ZN(n8860) );
  OAI21_X1 U10400 ( .B1(n8861), .B2(n9022), .A(n8860), .ZN(P2_U3204) );
  XNOR2_X1 U10401 ( .A(n8862), .B(n8868), .ZN(n8867) );
  INV_X1 U10402 ( .A(n9034), .ZN(n8874) );
  XNOR2_X1 U10403 ( .A(n8869), .B(n8868), .ZN(n9033) );
  AOI22_X1 U10404 ( .A1(n8870), .A2(n8999), .B1(n9000), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8871) );
  OAI21_X1 U10405 ( .B1(n9474), .B2(n9002), .A(n8871), .ZN(n8872) );
  AOI21_X1 U10406 ( .B1(n9033), .B2(n9004), .A(n8872), .ZN(n8873) );
  OAI21_X1 U10407 ( .B1(n8874), .B2(n9022), .A(n8873), .ZN(P2_U3205) );
  INV_X1 U10408 ( .A(n9037), .ZN(n8883) );
  XNOR2_X1 U10409 ( .A(n8878), .B(n8877), .ZN(n9038) );
  AOI22_X1 U10410 ( .A1(n8879), .A2(n8999), .B1(n9000), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8880) );
  OAI21_X1 U10411 ( .B1(n9477), .B2(n9002), .A(n8880), .ZN(n8881) );
  AOI21_X1 U10412 ( .B1(n9038), .B2(n9004), .A(n8881), .ZN(n8882) );
  OAI21_X1 U10413 ( .B1(n8883), .B2(n9022), .A(n8882), .ZN(P2_U3206) );
  XNOR2_X1 U10414 ( .A(n8885), .B(n8884), .ZN(n8886) );
  INV_X1 U10415 ( .A(n9039), .ZN(n8894) );
  XNOR2_X1 U10416 ( .A(n8889), .B(n8888), .ZN(n9040) );
  AOI22_X1 U10417 ( .A1(n8890), .A2(n8999), .B1(n9000), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8891) );
  OAI21_X1 U10418 ( .B1(n9481), .B2(n9002), .A(n8891), .ZN(n8892) );
  AOI21_X1 U10419 ( .B1(n9040), .B2(n9004), .A(n8892), .ZN(n8893) );
  OAI21_X1 U10420 ( .B1(n8894), .B2(n9022), .A(n8893), .ZN(P2_U3207) );
  XOR2_X1 U10421 ( .A(n8900), .B(n8895), .Z(n8896) );
  AOI21_X1 U10422 ( .B1(n8898), .B2(n9043), .A(n9044), .ZN(n8904) );
  AOI22_X1 U10423 ( .A1(n8899), .A2(n8999), .B1(n9022), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8903) );
  XNOR2_X1 U10424 ( .A(n8901), .B(n8900), .ZN(n9045) );
  NAND2_X1 U10425 ( .A1(n9045), .A2(n9004), .ZN(n8902) );
  OAI211_X1 U10426 ( .C1(n8904), .C2(n9022), .A(n8903), .B(n8902), .ZN(
        P2_U3208) );
  NOR2_X1 U10427 ( .A1(n9489), .A2(n8905), .ZN(n8909) );
  XNOR2_X1 U10428 ( .A(n8906), .B(n8914), .ZN(n8907) );
  OAI222_X1 U10429 ( .A1(n8953), .A2(n8908), .B1(n8929), .B2(n8993), .C1(n8907), .C2(n8990), .ZN(n9048) );
  AOI211_X1 U10430 ( .C1(n8999), .C2(n8910), .A(n8909), .B(n9048), .ZN(n8916)
         );
  NAND2_X1 U10431 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  XOR2_X1 U10432 ( .A(n8914), .B(n8913), .Z(n9049) );
  AOI22_X1 U10433 ( .A1(n9049), .A2(n9004), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9022), .ZN(n8915) );
  OAI21_X1 U10434 ( .B1(n8916), .B2(n9022), .A(n8915), .ZN(P2_U3209) );
  XNOR2_X1 U10435 ( .A(n8917), .B(n8920), .ZN(n8918) );
  OAI222_X1 U10436 ( .A1(n8953), .A2(n8919), .B1(n8993), .B2(n8939), .C1(n8990), .C2(n8918), .ZN(n9052) );
  INV_X1 U10437 ( .A(n9052), .ZN(n8926) );
  XNOR2_X1 U10438 ( .A(n8921), .B(n8920), .ZN(n9053) );
  AOI22_X1 U10439 ( .A1(n9000), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8922), .B2(
        n8999), .ZN(n8923) );
  OAI21_X1 U10440 ( .B1(n9493), .B2(n9002), .A(n8923), .ZN(n8924) );
  AOI21_X1 U10441 ( .B1(n9053), .B2(n9004), .A(n8924), .ZN(n8925) );
  OAI21_X1 U10442 ( .B1(n8926), .B2(n9022), .A(n8925), .ZN(P2_U3210) );
  XOR2_X1 U10443 ( .A(n8931), .B(n8927), .Z(n8928) );
  OAI222_X1 U10444 ( .A1(n8953), .A2(n8929), .B1(n8993), .B2(n8952), .C1(n8990), .C2(n8928), .ZN(n9056) );
  INV_X1 U10445 ( .A(n9056), .ZN(n8936) );
  XOR2_X1 U10446 ( .A(n8931), .B(n8930), .Z(n9057) );
  AOI22_X1 U10447 ( .A1(n9000), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8999), .B2(
        n8932), .ZN(n8933) );
  OAI21_X1 U10448 ( .B1(n9497), .B2(n9002), .A(n8933), .ZN(n8934) );
  AOI21_X1 U10449 ( .B1(n9057), .B2(n9004), .A(n8934), .ZN(n8935) );
  OAI21_X1 U10450 ( .B1(n8936), .B2(n9022), .A(n8935), .ZN(P2_U3211) );
  XNOR2_X1 U10451 ( .A(n8937), .B(n8940), .ZN(n8938) );
  OAI222_X1 U10452 ( .A1(n8953), .A2(n8939), .B1(n8993), .B2(n8964), .C1(n8990), .C2(n8938), .ZN(n9059) );
  INV_X1 U10453 ( .A(n9059), .ZN(n8946) );
  XNOR2_X1 U10454 ( .A(n8941), .B(n8940), .ZN(n9060) );
  AOI22_X1 U10455 ( .A1(n9000), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8999), .B2(
        n8942), .ZN(n8943) );
  OAI21_X1 U10456 ( .B1(n9501), .B2(n9002), .A(n8943), .ZN(n8944) );
  AOI21_X1 U10457 ( .B1(n9060), .B2(n9004), .A(n8944), .ZN(n8945) );
  OAI21_X1 U10458 ( .B1(n8946), .B2(n9022), .A(n8945), .ZN(P2_U3212) );
  OAI21_X1 U10459 ( .B1(n8948), .B2(n8955), .A(n8947), .ZN(n8949) );
  INV_X1 U10460 ( .A(n8949), .ZN(n8950) );
  OAI222_X1 U10461 ( .A1(n8953), .A2(n8952), .B1(n8993), .B2(n8951), .C1(n8990), .C2(n8950), .ZN(n9063) );
  AOI21_X1 U10462 ( .B1(n8999), .B2(n8954), .A(n9063), .ZN(n8959) );
  AOI22_X1 U10463 ( .A1(n9062), .A2(n9023), .B1(P2_REG2_REG_20__SCAN_IN), .B2(
        n9022), .ZN(n8958) );
  XNOR2_X1 U10464 ( .A(n8956), .B(n8955), .ZN(n9064) );
  NAND2_X1 U10465 ( .A1(n9064), .A2(n9004), .ZN(n8957) );
  OAI211_X1 U10466 ( .C1(n8959), .C2(n9000), .A(n8958), .B(n8957), .ZN(
        P2_U3213) );
  XNOR2_X1 U10467 ( .A(n8960), .B(n8963), .ZN(n9067) );
  INV_X1 U10468 ( .A(n9067), .ZN(n8972) );
  AOI211_X1 U10469 ( .C1(n8963), .C2(n8962), .A(n8990), .B(n8961), .ZN(n8966)
         );
  OAI22_X1 U10470 ( .A1(n8964), .A2(n8953), .B1(n8994), .B2(n8993), .ZN(n8965)
         );
  OR2_X1 U10471 ( .A1(n8966), .A2(n8965), .ZN(n9066) );
  INV_X1 U10472 ( .A(n8967), .ZN(n9509) );
  AOI22_X1 U10473 ( .A1(n9000), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8999), .B2(
        n8968), .ZN(n8969) );
  OAI21_X1 U10474 ( .B1(n9509), .B2(n9002), .A(n8969), .ZN(n8970) );
  AOI21_X1 U10475 ( .B1(n9066), .B2(n9020), .A(n8970), .ZN(n8971) );
  OAI21_X1 U10476 ( .B1(n8972), .B2(n9026), .A(n8971), .ZN(P2_U3214) );
  XNOR2_X1 U10477 ( .A(n8973), .B(n8980), .ZN(n8974) );
  NAND2_X1 U10478 ( .A1(n8974), .A2(n9017), .ZN(n8979) );
  NOR2_X1 U10479 ( .A1(n8975), .A2(n8993), .ZN(n8976) );
  AOI21_X1 U10480 ( .B1(n8977), .B2(n9014), .A(n8976), .ZN(n8978) );
  NAND2_X1 U10481 ( .A1(n8979), .A2(n8978), .ZN(n9075) );
  INV_X1 U10482 ( .A(n9073), .ZN(n8982) );
  NAND2_X1 U10483 ( .A1(n8981), .A2(n8980), .ZN(n9070) );
  NAND3_X1 U10484 ( .A1(n8982), .A2(n9004), .A3(n9070), .ZN(n8985) );
  AOI22_X1 U10485 ( .A1(n9000), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8999), .B2(
        n8983), .ZN(n8984) );
  OAI211_X1 U10486 ( .C1(n9071), .C2(n9002), .A(n8985), .B(n8984), .ZN(n8986)
         );
  AOI21_X1 U10487 ( .B1(n9075), .B2(n9020), .A(n8986), .ZN(n8987) );
  INV_X1 U10488 ( .A(n8987), .ZN(P2_U3215) );
  XNOR2_X1 U10489 ( .A(n8989), .B(n8988), .ZN(n8991) );
  OAI222_X1 U10490 ( .A1(n8953), .A2(n8994), .B1(n8993), .B2(n8992), .C1(n8991), .C2(n8990), .ZN(n9438) );
  INV_X1 U10491 ( .A(n9438), .ZN(n9006) );
  OAI21_X1 U10492 ( .B1(n5082), .B2(n8997), .A(n8996), .ZN(n9439) );
  AOI22_X1 U10493 ( .A1(n9000), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8999), .B2(
        n8998), .ZN(n9001) );
  OAI21_X1 U10494 ( .B1(n9515), .B2(n9002), .A(n9001), .ZN(n9003) );
  AOI21_X1 U10495 ( .B1(n9439), .B2(n9004), .A(n9003), .ZN(n9005) );
  OAI21_X1 U10496 ( .B1(n9006), .B2(n9022), .A(n9005), .ZN(P2_U3216) );
  OAI21_X1 U10497 ( .B1(n9008), .B2(n9010), .A(n9007), .ZN(n9447) );
  INV_X1 U10498 ( .A(n9009), .ZN(n9019) );
  XNOR2_X1 U10499 ( .A(n9011), .B(n9010), .ZN(n9016) );
  AOI222_X1 U10500 ( .A1(n9017), .A2(n9016), .B1(n9015), .B2(n9014), .C1(n9013), .C2(n9012), .ZN(n9446) );
  OAI21_X1 U10501 ( .B1(n9019), .B2(n9018), .A(n9446), .ZN(n9021) );
  NAND2_X1 U10502 ( .A1(n9021), .A2(n9020), .ZN(n9025) );
  AOI22_X1 U10503 ( .A1(n9444), .A2(n9023), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n9022), .ZN(n9024) );
  OAI211_X1 U10504 ( .C1(n9447), .C2(n9026), .A(n9025), .B(n9024), .ZN(
        P2_U3217) );
  NOR2_X1 U10505 ( .A1(n9457), .A2(n4671), .ZN(n9030) );
  AOI21_X1 U10506 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n4671), .A(n9030), .ZN(
        n9027) );
  OAI21_X1 U10507 ( .B1(n9459), .B2(n9442), .A(n9027), .ZN(P2_U3490) );
  NAND2_X1 U10508 ( .A1(n9029), .A2(n9028), .ZN(n9032) );
  INV_X1 U10509 ( .A(n9030), .ZN(n9031) );
  OAI211_X1 U10510 ( .C1(n9456), .C2(n6587), .A(n9032), .B(n9031), .ZN(
        P2_U3489) );
  INV_X1 U10511 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10512 ( .A(n9035), .B(n9471), .S(n9456), .Z(n9036) );
  OAI21_X1 U10513 ( .B1(n9474), .B2(n9442), .A(n9036), .ZN(P2_U3487) );
  INV_X1 U10514 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10515 ( .A(n9041), .B(n9478), .S(n9456), .Z(n9042) );
  OAI21_X1 U10516 ( .B1(n9481), .B2(n9442), .A(n9042), .ZN(P2_U3485) );
  INV_X1 U10517 ( .A(n9043), .ZN(n9485) );
  INV_X1 U10518 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9046) );
  MUX2_X1 U10519 ( .A(n9046), .B(n9482), .S(n9456), .Z(n9047) );
  OAI21_X1 U10520 ( .B1(n9485), .B2(n9442), .A(n9047), .ZN(P2_U3484) );
  INV_X1 U10521 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9050) );
  AOI21_X1 U10522 ( .B1(n9049), .B2(n9449), .A(n9048), .ZN(n9486) );
  MUX2_X1 U10523 ( .A(n9050), .B(n9486), .S(n9456), .Z(n9051) );
  OAI21_X1 U10524 ( .B1(n9489), .B2(n9442), .A(n9051), .ZN(P2_U3483) );
  INV_X1 U10525 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9054) );
  AOI21_X1 U10526 ( .B1(n9053), .B2(n9449), .A(n9052), .ZN(n9490) );
  MUX2_X1 U10527 ( .A(n9054), .B(n9490), .S(n9456), .Z(n9055) );
  OAI21_X1 U10528 ( .B1(n9493), .B2(n9442), .A(n9055), .ZN(P2_U3482) );
  AOI21_X1 U10529 ( .B1(n9449), .B2(n9057), .A(n9056), .ZN(n9494) );
  MUX2_X1 U10530 ( .A(n9409), .B(n9494), .S(n9456), .Z(n9058) );
  OAI21_X1 U10531 ( .B1(n9497), .B2(n9442), .A(n9058), .ZN(P2_U3481) );
  AOI21_X1 U10532 ( .B1(n9060), .B2(n9449), .A(n9059), .ZN(n9498) );
  MUX2_X1 U10533 ( .A(n9279), .B(n9498), .S(n9456), .Z(n9061) );
  OAI21_X1 U10534 ( .B1(n9501), .B2(n9442), .A(n9061), .ZN(P2_U3480) );
  INV_X1 U10535 ( .A(n9062), .ZN(n9505) );
  AOI21_X1 U10536 ( .B1(n9064), .B2(n9449), .A(n9063), .ZN(n9502) );
  MUX2_X1 U10537 ( .A(n9175), .B(n9502), .S(n9456), .Z(n9065) );
  OAI21_X1 U10538 ( .B1(n9505), .B2(n9442), .A(n9065), .ZN(P2_U3479) );
  INV_X1 U10539 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9068) );
  AOI21_X1 U10540 ( .B1(n9449), .B2(n9067), .A(n9066), .ZN(n9506) );
  MUX2_X1 U10541 ( .A(n9068), .B(n9506), .S(n9456), .Z(n9069) );
  OAI21_X1 U10542 ( .B1(n9509), .B2(n9442), .A(n9069), .ZN(P2_U3478) );
  NAND2_X1 U10543 ( .A1(n9070), .A2(n9449), .ZN(n9072) );
  OAI22_X1 U10544 ( .A1(n9073), .A2(n9072), .B1(n9071), .B2(n9454), .ZN(n9074)
         );
  MUX2_X1 U10545 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9510), .S(n9456), .Z(n9437) );
  AOI22_X1 U10546 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput249), .B1(
        P2_REG2_REG_8__SCAN_IN), .B2(keyinput143), .ZN(n9076) );
  OAI221_X1 U10547 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput249), .C1(
        P2_REG2_REG_8__SCAN_IN), .C2(keyinput143), .A(n9076), .ZN(n9083) );
  AOI22_X1 U10548 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput219), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput179), .ZN(n9077) );
  OAI221_X1 U10549 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput219), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput179), .A(n9077), .ZN(n9082) );
  AOI22_X1 U10550 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput145), .B1(
        P2_D_REG_25__SCAN_IN), .B2(keyinput168), .ZN(n9078) );
  OAI221_X1 U10551 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput145), .C1(
        P2_D_REG_25__SCAN_IN), .C2(keyinput168), .A(n9078), .ZN(n9081) );
  AOI22_X1 U10552 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput200), .B1(
        P2_REG0_REG_16__SCAN_IN), .B2(keyinput185), .ZN(n9079) );
  OAI221_X1 U10553 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput200), .C1(
        P2_REG0_REG_16__SCAN_IN), .C2(keyinput185), .A(n9079), .ZN(n9080) );
  NOR4_X1 U10554 ( .A1(n9083), .A2(n9082), .A3(n9081), .A4(n9080), .ZN(n9111)
         );
  AOI22_X1 U10555 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(keyinput195), .B1(
        P2_REG0_REG_7__SCAN_IN), .B2(keyinput189), .ZN(n9084) );
  OAI221_X1 U10556 ( .B1(P1_REG0_REG_24__SCAN_IN), .B2(keyinput195), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput189), .A(n9084), .ZN(n9091) );
  AOI22_X1 U10557 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput253), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput163), .ZN(n9085) );
  OAI221_X1 U10558 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput253), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput163), .A(n9085), .ZN(n9090) );
  AOI22_X1 U10559 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput182), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(keyinput131), .ZN(n9086) );
  OAI221_X1 U10560 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput182), .C1(
        P2_REG2_REG_0__SCAN_IN), .C2(keyinput131), .A(n9086), .ZN(n9089) );
  AOI22_X1 U10561 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(keyinput207), .B1(
        P2_REG0_REG_25__SCAN_IN), .B2(keyinput224), .ZN(n9087) );
  OAI221_X1 U10562 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(keyinput207), .C1(
        P2_REG0_REG_25__SCAN_IN), .C2(keyinput224), .A(n9087), .ZN(n9088) );
  NOR4_X1 U10563 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), .ZN(n9110)
         );
  AOI22_X1 U10564 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput218), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput241), .ZN(n9092) );
  OAI221_X1 U10565 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput218), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput241), .A(n9092), .ZN(n9099) );
  AOI22_X1 U10566 ( .A1(SI_30_), .A2(keyinput188), .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput231), .ZN(n9093) );
  OAI221_X1 U10567 ( .B1(SI_30_), .B2(keyinput188), .C1(
        P1_REG0_REG_21__SCAN_IN), .C2(keyinput231), .A(n9093), .ZN(n9098) );
  AOI22_X1 U10568 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput244), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput222), .ZN(n9094) );
  OAI221_X1 U10569 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput244), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput222), .A(n9094), .ZN(n9097) );
  AOI22_X1 U10570 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput159), .B1(
        P2_IR_REG_31__SCAN_IN), .B2(keyinput215), .ZN(n9095) );
  OAI221_X1 U10571 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput159), .C1(
        P2_IR_REG_31__SCAN_IN), .C2(keyinput215), .A(n9095), .ZN(n9096) );
  NOR4_X1 U10572 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), .ZN(n9109)
         );
  AOI22_X1 U10573 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(keyinput167), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput147), .ZN(n9100) );
  OAI221_X1 U10574 ( .B1(P2_IR_REG_4__SCAN_IN), .B2(keyinput167), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput147), .A(n9100), .ZN(n9107) );
  AOI22_X1 U10575 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput255), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput130), .ZN(n9101) );
  OAI221_X1 U10576 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput255), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput130), .A(n9101), .ZN(n9106) );
  AOI22_X1 U10577 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput171), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput176), .ZN(n9102) );
  OAI221_X1 U10578 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput171), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput176), .A(n9102), .ZN(n9105) );
  AOI22_X1 U10579 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(keyinput197), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput154), .ZN(n9103) );
  OAI221_X1 U10580 ( .B1(P1_REG0_REG_13__SCAN_IN), .B2(keyinput197), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput154), .A(n9103), .ZN(n9104) );
  NOR4_X1 U10581 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9108)
         );
  NAND4_X1 U10582 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n9244)
         );
  AOI22_X1 U10583 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput152), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput155), .ZN(n9112) );
  OAI221_X1 U10584 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput152), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput155), .A(n9112), .ZN(n9119) );
  AOI22_X1 U10585 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput151), .B1(
        P2_REG1_REG_18__SCAN_IN), .B2(keyinput129), .ZN(n9113) );
  OAI221_X1 U10586 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput151), .C1(
        P2_REG1_REG_18__SCAN_IN), .C2(keyinput129), .A(n9113), .ZN(n9118) );
  AOI22_X1 U10587 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput205), .B1(
        P2_REG2_REG_15__SCAN_IN), .B2(keyinput190), .ZN(n9114) );
  OAI221_X1 U10588 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput205), .C1(
        P2_REG2_REG_15__SCAN_IN), .C2(keyinput190), .A(n9114), .ZN(n9117) );
  AOI22_X1 U10589 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput138), .B1(
        P2_REG2_REG_13__SCAN_IN), .B2(keyinput184), .ZN(n9115) );
  OAI221_X1 U10590 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput138), .C1(
        P2_REG2_REG_13__SCAN_IN), .C2(keyinput184), .A(n9115), .ZN(n9116) );
  NOR4_X1 U10591 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(n9148)
         );
  AOI22_X1 U10592 ( .A1(P1_D_REG_9__SCAN_IN), .A2(keyinput194), .B1(
        P2_IR_REG_10__SCAN_IN), .B2(keyinput136), .ZN(n9120) );
  OAI221_X1 U10593 ( .B1(P1_D_REG_9__SCAN_IN), .B2(keyinput194), .C1(
        P2_IR_REG_10__SCAN_IN), .C2(keyinput136), .A(n9120), .ZN(n9127) );
  AOI22_X1 U10594 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(keyinput251), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput234), .ZN(n9121) );
  OAI221_X1 U10595 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(keyinput251), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput234), .A(n9121), .ZN(n9126) );
  AOI22_X1 U10596 ( .A1(SI_8_), .A2(keyinput209), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput237), .ZN(n9122) );
  OAI221_X1 U10597 ( .B1(SI_8_), .B2(keyinput209), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput237), .A(n9122), .ZN(n9125) );
  AOI22_X1 U10598 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput202), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput178), .ZN(n9123) );
  OAI221_X1 U10599 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput202), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput178), .A(n9123), .ZN(n9124) );
  NOR4_X1 U10600 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n9147)
         );
  AOI22_X1 U10601 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(keyinput212), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput146), .ZN(n9128) );
  OAI221_X1 U10602 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(keyinput212), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput146), .A(n9128), .ZN(n9135) );
  AOI22_X1 U10603 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(keyinput248), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput210), .ZN(n9129) );
  OAI221_X1 U10604 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(keyinput248), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput210), .A(n9129), .ZN(n9134) );
  AOI22_X1 U10605 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput225), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput160), .ZN(n9130) );
  OAI221_X1 U10606 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput225), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput160), .A(n9130), .ZN(n9133) );
  AOI22_X1 U10607 ( .A1(SI_4_), .A2(keyinput156), .B1(P2_DATAO_REG_5__SCAN_IN), 
        .B2(keyinput227), .ZN(n9131) );
  OAI221_X1 U10608 ( .B1(SI_4_), .B2(keyinput156), .C1(P2_DATAO_REG_5__SCAN_IN), .C2(keyinput227), .A(n9131), .ZN(n9132) );
  NOR4_X1 U10609 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n9146)
         );
  AOI22_X1 U10610 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput213), .B1(
        SI_16_), .B2(keyinput233), .ZN(n9136) );
  OAI221_X1 U10611 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput213), .C1(
        SI_16_), .C2(keyinput233), .A(n9136), .ZN(n9144) );
  AOI22_X1 U10612 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput186), .B1(
        P2_REG1_REG_21__SCAN_IN), .B2(keyinput238), .ZN(n9137) );
  OAI221_X1 U10613 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput186), .C1(
        P2_REG1_REG_21__SCAN_IN), .C2(keyinput238), .A(n9137), .ZN(n9143) );
  AOI22_X1 U10614 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput230), .B1(
        P1_REG2_REG_21__SCAN_IN), .B2(keyinput198), .ZN(n9138) );
  OAI221_X1 U10615 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput230), .C1(
        P1_REG2_REG_21__SCAN_IN), .C2(keyinput198), .A(n9138), .ZN(n9142) );
  AOI22_X1 U10616 ( .A1(P1_REG0_REG_25__SCAN_IN), .A2(keyinput201), .B1(n9140), 
        .B2(keyinput214), .ZN(n9139) );
  OAI221_X1 U10617 ( .B1(P1_REG0_REG_25__SCAN_IN), .B2(keyinput201), .C1(n9140), .C2(keyinput214), .A(n9139), .ZN(n9141) );
  NOR4_X1 U10618 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n9145)
         );
  NAND4_X1 U10619 ( .A1(n9148), .A2(n9147), .A3(n9146), .A4(n9145), .ZN(n9243)
         );
  AOI22_X1 U10620 ( .A1(n10015), .A2(keyinput157), .B1(n9600), .B2(keyinput134), .ZN(n9149) );
  OAI221_X1 U10621 ( .B1(n10015), .B2(keyinput157), .C1(n9600), .C2(
        keyinput134), .A(n9149), .ZN(n9158) );
  AOI22_X1 U10622 ( .A1(n9151), .A2(keyinput250), .B1(keyinput132), .B2(n9440), 
        .ZN(n9150) );
  OAI221_X1 U10623 ( .B1(n9151), .B2(keyinput250), .C1(n9440), .C2(keyinput132), .A(n9150), .ZN(n9157) );
  XNOR2_X1 U10624 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput254), .ZN(n9155)
         );
  XNOR2_X1 U10625 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput232), .ZN(n9154) );
  XNOR2_X1 U10626 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput172), .ZN(n9153) );
  XNOR2_X1 U10627 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput203), .ZN(n9152) );
  NAND4_X1 U10628 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), .ZN(n9156)
         );
  NOR3_X1 U10629 ( .A1(n9158), .A2(n9157), .A3(n9156), .ZN(n9196) );
  AOI22_X1 U10630 ( .A1(n6149), .A2(keyinput153), .B1(keyinput148), .B2(n9160), 
        .ZN(n9159) );
  OAI221_X1 U10631 ( .B1(n6149), .B2(keyinput153), .C1(n9160), .C2(keyinput148), .A(n9159), .ZN(n9169) );
  AOI22_X1 U10632 ( .A1(n10710), .A2(keyinput158), .B1(n9162), .B2(keyinput140), .ZN(n9161) );
  OAI221_X1 U10633 ( .B1(n10710), .B2(keyinput158), .C1(n9162), .C2(
        keyinput140), .A(n9161), .ZN(n9168) );
  AOI22_X1 U10634 ( .A1(n5365), .A2(keyinput220), .B1(n10592), .B2(keyinput183), .ZN(n9163) );
  OAI221_X1 U10635 ( .B1(n5365), .B2(keyinput220), .C1(n10592), .C2(
        keyinput183), .A(n9163), .ZN(n9167) );
  AOI22_X1 U10636 ( .A1(n10432), .A2(keyinput226), .B1(n9165), .B2(keyinput193), .ZN(n9164) );
  OAI221_X1 U10637 ( .B1(n10432), .B2(keyinput226), .C1(n9165), .C2(
        keyinput193), .A(n9164), .ZN(n9166) );
  NOR4_X1 U10638 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9195)
         );
  INV_X1 U10639 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10518) );
  AOI22_X1 U10640 ( .A1(n10518), .A2(keyinput246), .B1(keyinput208), .B2(n9255), .ZN(n9170) );
  OAI221_X1 U10641 ( .B1(n10518), .B2(keyinput246), .C1(n9255), .C2(
        keyinput208), .A(n9170), .ZN(n9181) );
  AOI22_X1 U10642 ( .A1(n9172), .A2(keyinput236), .B1(keyinput223), .B2(n7253), 
        .ZN(n9171) );
  OAI221_X1 U10643 ( .B1(n9172), .B2(keyinput236), .C1(n7253), .C2(keyinput223), .A(n9171), .ZN(n9180) );
  AOI22_X1 U10644 ( .A1(n9175), .A2(keyinput141), .B1(n9174), .B2(keyinput192), 
        .ZN(n9173) );
  OAI221_X1 U10645 ( .B1(n9175), .B2(keyinput141), .C1(n9174), .C2(keyinput192), .A(n9173), .ZN(n9179) );
  INV_X1 U10646 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10682) );
  XOR2_X1 U10647 ( .A(n10682), .B(keyinput173), .Z(n9177) );
  XNOR2_X1 U10648 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput174), .ZN(n9176) );
  NAND2_X1 U10649 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  NOR4_X1 U10650 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n9194)
         );
  INV_X1 U10651 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U10652 ( .A1(n10585), .A2(keyinput239), .B1(n6415), .B2(keyinput196), .ZN(n9182) );
  OAI221_X1 U10653 ( .B1(n10585), .B2(keyinput239), .C1(n6415), .C2(
        keyinput196), .A(n9182), .ZN(n9192) );
  AOI22_X1 U10654 ( .A1(n10729), .A2(keyinput216), .B1(n10636), .B2(
        keyinput169), .ZN(n9183) );
  OAI221_X1 U10655 ( .B1(n10729), .B2(keyinput216), .C1(n10636), .C2(
        keyinput169), .A(n9183), .ZN(n9191) );
  AOI22_X1 U10656 ( .A1(n9186), .A2(keyinput199), .B1(keyinput191), .B2(n9185), 
        .ZN(n9184) );
  OAI221_X1 U10657 ( .B1(n9186), .B2(keyinput199), .C1(n9185), .C2(keyinput191), .A(n9184), .ZN(n9190) );
  XNOR2_X1 U10658 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput206), .ZN(n9188)
         );
  XNOR2_X1 U10659 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput245), .ZN(n9187) );
  NAND2_X1 U10660 ( .A1(n9188), .A2(n9187), .ZN(n9189) );
  NOR4_X1 U10661 ( .A1(n9192), .A2(n9191), .A3(n9190), .A4(n9189), .ZN(n9193)
         );
  NAND4_X1 U10662 ( .A1(n9196), .A2(n9195), .A3(n9194), .A4(n9193), .ZN(n9242)
         );
  AOI22_X1 U10663 ( .A1(n9472), .A2(keyinput175), .B1(keyinput247), .B2(n9292), 
        .ZN(n9197) );
  OAI221_X1 U10664 ( .B1(n9472), .B2(keyinput175), .C1(n9292), .C2(keyinput247), .A(n9197), .ZN(n9206) );
  AOI22_X1 U10665 ( .A1(n9199), .A2(keyinput133), .B1(n9396), .B2(keyinput229), 
        .ZN(n9198) );
  OAI221_X1 U10666 ( .B1(n9199), .B2(keyinput133), .C1(n9396), .C2(keyinput229), .A(n9198), .ZN(n9205) );
  XNOR2_X1 U10667 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput139), .ZN(n9203) );
  XNOR2_X1 U10668 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput204), .ZN(n9202)
         );
  XNOR2_X1 U10669 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput221), .ZN(n9201) );
  XNOR2_X1 U10670 ( .A(keyinput217), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9200)
         );
  NAND4_X1 U10671 ( .A1(n9203), .A2(n9202), .A3(n9201), .A4(n9200), .ZN(n9204)
         );
  NOR3_X1 U10672 ( .A1(n9206), .A2(n9205), .A3(n9204), .ZN(n9240) );
  AOI22_X1 U10673 ( .A1(n6306), .A2(keyinput128), .B1(keyinput162), .B2(n5426), 
        .ZN(n9207) );
  OAI221_X1 U10674 ( .B1(n6306), .B2(keyinput128), .C1(n5426), .C2(keyinput162), .A(n9207), .ZN(n9215) );
  INV_X1 U10675 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9271) );
  AOI22_X1 U10676 ( .A1(n9668), .A2(keyinput240), .B1(keyinput243), .B2(n9271), 
        .ZN(n9208) );
  OAI221_X1 U10677 ( .B1(n9668), .B2(keyinput240), .C1(n9271), .C2(keyinput243), .A(n9208), .ZN(n9214) );
  INV_X1 U10678 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9262) );
  XOR2_X1 U10679 ( .A(n9262), .B(keyinput170), .Z(n9212) );
  INV_X1 U10680 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9420) );
  XOR2_X1 U10681 ( .A(n9420), .B(keyinput235), .Z(n9211) );
  XNOR2_X1 U10682 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput211), .ZN(n9210) );
  XNOR2_X1 U10683 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput161), .ZN(n9209) );
  NAND4_X1 U10684 ( .A1(n9212), .A2(n9211), .A3(n9210), .A4(n9209), .ZN(n9213)
         );
  NOR3_X1 U10685 ( .A1(n9215), .A2(n9214), .A3(n9213), .ZN(n9239) );
  INV_X1 U10686 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U10687 ( .A1(n10583), .A2(keyinput166), .B1(keyinput252), .B2(
        n10063), .ZN(n9216) );
  OAI221_X1 U10688 ( .B1(n10583), .B2(keyinput166), .C1(n10063), .C2(
        keyinput252), .A(n9216), .ZN(n9226) );
  AOI22_X1 U10689 ( .A1(n9218), .A2(keyinput181), .B1(keyinput164), .B2(n6990), 
        .ZN(n9217) );
  OAI221_X1 U10690 ( .B1(n9218), .B2(keyinput181), .C1(n6990), .C2(keyinput164), .A(n9217), .ZN(n9225) );
  AOI22_X1 U10691 ( .A1(n5199), .A2(keyinput180), .B1(n9220), .B2(keyinput135), 
        .ZN(n9219) );
  OAI221_X1 U10692 ( .B1(n5199), .B2(keyinput180), .C1(n9220), .C2(keyinput135), .A(n9219), .ZN(n9224) );
  INV_X1 U10693 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9222) );
  AOI22_X1 U10694 ( .A1(n9222), .A2(keyinput137), .B1(keyinput165), .B2(n9559), 
        .ZN(n9221) );
  OAI221_X1 U10695 ( .B1(n9222), .B2(keyinput137), .C1(n9559), .C2(keyinput165), .A(n9221), .ZN(n9223) );
  NOR4_X1 U10696 ( .A1(n9226), .A2(n9225), .A3(n9224), .A4(n9223), .ZN(n9238)
         );
  AOI22_X1 U10697 ( .A1(n9409), .A2(keyinput142), .B1(n9228), .B2(keyinput150), 
        .ZN(n9227) );
  OAI221_X1 U10698 ( .B1(n9409), .B2(keyinput142), .C1(n9228), .C2(keyinput150), .A(n9227), .ZN(n9236) );
  AOI22_X1 U10699 ( .A1(n5866), .A2(keyinput242), .B1(n10349), .B2(keyinput187), .ZN(n9229) );
  OAI221_X1 U10700 ( .B1(n5866), .B2(keyinput242), .C1(n10349), .C2(
        keyinput187), .A(n9229), .ZN(n9235) );
  XOR2_X1 U10701 ( .A(n9397), .B(keyinput228), .Z(n9233) );
  XNOR2_X1 U10702 ( .A(keyinput149), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n9232) );
  XNOR2_X1 U10703 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput144), .ZN(n9231) );
  XNOR2_X1 U10704 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput177), .ZN(n9230) );
  NAND4_X1 U10705 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n9234)
         );
  NOR3_X1 U10706 ( .A1(n9236), .A2(n9235), .A3(n9234), .ZN(n9237) );
  NAND4_X1 U10707 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n9241)
         );
  NOR4_X1 U10708 ( .A1(n9244), .A2(n9243), .A3(n9242), .A4(n9241), .ZN(n9435)
         );
  OAI22_X1 U10709 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(keyinput1), .B1(
        keyinput121), .B2(P1_D_REG_0__SCAN_IN), .ZN(n9245) );
  AOI221_X1 U10710 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(keyinput1), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput121), .A(n9245), .ZN(n9252) );
  OAI22_X1 U10711 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput54), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(keyinput88), .ZN(n9246) );
  AOI221_X1 U10712 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput54), .C1(
        keyinput88), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n9246), .ZN(n9251) );
  OAI22_X1 U10713 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput63), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput31), .ZN(n9247) );
  AOI221_X1 U10714 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput63), .C1(
        keyinput31), .C2(P1_REG2_REG_27__SCAN_IN), .A(n9247), .ZN(n9250) );
  OAI22_X1 U10715 ( .A1(P2_D_REG_24__SCAN_IN), .A2(keyinput108), .B1(
        P1_REG0_REG_21__SCAN_IN), .B2(keyinput103), .ZN(n9248) );
  AOI221_X1 U10716 ( .B1(P2_D_REG_24__SCAN_IN), .B2(keyinput108), .C1(
        keyinput103), .C2(P1_REG0_REG_21__SCAN_IN), .A(n9248), .ZN(n9249) );
  NAND4_X1 U10717 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n9258)
         );
  AOI22_X1 U10718 ( .A1(n5365), .A2(keyinput92), .B1(keyinput41), .B2(n10636), 
        .ZN(n9253) );
  OAI221_X1 U10719 ( .B1(n5365), .B2(keyinput92), .C1(n10636), .C2(keyinput41), 
        .A(n9253), .ZN(n9257) );
  AOI22_X1 U10720 ( .A1(n6149), .A2(keyinput25), .B1(keyinput80), .B2(n9255), 
        .ZN(n9254) );
  OAI221_X1 U10721 ( .B1(n6149), .B2(keyinput25), .C1(n9255), .C2(keyinput80), 
        .A(n9254), .ZN(n9256) );
  NOR3_X1 U10722 ( .A1(n9258), .A2(n9257), .A3(n9256), .ZN(n9301) );
  OAI22_X1 U10723 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput71), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput67), .ZN(n9259) );
  AOI221_X1 U10724 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput71), .C1(
        keyinput67), .C2(P1_REG0_REG_24__SCAN_IN), .A(n9259), .ZN(n9268) );
  OAI22_X1 U10725 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(keyinput70), .B1(
        keyinput24), .B2(P1_REG1_REG_22__SCAN_IN), .ZN(n9260) );
  AOI221_X1 U10726 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(keyinput70), .C1(
        P1_REG1_REG_22__SCAN_IN), .C2(keyinput24), .A(n9260), .ZN(n9267) );
  OAI22_X1 U10727 ( .A1(n9262), .A2(keyinput42), .B1(n5463), .B2(keyinput116), 
        .ZN(n9261) );
  AOI221_X1 U10728 ( .B1(n9262), .B2(keyinput42), .C1(keyinput116), .C2(n5463), 
        .A(n9261), .ZN(n9266) );
  OAI22_X1 U10729 ( .A1(n9264), .A2(keyinput51), .B1(keyinput48), .B2(
        P1_IR_REG_14__SCAN_IN), .ZN(n9263) );
  AOI221_X1 U10730 ( .B1(n9264), .B2(keyinput51), .C1(P1_IR_REG_14__SCAN_IN), 
        .C2(keyinput48), .A(n9263), .ZN(n9265) );
  NAND4_X1 U10731 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(n9285)
         );
  AOI22_X1 U10732 ( .A1(n9271), .A2(keyinput115), .B1(n9270), .B2(keyinput62), 
        .ZN(n9269) );
  OAI221_X1 U10733 ( .B1(n9271), .B2(keyinput115), .C1(n9270), .C2(keyinput62), 
        .A(n9269), .ZN(n9276) );
  AOI22_X1 U10734 ( .A1(n9274), .A2(keyinput126), .B1(n9273), .B2(keyinput105), 
        .ZN(n9272) );
  OAI221_X1 U10735 ( .B1(n9274), .B2(keyinput126), .C1(n9273), .C2(keyinput105), .A(n9272), .ZN(n9275) );
  NOR2_X1 U10736 ( .A1(n9276), .A2(n9275), .ZN(n9283) );
  INV_X1 U10737 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10587) );
  INV_X1 U10738 ( .A(keyinput66), .ZN(n9277) );
  XNOR2_X1 U10739 ( .A(n10587), .B(n9277), .ZN(n9282) );
  AOI22_X1 U10740 ( .A1(n10583), .A2(keyinput38), .B1(n9279), .B2(keyinput110), 
        .ZN(n9278) );
  OAI221_X1 U10741 ( .B1(n10583), .B2(keyinput38), .C1(n9279), .C2(keyinput110), .A(n9278), .ZN(n9280) );
  INV_X1 U10742 ( .A(n9280), .ZN(n9281) );
  NAND3_X1 U10743 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(n9284) );
  NOR2_X1 U10744 ( .A1(n9285), .A2(n9284), .ZN(n9300) );
  INV_X1 U10745 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U10746 ( .A1(n10584), .A2(keyinput94), .B1(n8702), .B2(keyinput89), 
        .ZN(n9286) );
  OAI221_X1 U10747 ( .B1(n10584), .B2(keyinput94), .C1(n8702), .C2(keyinput89), 
        .A(n9286), .ZN(n9290) );
  AOI22_X1 U10748 ( .A1(n9288), .A2(keyinput43), .B1(n5866), .B2(keyinput114), 
        .ZN(n9287) );
  OAI221_X1 U10749 ( .B1(n9288), .B2(keyinput43), .C1(n5866), .C2(keyinput114), 
        .A(n9287), .ZN(n9289) );
  NOR2_X1 U10750 ( .A1(n9290), .A2(n9289), .ZN(n9299) );
  AOI22_X1 U10751 ( .A1(n9293), .A2(keyinput76), .B1(keyinput119), .B2(n9292), 
        .ZN(n9291) );
  OAI221_X1 U10752 ( .B1(n9293), .B2(keyinput76), .C1(n9292), .C2(keyinput119), 
        .A(n9291), .ZN(n9297) );
  AOI22_X1 U10753 ( .A1(n9295), .A2(keyinput85), .B1(keyinput72), .B2(n10594), 
        .ZN(n9294) );
  OAI221_X1 U10754 ( .B1(n9295), .B2(keyinput85), .C1(n10594), .C2(keyinput72), 
        .A(n9294), .ZN(n9296) );
  NOR2_X1 U10755 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  NAND4_X1 U10756 ( .A1(n9301), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(n9394)
         );
  OAI22_X1 U10757 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput26), .B1(
        P1_REG0_REG_2__SCAN_IN), .B2(keyinput34), .ZN(n9302) );
  AOI221_X1 U10758 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput26), .C1(
        keyinput34), .C2(P1_REG0_REG_2__SCAN_IN), .A(n9302), .ZN(n9309) );
  OAI22_X1 U10759 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput13), .B1(
        keyinput5), .B2(P1_REG3_REG_7__SCAN_IN), .ZN(n9303) );
  AOI221_X1 U10760 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput13), .C1(
        P1_REG3_REG_7__SCAN_IN), .C2(keyinput5), .A(n9303), .ZN(n9308) );
  OAI22_X1 U10761 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput127), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput49), .ZN(n9304) );
  AOI221_X1 U10762 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput127), .C1(
        keyinput49), .C2(P1_IR_REG_10__SCAN_IN), .A(n9304), .ZN(n9307) );
  OAI22_X1 U10763 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput9), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput19), .ZN(n9305) );
  AOI221_X1 U10764 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput9), .C1(
        keyinput19), .C2(P2_IR_REG_9__SCAN_IN), .A(n9305), .ZN(n9306) );
  NAND4_X1 U10765 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n9319)
         );
  OAI22_X1 U10766 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput44), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput97), .ZN(n9310) );
  AOI221_X1 U10767 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput44), .C1(
        keyinput97), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n9310), .ZN(n9317) );
  OAI22_X1 U10768 ( .A1(P2_D_REG_5__SCAN_IN), .A2(keyinput86), .B1(keyinput60), 
        .B2(SI_30_), .ZN(n9311) );
  AOI221_X1 U10769 ( .B1(P2_D_REG_5__SCAN_IN), .B2(keyinput86), .C1(SI_30_), 
        .C2(keyinput60), .A(n9311), .ZN(n9316) );
  OAI22_X1 U10770 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput27), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(keyinput3), .ZN(n9312) );
  AOI221_X1 U10771 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput27), .C1(
        keyinput3), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9312), .ZN(n9315) );
  OAI22_X1 U10772 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(keyinput7), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput113), .ZN(n9313) );
  AOI221_X1 U10773 ( .B1(P2_IR_REG_11__SCAN_IN), .B2(keyinput7), .C1(
        keyinput113), .C2(P2_D_REG_31__SCAN_IN), .A(n9313), .ZN(n9314) );
  NAND4_X1 U10774 ( .A1(n9317), .A2(n9316), .A3(n9315), .A4(n9314), .ZN(n9318)
         );
  NOR2_X1 U10775 ( .A1(n9319), .A2(n9318), .ZN(n9392) );
  OAI22_X1 U10776 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput65), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput104), .ZN(n9320) );
  AOI221_X1 U10777 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput65), .C1(
        keyinput104), .C2(P2_REG2_REG_2__SCAN_IN), .A(n9320), .ZN(n9327) );
  OAI22_X1 U10778 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput112), .B1(
        keyinput52), .B2(P1_REG2_REG_28__SCAN_IN), .ZN(n9321) );
  AOI221_X1 U10779 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput112), .C1(
        P1_REG2_REG_28__SCAN_IN), .C2(keyinput52), .A(n9321), .ZN(n9326) );
  OAI22_X1 U10780 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput78), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(keyinput122), .ZN(n9322) );
  AOI221_X1 U10781 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput78), .C1(
        keyinput122), .C2(P1_DATAO_REG_9__SCAN_IN), .A(n9322), .ZN(n9325) );
  OAI22_X1 U10782 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(keyinput99), .B1(
        keyinput32), .B2(P1_IR_REG_31__SCAN_IN), .ZN(n9323) );
  AOI221_X1 U10783 ( .B1(P2_DATAO_REG_5__SCAN_IN), .B2(keyinput99), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput32), .A(n9323), .ZN(n9324) );
  NAND4_X1 U10784 ( .A1(n9327), .A2(n9326), .A3(n9325), .A4(n9324), .ZN(n9338)
         );
  AOI22_X1 U10785 ( .A1(n6990), .A2(keyinput36), .B1(keyinput73), .B2(n9329), 
        .ZN(n9328) );
  OAI221_X1 U10786 ( .B1(n6990), .B2(keyinput36), .C1(n9329), .C2(keyinput73), 
        .A(n9328), .ZN(n9330) );
  INV_X1 U10787 ( .A(n9330), .ZN(n9336) );
  AOI22_X1 U10788 ( .A1(n7666), .A2(keyinput15), .B1(keyinput6), .B2(n9600), 
        .ZN(n9331) );
  OAI221_X1 U10789 ( .B1(n7666), .B2(keyinput15), .C1(n9600), .C2(keyinput6), 
        .A(n9331), .ZN(n9332) );
  INV_X1 U10790 ( .A(n9332), .ZN(n9335) );
  INV_X1 U10791 ( .A(keyinput111), .ZN(n9333) );
  XNOR2_X1 U10792 ( .A(n10585), .B(n9333), .ZN(n9334) );
  NAND3_X1 U10793 ( .A1(n9336), .A2(n9335), .A3(n9334), .ZN(n9337) );
  NOR2_X1 U10794 ( .A1(n9338), .A2(n9337), .ZN(n9391) );
  OAI22_X1 U10795 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput64), .B1(
        P1_REG2_REG_10__SCAN_IN), .B2(keyinput95), .ZN(n9339) );
  AOI221_X1 U10796 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput64), .C1(
        keyinput95), .C2(P1_REG2_REG_10__SCAN_IN), .A(n9339), .ZN(n9346) );
  OAI22_X1 U10797 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput35), .B1(
        P1_REG2_REG_8__SCAN_IN), .B2(keyinput91), .ZN(n9340) );
  AOI221_X1 U10798 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput35), .C1(
        keyinput91), .C2(P1_REG2_REG_8__SCAN_IN), .A(n9340), .ZN(n9345) );
  OAI22_X1 U10799 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(keyinput4), .B1(
        keyinput58), .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9341) );
  AOI221_X1 U10800 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(keyinput4), .C1(
        P1_ADDR_REG_2__SCAN_IN), .C2(keyinput58), .A(n9341), .ZN(n9344) );
  OAI22_X1 U10801 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput18), .B1(
        P2_ADDR_REG_0__SCAN_IN), .B2(keyinput102), .ZN(n9342) );
  AOI221_X1 U10802 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput18), .C1(
        keyinput102), .C2(P2_ADDR_REG_0__SCAN_IN), .A(n9342), .ZN(n9343) );
  NAND4_X1 U10803 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n9356)
         );
  OAI22_X1 U10804 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput53), .B1(keyinput84), 
        .B2(P2_REG2_REG_19__SCAN_IN), .ZN(n9347) );
  AOI221_X1 U10805 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput53), .C1(
        P2_REG2_REG_19__SCAN_IN), .C2(keyinput84), .A(n9347), .ZN(n9354) );
  OAI22_X1 U10806 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(keyinput39), .B1(keyinput22), .B2(P2_D_REG_6__SCAN_IN), .ZN(n9348) );
  AOI221_X1 U10807 ( .B1(P2_IR_REG_4__SCAN_IN), .B2(keyinput39), .C1(
        P2_D_REG_6__SCAN_IN), .C2(keyinput22), .A(n9348), .ZN(n9353) );
  OAI22_X1 U10808 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput56), .B1(
        keyinput12), .B2(P1_REG2_REG_22__SCAN_IN), .ZN(n9349) );
  AOI221_X1 U10809 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput56), .C1(
        P1_REG2_REG_22__SCAN_IN), .C2(keyinput12), .A(n9349), .ZN(n9352) );
  OAI22_X1 U10810 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput87), .B1(
        P2_IR_REG_3__SCAN_IN), .B2(keyinput16), .ZN(n9350) );
  AOI221_X1 U10811 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput87), .C1(
        keyinput16), .C2(P2_IR_REG_3__SCAN_IN), .A(n9350), .ZN(n9351) );
  NAND4_X1 U10812 ( .A1(n9354), .A2(n9353), .A3(n9352), .A4(n9351), .ZN(n9355)
         );
  NOR2_X1 U10813 ( .A1(n9356), .A2(n9355), .ZN(n9390) );
  OAI22_X1 U10814 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput90), .B1(
        keyinput57), .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n9357) );
  AOI221_X1 U10815 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput90), .C1(
        P2_REG0_REG_16__SCAN_IN), .C2(keyinput57), .A(n9357), .ZN(n9364) );
  OAI22_X1 U10816 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput117), .B1(
        keyinput21), .B2(P1_REG1_REG_9__SCAN_IN), .ZN(n9358) );
  AOI221_X1 U10817 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput117), .C1(
        P1_REG1_REG_9__SCAN_IN), .C2(keyinput21), .A(n9358), .ZN(n9363) );
  OAI22_X1 U10818 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput82), .B1(
        P1_REG3_REG_19__SCAN_IN), .B2(keyinput37), .ZN(n9359) );
  AOI221_X1 U10819 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput82), .C1(
        keyinput37), .C2(P1_REG3_REG_19__SCAN_IN), .A(n9359), .ZN(n9362) );
  OAI22_X1 U10820 ( .A1(P1_D_REG_31__SCAN_IN), .A2(keyinput50), .B1(
        P1_REG1_REG_23__SCAN_IN), .B2(keyinput59), .ZN(n9360) );
  AOI221_X1 U10821 ( .B1(P1_D_REG_31__SCAN_IN), .B2(keyinput50), .C1(
        keyinput59), .C2(P1_REG1_REG_23__SCAN_IN), .A(n9360), .ZN(n9361) );
  NAND4_X1 U10822 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9388)
         );
  XNOR2_X1 U10823 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput109), .ZN(n9368)
         );
  XNOR2_X1 U10824 ( .A(SI_4_), .B(keyinput28), .ZN(n9367) );
  XNOR2_X1 U10825 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput77), .ZN(n9366) );
  XNOR2_X1 U10826 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput98), .ZN(n9365) );
  NAND4_X1 U10827 ( .A1(n9368), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n9374)
         );
  XNOR2_X1 U10828 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput83), .ZN(n9372) );
  XNOR2_X1 U10829 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput11), .ZN(n9371) );
  XNOR2_X1 U10830 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput2), .ZN(n9370) );
  XNOR2_X1 U10831 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput46), .ZN(n9369) );
  NAND4_X1 U10832 ( .A1(n9372), .A2(n9371), .A3(n9370), .A4(n9369), .ZN(n9373)
         );
  NOR2_X1 U10833 ( .A1(n9374), .A2(n9373), .ZN(n9386) );
  XNOR2_X1 U10834 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput75), .ZN(n9378) );
  XNOR2_X1 U10835 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput8), .ZN(n9377) );
  XNOR2_X1 U10836 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput93), .ZN(n9376) );
  XNOR2_X1 U10837 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput33), .ZN(n9375) );
  NAND4_X1 U10838 ( .A1(n9378), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n9384)
         );
  XNOR2_X1 U10839 ( .A(keyinput123), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9382) );
  XNOR2_X1 U10840 ( .A(keyinput30), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n9381) );
  XNOR2_X1 U10841 ( .A(keyinput20), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U10842 ( .A(keyinput23), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n9379) );
  NAND4_X1 U10843 ( .A1(n9382), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9383)
         );
  NOR2_X1 U10844 ( .A1(n9384), .A2(n9383), .ZN(n9385) );
  NAND2_X1 U10845 ( .A1(n9386), .A2(n9385), .ZN(n9387) );
  NOR2_X1 U10846 ( .A1(n9388), .A2(n9387), .ZN(n9389) );
  NAND4_X1 U10847 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), .ZN(n9393)
         );
  NOR2_X1 U10848 ( .A1(n9394), .A2(n9393), .ZN(n9433) );
  AOI22_X1 U10849 ( .A1(n9397), .A2(keyinput100), .B1(n9396), .B2(keyinput101), 
        .ZN(n9395) );
  OAI221_X1 U10850 ( .B1(n9397), .B2(keyinput100), .C1(n9396), .C2(keyinput101), .A(n9395), .ZN(n9406) );
  AOI22_X1 U10851 ( .A1(n10682), .A2(keyinput45), .B1(n9483), .B2(keyinput96), 
        .ZN(n9398) );
  OAI221_X1 U10852 ( .B1(n10682), .B2(keyinput45), .C1(n9483), .C2(keyinput96), 
        .A(n9398), .ZN(n9405) );
  AOI22_X1 U10853 ( .A1(n6415), .A2(keyinput68), .B1(n9400), .B2(keyinput17), 
        .ZN(n9399) );
  OAI221_X1 U10854 ( .B1(n6415), .B2(keyinput68), .C1(n9400), .C2(keyinput17), 
        .A(n9399), .ZN(n9404) );
  AOI22_X1 U10855 ( .A1(n10015), .A2(keyinput29), .B1(n9402), .B2(keyinput79), 
        .ZN(n9401) );
  OAI221_X1 U10856 ( .B1(n10015), .B2(keyinput29), .C1(n9402), .C2(keyinput79), 
        .A(n9401), .ZN(n9403) );
  NOR4_X1 U10857 ( .A1(n9406), .A2(n9405), .A3(n9404), .A4(n9403), .ZN(n9432)
         );
  AOI22_X1 U10858 ( .A1(n9409), .A2(keyinput14), .B1(keyinput69), .B2(n9408), 
        .ZN(n9407) );
  OAI221_X1 U10859 ( .B1(n9409), .B2(keyinput14), .C1(n9408), .C2(keyinput69), 
        .A(n9407), .ZN(n9418) );
  AOI22_X1 U10860 ( .A1(n9472), .A2(keyinput47), .B1(keyinput118), .B2(n10518), 
        .ZN(n9410) );
  OAI221_X1 U10861 ( .B1(n9472), .B2(keyinput47), .C1(n10518), .C2(keyinput118), .A(n9410), .ZN(n9417) );
  AOI22_X1 U10862 ( .A1(n10063), .A2(keyinput124), .B1(n9412), .B2(keyinput120), .ZN(n9411) );
  OAI221_X1 U10863 ( .B1(n10063), .B2(keyinput124), .C1(n9412), .C2(
        keyinput120), .A(n9411), .ZN(n9416) );
  INV_X1 U10864 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10436) );
  INV_X1 U10865 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9414) );
  AOI22_X1 U10866 ( .A1(n10436), .A2(keyinput125), .B1(n9414), .B2(keyinput106), .ZN(n9413) );
  OAI221_X1 U10867 ( .B1(n10436), .B2(keyinput125), .C1(n9414), .C2(
        keyinput106), .A(n9413), .ZN(n9415) );
  NOR4_X1 U10868 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n9415), .ZN(n9431)
         );
  AOI22_X1 U10869 ( .A1(n10586), .A2(keyinput74), .B1(n9420), .B2(keyinput107), 
        .ZN(n9419) );
  OAI221_X1 U10870 ( .B1(n10586), .B2(keyinput74), .C1(n9420), .C2(keyinput107), .A(n9419), .ZN(n9429) );
  AOI22_X1 U10871 ( .A1(n9422), .A2(keyinput81), .B1(keyinput0), .B2(n6306), 
        .ZN(n9421) );
  OAI221_X1 U10872 ( .B1(n9422), .B2(keyinput81), .C1(n6306), .C2(keyinput0), 
        .A(n9421), .ZN(n9428) );
  AOI22_X1 U10873 ( .A1(n10592), .A2(keyinput55), .B1(keyinput10), .B2(n10233), 
        .ZN(n9423) );
  OAI221_X1 U10874 ( .B1(n10592), .B2(keyinput55), .C1(n10233), .C2(keyinput10), .A(n9423), .ZN(n9427) );
  AOI22_X1 U10875 ( .A1(n6356), .A2(keyinput61), .B1(n9425), .B2(keyinput40), 
        .ZN(n9424) );
  OAI221_X1 U10876 ( .B1(n6356), .B2(keyinput61), .C1(n9425), .C2(keyinput40), 
        .A(n9424), .ZN(n9426) );
  NOR4_X1 U10877 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n9430)
         );
  NAND4_X1 U10878 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(n9430), .ZN(n9434)
         );
  OR2_X1 U10879 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  XNOR2_X1 U10880 ( .A(n9437), .B(n9436), .ZN(P2_U3477) );
  AOI21_X1 U10881 ( .B1(n9449), .B2(n9439), .A(n9438), .ZN(n9511) );
  MUX2_X1 U10882 ( .A(n9440), .B(n9511), .S(n9456), .Z(n9441) );
  OAI21_X1 U10883 ( .B1(n9515), .B2(n9442), .A(n9441), .ZN(P2_U3476) );
  NAND2_X1 U10884 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  OAI211_X1 U10885 ( .C1(n9448), .C2(n9447), .A(n9446), .B(n9445), .ZN(n9516)
         );
  MUX2_X1 U10886 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9516), .S(n9456), .Z(
        P2_U3475) );
  NAND3_X1 U10887 ( .A1(n9451), .A2(n9450), .A3(n9449), .ZN(n9452) );
  OAI211_X1 U10888 ( .C1(n9455), .C2(n9454), .A(n9453), .B(n9452), .ZN(n9517)
         );
  MUX2_X1 U10889 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9517), .S(n9456), .Z(
        P2_U3474) );
  NOR2_X1 U10890 ( .A1(n9457), .A2(n10685), .ZN(n9460) );
  AOI21_X1 U10891 ( .B1(n10685), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9460), .ZN(
        n9458) );
  OAI21_X1 U10892 ( .B1(n9459), .B2(n9514), .A(n9458), .ZN(P2_U3458) );
  AOI21_X1 U10893 ( .B1(n10685), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9460), .ZN(
        n9461) );
  OAI21_X1 U10894 ( .B1(n9462), .B2(n9514), .A(n9461), .ZN(P2_U3457) );
  NAND2_X1 U10895 ( .A1(n9463), .A2(n10683), .ZN(n9466) );
  INV_X1 U10896 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U10897 ( .A1(n9466), .A2(n9465), .ZN(n9470) );
  NAND2_X1 U10898 ( .A1(n9468), .A2(n9467), .ZN(n9469) );
  NAND2_X1 U10899 ( .A1(n9470), .A2(n9469), .ZN(P2_U3456) );
  MUX2_X1 U10900 ( .A(n9472), .B(n9471), .S(n10683), .Z(n9473) );
  OAI21_X1 U10901 ( .B1(n9474), .B2(n9514), .A(n9473), .ZN(P2_U3455) );
  INV_X1 U10902 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U10903 ( .A(n9479), .B(n9478), .S(n10683), .Z(n9480) );
  OAI21_X1 U10904 ( .B1(n9481), .B2(n9514), .A(n9480), .ZN(P2_U3453) );
  MUX2_X1 U10905 ( .A(n9483), .B(n9482), .S(n10683), .Z(n9484) );
  OAI21_X1 U10906 ( .B1(n9485), .B2(n9514), .A(n9484), .ZN(P2_U3452) );
  INV_X1 U10907 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9487) );
  MUX2_X1 U10908 ( .A(n9487), .B(n9486), .S(n10683), .Z(n9488) );
  OAI21_X1 U10909 ( .B1(n9489), .B2(n9514), .A(n9488), .ZN(P2_U3451) );
  INV_X1 U10910 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9491) );
  MUX2_X1 U10911 ( .A(n9491), .B(n9490), .S(n10683), .Z(n9492) );
  OAI21_X1 U10912 ( .B1(n9493), .B2(n9514), .A(n9492), .ZN(P2_U3450) );
  INV_X1 U10913 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U10914 ( .A(n9495), .B(n9494), .S(n10683), .Z(n9496) );
  OAI21_X1 U10915 ( .B1(n9497), .B2(n9514), .A(n9496), .ZN(P2_U3449) );
  INV_X1 U10916 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9499) );
  MUX2_X1 U10917 ( .A(n9499), .B(n9498), .S(n10683), .Z(n9500) );
  OAI21_X1 U10918 ( .B1(n9501), .B2(n9514), .A(n9500), .ZN(P2_U3448) );
  INV_X1 U10919 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9503) );
  MUX2_X1 U10920 ( .A(n9503), .B(n9502), .S(n10683), .Z(n9504) );
  OAI21_X1 U10921 ( .B1(n9505), .B2(n9514), .A(n9504), .ZN(P2_U3447) );
  INV_X1 U10922 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9507) );
  MUX2_X1 U10923 ( .A(n9507), .B(n9506), .S(n10683), .Z(n9508) );
  OAI21_X1 U10924 ( .B1(n9509), .B2(n9514), .A(n9508), .ZN(P2_U3446) );
  MUX2_X1 U10925 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9510), .S(n10683), .Z(
        P2_U3444) );
  INV_X1 U10926 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9512) );
  MUX2_X1 U10927 ( .A(n9512), .B(n9511), .S(n10683), .Z(n9513) );
  OAI21_X1 U10928 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(P2_U3441) );
  MUX2_X1 U10929 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9516), .S(n10683), .Z(
        P2_U3438) );
  MUX2_X1 U10930 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9517), .S(n10683), .Z(
        P2_U3435) );
  INV_X1 U10931 ( .A(n9673), .ZN(n10466) );
  NOR4_X1 U10932 ( .A1(n9520), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9518), .ZN(n9521) );
  AOI21_X1 U10933 ( .B1(n9522), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9521), .ZN(
        n9523) );
  OAI21_X1 U10934 ( .B1(n10466), .B2(n9524), .A(n9523), .ZN(P2_U3264) );
  MUX2_X1 U10935 ( .A(n9525), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10936 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  XOR2_X1 U10937 ( .A(n9529), .B(n9528), .Z(n9536) );
  AOI22_X1 U10938 ( .A1(n10541), .A2(n9530), .B1(P1_REG3_REG_14__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9531) );
  OAI21_X1 U10939 ( .B1(n9532), .B2(n10547), .A(n9531), .ZN(n9533) );
  AOI21_X1 U10940 ( .B1(n9534), .B2(n10502), .A(n9533), .ZN(n9535) );
  OAI21_X1 U10941 ( .B1(n9536), .B2(n10535), .A(n9535), .ZN(P1_U3215) );
  AOI21_X1 U10942 ( .B1(n9539), .B2(n9537), .A(n9538), .ZN(n9545) );
  AND2_X1 U10943 ( .A1(n9965), .A2(n9666), .ZN(n9540) );
  AOI21_X1 U10944 ( .B1(n9963), .B2(n9667), .A(n9540), .ZN(n10344) );
  INV_X1 U10945 ( .A(n9541), .ZN(n10182) );
  AOI22_X1 U10946 ( .A1(n10182), .A2(n9638), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9542) );
  OAI21_X1 U10947 ( .B1(n10344), .B2(n10492), .A(n9542), .ZN(n9543) );
  AOI21_X1 U10948 ( .B1(n10179), .B2(n10515), .A(n9543), .ZN(n9544) );
  OAI21_X1 U10949 ( .B1(n9545), .B2(n10535), .A(n9544), .ZN(P1_U3216) );
  OAI21_X1 U10950 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9549) );
  NAND2_X1 U10951 ( .A1(n9549), .A2(n10527), .ZN(n9555) );
  AOI22_X1 U10952 ( .A1(n10541), .A2(n9550), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n9554) );
  NAND2_X1 U10953 ( .A1(n9638), .A2(n5460), .ZN(n9553) );
  NAND2_X1 U10954 ( .A1(n10502), .A2(n4561), .ZN(n9552) );
  NAND4_X1 U10955 ( .A1(n9555), .A2(n9554), .A3(n9553), .A4(n9552), .ZN(
        P1_U3218) );
  XOR2_X1 U10956 ( .A(n9556), .B(n9557), .Z(n9563) );
  NOR2_X1 U10957 ( .A1(n10547), .A2(n10232), .ZN(n9561) );
  AND2_X1 U10958 ( .A1(n9969), .A2(n9666), .ZN(n9558) );
  AOI21_X1 U10959 ( .B1(n9967), .B2(n9667), .A(n9558), .ZN(n10239) );
  OAI22_X1 U10960 ( .A1(n10239), .A2(n10492), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9559), .ZN(n9560) );
  AOI211_X1 U10961 ( .C1(n10369), .C2(n10515), .A(n9561), .B(n9560), .ZN(n9562) );
  OAI21_X1 U10962 ( .B1(n9563), .B2(n10535), .A(n9562), .ZN(P1_U3219) );
  NAND2_X1 U10963 ( .A1(n9565), .A2(n9564), .ZN(n9571) );
  OR2_X1 U10964 ( .A1(n9566), .A2(n9567), .ZN(n9569) );
  NAND2_X1 U10965 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  XOR2_X1 U10966 ( .A(n9571), .B(n9570), .Z(n9577) );
  NAND2_X1 U10967 ( .A1(n9965), .A2(n9667), .ZN(n9573) );
  NAND2_X1 U10968 ( .A1(n9967), .A2(n9666), .ZN(n9572) );
  NAND2_X1 U10969 ( .A1(n9573), .A2(n9572), .ZN(n10205) );
  AOI22_X1 U10970 ( .A1(n10205), .A2(n10541), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9574) );
  OAI21_X1 U10971 ( .B1(n10210), .B2(n10547), .A(n9574), .ZN(n9575) );
  AOI21_X1 U10972 ( .B1(n10428), .B2(n10515), .A(n9575), .ZN(n9576) );
  OAI21_X1 U10973 ( .B1(n9577), .B2(n10535), .A(n9576), .ZN(P1_U3223) );
  XOR2_X1 U10974 ( .A(n9579), .B(n9578), .Z(n9583) );
  AOI22_X1 U10975 ( .A1(n9961), .A2(n9667), .B1(n9666), .B2(n9963), .ZN(n10148) );
  AOI22_X1 U10976 ( .A1(n10153), .A2(n9638), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9580) );
  OAI21_X1 U10977 ( .B1(n10148), .B2(n10492), .A(n9580), .ZN(n9581) );
  AOI21_X1 U10978 ( .B1(n10411), .B2(n10515), .A(n9581), .ZN(n9582) );
  OAI21_X1 U10979 ( .B1(n9583), .B2(n10535), .A(n9582), .ZN(P1_U3225) );
  INV_X1 U10980 ( .A(n9587), .ZN(n9584) );
  NOR2_X1 U10981 ( .A1(n9585), .A2(n9584), .ZN(n9590) );
  AOI21_X1 U10982 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n9589) );
  OAI21_X1 U10983 ( .B1(n9590), .B2(n9589), .A(n10527), .ZN(n9593) );
  AOI22_X1 U10984 ( .A1(n9970), .A2(n9667), .B1(n9972), .B2(n9666), .ZN(n10283) );
  NAND2_X1 U10985 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10027)
         );
  OAI21_X1 U10986 ( .B1(n10492), .B2(n10283), .A(n10027), .ZN(n9591) );
  AOI21_X1 U10987 ( .B1(n10291), .B2(n9638), .A(n9591), .ZN(n9592) );
  OAI211_X1 U10988 ( .C1(n10293), .C2(n10543), .A(n9593), .B(n9592), .ZN(
        P1_U3226) );
  OAI21_X1 U10989 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9597) );
  NAND2_X1 U10990 ( .A1(n9597), .A2(n10527), .ZN(n9603) );
  NAND2_X1 U10991 ( .A1(n9969), .A2(n9667), .ZN(n9599) );
  NAND2_X1 U10992 ( .A1(n9971), .A2(n9666), .ZN(n9598) );
  NAND2_X1 U10993 ( .A1(n9599), .A2(n9598), .ZN(n10265) );
  NOR2_X1 U10994 ( .A1(n9600), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10054) );
  NOR2_X1 U10995 ( .A1(n10547), .A2(n10271), .ZN(n9601) );
  AOI211_X1 U10996 ( .C1(n10541), .C2(n10265), .A(n10054), .B(n9601), .ZN(
        n9602) );
  OAI211_X1 U10997 ( .C1(n10274), .C2(n10543), .A(n9603), .B(n9602), .ZN(
        P1_U3228) );
  XOR2_X1 U10998 ( .A(n9604), .B(n4584), .Z(n9608) );
  AOI22_X1 U10999 ( .A1(n9962), .A2(n9667), .B1(n9666), .B2(n9964), .ZN(n10164) );
  AOI22_X1 U11000 ( .A1(n10167), .A2(n9638), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9605) );
  OAI21_X1 U11001 ( .B1(n10164), .B2(n10492), .A(n9605), .ZN(n9606) );
  AOI21_X1 U11002 ( .B1(n10341), .B2(n10515), .A(n9606), .ZN(n9607) );
  OAI21_X1 U11003 ( .B1(n9608), .B2(n10535), .A(n9607), .ZN(P1_U3229) );
  XNOR2_X1 U11004 ( .A(n9610), .B(n9609), .ZN(n9611) );
  XNOR2_X1 U11005 ( .A(n9566), .B(n9611), .ZN(n9617) );
  AND2_X1 U11006 ( .A1(n9968), .A2(n9666), .ZN(n9612) );
  AOI21_X1 U11007 ( .B1(n9966), .B2(n9667), .A(n9612), .ZN(n10219) );
  OAI22_X1 U11008 ( .A1(n10219), .A2(n10492), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9613), .ZN(n9615) );
  NOR2_X1 U11009 ( .A1(n10225), .A2(n10543), .ZN(n9614) );
  AOI211_X1 U11010 ( .C1(n9638), .C2(n10222), .A(n9615), .B(n9614), .ZN(n9616)
         );
  OAI21_X1 U11011 ( .B1(n9617), .B2(n10535), .A(n9616), .ZN(P1_U3233) );
  OAI21_X1 U11012 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9621) );
  NAND2_X1 U11013 ( .A1(n9621), .A2(n10527), .ZN(n9628) );
  INV_X1 U11014 ( .A(n9622), .ZN(n9626) );
  OAI22_X1 U11015 ( .A1(n10492), .A2(n9624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9623), .ZN(n9625) );
  AOI21_X1 U11016 ( .B1(n9626), .B2(n9638), .A(n9625), .ZN(n9627) );
  OAI211_X1 U11017 ( .C1(n9629), .C2(n10543), .A(n9628), .B(n9627), .ZN(
        P1_U3234) );
  INV_X1 U11018 ( .A(n9537), .ZN(n9636) );
  INV_X1 U11019 ( .A(n9630), .ZN(n9632) );
  NAND2_X1 U11020 ( .A1(n9632), .A2(n9631), .ZN(n9634) );
  AOI22_X1 U11021 ( .A1(n9636), .A2(n9635), .B1(n9634), .B2(n9633), .ZN(n9642)
         );
  AND2_X1 U11022 ( .A1(n9966), .A2(n9666), .ZN(n9637) );
  AOI21_X1 U11023 ( .B1(n9964), .B2(n9667), .A(n9637), .ZN(n10191) );
  AOI22_X1 U11024 ( .A1(n9638), .A2(n10195), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9639) );
  OAI21_X1 U11025 ( .B1(n10191), .B2(n10492), .A(n9639), .ZN(n9640) );
  AOI21_X1 U11026 ( .B1(n10194), .B2(n10515), .A(n9640), .ZN(n9641) );
  OAI21_X1 U11027 ( .B1(n9642), .B2(n10535), .A(n9641), .ZN(P1_U3235) );
  XNOR2_X1 U11028 ( .A(n9644), .B(n9643), .ZN(n9645) );
  XNOR2_X1 U11029 ( .A(n9646), .B(n9645), .ZN(n9652) );
  NOR2_X1 U11030 ( .A1(n10547), .A2(n10252), .ZN(n9650) );
  AND2_X1 U11031 ( .A1(n9970), .A2(n9666), .ZN(n9647) );
  AOI21_X1 U11032 ( .B1(n9968), .B2(n9667), .A(n9647), .ZN(n10248) );
  OAI22_X1 U11033 ( .A1(n10248), .A2(n10492), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9648), .ZN(n9649) );
  AOI211_X1 U11034 ( .C1(n10374), .C2(n10502), .A(n9650), .B(n9649), .ZN(n9651) );
  OAI21_X1 U11035 ( .B1(n9652), .B2(n10535), .A(n9651), .ZN(P1_U3238) );
  OAI211_X1 U11036 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n10527), .ZN(n9661)
         );
  NAND2_X1 U11037 ( .A1(n9960), .A2(n9667), .ZN(n9657) );
  NAND2_X1 U11038 ( .A1(n9962), .A2(n9666), .ZN(n9656) );
  NAND2_X1 U11039 ( .A1(n9657), .A2(n9656), .ZN(n10134) );
  OAI22_X1 U11040 ( .A1(n10138), .A2(n10547), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9658), .ZN(n9659) );
  AOI21_X1 U11041 ( .B1(n10134), .B2(n10541), .A(n9659), .ZN(n9660) );
  OAI211_X1 U11042 ( .C1(n10142), .C2(n10543), .A(n9661), .B(n9660), .ZN(
        P1_U3240) );
  NAND2_X1 U11043 ( .A1(n9663), .A2(n9662), .ZN(n9665) );
  XNOR2_X1 U11044 ( .A(n9665), .B(n9664), .ZN(n9672) );
  NOR2_X1 U11045 ( .A1(n10547), .A2(n10297), .ZN(n9670) );
  AOI22_X1 U11046 ( .A1(n9667), .A2(n9971), .B1(n9973), .B2(n9666), .ZN(n10301) );
  OAI22_X1 U11047 ( .A1(n10492), .A2(n10301), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9668), .ZN(n9669) );
  AOI211_X1 U11048 ( .C1(n10454), .C2(n10502), .A(n9670), .B(n9669), .ZN(n9671) );
  OAI21_X1 U11049 ( .B1(n9672), .B2(n10535), .A(n9671), .ZN(P1_U3241) );
  NAND2_X1 U11050 ( .A1(n9673), .A2(n5337), .ZN(n9676) );
  OR2_X1 U11051 ( .A1(n5420), .A2(n9674), .ZN(n9675) );
  INV_X1 U11052 ( .A(n10398), .ZN(n9792) );
  NAND2_X1 U11053 ( .A1(n9792), .A2(n10104), .ZN(n9931) );
  INV_X1 U11054 ( .A(n9931), .ZN(n9800) );
  AND2_X1 U11055 ( .A1(n9770), .A2(n9677), .ZN(n9842) );
  INV_X1 U11056 ( .A(n10217), .ZN(n9679) );
  NAND2_X1 U11057 ( .A1(n10202), .A2(n9941), .ZN(n9678) );
  OAI21_X1 U11058 ( .B1(n9679), .B2(n10369), .A(n9678), .ZN(n9680) );
  NAND2_X1 U11059 ( .A1(n9680), .A2(n9906), .ZN(n9683) );
  NAND3_X1 U11060 ( .A1(n9681), .A2(n9968), .A3(n9795), .ZN(n9682) );
  NAND2_X1 U11061 ( .A1(n9683), .A2(n9682), .ZN(n9756) );
  INV_X1 U11062 ( .A(n9743), .ZN(n9825) );
  INV_X1 U11063 ( .A(n9809), .ZN(n9877) );
  OAI211_X1 U11064 ( .C1(n9684), .C2(n9877), .A(n9813), .B(n9703), .ZN(n9686)
         );
  AND4_X1 U11065 ( .A1(n9882), .A2(n9880), .A3(n9879), .A4(n9795), .ZN(n9685)
         );
  NAND2_X1 U11066 ( .A1(n9686), .A2(n9685), .ZN(n9712) );
  NAND2_X1 U11067 ( .A1(n9982), .A2(n9795), .ZN(n9692) );
  INV_X1 U11068 ( .A(n9692), .ZN(n9687) );
  AOI22_X1 U11069 ( .A1(n9687), .A2(n10602), .B1(n9981), .B2(n9795), .ZN(n9699) );
  NAND2_X1 U11070 ( .A1(n9688), .A2(n9941), .ZN(n9691) );
  OAI22_X1 U11071 ( .A1(n9691), .A2(n10602), .B1(n9981), .B2(n9795), .ZN(n9689) );
  NAND2_X1 U11072 ( .A1(n9689), .A2(n9698), .ZN(n9697) );
  OAI21_X1 U11073 ( .B1(n9691), .B2(n9981), .A(n9690), .ZN(n9695) );
  OAI21_X1 U11074 ( .B1(n9693), .B2(n9692), .A(n10602), .ZN(n9694) );
  NAND2_X1 U11075 ( .A1(n9695), .A2(n9694), .ZN(n9696) );
  OAI211_X1 U11076 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9700)
         );
  INV_X1 U11077 ( .A(n9700), .ZN(n9710) );
  INV_X1 U11078 ( .A(n9701), .ZN(n9702) );
  NAND2_X1 U11079 ( .A1(n9702), .A2(n9808), .ZN(n9870) );
  AND2_X1 U11080 ( .A1(n9704), .A2(n9703), .ZN(n9872) );
  NAND2_X1 U11081 ( .A1(n9809), .A2(n9879), .ZN(n9705) );
  AOI21_X1 U11082 ( .B1(n9870), .B2(n9872), .A(n9705), .ZN(n9708) );
  NAND4_X1 U11083 ( .A1(n9706), .A2(n9884), .A3(n9876), .A4(n9941), .ZN(n9707)
         );
  OR2_X1 U11084 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  NAND4_X1 U11085 ( .A1(n9712), .A2(n9711), .A3(n9710), .A4(n9709), .ZN(n9719)
         );
  NAND2_X1 U11086 ( .A1(n9714), .A2(n9713), .ZN(n9716) );
  MUX2_X1 U11087 ( .A(n9716), .B(n9715), .S(n9795), .Z(n9717) );
  INV_X1 U11088 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U11089 ( .A1(n9719), .A2(n9718), .ZN(n9724) );
  INV_X1 U11090 ( .A(n9720), .ZN(n9721) );
  MUX2_X1 U11091 ( .A(n9722), .B(n9721), .S(n9795), .Z(n9723) );
  NAND2_X1 U11092 ( .A1(n9724), .A2(n9723), .ZN(n9735) );
  NAND2_X1 U11093 ( .A1(n9735), .A2(n9732), .ZN(n9725) );
  NAND2_X1 U11094 ( .A1(n9738), .A2(n9736), .ZN(n9890) );
  AOI21_X1 U11095 ( .B1(n9725), .B2(n9891), .A(n9890), .ZN(n9726) );
  NAND2_X1 U11096 ( .A1(n9739), .A2(n9737), .ZN(n9895) );
  OAI21_X1 U11097 ( .B1(n9726), .B2(n9895), .A(n9893), .ZN(n9727) );
  NAND2_X1 U11098 ( .A1(n9727), .A2(n9897), .ZN(n9728) );
  NAND3_X1 U11099 ( .A1(n9825), .A2(n9894), .A3(n9728), .ZN(n9729) );
  NAND4_X1 U11100 ( .A1(n9900), .A2(n10298), .A3(n9899), .A4(n9729), .ZN(n9745) );
  NAND2_X1 U11101 ( .A1(n10260), .A2(n9972), .ZN(n9730) );
  NAND2_X1 U11102 ( .A1(n9730), .A2(n9941), .ZN(n9749) );
  AND2_X1 U11103 ( .A1(n9746), .A2(n9731), .ZN(n9903) );
  INV_X1 U11104 ( .A(n9732), .ZN(n9734) );
  AOI21_X1 U11105 ( .B1(n9740), .B2(n9739), .A(n4857), .ZN(n9742) );
  INV_X1 U11106 ( .A(n9897), .ZN(n9741) );
  NAND2_X1 U11107 ( .A1(n9900), .A2(n4853), .ZN(n9747) );
  NAND2_X1 U11108 ( .A1(n9747), .A2(n10260), .ZN(n9748) );
  NAND2_X1 U11109 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  NAND2_X1 U11110 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U11111 ( .A1(n9752), .A2(n10268), .ZN(n9759) );
  NAND2_X1 U11112 ( .A1(n9760), .A2(n9753), .ZN(n9828) );
  INV_X1 U11113 ( .A(n9828), .ZN(n9910) );
  NAND2_X1 U11114 ( .A1(n9759), .A2(n9910), .ZN(n9754) );
  NAND4_X1 U11115 ( .A1(n9754), .A2(n9905), .A3(n9906), .A4(n9795), .ZN(n9755)
         );
  NAND2_X1 U11116 ( .A1(n9756), .A2(n9755), .ZN(n9758) );
  NAND2_X1 U11117 ( .A1(n9861), .A2(n9795), .ZN(n9757) );
  NAND2_X1 U11118 ( .A1(n9758), .A2(n9757), .ZN(n9767) );
  NAND3_X1 U11119 ( .A1(n9759), .A2(n10245), .A3(n9905), .ZN(n9761) );
  INV_X1 U11120 ( .A(n9763), .ZN(n9764) );
  AOI21_X1 U11121 ( .B1(n9941), .B2(n9765), .A(n9764), .ZN(n9766) );
  OAI21_X1 U11122 ( .B1(n9768), .B2(n10160), .A(n9841), .ZN(n9773) );
  NOR2_X1 U11123 ( .A1(n9771), .A2(n10160), .ZN(n9772) );
  INV_X1 U11124 ( .A(n9848), .ZN(n9774) );
  NAND2_X1 U11125 ( .A1(n9847), .A2(n9805), .ZN(n9845) );
  INV_X1 U11126 ( .A(n9845), .ZN(n9776) );
  INV_X1 U11127 ( .A(n9854), .ZN(n9864) );
  AND2_X1 U11128 ( .A1(n9778), .A2(n9777), .ZN(n9857) );
  NAND2_X1 U11129 ( .A1(n9780), .A2(n9779), .ZN(n9784) );
  NAND2_X1 U11130 ( .A1(n9781), .A2(n9854), .ZN(n9782) );
  AOI21_X1 U11131 ( .B1(n9782), .B2(n9857), .A(n9863), .ZN(n9783) );
  MUX2_X1 U11132 ( .A(n9784), .B(n9783), .S(n9941), .Z(n9788) );
  INV_X1 U11133 ( .A(n9913), .ZN(n9786) );
  INV_X1 U11134 ( .A(n9866), .ZN(n9785) );
  MUX2_X1 U11135 ( .A(n9786), .B(n9785), .S(n9795), .Z(n9787) );
  NAND2_X1 U11136 ( .A1(n9789), .A2(n5337), .ZN(n9791) );
  INV_X1 U11137 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10469) );
  OR2_X1 U11138 ( .A1(n5420), .A2(n10469), .ZN(n9790) );
  MUX2_X1 U11139 ( .A(n9941), .B(n9796), .S(n10108), .Z(n9794) );
  INV_X1 U11140 ( .A(n9804), .ZN(n9957) );
  NAND2_X1 U11141 ( .A1(n9792), .A2(n9957), .ZN(n9793) );
  MUX2_X1 U11142 ( .A(n9796), .B(n9795), .S(n10108), .Z(n9799) );
  NAND2_X1 U11143 ( .A1(n9929), .A2(n9957), .ZN(n9797) );
  NAND2_X1 U11144 ( .A1(n9943), .A2(n9797), .ZN(n9798) );
  AOI21_X1 U11145 ( .B1(n9941), .B2(n9800), .A(n9922), .ZN(n9956) );
  INV_X1 U11146 ( .A(n9801), .ZN(n9942) );
  NOR2_X1 U11147 ( .A1(n9940), .A2(n9802), .ZN(n9950) );
  OAI211_X1 U11148 ( .C1(n9943), .C2(n9938), .A(n9942), .B(n9950), .ZN(n9955)
         );
  NOR2_X1 U11149 ( .A1(n10108), .A2(n9804), .ZN(n9930) );
  INV_X1 U11150 ( .A(n9930), .ZN(n9803) );
  NAND2_X1 U11151 ( .A1(n9931), .A2(n9803), .ZN(n9915) );
  NAND2_X1 U11152 ( .A1(n10108), .A2(n9804), .ZN(n9914) );
  NAND2_X1 U11153 ( .A1(n9805), .A2(n9848), .ZN(n10146) );
  XNOR2_X1 U11154 ( .A(n10428), .B(n9806), .ZN(n10204) );
  NAND3_X1 U11155 ( .A1(n9809), .A2(n9808), .A3(n9807), .ZN(n9810) );
  NOR2_X1 U11156 ( .A1(n9811), .A2(n9810), .ZN(n9814) );
  NAND4_X1 U11157 ( .A1(n9814), .A2(n9813), .A3(n9872), .A4(n9812), .ZN(n9816)
         );
  NOR2_X1 U11158 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  AND4_X1 U11159 ( .A1(n9887), .A2(n9886), .A3(n9817), .A4(n9882), .ZN(n9818)
         );
  NAND4_X1 U11160 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9822)
         );
  NOR2_X1 U11161 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  NAND2_X1 U11162 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  NOR2_X1 U11163 ( .A1(n10305), .A2(n9826), .ZN(n9827) );
  NAND4_X1 U11164 ( .A1(n9905), .A2(n10287), .A3(n9827), .A4(n10245), .ZN(
        n9829) );
  NOR2_X1 U11165 ( .A1(n9829), .A2(n9828), .ZN(n9830) );
  NAND3_X1 U11166 ( .A1(n10217), .A2(n10236), .A3(n9830), .ZN(n9831) );
  NOR3_X1 U11167 ( .A1(n9832), .A2(n10204), .A3(n9831), .ZN(n9833) );
  NAND2_X1 U11168 ( .A1(n10176), .A2(n9833), .ZN(n9834) );
  OR4_X1 U11169 ( .A1(n10128), .A2(n10146), .A3(n9834), .A4(n10160), .ZN(n9835) );
  NOR2_X1 U11170 ( .A1(n9836), .A2(n9835), .ZN(n9837) );
  NAND4_X1 U11171 ( .A1(n9914), .A2(n9838), .A3(n10116), .A4(n9837), .ZN(n9839) );
  OR3_X1 U11172 ( .A1(n9933), .A2(n9915), .A3(n9839), .ZN(n9935) );
  INV_X1 U11173 ( .A(n9935), .ZN(n9920) );
  NAND2_X1 U11174 ( .A1(n9841), .A2(n9840), .ZN(n9846) );
  NOR2_X1 U11175 ( .A1(n9846), .A2(n9842), .ZN(n9843) );
  OR3_X1 U11176 ( .A1(n9845), .A2(n9844), .A3(n9843), .ZN(n9862) );
  INV_X1 U11177 ( .A(n9846), .ZN(n9850) );
  INV_X1 U11178 ( .A(n9847), .ZN(n9849) );
  OAI22_X1 U11179 ( .A1(n9862), .A2(n9850), .B1(n9849), .B2(n9848), .ZN(n9856)
         );
  AND2_X1 U11180 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NOR2_X1 U11181 ( .A1(n9862), .A2(n9853), .ZN(n9855) );
  OAI21_X1 U11182 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9858) );
  AND2_X1 U11183 ( .A1(n9858), .A2(n9857), .ZN(n9865) );
  INV_X1 U11184 ( .A(n9865), .ZN(n9860) );
  NOR2_X1 U11185 ( .A1(n9862), .A2(n9861), .ZN(n9868) );
  AOI21_X1 U11186 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9867) );
  INV_X1 U11187 ( .A(n9870), .ZN(n9875) );
  OAI211_X1 U11188 ( .C1(n4688), .C2(n5897), .A(n9871), .B(n5820), .ZN(n9874)
         );
  INV_X1 U11189 ( .A(n9872), .ZN(n9873) );
  AOI21_X1 U11190 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(n9878) );
  OAI21_X1 U11191 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(n9881) );
  NAND3_X1 U11192 ( .A1(n9881), .A2(n9880), .A3(n9879), .ZN(n9885) );
  INV_X1 U11193 ( .A(n9882), .ZN(n9883) );
  AOI21_X1 U11194 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9889) );
  INV_X1 U11195 ( .A(n9886), .ZN(n9888) );
  OAI21_X1 U11196 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9892) );
  AOI21_X1 U11197 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9896) );
  OAI211_X1 U11198 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9898)
         );
  NAND3_X1 U11199 ( .A1(n9898), .A2(n9897), .A3(n10298), .ZN(n9902) );
  INV_X1 U11200 ( .A(n9899), .ZN(n9901) );
  AOI211_X1 U11201 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n4800), .ZN(n9904)
         );
  OAI21_X1 U11202 ( .B1(n9904), .B2(n4804), .A(n10245), .ZN(n9909) );
  INV_X1 U11203 ( .A(n9905), .ZN(n9908) );
  INV_X1 U11204 ( .A(n9906), .ZN(n9907) );
  AOI211_X1 U11205 ( .C1(n9910), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9911)
         );
  NOR3_X1 U11206 ( .A1(n9923), .A2(n4851), .A3(n9911), .ZN(n9912) );
  NOR2_X1 U11207 ( .A1(n9924), .A2(n9912), .ZN(n9917) );
  NAND2_X1 U11208 ( .A1(n9914), .A2(n9913), .ZN(n9927) );
  INV_X1 U11209 ( .A(n9915), .ZN(n9916) );
  OAI21_X1 U11210 ( .B1(n9917), .B2(n9927), .A(n9916), .ZN(n9944) );
  NAND2_X1 U11211 ( .A1(n9944), .A2(n9943), .ZN(n9919) );
  MUX2_X1 U11212 ( .A(n9920), .B(n9919), .S(n4549), .Z(n9921) );
  INV_X1 U11213 ( .A(n9923), .ZN(n9925) );
  AOI21_X1 U11214 ( .B1(n4687), .B2(n9925), .A(n9924), .ZN(n9926) );
  AOI21_X1 U11215 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n9934) );
  OAI211_X1 U11216 ( .C1(n9934), .C2(n9933), .A(n9932), .B(n9931), .ZN(n9937)
         );
  NAND3_X1 U11217 ( .A1(n9937), .A2(n9936), .A3(n9935), .ZN(n9939) );
  AOI21_X1 U11218 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(n9946) );
  NAND3_X1 U11219 ( .A1(n9944), .A2(n9949), .A3(n9943), .ZN(n9945) );
  NAND3_X1 U11220 ( .A1(n9947), .A2(n9946), .A3(n9945), .ZN(n9954) );
  NAND3_X1 U11221 ( .A1(n9666), .A2(n9949), .A3(n9948), .ZN(n9952) );
  INV_X1 U11222 ( .A(n9950), .ZN(n9951) );
  OAI211_X1 U11223 ( .C1(n9952), .C2(n10458), .A(P1_B_REG_SCAN_IN), .B(n9951), 
        .ZN(n9953) );
  OAI211_X1 U11224 ( .C1(n9956), .C2(n9955), .A(n9954), .B(n9953), .ZN(
        P1_U3242) );
  MUX2_X1 U11225 ( .A(n9957), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9985), .Z(
        P1_U3584) );
  MUX2_X1 U11226 ( .A(n9958), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9985), .Z(
        P1_U3583) );
  MUX2_X1 U11227 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9959), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11228 ( .A(n9960), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9985), .Z(
        P1_U3581) );
  MUX2_X1 U11229 ( .A(n9961), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9985), .Z(
        P1_U3580) );
  MUX2_X1 U11230 ( .A(n9962), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9985), .Z(
        P1_U3579) );
  MUX2_X1 U11231 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9963), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11232 ( .A(n9964), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9985), .Z(
        P1_U3577) );
  MUX2_X1 U11233 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9965), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11234 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9966), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11235 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9967), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11236 ( .A(n9968), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9985), .Z(
        P1_U3573) );
  MUX2_X1 U11237 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9969), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11238 ( .A(n9970), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9985), .Z(
        P1_U3571) );
  MUX2_X1 U11239 ( .A(n9971), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9985), .Z(
        P1_U3570) );
  MUX2_X1 U11240 ( .A(n9972), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9985), .Z(
        P1_U3569) );
  MUX2_X1 U11241 ( .A(n9973), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9985), .Z(
        P1_U3568) );
  MUX2_X1 U11242 ( .A(n9974), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9985), .Z(
        P1_U3567) );
  MUX2_X1 U11243 ( .A(n9975), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9985), .Z(
        P1_U3566) );
  MUX2_X1 U11244 ( .A(n9976), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9985), .Z(
        P1_U3565) );
  MUX2_X1 U11245 ( .A(n9977), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9985), .Z(
        P1_U3564) );
  MUX2_X1 U11246 ( .A(n9978), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9985), .Z(
        P1_U3563) );
  MUX2_X1 U11247 ( .A(n9979), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9985), .Z(
        P1_U3562) );
  MUX2_X1 U11248 ( .A(n9980), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9985), .Z(
        P1_U3561) );
  MUX2_X1 U11249 ( .A(n9981), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9985), .Z(
        P1_U3560) );
  MUX2_X1 U11250 ( .A(n9982), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9985), .Z(
        P1_U3559) );
  MUX2_X1 U11251 ( .A(n9983), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9985), .Z(
        P1_U3558) );
  MUX2_X1 U11252 ( .A(n9984), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9985), .Z(
        P1_U3557) );
  MUX2_X1 U11253 ( .A(n9986), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9985), .Z(
        P1_U3556) );
  MUX2_X1 U11254 ( .A(n9987), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9985), .Z(
        P1_U3555) );
  OAI211_X1 U11255 ( .C1(n9990), .C2(n9989), .A(n10087), .B(n9988), .ZN(n9997)
         );
  AOI22_X1 U11256 ( .A1(n10055), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9996) );
  NAND2_X1 U11257 ( .A1(n10072), .A2(n5400), .ZN(n9995) );
  OAI211_X1 U11258 ( .C1(n9993), .C2(n9992), .A(n10093), .B(n9991), .ZN(n9994)
         );
  NAND4_X1 U11259 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(
        P1_U3244) );
  NAND2_X1 U11260 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9998) );
  OAI21_X1 U11261 ( .B1(n10099), .B2(n9999), .A(n9998), .ZN(n10000) );
  AOI21_X1 U11262 ( .B1(n10072), .B2(n4690), .A(n10000), .ZN(n10010) );
  INV_X1 U11263 ( .A(n10001), .ZN(n10002) );
  OAI211_X1 U11264 ( .C1(n10004), .C2(n10003), .A(n10093), .B(n10002), .ZN(
        n10009) );
  OAI211_X1 U11265 ( .C1(n10007), .C2(n10006), .A(n10087), .B(n10005), .ZN(
        n10008) );
  NAND3_X1 U11266 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(P1_U3246) );
  AOI211_X1 U11267 ( .C1(n10013), .C2(n10012), .A(n10090), .B(n10011), .ZN(
        n10014) );
  INV_X1 U11268 ( .A(n10014), .ZN(n10023) );
  NAND2_X1 U11269 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10521) );
  OAI21_X1 U11270 ( .B1(n10099), .B2(n10015), .A(n10521), .ZN(n10016) );
  AOI21_X1 U11271 ( .B1(n10072), .B2(n10017), .A(n10016), .ZN(n10022) );
  OAI211_X1 U11272 ( .C1(n10020), .C2(n10019), .A(n10018), .B(n10093), .ZN(
        n10021) );
  NAND3_X1 U11273 ( .A1(n10023), .A2(n10022), .A3(n10021), .ZN(P1_U3251) );
  XNOR2_X1 U11274 ( .A(n10049), .B(n10044), .ZN(n10046) );
  NOR2_X1 U11275 ( .A1(n10024), .A2(n10032), .ZN(n10026) );
  XOR2_X1 U11276 ( .A(n10046), .B(n10047), .Z(n10043) );
  INV_X1 U11277 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10028) );
  OAI21_X1 U11278 ( .B1(n10099), .B2(n10028), .A(n10027), .ZN(n10041) );
  OR2_X1 U11279 ( .A1(n10049), .A2(n10029), .ZN(n10031) );
  NAND2_X1 U11280 ( .A1(n10049), .A2(n10029), .ZN(n10030) );
  AND2_X1 U11281 ( .A1(n10031), .A2(n10030), .ZN(n10039) );
  NOR2_X1 U11282 ( .A1(n10033), .A2(n10032), .ZN(n10035) );
  INV_X1 U11283 ( .A(n10051), .ZN(n10036) );
  AOI211_X1 U11284 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10040) );
  AOI211_X1 U11285 ( .C1(n10072), .C2(n10049), .A(n10041), .B(n10040), .ZN(
        n10042) );
  OAI21_X1 U11286 ( .B1(n10043), .B2(n10090), .A(n10042), .ZN(P1_U3259) );
  XNOR2_X1 U11287 ( .A(n10064), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10065) );
  XOR2_X1 U11288 ( .A(n10065), .B(n10066), .Z(n10061) );
  OR2_X1 U11289 ( .A1(n10064), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U11290 ( .A1(n10064), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10048) );
  AND2_X1 U11291 ( .A1(n10073), .A2(n10048), .ZN(n10053) );
  NAND2_X1 U11292 ( .A1(n10049), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U11293 ( .A1(n10052), .A2(n10053), .ZN(n10074) );
  OAI21_X1 U11294 ( .B1(n10053), .B2(n10052), .A(n10074), .ZN(n10059) );
  AOI21_X1 U11295 ( .B1(n10055), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10054), 
        .ZN(n10056) );
  OAI21_X1 U11296 ( .B1(n10057), .B2(n10089), .A(n10056), .ZN(n10058) );
  AOI21_X1 U11297 ( .B1(n10059), .B2(n10093), .A(n10058), .ZN(n10060) );
  OAI21_X1 U11298 ( .B1(n10061), .B2(n10090), .A(n10060), .ZN(P1_U3260) );
  NAND2_X1 U11299 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n10062)
         );
  OAI21_X1 U11300 ( .B1(n10099), .B2(n10063), .A(n10062), .ZN(n10071) );
  OAI22_X1 U11301 ( .A1(n10066), .A2(n10065), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n10064), .ZN(n10069) );
  NAND2_X1 U11302 ( .A1(n10075), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10084) );
  OAI21_X1 U11303 ( .B1(n10075), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10084), 
        .ZN(n10068) );
  INV_X1 U11304 ( .A(n10085), .ZN(n10067) );
  AOI211_X1 U11305 ( .C1(n10069), .C2(n10068), .A(n10090), .B(n10067), .ZN(
        n10070) );
  AOI211_X1 U11306 ( .C1(n10072), .C2(n10075), .A(n10071), .B(n10070), .ZN(
        n10080) );
  AND2_X1 U11307 ( .A1(n10074), .A2(n10073), .ZN(n10078) );
  OR2_X1 U11308 ( .A1(n10075), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U11309 ( .A1(n10075), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10081) );
  AND2_X1 U11310 ( .A1(n10076), .A2(n10081), .ZN(n10077) );
  NAND2_X1 U11311 ( .A1(n10078), .A2(n10077), .ZN(n10082) );
  OAI211_X1 U11312 ( .C1(n10078), .C2(n10077), .A(n10082), .B(n10093), .ZN(
        n10079) );
  NAND2_X1 U11313 ( .A1(n10080), .A2(n10079), .ZN(P1_U3261) );
  INV_X1 U11314 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U11315 ( .A1(n10082), .A2(n10081), .ZN(n10083) );
  XNOR2_X1 U11316 ( .A(n10083), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n10094) );
  INV_X1 U11317 ( .A(n10094), .ZN(n10088) );
  NAND2_X1 U11318 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  INV_X1 U11319 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10370) );
  XNOR2_X1 U11320 ( .A(n10086), .B(n10370), .ZN(n10091) );
  AOI22_X1 U11321 ( .A1(n10088), .A2(n10093), .B1(n10091), .B2(n10087), .ZN(
        n10096) );
  OAI21_X1 U11322 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(n10092) );
  AOI21_X1 U11323 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(n10095) );
  MUX2_X1 U11324 ( .A(n10096), .B(n10095), .S(n10211), .Z(n10098) );
  NAND2_X1 U11325 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n10097)
         );
  OAI211_X1 U11326 ( .C1(n10100), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        P1_U3262) );
  XNOR2_X1 U11327 ( .A(n10398), .B(n10101), .ZN(n10102) );
  NAND2_X1 U11328 ( .A1(n10315), .A2(n10548), .ZN(n10107) );
  NOR2_X1 U11329 ( .A1(n10104), .A2(n10103), .ZN(n10318) );
  INV_X1 U11330 ( .A(n10318), .ZN(n10105) );
  NOR2_X1 U11331 ( .A1(n10563), .A2(n10105), .ZN(n10111) );
  AOI21_X1 U11332 ( .B1(n10553), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10111), 
        .ZN(n10106) );
  OAI211_X1 U11333 ( .C1(n10398), .C2(n10556), .A(n10107), .B(n10106), .ZN(
        P1_U3263) );
  XOR2_X1 U11334 ( .A(n10109), .B(n10108), .Z(n10320) );
  NAND2_X1 U11335 ( .A1(n10320), .A2(n10110), .ZN(n10113) );
  AOI21_X1 U11336 ( .B1(n10553), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10111), 
        .ZN(n10112) );
  OAI211_X1 U11337 ( .C1(n4848), .C2(n10556), .A(n10113), .B(n10112), .ZN(
        P1_U3264) );
  OAI21_X1 U11338 ( .B1(n10116), .B2(n10115), .A(n10114), .ZN(n10119) );
  INV_X1 U11339 ( .A(n10117), .ZN(n10118) );
  AOI21_X1 U11340 ( .B1(n10119), .B2(n10285), .A(n10118), .ZN(n10328) );
  NAND3_X1 U11341 ( .A1(n10324), .A2(n10323), .A3(n10560), .ZN(n10127) );
  AOI211_X1 U11342 ( .C1(n10326), .C2(n10121), .A(n10308), .B(n10120), .ZN(
        n10325) );
  AOI22_X1 U11343 ( .A1(n10122), .A2(n10551), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10563), .ZN(n10123) );
  OAI21_X1 U11344 ( .B1(n10124), .B2(n10556), .A(n10123), .ZN(n10125) );
  AOI21_X1 U11345 ( .B1(n10325), .B2(n10548), .A(n10125), .ZN(n10126) );
  OAI211_X1 U11346 ( .C1(n10553), .C2(n10328), .A(n10127), .B(n10126), .ZN(
        P1_U3265) );
  XNOR2_X1 U11347 ( .A(n10129), .B(n10128), .ZN(n10408) );
  OAI21_X1 U11348 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10133) );
  NAND2_X1 U11349 ( .A1(n10133), .A2(n10285), .ZN(n10136) );
  INV_X1 U11350 ( .A(n10134), .ZN(n10135) );
  NAND2_X1 U11351 ( .A1(n10136), .A2(n10135), .ZN(n10331) );
  AOI211_X1 U11352 ( .C1(n10406), .C2(n10151), .A(n10308), .B(n10137), .ZN(
        n10330) );
  NAND2_X1 U11353 ( .A1(n10330), .A2(n10548), .ZN(n10141) );
  INV_X1 U11354 ( .A(n10138), .ZN(n10139) );
  AOI22_X1 U11355 ( .A1(n10139), .A2(n10551), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10563), .ZN(n10140) );
  OAI211_X1 U11356 ( .C1(n10142), .C2(n10556), .A(n10141), .B(n10140), .ZN(
        n10143) );
  AOI21_X1 U11357 ( .B1(n5878), .B2(n10331), .A(n10143), .ZN(n10144) );
  OAI21_X1 U11358 ( .B1(n10408), .B2(n10259), .A(n10144), .ZN(P1_U3267) );
  XOR2_X1 U11359 ( .A(n10146), .B(n10145), .Z(n10413) );
  XNOR2_X1 U11360 ( .A(n10147), .B(n10146), .ZN(n10150) );
  INV_X1 U11361 ( .A(n10148), .ZN(n10149) );
  AOI21_X1 U11362 ( .B1(n10150), .B2(n10285), .A(n10149), .ZN(n10336) );
  INV_X1 U11363 ( .A(n10336), .ZN(n10157) );
  OAI211_X1 U11364 ( .C1(n10152), .C2(n10166), .A(n10151), .B(n10319), .ZN(
        n10335) );
  AOI22_X1 U11365 ( .A1(n10153), .A2(n10551), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10563), .ZN(n10155) );
  NAND2_X1 U11366 ( .A1(n10411), .A2(n10278), .ZN(n10154) );
  OAI211_X1 U11367 ( .C1(n10335), .C2(n10275), .A(n10155), .B(n10154), .ZN(
        n10156) );
  AOI21_X1 U11368 ( .B1(n10157), .B2(n10241), .A(n10156), .ZN(n10158) );
  OAI21_X1 U11369 ( .B1(n10413), .B2(n10259), .A(n10158), .ZN(P1_U3268) );
  XNOR2_X1 U11370 ( .A(n10159), .B(n10160), .ZN(n10417) );
  INV_X1 U11371 ( .A(n10160), .ZN(n10161) );
  XNOR2_X1 U11372 ( .A(n10162), .B(n10161), .ZN(n10163) );
  NAND2_X1 U11373 ( .A1(n10163), .A2(n10285), .ZN(n10165) );
  NAND2_X1 U11374 ( .A1(n10165), .A2(n10164), .ZN(n10340) );
  AOI211_X1 U11375 ( .C1(n10341), .C2(n10180), .A(n10308), .B(n10166), .ZN(
        n10339) );
  NAND2_X1 U11376 ( .A1(n10339), .A2(n10548), .ZN(n10169) );
  AOI22_X1 U11377 ( .A1(n10167), .A2(n10551), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10563), .ZN(n10168) );
  OAI211_X1 U11378 ( .C1(n10170), .C2(n10556), .A(n10169), .B(n10168), .ZN(
        n10171) );
  AOI21_X1 U11379 ( .B1(n10241), .B2(n10340), .A(n10171), .ZN(n10172) );
  OAI21_X1 U11380 ( .B1(n10417), .B2(n10259), .A(n10172), .ZN(P1_U3269) );
  XNOR2_X1 U11381 ( .A(n10173), .B(n10176), .ZN(n10421) );
  AOI22_X1 U11382 ( .A1(n10179), .A2(n10278), .B1(n10553), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n10186) );
  OAI21_X1 U11383 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10177) );
  AND2_X1 U11384 ( .A1(n10177), .A2(n10285), .ZN(n10348) );
  AOI21_X1 U11385 ( .B1(n10179), .B2(n10193), .A(n10308), .ZN(n10181) );
  NAND2_X1 U11386 ( .A1(n10181), .A2(n10180), .ZN(n10345) );
  NAND2_X1 U11387 ( .A1(n10182), .A2(n10551), .ZN(n10183) );
  OAI211_X1 U11388 ( .C1(n10345), .C2(n10211), .A(n10344), .B(n10183), .ZN(
        n10184) );
  OAI21_X1 U11389 ( .B1(n10348), .B2(n10184), .A(n5878), .ZN(n10185) );
  OAI211_X1 U11390 ( .C1(n10421), .C2(n10259), .A(n10186), .B(n10185), .ZN(
        P1_U3270) );
  XNOR2_X1 U11391 ( .A(n10187), .B(n10190), .ZN(n10353) );
  INV_X1 U11392 ( .A(n10353), .ZN(n10200) );
  OAI211_X1 U11393 ( .C1(n10190), .C2(n10189), .A(n10188), .B(n10285), .ZN(
        n10192) );
  NAND2_X1 U11394 ( .A1(n10192), .A2(n10191), .ZN(n10351) );
  AOI211_X1 U11395 ( .C1(n10194), .C2(n10208), .A(n10308), .B(n10178), .ZN(
        n10352) );
  NAND2_X1 U11396 ( .A1(n10352), .A2(n10548), .ZN(n10197) );
  AOI22_X1 U11397 ( .A1(n10195), .A2(n10551), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10563), .ZN(n10196) );
  OAI211_X1 U11398 ( .C1(n4942), .C2(n10556), .A(n10197), .B(n10196), .ZN(
        n10198) );
  AOI21_X1 U11399 ( .B1(n5878), .B2(n10351), .A(n10198), .ZN(n10199) );
  OAI21_X1 U11400 ( .B1(n10200), .B2(n10259), .A(n10199), .ZN(P1_U3271) );
  XOR2_X1 U11401 ( .A(n10201), .B(n10204), .Z(n10430) );
  AOI22_X1 U11402 ( .A1(n10428), .A2(n10278), .B1(n10553), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U11403 ( .A1(n10217), .A2(n4687), .ZN(n10216) );
  NAND2_X1 U11404 ( .A1(n10216), .A2(n10202), .ZN(n10203) );
  XOR2_X1 U11405 ( .A(n10204), .B(n10203), .Z(n10207) );
  INV_X1 U11406 ( .A(n10205), .ZN(n10206) );
  OAI21_X1 U11407 ( .B1(n10207), .B2(n10302), .A(n10206), .ZN(n10357) );
  OAI211_X1 U11408 ( .C1(n10209), .C2(n10221), .A(n10319), .B(n10208), .ZN(
        n10358) );
  OAI22_X1 U11409 ( .A1(n10358), .A2(n10211), .B1(n10270), .B2(n10210), .ZN(
        n10212) );
  OAI21_X1 U11410 ( .B1(n10357), .B2(n10212), .A(n10241), .ZN(n10213) );
  OAI211_X1 U11411 ( .C1(n10430), .C2(n10259), .A(n10214), .B(n10213), .ZN(
        P1_U3272) );
  XNOR2_X1 U11412 ( .A(n10215), .B(n10217), .ZN(n10434) );
  OAI211_X1 U11413 ( .C1(n4687), .C2(n10217), .A(n10216), .B(n10285), .ZN(
        n10220) );
  NAND2_X1 U11414 ( .A1(n10220), .A2(n10219), .ZN(n10363) );
  AOI211_X1 U11415 ( .C1(n10364), .C2(n4847), .A(n10308), .B(n10221), .ZN(
        n10362) );
  NAND2_X1 U11416 ( .A1(n10362), .A2(n10548), .ZN(n10224) );
  AOI22_X1 U11417 ( .A1(n10553), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10222), 
        .B2(n10551), .ZN(n10223) );
  OAI211_X1 U11418 ( .C1(n10225), .C2(n10556), .A(n10224), .B(n10223), .ZN(
        n10226) );
  AOI21_X1 U11419 ( .B1(n5878), .B2(n10363), .A(n10226), .ZN(n10227) );
  OAI21_X1 U11420 ( .B1(n10434), .B2(n10259), .A(n10227), .ZN(P1_U3273) );
  XOR2_X1 U11421 ( .A(n10236), .B(n10228), .Z(n10438) );
  NAND2_X1 U11422 ( .A1(n10250), .A2(n10369), .ZN(n10229) );
  NAND2_X1 U11423 ( .A1(n10229), .A2(n10319), .ZN(n10230) );
  NOR2_X1 U11424 ( .A1(n10231), .A2(n10230), .ZN(n10368) );
  NOR2_X1 U11425 ( .A1(n4845), .A2(n10556), .ZN(n10235) );
  OAI22_X1 U11426 ( .A1(n10241), .A2(n10233), .B1(n10232), .B2(n10270), .ZN(
        n10234) );
  AOI211_X1 U11427 ( .C1(n10368), .C2(n10548), .A(n10235), .B(n10234), .ZN(
        n10243) );
  XNOR2_X1 U11428 ( .A(n10237), .B(n10236), .ZN(n10238) );
  NAND2_X1 U11429 ( .A1(n10238), .A2(n10285), .ZN(n10240) );
  NAND2_X1 U11430 ( .A1(n10240), .A2(n10239), .ZN(n10367) );
  NAND2_X1 U11431 ( .A1(n10367), .A2(n10241), .ZN(n10242) );
  OAI211_X1 U11432 ( .C1(n10438), .C2(n10259), .A(n10243), .B(n10242), .ZN(
        P1_U3274) );
  XOR2_X1 U11433 ( .A(n10246), .B(n10244), .Z(n10442) );
  NAND2_X1 U11434 ( .A1(n10263), .A2(n10245), .ZN(n10247) );
  XNOR2_X1 U11435 ( .A(n10247), .B(n10246), .ZN(n10249) );
  OAI21_X1 U11436 ( .B1(n10249), .B2(n10302), .A(n10248), .ZN(n10373) );
  INV_X1 U11437 ( .A(n10250), .ZN(n10251) );
  AOI211_X1 U11438 ( .C1(n10374), .C2(n10273), .A(n10308), .B(n10251), .ZN(
        n10372) );
  NAND2_X1 U11439 ( .A1(n10372), .A2(n10548), .ZN(n10255) );
  INV_X1 U11440 ( .A(n10252), .ZN(n10253) );
  AOI22_X1 U11441 ( .A1(n10553), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10253), 
        .B2(n10551), .ZN(n10254) );
  OAI211_X1 U11442 ( .C1(n10256), .C2(n10556), .A(n10255), .B(n10254), .ZN(
        n10257) );
  AOI21_X1 U11443 ( .B1(n5878), .B2(n10373), .A(n10257), .ZN(n10258) );
  OAI21_X1 U11444 ( .B1(n10442), .B2(n10259), .A(n10258), .ZN(P1_U3275) );
  NAND2_X1 U11445 ( .A1(n10281), .A2(n10260), .ZN(n10262) );
  INV_X1 U11446 ( .A(n10268), .ZN(n10261) );
  NAND2_X1 U11447 ( .A1(n10262), .A2(n10261), .ZN(n10264) );
  NAND3_X1 U11448 ( .A1(n10264), .A2(n10263), .A3(n10285), .ZN(n10267) );
  INV_X1 U11449 ( .A(n10265), .ZN(n10266) );
  XNOR2_X1 U11450 ( .A(n4637), .B(n10268), .ZN(n10448) );
  INV_X1 U11451 ( .A(n10448), .ZN(n10269) );
  NAND2_X1 U11452 ( .A1(n10269), .A2(n10560), .ZN(n10280) );
  OAI22_X1 U11453 ( .A1(n5878), .A2(n10272), .B1(n10271), .B2(n10270), .ZN(
        n10277) );
  OAI211_X1 U11454 ( .C1(n10289), .C2(n10274), .A(n10319), .B(n10273), .ZN(
        n10377) );
  NOR2_X1 U11455 ( .A1(n10377), .A2(n10275), .ZN(n10276) );
  AOI211_X1 U11456 ( .C1(n10278), .C2(n10443), .A(n10277), .B(n10276), .ZN(
        n10279) );
  OAI211_X1 U11457 ( .C1(n10563), .C2(n10378), .A(n10280), .B(n10279), .ZN(
        P1_U3276) );
  OAI21_X1 U11458 ( .B1(n10287), .B2(n10282), .A(n10281), .ZN(n10286) );
  INV_X1 U11459 ( .A(n10283), .ZN(n10284) );
  AOI21_X1 U11460 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(n10386) );
  NAND2_X1 U11461 ( .A1(n10288), .A2(n10287), .ZN(n10382) );
  NAND3_X1 U11462 ( .A1(n4922), .A2(n10560), .A3(n10382), .ZN(n10296) );
  INV_X1 U11463 ( .A(n10307), .ZN(n10290) );
  AOI211_X1 U11464 ( .C1(n10384), .C2(n10290), .A(n10308), .B(n10289), .ZN(
        n10383) );
  AOI22_X1 U11465 ( .A1(n10553), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10291), 
        .B2(n10551), .ZN(n10292) );
  OAI21_X1 U11466 ( .B1(n10293), .B2(n10556), .A(n10292), .ZN(n10294) );
  AOI21_X1 U11467 ( .B1(n10383), .B2(n10548), .A(n10294), .ZN(n10295) );
  OAI211_X1 U11468 ( .C1(n10563), .C2(n10386), .A(n10296), .B(n10295), .ZN(
        P1_U3277) );
  INV_X1 U11469 ( .A(n10297), .ZN(n10304) );
  NAND2_X1 U11470 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  XOR2_X1 U11471 ( .A(n10305), .B(n10300), .Z(n10303) );
  OAI21_X1 U11472 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10390) );
  AOI21_X1 U11473 ( .B1(n10304), .B2(n10551), .A(n10390), .ZN(n10314) );
  XNOR2_X1 U11474 ( .A(n10306), .B(n10305), .ZN(n10452) );
  NAND2_X1 U11475 ( .A1(n10452), .A2(n10560), .ZN(n10313) );
  AOI211_X1 U11476 ( .C1(n10454), .C2(n10309), .A(n10308), .B(n10307), .ZN(
        n10389) );
  OAI22_X1 U11477 ( .A1(n10310), .A2(n10556), .B1(n5878), .B2(n8051), .ZN(
        n10311) );
  AOI21_X1 U11478 ( .B1(n10389), .B2(n10548), .A(n10311), .ZN(n10312) );
  OAI211_X1 U11479 ( .C1(n10553), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        P1_U3278) );
  INV_X1 U11480 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U11481 ( .A1(n10315), .A2(n10318), .ZN(n10395) );
  MUX2_X1 U11482 ( .A(n10316), .B(n10395), .S(n10643), .Z(n10317) );
  OAI21_X1 U11483 ( .B1(n10398), .B2(n10356), .A(n10317), .ZN(P1_U3553) );
  INV_X1 U11484 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10321) );
  AOI21_X1 U11485 ( .B1(n10320), .B2(n10319), .A(n10318), .ZN(n10399) );
  MUX2_X1 U11486 ( .A(n10321), .B(n10399), .S(n10643), .Z(n10322) );
  OAI21_X1 U11487 ( .B1(n4848), .B2(n10356), .A(n10322), .ZN(P1_U3552) );
  AOI21_X1 U11488 ( .B1(n10626), .B2(n10326), .A(n10325), .ZN(n10327) );
  NAND3_X1 U11489 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10402) );
  MUX2_X1 U11490 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10402), .S(n10643), .Z(
        P1_U3550) );
  NOR2_X1 U11491 ( .A1(n10331), .A2(n10330), .ZN(n10403) );
  MUX2_X1 U11492 ( .A(n10332), .B(n10403), .S(n10643), .Z(n10334) );
  NAND2_X1 U11493 ( .A1(n10406), .A2(n10392), .ZN(n10333) );
  OAI211_X1 U11494 ( .C1(n10408), .C2(n10381), .A(n10334), .B(n10333), .ZN(
        P1_U3548) );
  NAND2_X1 U11495 ( .A1(n10336), .A2(n10335), .ZN(n10409) );
  MUX2_X1 U11496 ( .A(n10409), .B(P1_REG1_REG_25__SCAN_IN), .S(n10641), .Z(
        n10337) );
  AOI21_X1 U11497 ( .B1(n10392), .B2(n10411), .A(n10337), .ZN(n10338) );
  OAI21_X1 U11498 ( .B1(n10413), .B2(n10381), .A(n10338), .ZN(P1_U3547) );
  INV_X1 U11499 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10342) );
  AOI211_X1 U11500 ( .C1(n10626), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        n10414) );
  MUX2_X1 U11501 ( .A(n10342), .B(n10414), .S(n10643), .Z(n10343) );
  OAI21_X1 U11502 ( .B1(n10417), .B2(n10381), .A(n10343), .ZN(P1_U3546) );
  OAI211_X1 U11503 ( .C1(n10346), .C2(n10617), .A(n10345), .B(n10344), .ZN(
        n10347) );
  NOR2_X1 U11504 ( .A1(n10348), .A2(n10347), .ZN(n10418) );
  MUX2_X1 U11505 ( .A(n10349), .B(n10418), .S(n10643), .Z(n10350) );
  OAI21_X1 U11506 ( .B1(n10421), .B2(n10381), .A(n10350), .ZN(P1_U3545) );
  AOI211_X1 U11507 ( .C1(n10353), .C2(n10622), .A(n10352), .B(n10351), .ZN(
        n10422) );
  MUX2_X1 U11508 ( .A(n10354), .B(n10422), .S(n10643), .Z(n10355) );
  OAI21_X1 U11509 ( .B1(n4942), .B2(n10356), .A(n10355), .ZN(P1_U3544) );
  INV_X1 U11510 ( .A(n10357), .ZN(n10359) );
  NAND2_X1 U11511 ( .A1(n10359), .A2(n10358), .ZN(n10426) );
  MUX2_X1 U11512 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10426), .S(n10643), .Z(
        n10360) );
  AOI21_X1 U11513 ( .B1(n10392), .B2(n10428), .A(n10360), .ZN(n10361) );
  OAI21_X1 U11514 ( .B1(n10430), .B2(n10381), .A(n10361), .ZN(P1_U3543) );
  INV_X1 U11515 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10365) );
  AOI211_X1 U11516 ( .C1(n10626), .C2(n10364), .A(n10363), .B(n10362), .ZN(
        n10431) );
  MUX2_X1 U11517 ( .A(n10365), .B(n10431), .S(n10643), .Z(n10366) );
  OAI21_X1 U11518 ( .B1(n10434), .B2(n10381), .A(n10366), .ZN(P1_U3542) );
  AOI211_X1 U11519 ( .C1(n10626), .C2(n10369), .A(n10368), .B(n10367), .ZN(
        n10435) );
  MUX2_X1 U11520 ( .A(n10370), .B(n10435), .S(n10643), .Z(n10371) );
  OAI21_X1 U11521 ( .B1(n10438), .B2(n10381), .A(n10371), .ZN(P1_U3541) );
  INV_X1 U11522 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10375) );
  AOI211_X1 U11523 ( .C1(n10626), .C2(n10374), .A(n10373), .B(n10372), .ZN(
        n10439) );
  MUX2_X1 U11524 ( .A(n10375), .B(n10439), .S(n10643), .Z(n10376) );
  OAI21_X1 U11525 ( .B1(n10442), .B2(n10381), .A(n10376), .ZN(P1_U3540) );
  AOI22_X1 U11526 ( .A1(n10443), .A2(n10392), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n10641), .ZN(n10380) );
  NAND2_X1 U11527 ( .A1(n10378), .A2(n10377), .ZN(n10444) );
  NAND2_X1 U11528 ( .A1(n10444), .A2(n10643), .ZN(n10379) );
  OAI211_X1 U11529 ( .C1(n10448), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        P1_U3539) );
  NAND2_X1 U11530 ( .A1(n10382), .A2(n10622), .ZN(n10387) );
  AOI21_X1 U11531 ( .B1(n10626), .B2(n10384), .A(n10383), .ZN(n10385) );
  OAI211_X1 U11532 ( .C1(n10388), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        n10450) );
  MUX2_X1 U11533 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10450), .S(n10643), .Z(
        P1_U3538) );
  NOR2_X1 U11534 ( .A1(n10390), .A2(n10389), .ZN(n10457) );
  NAND2_X1 U11535 ( .A1(n10452), .A2(n10391), .ZN(n10394) );
  AOI22_X1 U11536 ( .A1(n10454), .A2(n10392), .B1(P1_REG1_REG_15__SCAN_IN), 
        .B2(n10641), .ZN(n10393) );
  OAI211_X1 U11537 ( .C1(n10457), .C2(n10641), .A(n10394), .B(n10393), .ZN(
        P1_U3537) );
  MUX2_X1 U11538 ( .A(n10396), .B(n10395), .S(n10449), .Z(n10397) );
  OAI21_X1 U11539 ( .B1(n10398), .B2(n10425), .A(n10397), .ZN(P1_U3521) );
  MUX2_X1 U11540 ( .A(n10400), .B(n10399), .S(n10449), .Z(n10401) );
  OAI21_X1 U11541 ( .B1(n4848), .B2(n10425), .A(n10401), .ZN(P1_U3520) );
  MUX2_X1 U11542 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10402), .S(n10449), .Z(
        P1_U3518) );
  INV_X1 U11543 ( .A(n10403), .ZN(n10404) );
  MUX2_X1 U11544 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10404), .S(n10449), .Z(
        n10405) );
  AOI21_X1 U11545 ( .B1(n10453), .B2(n10406), .A(n10405), .ZN(n10407) );
  OAI21_X1 U11546 ( .B1(n10408), .B2(n10447), .A(n10407), .ZN(P1_U3516) );
  MUX2_X1 U11547 ( .A(n10409), .B(P1_REG0_REG_25__SCAN_IN), .S(n10634), .Z(
        n10410) );
  AOI21_X1 U11548 ( .B1(n10453), .B2(n10411), .A(n10410), .ZN(n10412) );
  OAI21_X1 U11549 ( .B1(n10413), .B2(n10447), .A(n10412), .ZN(P1_U3515) );
  MUX2_X1 U11550 ( .A(n10415), .B(n10414), .S(n10449), .Z(n10416) );
  OAI21_X1 U11551 ( .B1(n10417), .B2(n10447), .A(n10416), .ZN(P1_U3514) );
  INV_X1 U11552 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10419) );
  MUX2_X1 U11553 ( .A(n10419), .B(n10418), .S(n10449), .Z(n10420) );
  OAI21_X1 U11554 ( .B1(n10421), .B2(n10447), .A(n10420), .ZN(P1_U3513) );
  INV_X1 U11555 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10423) );
  MUX2_X1 U11556 ( .A(n10423), .B(n10422), .S(n10449), .Z(n10424) );
  OAI21_X1 U11557 ( .B1(n4942), .B2(n10425), .A(n10424), .ZN(P1_U3512) );
  MUX2_X1 U11558 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10426), .S(n10449), .Z(
        n10427) );
  AOI21_X1 U11559 ( .B1(n10453), .B2(n10428), .A(n10427), .ZN(n10429) );
  OAI21_X1 U11560 ( .B1(n10430), .B2(n10447), .A(n10429), .ZN(P1_U3511) );
  MUX2_X1 U11561 ( .A(n10432), .B(n10431), .S(n10449), .Z(n10433) );
  OAI21_X1 U11562 ( .B1(n10434), .B2(n10447), .A(n10433), .ZN(P1_U3510) );
  MUX2_X1 U11563 ( .A(n10436), .B(n10435), .S(n10449), .Z(n10437) );
  OAI21_X1 U11564 ( .B1(n10438), .B2(n10447), .A(n10437), .ZN(P1_U3509) );
  INV_X1 U11565 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10440) );
  MUX2_X1 U11566 ( .A(n10440), .B(n10439), .S(n10449), .Z(n10441) );
  OAI21_X1 U11567 ( .B1(n10442), .B2(n10447), .A(n10441), .ZN(P1_U3507) );
  AOI22_X1 U11568 ( .A1(n10443), .A2(n10453), .B1(P1_REG0_REG_17__SCAN_IN), 
        .B2(n10634), .ZN(n10446) );
  NAND2_X1 U11569 ( .A1(n10444), .A2(n10449), .ZN(n10445) );
  OAI211_X1 U11570 ( .C1(n10448), .C2(n10447), .A(n10446), .B(n10445), .ZN(
        P1_U3504) );
  MUX2_X1 U11571 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10450), .S(n10449), .Z(
        P1_U3501) );
  NAND2_X1 U11572 ( .A1(n10452), .A2(n10451), .ZN(n10456) );
  AOI22_X1 U11573 ( .A1(n10454), .A2(n10453), .B1(P1_REG0_REG_15__SCAN_IN), 
        .B2(n10634), .ZN(n10455) );
  OAI211_X1 U11574 ( .C1(n10457), .C2(n10634), .A(n10456), .B(n10455), .ZN(
        P1_U3498) );
  MUX2_X1 U11575 ( .A(n10459), .B(P1_D_REG_0__SCAN_IN), .S(n10458), .Z(
        P1_U3439) );
  NOR4_X1 U11576 ( .A1(n10462), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10461), .A4(
        P1_U3086), .ZN(n10463) );
  AOI21_X1 U11577 ( .B1(n10464), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10463), 
        .ZN(n10465) );
  OAI21_X1 U11578 ( .B1(n10466), .B2(n10472), .A(n10465), .ZN(P1_U3324) );
  OAI222_X1 U11579 ( .A1(n10470), .A2(n10469), .B1(n10472), .B2(n10468), .C1(
        n10467), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U11580 ( .A1(n10470), .A2(n10474), .B1(P1_U3086), .B2(n10473), 
        .C1(n10472), .C2(n10471), .ZN(P1_U3326) );
  MUX2_X1 U11581 ( .A(n10475), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11582 ( .A(n10476), .ZN(n10477) );
  AOI21_X1 U11583 ( .B1(n10541), .B2(n10478), .A(n10477), .ZN(n10479) );
  INV_X1 U11584 ( .A(n10479), .ZN(n10485) );
  NAND2_X1 U11585 ( .A1(n10481), .A2(n10482), .ZN(n10483) );
  AOI21_X1 U11586 ( .B1(n10480), .B2(n10483), .A(n10535), .ZN(n10484) );
  AOI211_X1 U11587 ( .C1(n10486), .C2(n10502), .A(n10485), .B(n10484), .ZN(
        n10487) );
  OAI21_X1 U11588 ( .B1(n10488), .B2(n10547), .A(n10487), .ZN(P1_U3217) );
  INV_X1 U11589 ( .A(n10489), .ZN(n10490) );
  OAI21_X1 U11590 ( .B1(n10492), .B2(n10491), .A(n10490), .ZN(n10501) );
  INV_X1 U11591 ( .A(n10495), .ZN(n10496) );
  NAND3_X1 U11592 ( .A1(n10494), .A2(n10497), .A3(n10496), .ZN(n10498) );
  AOI21_X1 U11593 ( .B1(n10499), .B2(n10498), .A(n10535), .ZN(n10500) );
  AOI211_X1 U11594 ( .C1(n10503), .C2(n10502), .A(n10501), .B(n10500), .ZN(
        n10504) );
  OAI21_X1 U11595 ( .B1(n10505), .B2(n10547), .A(n10504), .ZN(P1_U3224) );
  INV_X1 U11596 ( .A(n10506), .ZN(n10507) );
  AOI21_X1 U11597 ( .B1(n10541), .B2(n10508), .A(n10507), .ZN(n10509) );
  INV_X1 U11598 ( .A(n10509), .ZN(n10514) );
  INV_X1 U11599 ( .A(n10510), .ZN(n10511) );
  AOI21_X1 U11600 ( .B1(n10494), .B2(n10512), .A(n10535), .ZN(n10513) );
  AOI211_X1 U11601 ( .C1(n10625), .C2(n10515), .A(n10514), .B(n10513), .ZN(
        n10516) );
  OAI21_X1 U11602 ( .B1(n10517), .B2(n10547), .A(n10516), .ZN(P1_U3236) );
  XOR2_X1 U11603 ( .A(n10518), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11604 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11605 ( .B1(n10520), .B2(n10519), .A(n7737), .ZN(n10528) );
  INV_X1 U11606 ( .A(n10521), .ZN(n10522) );
  AOI21_X1 U11607 ( .B1(n10541), .B2(n10523), .A(n10522), .ZN(n10524) );
  OAI21_X1 U11608 ( .B1(n10525), .B2(n10543), .A(n10524), .ZN(n10526) );
  AOI21_X1 U11609 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(n10529) );
  OAI21_X1 U11610 ( .B1(n10530), .B2(n10547), .A(n10529), .ZN(P1_U3221) );
  INV_X1 U11611 ( .A(n10531), .ZN(n10532) );
  NAND3_X1 U11612 ( .A1(n10534), .A2(n10533), .A3(n10532), .ZN(n10537) );
  AOI21_X1 U11613 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(n10545) );
  INV_X1 U11614 ( .A(n10538), .ZN(n10539) );
  AOI21_X1 U11615 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(n10542) );
  OAI21_X1 U11616 ( .B1(n10557), .B2(n10543), .A(n10542), .ZN(n10544) );
  NOR2_X1 U11617 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  OAI21_X1 U11618 ( .B1(n10550), .B2(n10547), .A(n10546), .ZN(P1_U3239) );
  NAND2_X1 U11619 ( .A1(n10549), .A2(n10548), .ZN(n10555) );
  INV_X1 U11620 ( .A(n10550), .ZN(n10552) );
  AOI22_X1 U11621 ( .A1(n10553), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10552), 
        .B2(n10551), .ZN(n10554) );
  OAI211_X1 U11622 ( .C1(n10557), .C2(n10556), .A(n10555), .B(n10554), .ZN(
        n10558) );
  AOI21_X1 U11623 ( .B1(n10560), .B2(n10559), .A(n10558), .ZN(n10561) );
  OAI21_X1 U11624 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(P1_U3287) );
  NOR2_X1 U11625 ( .A1(n4550), .A2(n10564), .ZN(P1_U3294) );
  INV_X1 U11626 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U11627 ( .A1(n4550), .A2(n10566), .ZN(P1_U3295) );
  INV_X1 U11628 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10567) );
  NOR2_X1 U11629 ( .A1(n4550), .A2(n10567), .ZN(P1_U3296) );
  INV_X1 U11630 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U11631 ( .A1(n4550), .A2(n10568), .ZN(P1_U3297) );
  INV_X1 U11632 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U11633 ( .A1(n4550), .A2(n10569), .ZN(P1_U3298) );
  INV_X1 U11634 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U11635 ( .A1(n4550), .A2(n10570), .ZN(P1_U3299) );
  INV_X1 U11636 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U11637 ( .A1(n4550), .A2(n10571), .ZN(P1_U3300) );
  INV_X1 U11638 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U11639 ( .A1(n4550), .A2(n10572), .ZN(P1_U3301) );
  INV_X1 U11640 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10573) );
  NOR2_X1 U11641 ( .A1(n4550), .A2(n10573), .ZN(P1_U3302) );
  INV_X1 U11642 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10574) );
  NOR2_X1 U11643 ( .A1(n4550), .A2(n10574), .ZN(P1_U3303) );
  INV_X1 U11644 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U11645 ( .A1(n4550), .A2(n10575), .ZN(P1_U3304) );
  INV_X1 U11646 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U11647 ( .A1(n4550), .A2(n10576), .ZN(P1_U3305) );
  INV_X1 U11648 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10577) );
  NOR2_X1 U11649 ( .A1(n4550), .A2(n10577), .ZN(P1_U3306) );
  INV_X1 U11650 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10578) );
  NOR2_X1 U11651 ( .A1(n4550), .A2(n10578), .ZN(P1_U3307) );
  INV_X1 U11652 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10579) );
  NOR2_X1 U11653 ( .A1(n4550), .A2(n10579), .ZN(P1_U3308) );
  INV_X1 U11654 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10580) );
  NOR2_X1 U11655 ( .A1(n4550), .A2(n10580), .ZN(P1_U3309) );
  INV_X1 U11656 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10581) );
  NOR2_X1 U11657 ( .A1(n4550), .A2(n10581), .ZN(P1_U3310) );
  INV_X1 U11658 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10582) );
  NOR2_X1 U11659 ( .A1(n4550), .A2(n10582), .ZN(P1_U3311) );
  NOR2_X1 U11660 ( .A1(n4550), .A2(n10583), .ZN(P1_U3312) );
  NOR2_X1 U11661 ( .A1(n4550), .A2(n10584), .ZN(P1_U3313) );
  NOR2_X1 U11662 ( .A1(n4550), .A2(n10585), .ZN(P1_U3314) );
  NOR2_X1 U11663 ( .A1(n4550), .A2(n10586), .ZN(P1_U3315) );
  NOR2_X1 U11664 ( .A1(n4550), .A2(n10587), .ZN(P1_U3316) );
  INV_X1 U11665 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10588) );
  NOR2_X1 U11666 ( .A1(n4550), .A2(n10588), .ZN(P1_U3317) );
  INV_X1 U11667 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10589) );
  NOR2_X1 U11668 ( .A1(n4550), .A2(n10589), .ZN(P1_U3318) );
  INV_X1 U11669 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10590) );
  NOR2_X1 U11670 ( .A1(n4550), .A2(n10590), .ZN(P1_U3319) );
  INV_X1 U11671 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U11672 ( .A1(n4550), .A2(n10591), .ZN(P1_U3320) );
  NOR2_X1 U11673 ( .A1(n4550), .A2(n10592), .ZN(P1_U3321) );
  INV_X1 U11674 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10593) );
  NOR2_X1 U11675 ( .A1(n4550), .A2(n10593), .ZN(P1_U3322) );
  NOR2_X1 U11676 ( .A1(n4550), .A2(n10594), .ZN(P1_U3323) );
  AOI21_X1 U11677 ( .B1(n10626), .B2(n5897), .A(n10595), .ZN(n10596) );
  OAI21_X1 U11678 ( .B1(n10597), .B2(n10629), .A(n10596), .ZN(n10598) );
  AOI211_X1 U11679 ( .C1(n10633), .C2(n10600), .A(n10599), .B(n10598), .ZN(
        n10637) );
  AOI22_X1 U11680 ( .A1(n10449), .A2(n10637), .B1(n5403), .B2(n10634), .ZN(
        P1_U3456) );
  OAI21_X1 U11681 ( .B1(n10602), .B2(n10617), .A(n10601), .ZN(n10604) );
  AOI211_X1 U11682 ( .C1(n10622), .C2(n10605), .A(n10604), .B(n10603), .ZN(
        n10638) );
  INV_X1 U11683 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U11684 ( .A1(n10449), .A2(n10638), .B1(n10606), .B2(n10634), .ZN(
        P1_U3468) );
  INV_X1 U11685 ( .A(n10629), .ZN(n10611) );
  AND2_X1 U11686 ( .A1(n10607), .A2(n10626), .ZN(n10608) );
  OR2_X1 U11687 ( .A1(n10609), .A2(n10608), .ZN(n10610) );
  AOI21_X1 U11688 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10613) );
  INV_X1 U11689 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U11690 ( .A1(n10449), .A2(n10639), .B1(n10615), .B2(n10634), .ZN(
        P1_U3474) );
  OAI21_X1 U11691 ( .B1(n10618), .B2(n10617), .A(n10616), .ZN(n10620) );
  AOI211_X1 U11692 ( .C1(n10622), .C2(n10621), .A(n10620), .B(n10619), .ZN(
        n10640) );
  INV_X1 U11693 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U11694 ( .A1(n10449), .A2(n10640), .B1(n10623), .B2(n10634), .ZN(
        P1_U3480) );
  INV_X1 U11695 ( .A(n10632), .ZN(n10630) );
  AOI21_X1 U11696 ( .B1(n10626), .B2(n10625), .A(n10624), .ZN(n10627) );
  OAI211_X1 U11697 ( .C1(n10630), .C2(n10629), .A(n10628), .B(n10627), .ZN(
        n10631) );
  AOI21_X1 U11698 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(n10642) );
  INV_X1 U11699 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U11700 ( .A1(n10449), .A2(n10642), .B1(n10635), .B2(n10634), .ZN(
        P1_U3486) );
  AOI22_X1 U11701 ( .A1(n10643), .A2(n10637), .B1(n10636), .B2(n10641), .ZN(
        P1_U3523) );
  AOI22_X1 U11702 ( .A1(n10643), .A2(n10638), .B1(n6960), .B2(n10641), .ZN(
        P1_U3527) );
  AOI22_X1 U11703 ( .A1(n10643), .A2(n10639), .B1(n6997), .B2(n10641), .ZN(
        P1_U3529) );
  AOI22_X1 U11704 ( .A1(n10643), .A2(n10640), .B1(n7117), .B2(n10641), .ZN(
        P1_U3531) );
  AOI22_X1 U11705 ( .A1(n10643), .A2(n10642), .B1(n7352), .B2(n10641), .ZN(
        P1_U3533) );
  INV_X1 U11706 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10658) );
  OAI21_X1 U11707 ( .B1(n10646), .B2(n10645), .A(n10644), .ZN(n10647) );
  AOI22_X1 U11708 ( .A1(n10650), .A2(n10649), .B1(n10648), .B2(n10647), .ZN(
        n10656) );
  OAI211_X1 U11709 ( .C1(n10654), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        n10655) );
  OAI211_X1 U11710 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        n10659) );
  INV_X1 U11711 ( .A(n10659), .ZN(n10666) );
  OAI21_X1 U11712 ( .B1(n10662), .B2(n10661), .A(n10660), .ZN(n10663) );
  NAND2_X1 U11713 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  OAI211_X1 U11714 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6939), .A(n10666), .B(
        n10665), .ZN(P2_U3184) );
  INV_X1 U11715 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U11716 ( .A1(n10685), .A2(n10668), .B1(n10667), .B2(n10683), .ZN(
        P2_U3393) );
  AOI22_X1 U11717 ( .A1(n10685), .A2(n6254), .B1(n10669), .B2(n10683), .ZN(
        P2_U3396) );
  INV_X1 U11718 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U11719 ( .A1(n10685), .A2(n10671), .B1(n10670), .B2(n10683), .ZN(
        P2_U3399) );
  AOI22_X1 U11720 ( .A1(n10685), .A2(n6306), .B1(n10672), .B2(n10683), .ZN(
        P2_U3402) );
  INV_X1 U11721 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U11722 ( .A1(n10685), .A2(n10674), .B1(n10673), .B2(n10683), .ZN(
        P2_U3405) );
  INV_X1 U11723 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U11724 ( .A1(n10685), .A2(n10676), .B1(n10675), .B2(n10683), .ZN(
        P2_U3408) );
  AOI22_X1 U11725 ( .A1(n10685), .A2(n6356), .B1(n10677), .B2(n10683), .ZN(
        P2_U3411) );
  AOI22_X1 U11726 ( .A1(n10685), .A2(n6367), .B1(n10678), .B2(n10683), .ZN(
        P2_U3414) );
  INV_X1 U11727 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U11728 ( .A1(n10685), .A2(n10680), .B1(n10679), .B2(n10683), .ZN(
        P2_U3417) );
  AOI22_X1 U11729 ( .A1(n10685), .A2(n10682), .B1(n10681), .B2(n10683), .ZN(
        P2_U3420) );
  AOI22_X1 U11730 ( .A1(n10685), .A2(n6413), .B1(n10684), .B2(n10683), .ZN(
        P2_U3423) );
  INV_X1 U11731 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U11732 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  XOR2_X1 U11733 ( .A(n10690), .B(n10689), .Z(ADD_1068_U5) );
  XOR2_X1 U11734 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11735 ( .B1(n10693), .B2(n10692), .A(n10691), .ZN(ADD_1068_U55) );
  AOI21_X1 U11736 ( .B1(n10696), .B2(n10695), .A(n10694), .ZN(ADD_1068_U56) );
  AOI21_X1 U11737 ( .B1(n10699), .B2(n10698), .A(n10697), .ZN(ADD_1068_U57) );
  AOI21_X1 U11738 ( .B1(n10702), .B2(n10701), .A(n10700), .ZN(ADD_1068_U58) );
  AOI21_X1 U11739 ( .B1(n10705), .B2(n10704), .A(n10703), .ZN(ADD_1068_U59) );
  AOI21_X1 U11740 ( .B1(n10708), .B2(n10707), .A(n10706), .ZN(ADD_1068_U60) );
  OAI21_X1 U11741 ( .B1(n10711), .B2(n10710), .A(n10709), .ZN(n10713) );
  XNOR2_X1 U11742 ( .A(n10713), .B(n10712), .ZN(ADD_1068_U61) );
  XOR2_X1 U11743 ( .A(n10715), .B(n10714), .Z(ADD_1068_U62) );
  NOR2_X1 U11744 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  XNOR2_X1 U11745 ( .A(n10719), .B(n10718), .ZN(ADD_1068_U63) );
  XOR2_X1 U11746 ( .A(n10720), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11747 ( .A1(n10722), .A2(n10721), .ZN(n10723) );
  XOR2_X1 U11748 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10723), .Z(ADD_1068_U51) );
  AOI21_X1 U11749 ( .B1(n10726), .B2(n10725), .A(n10724), .ZN(ADD_1068_U47) );
  AOI21_X1 U11750 ( .B1(n10729), .B2(n10728), .A(n10727), .ZN(ADD_1068_U49) );
  AOI21_X1 U11751 ( .B1(n10732), .B2(n10731), .A(n10730), .ZN(ADD_1068_U48) );
  XOR2_X1 U11752 ( .A(n10734), .B(n10733), .Z(ADD_1068_U54) );
  XOR2_X1 U11753 ( .A(n10736), .B(n10735), .Z(ADD_1068_U53) );
  XNOR2_X1 U11754 ( .A(n10738), .B(n10737), .ZN(ADD_1068_U52) );
  INV_X1 U5103 ( .A(n6117), .ZN(n4542) );
  CLKBUF_X2 U5051 ( .A(n5936), .Z(n6112) );
  CLKBUF_X1 U5067 ( .A(n6110), .Z(n6115) );
  INV_X4 U5068 ( .A(n4542), .ZN(n4543) );
  CLKBUF_X1 U5070 ( .A(n9551), .Z(n4560) );
  CLKBUF_X1 U5104 ( .A(n5427), .Z(n4552) );
  CLKBUF_X1 U5125 ( .A(n7763), .Z(n4559) );
  CLKBUF_X1 U5143 ( .A(n5425), .Z(n5766) );
  CLKBUF_X1 U5199 ( .A(n5889), .Z(n6685) );
  CLKBUF_X1 U5203 ( .A(n9918), .Z(n4549) );
  CLKBUF_X1 U5252 ( .A(n6798), .Z(n4548) );
  CLKBUF_X2 U6148 ( .A(n5822), .Z(n9938) );
  CLKBUF_X2 U6572 ( .A(n6721), .Z(n4554) );
endmodule

