

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4295, n4296, n4297, n4298, n4299, n4300, n4302, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066;

  NAND2_X2 U4801 ( .A1(n8658), .A2(n8902), .ZN(n8981) );
  INV_X1 U4802 ( .A(n9052), .ZN(n9213) );
  NAND2_X1 U4803 ( .A1(n4838), .A2(n4836), .ZN(n7071) );
  INV_X1 U4804 ( .A(n9377), .ZN(n9165) );
  INV_X1 U4806 ( .A(n5548), .ZN(n5602) );
  CLKBUF_X2 U4807 ( .A(n5789), .Z(n6589) );
  INV_X2 U4808 ( .A(n5744), .ZN(n6103) );
  NAND2_X4 U4809 ( .A1(n6299), .A2(n4942), .ZN(n5550) );
  INV_X1 U4810 ( .A(n6756), .ZN(n6755) );
  NOR2_X1 U4811 ( .A1(n7232), .A2(n5615), .ZN(n4900) );
  NAND2_X1 U4812 ( .A1(n4881), .A2(n4862), .ZN(n5062) );
  CLKBUF_X1 U4813 ( .A(n8499), .Z(n4295) );
  OAI21_X1 U4814 ( .B1(n5648), .B2(n9534), .A(n9602), .ZN(n8499) );
  INV_X2 U4815 ( .A(n4982), .ZN(n5567) );
  NAND2_X1 U4816 ( .A1(n6430), .A2(n6605), .ZN(n6433) );
  OAI21_X1 U4817 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5470) );
  CLKBUF_X2 U4818 ( .A(n5739), .Z(n7622) );
  NAND2_X1 U4819 ( .A1(n6055), .A2(n6056), .ZN(n6068) );
  OAI21_X1 U4820 ( .B1(n7725), .B2(n7724), .A(n7723), .ZN(n7722) );
  CLKBUF_X2 U4821 ( .A(n5891), .Z(n4307) );
  INV_X1 U4822 ( .A(n7588), .ZN(n7389) );
  INV_X1 U4823 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5904) );
  CLKBUF_X2 U4824 ( .A(n5548), .Z(n4297) );
  INV_X1 U4825 ( .A(n8620), .ZN(n5372) );
  AND2_X1 U4826 ( .A1(n5593), .A2(n5592), .ZN(n8974) );
  INV_X1 U4827 ( .A(n9032), .ZN(n9204) );
  NAND2_X1 U4828 ( .A1(n8649), .A2(n8667), .ZN(n9156) );
  INV_X1 U4829 ( .A(n6796), .ZN(n9637) );
  AND4_X1 U4830 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n8119)
         );
  INV_X1 U4831 ( .A(n9096), .ZN(n9228) );
  NAND2_X1 U4832 ( .A1(n5299), .A2(n5298), .ZN(n9244) );
  INV_X1 U4833 ( .A(n9194), .ZN(n9004) );
  AOI21_X1 U4834 ( .B1(n8977), .B2(n8981), .A(n8948), .ZN(n8963) );
  OR2_X1 U4835 ( .A1(n7525), .A2(n7527), .ZN(n4296) );
  XNOR2_X1 U4836 ( .A(n4904), .B(n4903), .ZN(n8873) );
  INV_X4 U4837 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5794) );
  NAND2_X2 U4839 ( .A1(n8287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  NOR2_X2 U4840 ( .A1(n5996), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5721) );
  XNOR2_X2 U4842 ( .A(n4998), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9350) );
  XNOR2_X2 U4843 ( .A(n4407), .B(n4406), .ZN(n7804) );
  OR2_X2 U4844 ( .A1(n7803), .A2(n4386), .ZN(n4407) );
  OAI22_X2 U4845 ( .A1(n7955), .A2(n6215), .B1(n6110), .B2(n7738), .ZN(n7945)
         );
  NAND2_X2 U4846 ( .A1(n4823), .A2(n4822), .ZN(n7955) );
  OAI21_X2 U4847 ( .B1(n8050), .B2(n7559), .A(n7557), .ZN(n8035) );
  NOR2_X2 U4848 ( .A1(n7765), .A2(n7764), .ZN(n7774) );
  XNOR2_X2 U4849 ( .A(n7773), .B(n7789), .ZN(n7765) );
  XNOR2_X2 U4850 ( .A(n5689), .B(n5688), .ZN(n6155) );
  BUF_X8 U4851 ( .A(n4975), .Z(n4298) );
  NOR2_X2 U4852 ( .A1(n6850), .A2(n4400), .ZN(n9758) );
  NOR2_X2 U4853 ( .A1(n6461), .A2(n6470), .ZN(n6850) );
  NAND2_X1 U4854 ( .A1(n8616), .A2(n8615), .ZN(n9172) );
  NAND2_X1 U4855 ( .A1(n6255), .A2(n7500), .ZN(n7984) );
  AOI21_X1 U4856 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n8595) );
  NAND2_X1 U4857 ( .A1(n6228), .A2(n6227), .ZN(n6286) );
  OAI21_X1 U4858 ( .B1(n8018), .B2(n6252), .A(n7487), .ZN(n8006) );
  NAND2_X1 U4859 ( .A1(n4568), .A2(n7480), .ZN(n8018) );
  XNOR2_X1 U4860 ( .A(n7360), .B(SI_29_), .ZN(n8602) );
  AND2_X1 U4861 ( .A1(n5538), .A2(n5537), .ZN(n9194) );
  NAND2_X1 U4862 ( .A1(n5694), .A2(n5693), .ZN(n8213) );
  AND2_X1 U4863 ( .A1(n8898), .A2(n8680), .ZN(n9023) );
  XNOR2_X1 U4864 ( .A(n7655), .B(n7979), .ZN(n7972) );
  NAND2_X1 U4865 ( .A1(n6763), .A2(n7566), .ZN(n6874) );
  OAI21_X1 U4866 ( .B1(n6811), .B2(n7404), .A(n7414), .ZN(n6763) );
  AND2_X1 U4867 ( .A1(n4674), .A2(n4672), .ZN(n4671) );
  OR2_X1 U4868 ( .A1(n8910), .A2(n7195), .ZN(n8663) );
  AND2_X1 U4869 ( .A1(n4563), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7029) );
  OAI21_X1 U4870 ( .B1(n5235), .B2(n4807), .A(n4805), .ZN(n5283) );
  INV_X1 U4871 ( .A(n6919), .ZN(n9655) );
  INV_X16 U4872 ( .A(n9138), .ZN(n9616) );
  NAND2_X1 U4873 ( .A1(n7412), .A2(n7409), .ZN(n7561) );
  INV_X1 U4874 ( .A(n9837), .ZN(n6966) );
  NOR2_X2 U4875 ( .A1(n6751), .A2(n6755), .ZN(n6780) );
  AND2_X1 U4876 ( .A1(n6431), .A2(n6433), .ZN(n6607) );
  XNOR2_X1 U4877 ( .A(n5704), .B(n5703), .ZN(n7277) );
  AOI21_X1 U4878 ( .B1(n6433), .B2(n4559), .A(n4391), .ZN(n4558) );
  INV_X1 U4879 ( .A(n6188), .ZN(n4595) );
  NAND2_X1 U4880 ( .A1(n5701), .A2(n5702), .ZN(n5712) );
  NAND2_X1 U4881 ( .A1(n5702), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  INV_X2 U4882 ( .A(n5550), .ZN(n4943) );
  INV_X1 U4883 ( .A(n5891), .ZN(n4306) );
  CLKBUF_X1 U4885 ( .A(n8873), .Z(n4305) );
  XNOR2_X1 U4886 ( .A(n5677), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U4887 ( .A1(n8708), .A2(n6955), .ZN(n6749) );
  OAI21_X1 U4888 ( .B1(n4905), .B2(n4312), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4915) );
  OR2_X1 U4889 ( .A1(n4905), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4906) );
  INV_X2 U4890 ( .A(n4298), .ZN(n8613) );
  NAND2_X2 U4891 ( .A1(n5771), .A2(n5770), .ZN(n6411) );
  XNOR2_X1 U4892 ( .A(n5827), .B(n5826), .ZN(n6459) );
  CLKBUF_X1 U4893 ( .A(n8799), .Z(n4300) );
  INV_X1 U4894 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5665) );
  XNOR2_X1 U4895 ( .A(n7548), .B(n7526), .ZN(n7931) );
  NAND2_X1 U4896 ( .A1(n8366), .A2(n5556), .ZN(n8494) );
  AOI21_X1 U4897 ( .B1(n4435), .B2(n4336), .A(n4429), .ZN(n4428) );
  NAND2_X1 U4898 ( .A1(n8627), .A2(n8881), .ZN(n8767) );
  INV_X1 U4899 ( .A(n9172), .ZN(n8627) );
  NAND2_X1 U4900 ( .A1(n7545), .A2(n7544), .ZN(n8203) );
  NAND2_X1 U4901 ( .A1(n8611), .A2(n8610), .ZN(n8876) );
  NOR2_X1 U4902 ( .A1(n4549), .A2(n4546), .ZN(n4545) );
  AND2_X1 U4903 ( .A1(n4554), .A2(n4553), .ZN(n4549) );
  AOI21_X1 U4904 ( .B1(n4575), .B2(n4577), .A(n7935), .ZN(n4573) );
  AOI21_X1 U4905 ( .B1(n4359), .B2(n4746), .A(n4744), .ZN(n4743) );
  NAND2_X2 U4906 ( .A1(n5566), .A2(n5565), .ZN(n9190) );
  XNOR2_X1 U4907 ( .A(n6222), .B(n6221), .ZN(n7600) );
  NAND2_X1 U4908 ( .A1(n6099), .A2(n6098), .ZN(n8219) );
  NAND2_X1 U4909 ( .A1(n8937), .A2(n8936), .ZN(n9035) );
  INV_X1 U4910 ( .A(n4779), .ZN(n6222) );
  NAND2_X1 U4911 ( .A1(n6085), .A2(n6084), .ZN(n7655) );
  XNOR2_X1 U4912 ( .A(n5558), .B(n5557), .ZN(n8299) );
  OR2_X1 U4913 ( .A1(n9204), .A2(n8940), .ZN(n8898) );
  NAND2_X1 U4914 ( .A1(n6070), .A2(n6069), .ZN(n8226) );
  NAND2_X1 U4915 ( .A1(n5473), .A2(n5472), .ZN(n9209) );
  OR2_X1 U4916 ( .A1(n9213), .A2(n8934), .ZN(n9036) );
  OR2_X1 U4917 ( .A1(n8553), .A2(n8612), .ZN(n4489) );
  NAND2_X1 U4918 ( .A1(n5728), .A2(n5727), .ZN(n7997) );
  OR4_X1 U4919 ( .A1(n9066), .A2(n9101), .A3(n9113), .A4(n8652), .ZN(n8653) );
  AOI21_X1 U4920 ( .B1(n4585), .B2(n4584), .A(n4583), .ZN(n4582) );
  AND2_X1 U4921 ( .A1(n4608), .A2(n7458), .ZN(n4606) );
  NAND2_X1 U4922 ( .A1(n5407), .A2(n5406), .ZN(n9223) );
  AND2_X1 U4923 ( .A1(n4609), .A2(n7459), .ZN(n4608) );
  AND2_X1 U4924 ( .A1(n5390), .A2(n5389), .ZN(n9096) );
  NAND2_X1 U4925 ( .A1(n6011), .A2(n6010), .ZN(n8255) );
  AOI21_X1 U4926 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8833), .A(n9465), .ZN(
        n8822) );
  NAND2_X1 U4927 ( .A1(n4530), .A2(n4330), .ZN(n9510) );
  NAND2_X1 U4928 ( .A1(n6971), .A2(n6975), .ZN(n7061) );
  OAI21_X1 U4929 ( .B1(n5405), .B2(n5404), .A(n5403), .ZN(n5420) );
  OR2_X1 U4930 ( .A1(n9239), .A2(n8560), .ZN(n9109) );
  OR2_X1 U4931 ( .A1(n7196), .A2(n4534), .ZN(n4530) );
  NAND2_X1 U4932 ( .A1(n5985), .A2(n5984), .ZN(n8179) );
  NAND2_X1 U4933 ( .A1(n5999), .A2(n5998), .ZN(n8261) );
  AOI21_X1 U4934 ( .B1(n4671), .B2(n4676), .A(n4669), .ZN(n4668) );
  NAND2_X1 U4935 ( .A1(n4784), .A2(n5386), .ZN(n5405) );
  NAND2_X1 U4936 ( .A1(n6243), .A2(n7412), .ZN(n6811) );
  AOI21_X1 U4937 ( .B1(n4536), .B2(n4533), .A(n4532), .ZN(n4531) );
  AND2_X1 U4938 ( .A1(n9155), .A2(n8550), .ZN(n9511) );
  AND2_X1 U4939 ( .A1(n8911), .A2(n4537), .ZN(n4536) );
  OR2_X1 U4940 ( .A1(n9520), .A2(n8543), .ZN(n9155) );
  AOI21_X1 U4941 ( .B1(n4677), .B2(n4675), .A(n5155), .ZN(n4674) );
  NAND2_X1 U4942 ( .A1(n5938), .A2(n5937), .ZN(n8110) );
  NAND2_X1 U4943 ( .A1(n5268), .A2(n5267), .ZN(n9520) );
  NAND2_X1 U4944 ( .A1(n5955), .A2(n5954), .ZN(n8279) );
  AND2_X1 U4945 ( .A1(n4763), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U4946 ( .A1(n5218), .A2(n5217), .ZN(n8910) );
  AND2_X1 U4947 ( .A1(n5151), .A2(n4327), .ZN(n4677) );
  NAND2_X1 U4948 ( .A1(n6685), .A2(n5033), .ZN(n6716) );
  NAND2_X1 U4949 ( .A1(n5210), .A2(n5209), .ZN(n5235) );
  NAND2_X1 U4950 ( .A1(n6788), .A2(n6787), .ZN(n6893) );
  NAND2_X1 U4951 ( .A1(n7386), .A2(n6179), .ZN(n6728) );
  NAND2_X1 U4952 ( .A1(n4544), .A2(n4542), .ZN(n8431) );
  XNOR2_X1 U4953 ( .A(n4440), .B(n5187), .ZN(n6340) );
  INV_X1 U4954 ( .A(n6920), .ZN(n9662) );
  NAND2_X1 U4955 ( .A1(n4851), .A2(n9783), .ZN(n7391) );
  NAND2_X1 U4956 ( .A1(n6440), .A2(n4403), .ZN(n6604) );
  NAND4_X1 U4957 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n7751)
         );
  NAND4_X1 U4958 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n6751)
         );
  NAND4_X1 U4959 ( .A1(n4967), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n8791)
         );
  AND2_X2 U4960 ( .A1(n7596), .A2(n7389), .ZN(n7519) );
  CLKBUF_X1 U4961 ( .A(n5131), .Z(n5642) );
  NAND2_X1 U4962 ( .A1(n8873), .A2(n8769), .ZN(n6509) );
  INV_X2 U4963 ( .A(n4992), .ZN(n4723) );
  INV_X2 U4964 ( .A(n5131), .ZN(n5594) );
  NAND2_X1 U4965 ( .A1(n5065), .A2(n5064), .ZN(n4515) );
  CLKBUF_X3 U4966 ( .A(n5741), .Z(n6594) );
  NAND2_X1 U4967 ( .A1(n5716), .A2(n6132), .ZN(n7588) );
  AND2_X2 U4968 ( .A1(n9306), .A2(n4937), .ZN(n5040) );
  AND2_X2 U4969 ( .A1(n4936), .A2(n4937), .ZN(n8620) );
  CLKBUF_X1 U4970 ( .A(n4999), .Z(n8603) );
  XNOR2_X1 U4971 ( .A(n5720), .B(n5719), .ZN(n7586) );
  CLKBUF_X1 U4972 ( .A(n5120), .Z(n5387) );
  NAND2_X1 U4973 ( .A1(n4639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U4974 ( .A1(n6394), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U4975 ( .A1(n5369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4904) );
  OR2_X1 U4976 ( .A1(n6393), .A2(n6494), .ZN(n6394) );
  NAND2_X1 U4977 ( .A1(n5640), .A2(n6540), .ZN(n4952) );
  BUF_X4 U4978 ( .A(n6155), .Z(n6156) );
  NAND2_X1 U4979 ( .A1(n4895), .A2(n4898), .ZN(n7232) );
  AOI21_X1 U4980 ( .B1(n5087), .B2(n4419), .A(n4358), .ZN(n4418) );
  XNOR2_X1 U4981 ( .A(n5622), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8769) );
  MUX2_X1 U4982 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4892), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4895) );
  AOI21_X1 U4983 ( .B1(n4413), .B2(n5019), .A(n4357), .ZN(n4412) );
  XNOR2_X1 U4984 ( .A(n4916), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6540) );
  XNOR2_X1 U4985 ( .A(n4934), .B(n4933), .ZN(n4936) );
  OAI21_X1 U4986 ( .B1(n4934), .B2(n4924), .A(P1_IR_REG_30__SCAN_IN), .ZN(
        n4932) );
  XNOR2_X1 U4987 ( .A(n4915), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5620) );
  OR2_X1 U4988 ( .A1(n6502), .A2(n5740), .ZN(n6500) );
  NOR2_X1 U4989 ( .A1(n4774), .A2(n4772), .ZN(n4771) );
  NOR2_X1 U4990 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  AND2_X1 U4991 ( .A1(n4887), .A2(n4888), .ZN(n4773) );
  AND2_X1 U4992 ( .A1(n5665), .A2(n5805), .ZN(n4570) );
  NAND2_X1 U4993 ( .A1(n6682), .A2(n4918), .ZN(n4411) );
  AND2_X1 U4994 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6682) );
  INV_X1 U4995 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4903) );
  INV_X1 U4996 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4516) );
  NOR3_X1 U4997 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n4889) );
  INV_X4 U4998 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4999 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4918) );
  NOR2_X1 U5000 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4884) );
  NOR2_X1 U5001 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4883) );
  NOR2_X1 U5002 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4882) );
  INV_X1 U5003 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4887) );
  INV_X1 U5004 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5016) );
  OR2_X1 U5005 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4890) );
  INV_X1 U5006 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6129) );
  INV_X1 U5007 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5723) );
  INV_X1 U5008 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5948) );
  INV_X1 U5009 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5951) );
  INV_X1 U5010 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5914) );
  INV_X1 U5011 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5699) );
  INV_X1 U5012 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5859) );
  INV_X4 U5013 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AND2_X1 U5014 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4924) );
  NAND2_X1 U5015 ( .A1(n7071), .A2(n6202), .ZN(n7206) );
  NAND2_X1 U5016 ( .A1(n5736), .A2(n5665), .ZN(n5770) );
  INV_X2 U5017 ( .A(n5772), .ZN(n7542) );
  OR2_X1 U5018 ( .A1(n5772), .A2(n6317), .ZN(n4850) );
  OAI22_X1 U5019 ( .A1(n7936), .A2(n6220), .B1(n7524), .B2(n7528), .ZN(n6235)
         );
  OAI22_X2 U5020 ( .A1(n8001), .A2(n8005), .B1(n8159), .B2(n7741), .ZN(n7991)
         );
  NOR2_X2 U5021 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  NOR2_X2 U5022 ( .A1(n6621), .A2(n6620), .ZN(n6619) );
  AND2_X2 U5023 ( .A1(n4411), .A2(n4410), .ZN(n4975) );
  NOR2_X2 U5024 ( .A1(n9756), .A2(n4404), .ZN(n7027) );
  XNOR2_X2 U5025 ( .A(n4978), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6646) );
  NAND2_X2 U5026 ( .A1(n6194), .A2(n6193), .ZN(n6816) );
  NAND2_X1 U5027 ( .A1(n4911), .A2(n6299), .ZN(n4299) );
  INV_X4 U5028 ( .A(n5601), .ZN(n5551) );
  OR2_X1 U5029 ( .A1(n5679), .A2(n5904), .ZN(n5677) );
  NOR2_X2 U5030 ( .A1(n7030), .A2(n7029), .ZN(n7033) );
  XNOR2_X1 U5031 ( .A(n4493), .B(P1_IR_REG_1__SCAN_IN), .ZN(n8799) );
  OAI21_X2 U5032 ( .B1(n8615), .B2(n6526), .A(n4920), .ZN(n6756) );
  BUF_X1 U5033 ( .A(n5695), .Z(n5996) );
  NAND2_X2 U5034 ( .A1(n7391), .A2(n7390), .ZN(n7386) );
  INV_X1 U5036 ( .A(n4298), .ZN(n4302) );
  OR2_X1 U5037 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  NAND3_X1 U5038 ( .A1(n6749), .A2(n6299), .A3(n6509), .ZN(n5548) );
  NAND2_X2 U5039 ( .A1(n8873), .A2(n6955), .ZN(n5626) );
  OR2_X1 U5040 ( .A1(n5707), .A2(n5904), .ZN(n5689) );
  INV_X2 U5041 ( .A(n6178), .ZN(n4851) );
  AND4_X4 U5042 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(n6178)
         );
  NOR2_X2 U5044 ( .A1(n5838), .A2(n5670), .ZN(n5980) );
  OAI21_X2 U5045 ( .B1(n7206), .B2(n4854), .A(n4852), .ZN(n7280) );
  NAND2_X1 U5046 ( .A1(n5681), .A2(n5682), .ZN(n5891) );
  AOI22_X2 U5047 ( .A1(n8014), .A2(n8017), .B1(n8004), .B2(n7639), .ZN(n8001)
         );
  NAND2_X1 U5048 ( .A1(n6383), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5049 ( .A1(n4719), .A2(n4322), .ZN(n4715) );
  AOI21_X1 U5050 ( .B1(n4311), .B2(n4737), .A(n4736), .ZN(n4735) );
  NOR2_X1 U5051 ( .A1(n9228), .A2(n8926), .ZN(n4736) );
  NOR2_X1 U5052 ( .A1(n4740), .A2(n8927), .ZN(n4737) );
  NAND2_X1 U5053 ( .A1(n8600), .A2(n8601), .ZN(n4486) );
  INV_X1 U5054 ( .A(n8599), .ZN(n4485) );
  INV_X1 U5055 ( .A(n4781), .ZN(n4780) );
  OAI21_X1 U5056 ( .B1(n5589), .B2(n4782), .A(n6221), .ZN(n4781) );
  AND2_X1 U5057 ( .A1(n7522), .A2(n7532), .ZN(n4809) );
  INV_X1 U5058 ( .A(n4803), .ZN(n4798) );
  INV_X1 U5059 ( .A(n5309), .ZN(n5293) );
  NAND2_X1 U5060 ( .A1(n7632), .A2(n6052), .ZN(n6055) );
  AND2_X1 U5061 ( .A1(n7533), .A2(n7532), .ZN(n7549) );
  OR2_X1 U5062 ( .A1(n6442), .A2(n6421), .ZN(n4865) );
  INV_X1 U5063 ( .A(n6425), .ZN(n4722) );
  INV_X1 U5064 ( .A(n9760), .ZN(n4693) );
  INV_X1 U5065 ( .A(n6832), .ZN(n4694) );
  NAND2_X1 U5066 ( .A1(n4589), .A2(n4594), .ZN(n7402) );
  NAND2_X1 U5067 ( .A1(n5756), .A2(n5681), .ZN(n5789) );
  NOR2_X1 U5068 ( .A1(n4831), .A2(n4828), .ZN(n4827) );
  NOR2_X1 U5069 ( .A1(n4332), .A2(n4835), .ZN(n4831) );
  INV_X1 U5070 ( .A(n4833), .ZN(n4828) );
  OR2_X1 U5071 ( .A1(n7991), .A2(n4829), .ZN(n4825) );
  INV_X1 U5072 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5671) );
  INV_X1 U5073 ( .A(n7060), .ZN(n4675) );
  AND2_X1 U5074 ( .A1(n9143), .A2(n8667), .ZN(n4541) );
  NAND2_X1 U5075 ( .A1(n9675), .A2(n7116), .ZN(n4768) );
  OR2_X1 U5076 ( .A1(n9190), .A2(n8596), .ZN(n8658) );
  AND2_X1 U5077 ( .A1(n4751), .A2(n4353), .ZN(n4749) );
  INV_X1 U5078 ( .A(n8780), .ZN(n8920) );
  INV_X1 U5079 ( .A(n4815), .ZN(n4814) );
  INV_X1 U5080 ( .A(n4773), .ZN(n4772) );
  NAND2_X1 U5081 ( .A1(n4889), .A2(n4775), .ZN(n4774) );
  INV_X1 U5082 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U5083 ( .A1(n4787), .A2(n4786), .ZN(n4785) );
  INV_X1 U5084 ( .A(n5360), .ZN(n4786) );
  NOR2_X1 U5085 ( .A1(n5141), .A2(n4792), .ZN(n4791) );
  INV_X1 U5086 ( .A(n5109), .ZN(n4792) );
  AND2_X1 U5087 ( .A1(n5158), .A2(n5119), .ZN(n5156) );
  AND2_X1 U5088 ( .A1(n7675), .A2(n4866), .ZN(n6081) );
  OR2_X1 U5089 ( .A1(n7603), .A2(n8003), .ZN(n4866) );
  AND2_X1 U5090 ( .A1(n6093), .A2(n6092), .ZN(n7509) );
  INV_X1 U5091 ( .A(n4307), .ZN(n6229) );
  OAI211_X1 U5092 ( .C1(n5771), .C2(n5777), .A(n4686), .B(n4685), .ZN(n9740)
         );
  NAND2_X1 U5093 ( .A1(n4687), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4686) );
  OAI211_X1 U5094 ( .C1(n6456), .C2(n4718), .A(n4716), .B(n4714), .ZN(n6457)
         );
  NAND2_X1 U5095 ( .A1(n4715), .A2(n6852), .ZN(n4714) );
  NAND2_X1 U5096 ( .A1(n4718), .A2(n4339), .ZN(n4716) );
  NAND2_X1 U5097 ( .A1(n4395), .A2(n4380), .ZN(n4700) );
  NAND2_X1 U5098 ( .A1(n7791), .A2(n4702), .ZN(n4701) );
  INV_X1 U5099 ( .A(n7793), .ZN(n4702) );
  INV_X1 U5100 ( .A(n7835), .ZN(n4406) );
  AND2_X1 U5101 ( .A1(n4846), .A2(n4338), .ZN(n4845) );
  NAND2_X1 U5102 ( .A1(n6874), .A2(n7427), .ZN(n6246) );
  INV_X1 U5103 ( .A(n4844), .ZN(n4843) );
  AND2_X1 U5104 ( .A1(n6276), .A2(n6275), .ZN(n6704) );
  OR2_X1 U5105 ( .A1(n7991), .A2(n6214), .ZN(n4832) );
  INV_X1 U5106 ( .A(n7543), .ZN(n6020) );
  AND2_X1 U5107 ( .A1(n6267), .A2(n7519), .ZN(n8096) );
  INV_X1 U5108 ( .A(n4655), .ZN(n4654) );
  OAI21_X1 U5109 ( .B1(n8357), .B2(n4656), .A(n5458), .ZN(n4655) );
  INV_X1 U5110 ( .A(n5439), .ZN(n4656) );
  AND2_X1 U5111 ( .A1(n8769), .A2(n8708), .ZN(n8697) );
  INV_X1 U5112 ( .A(n5040), .ZN(n5476) );
  NAND2_X1 U5114 ( .A1(n4935), .A2(n4936), .ZN(n5131) );
  OAI21_X1 U5115 ( .B1(n6893), .B2(n4487), .A(n8712), .ZN(n9576) );
  INV_X1 U5116 ( .A(n6894), .ZN(n4487) );
  OR2_X1 U5117 ( .A1(n9213), .A2(n8935), .ZN(n8936) );
  NAND2_X1 U5118 ( .A1(n9048), .A2(n4876), .ZN(n8937) );
  INV_X1 U5119 ( .A(n8927), .ZN(n4738) );
  NOR2_X1 U5120 ( .A1(n4741), .A2(n8924), .ZN(n4740) );
  NOR2_X1 U5121 ( .A1(n9124), .A2(n4742), .ZN(n4741) );
  AND2_X1 U5122 ( .A1(n8630), .A2(n8768), .ZN(n9596) );
  INV_X1 U5123 ( .A(n6378), .ZN(n6303) );
  NAND2_X1 U5124 ( .A1(n4817), .A2(n7583), .ZN(n7546) );
  NAND2_X1 U5125 ( .A1(n4443), .A2(n7535), .ZN(n4442) );
  NAND2_X1 U5126 ( .A1(n7434), .A2(n7519), .ZN(n4441) );
  NAND2_X1 U5127 ( .A1(n4427), .A2(n7535), .ZN(n4426) );
  NOR2_X1 U5128 ( .A1(n4472), .A2(n4471), .ZN(n4470) );
  INV_X1 U5129 ( .A(n8728), .ZN(n4472) );
  NAND2_X1 U5130 ( .A1(n8540), .A2(n8612), .ZN(n4471) );
  NAND2_X1 U5131 ( .A1(n7467), .A2(n7468), .ZN(n7475) );
  NAND2_X1 U5132 ( .A1(n4780), .A2(n4782), .ZN(n4778) );
  NAND2_X1 U5133 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  NAND2_X1 U5134 ( .A1(n4482), .A2(n8607), .ZN(n8625) );
  NAND2_X1 U5135 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  OAI211_X1 U5136 ( .C1(n8598), .C2(n8597), .A(n4486), .B(n4485), .ZN(n4484)
         );
  NAND2_X1 U5137 ( .A1(n8646), .A2(n8537), .ZN(n4537) );
  NAND2_X1 U5138 ( .A1(n4492), .A2(n4871), .ZN(n4491) );
  INV_X1 U5139 ( .A(n4890), .ZN(n4492) );
  INV_X1 U5140 ( .A(n5385), .ZN(n4787) );
  NAND2_X1 U5141 ( .A1(n4808), .A2(n5258), .ZN(n4807) );
  NAND2_X1 U5142 ( .A1(n5234), .A2(n5233), .ZN(n4808) );
  INV_X1 U5143 ( .A(n5158), .ZN(n4796) );
  INV_X1 U5144 ( .A(SI_11_), .ZN(n5163) );
  NAND2_X1 U5145 ( .A1(n4418), .A2(n4420), .ZN(n4417) );
  OAI21_X1 U5146 ( .B1(n4431), .B2(n4430), .A(n4428), .ZN(n4819) );
  NAND2_X1 U5147 ( .A1(n4435), .A2(n4432), .ZN(n4430) );
  NAND2_X1 U5148 ( .A1(n6411), .A2(n9946), .ZN(n4405) );
  NOR2_X1 U5149 ( .A1(n4712), .A2(n6852), .ZN(n4711) );
  NAND2_X1 U5150 ( .A1(n4718), .A2(n4717), .ZN(n4713) );
  INV_X1 U5151 ( .A(n4715), .ZN(n4717) );
  AND2_X1 U5152 ( .A1(n6854), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4404) );
  NOR2_X1 U5153 ( .A1(n7133), .A2(n4408), .ZN(n7135) );
  AND2_X1 U5154 ( .A1(n7134), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5155 ( .A1(n6024), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5156 ( .A1(n4855), .A2(n6205), .ZN(n4854) );
  NOR2_X1 U5157 ( .A1(n5845), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5844) );
  OR2_X1 U5158 ( .A1(n8226), .A2(n7993), .ZN(n7502) );
  OR2_X1 U5159 ( .A1(n8249), .A2(n7717), .ZN(n7478) );
  INV_X1 U5160 ( .A(n4611), .ZN(n4604) );
  OR2_X1 U5161 ( .A1(n8261), .A2(n7338), .ZN(n7471) );
  AOI21_X1 U5162 ( .B1(n4618), .B2(n7568), .A(n4616), .ZN(n4615) );
  INV_X1 U5163 ( .A(n7436), .ZN(n4616) );
  NAND2_X1 U5164 ( .A1(n5763), .A2(n6730), .ZN(n7388) );
  INV_X1 U5165 ( .A(n7277), .ZN(n6128) );
  INV_X1 U5166 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5688) );
  NOR2_X1 U5167 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4641) );
  OR2_X1 U5168 ( .A1(n5874), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5903) );
  INV_X1 U5169 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5666) );
  INV_X1 U5170 ( .A(n4319), .ZN(n4651) );
  NAND2_X1 U5171 ( .A1(n8625), .A2(n8876), .ZN(n4481) );
  OR2_X1 U5172 ( .A1(n8876), .A2(n8612), .ZN(n4480) );
  INV_X1 U5173 ( .A(n4937), .ZN(n4935) );
  INV_X1 U5174 ( .A(n8964), .ZN(n4554) );
  INV_X1 U5175 ( .A(n8981), .ZN(n4551) );
  OR2_X1 U5176 ( .A1(n7119), .A2(n8473), .ZN(n4451) );
  AND2_X1 U5177 ( .A1(n8634), .A2(n8744), .ZN(n8674) );
  INV_X1 U5178 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4913) );
  INV_X1 U5179 ( .A(n5591), .ZN(n4782) );
  AND2_X1 U5180 ( .A1(n5591), .A2(n5564), .ZN(n5589) );
  AND2_X1 U5181 ( .A1(n5559), .A2(n5536), .ZN(n5557) );
  INV_X1 U5182 ( .A(n5532), .ZN(n4816) );
  AND2_X1 U5183 ( .A1(n5532), .A2(n5518), .ZN(n5530) );
  INV_X1 U5184 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4893) );
  INV_X1 U5185 ( .A(n4491), .ZN(n4457) );
  INV_X1 U5186 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5624) );
  INV_X1 U5187 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5621) );
  INV_X1 U5188 ( .A(n4800), .ZN(n4799) );
  AOI21_X1 U5189 ( .B1(n4798), .B2(n4800), .A(n4356), .ZN(n4797) );
  NOR2_X1 U5190 ( .A1(n4801), .A2(n5338), .ZN(n4800) );
  INV_X1 U5191 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5291) );
  INV_X1 U5192 ( .A(SI_14_), .ZN(n5287) );
  INV_X1 U5193 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U5194 ( .A1(n7337), .A2(n7336), .ZN(n4587) );
  NAND2_X1 U5195 ( .A1(n7086), .A2(n4341), .ZN(n7239) );
  NAND2_X1 U5196 ( .A1(n6058), .A2(n6057), .ZN(n4638) );
  NAND2_X1 U5197 ( .A1(n4587), .A2(n4585), .ZN(n7709) );
  NAND2_X1 U5198 ( .A1(n4581), .A2(n4334), .ZN(n7713) );
  NAND2_X1 U5199 ( .A1(n4582), .A2(n4586), .ZN(n4580) );
  NOR2_X1 U5200 ( .A1(n4350), .A2(n4624), .ZN(n4623) );
  INV_X1 U5201 ( .A(n4626), .ZN(n4624) );
  OR2_X1 U5202 ( .A1(n6283), .A2(n6280), .ZN(n6168) );
  AOI21_X1 U5203 ( .B1(n4869), .B2(n7588), .A(n7586), .ZN(n7587) );
  AND4_X1 U5204 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n6989)
         );
  NAND2_X1 U5205 ( .A1(n5800), .A2(n5802), .ZN(n4593) );
  NAND2_X1 U5206 ( .A1(n6381), .A2(n4688), .ZN(n4690) );
  NOR2_X1 U5207 ( .A1(n4689), .A2(n6499), .ZN(n4688) );
  AOI21_X1 U5208 ( .B1(n4690), .B2(n6382), .A(n9740), .ZN(n9739) );
  AND2_X1 U5209 ( .A1(n6385), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U5210 ( .A1(n6386), .A2(n6385), .ZN(n4697) );
  NAND2_X1 U5211 ( .A1(n4567), .A2(n6395), .ZN(n6429) );
  NAND2_X1 U5212 ( .A1(n6458), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6833) );
  AND2_X1 U5213 ( .A1(n5903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5875) );
  AND3_X1 U5214 ( .A1(n4691), .A2(n4692), .A3(n4384), .ZN(n7010) );
  OR2_X1 U5215 ( .A1(n7138), .A2(n7137), .ZN(n4561) );
  NAND2_X1 U5216 ( .A1(n4396), .A2(n4381), .ZN(n4706) );
  INV_X1 U5217 ( .A(n7158), .ZN(n4396) );
  NAND2_X1 U5218 ( .A1(n7128), .A2(n4708), .ZN(n4707) );
  INV_X1 U5219 ( .A(n7129), .ZN(n4708) );
  OR2_X1 U5220 ( .A1(n7754), .A2(n7755), .ZN(n4705) );
  AND3_X1 U5221 ( .A1(n4701), .A2(n4703), .A3(n4700), .ZN(n7834) );
  OR2_X1 U5222 ( .A1(n7848), .A2(n7847), .ZN(n7882) );
  NAND2_X1 U5223 ( .A1(n7375), .A2(n4872), .ZN(n7531) );
  NAND2_X1 U5224 ( .A1(n8609), .A2(n7542), .ZN(n7375) );
  AND2_X1 U5225 ( .A1(n8025), .A2(n4363), .ZN(n4848) );
  OR2_X1 U5226 ( .A1(n8037), .A2(n8036), .ZN(n4849) );
  AND4_X1 U5227 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n7345)
         );
  INV_X1 U5228 ( .A(n7388), .ZN(n6726) );
  OR3_X1 U5229 ( .A1(n6280), .A2(n6279), .A3(n6278), .ZN(n6705) );
  OR2_X1 U5230 ( .A1(n7944), .A2(n7516), .ZN(n4577) );
  INV_X1 U5231 ( .A(n4576), .ZN(n4575) );
  OAI21_X1 U5232 ( .B1(n4578), .B2(n4577), .A(n7521), .ZN(n4576) );
  NOR2_X1 U5233 ( .A1(n7515), .A2(n4579), .ZN(n4578) );
  INV_X1 U5234 ( .A(n7510), .ZN(n4579) );
  XNOR2_X1 U5235 ( .A(n8213), .B(n7732), .ZN(n7944) );
  OR2_X1 U5236 ( .A1(n7515), .A2(n7516), .ZN(n7954) );
  AOI21_X1 U5237 ( .B1(n4824), .B2(n4829), .A(n4355), .ZN(n4822) );
  INV_X1 U5238 ( .A(n7954), .ZN(n7952) );
  NAND2_X1 U5239 ( .A1(n4825), .A2(n4826), .ZN(n7962) );
  INV_X1 U5240 ( .A(n4827), .ZN(n4826) );
  AND2_X1 U5241 ( .A1(n7504), .A2(n7502), .ZN(n7985) );
  NAND2_X1 U5242 ( .A1(n6045), .A2(n6044), .ZN(n8163) );
  AND3_X1 U5243 ( .A1(n6038), .A2(n6037), .A3(n6036), .ZN(n8042) );
  INV_X1 U5244 ( .A(n8096), .ZN(n8120) );
  NAND2_X1 U5245 ( .A1(n7519), .A2(n6266), .ZN(n8118) );
  AND2_X1 U5246 ( .A1(n7478), .A2(n7477), .ZN(n8036) );
  NOR2_X1 U5247 ( .A1(n6250), .A2(n7450), .ZN(n4611) );
  NOR2_X1 U5248 ( .A1(n7425), .A2(n4619), .ZN(n4618) );
  INV_X1 U5249 ( .A(n7426), .ZN(n4619) );
  NAND2_X1 U5250 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  INV_X1 U5251 ( .A(n6935), .ZN(n4622) );
  AND2_X1 U5252 ( .A1(n5879), .A2(n5878), .ZN(n9819) );
  OR2_X1 U5253 ( .A1(n6237), .A2(n6136), .ZN(n6287) );
  AND2_X1 U5254 ( .A1(n6131), .A2(n8285), .ZN(n6290) );
  NAND2_X1 U5255 ( .A1(n6114), .A2(n6113), .ZN(n6273) );
  NAND2_X1 U5256 ( .A1(n5676), .A2(n4860), .ZN(n4859) );
  INV_X1 U5257 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4860) );
  NAND2_X1 U5258 ( .A1(n5698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U5259 ( .A1(n5700), .A2(n5699), .ZN(n5702) );
  NAND2_X1 U5260 ( .A1(n5717), .A2(n4641), .ZN(n6132) );
  INV_X1 U5261 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5719) );
  XNOR2_X1 U5262 ( .A(n5725), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7896) );
  OR2_X1 U5263 ( .A1(n5858), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5874) );
  CLKBUF_X1 U5264 ( .A(n5838), .Z(n5858) );
  NAND2_X1 U5265 ( .A1(n5666), .A2(n5794), .ZN(n4857) );
  INV_X1 U5266 ( .A(n5769), .ZN(n5771) );
  NAND2_X1 U5267 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5768) );
  NAND2_X1 U5268 ( .A1(n5904), .A2(n5665), .ZN(n5767) );
  NAND2_X1 U5269 ( .A1(n5738), .A2(n5737), .ZN(n6380) );
  INV_X1 U5270 ( .A(n4663), .ZN(n4662) );
  OAI21_X1 U5271 ( .B1(n4666), .B2(n4664), .A(n8480), .ZN(n4663) );
  INV_X1 U5272 ( .A(n4665), .ZN(n4664) );
  AND2_X1 U5273 ( .A1(n5581), .A2(n5580), .ZN(n5631) );
  INV_X1 U5274 ( .A(n4677), .ZN(n4676) );
  INV_X1 U5275 ( .A(n5204), .ZN(n4672) );
  NAND2_X1 U5276 ( .A1(n4646), .A2(n4651), .ZN(n4650) );
  INV_X1 U5277 ( .A(n6716), .ZN(n4646) );
  NAND2_X1 U5278 ( .A1(n4651), .A2(n4649), .ZN(n4648) );
  INV_X1 U5279 ( .A(n5037), .ZN(n4649) );
  NAND2_X1 U5280 ( .A1(n8356), .A2(n8357), .ZN(n8355) );
  INV_X1 U5281 ( .A(n8457), .ZN(n5460) );
  INV_X1 U5282 ( .A(n8935), .ZN(n8934) );
  XNOR2_X1 U5283 ( .A(n4679), .B(n5602), .ZN(n4984) );
  OAI21_X1 U5284 ( .B1(n4982), .B2(n9629), .A(n4983), .ZN(n4679) );
  OR2_X1 U5285 ( .A1(n8398), .A2(n8399), .ZN(n4665) );
  AND2_X1 U5286 ( .A1(n8697), .A2(n5626), .ZN(n6515) );
  NAND2_X1 U5287 ( .A1(n4361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5622) );
  INV_X1 U5288 ( .A(n6955), .ZN(n8756) );
  NAND2_X1 U5289 ( .A1(n8758), .A2(n8757), .ZN(n8760) );
  AND2_X1 U5290 ( .A1(n5575), .A2(n5574), .ZN(n8596) );
  AND2_X1 U5291 ( .A1(n5547), .A2(n5546), .ZN(n8945) );
  NAND2_X1 U5292 ( .A1(n9340), .A2(n6529), .ZN(n4506) );
  NAND2_X1 U5293 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  INV_X1 U5294 ( .A(n9394), .ZN(n4503) );
  NAND2_X1 U5295 ( .A1(n4506), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U5296 ( .A1(n9350), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5297 ( .A1(n8805), .A2(n8806), .ZN(n8804) );
  OR2_X1 U5298 ( .A1(n9318), .A2(n9317), .ZN(n4497) );
  OR2_X1 U5299 ( .A1(n5569), .A2(n5568), .ZN(n5641) );
  OR2_X1 U5300 ( .A1(n9199), .A2(n8944), .ZN(n8992) );
  NAND2_X1 U5301 ( .A1(n5451), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5474) );
  INV_X1 U5302 ( .A(n5410), .ZN(n5408) );
  INV_X1 U5303 ( .A(n4539), .ZN(n4538) );
  OAI21_X1 U5304 ( .B1(n4541), .B2(n4540), .A(n9134), .ZN(n4539) );
  INV_X1 U5305 ( .A(n8669), .ZN(n4540) );
  NAND2_X1 U5306 ( .A1(n8668), .A2(n4541), .ZN(n9142) );
  OAI21_X1 U5307 ( .B1(n9507), .B2(n9511), .A(n8916), .ZN(n9154) );
  NAND2_X1 U5308 ( .A1(n9522), .A2(n9706), .ZN(n9523) );
  INV_X2 U5309 ( .A(n5000), .ZN(n8608) );
  NAND2_X1 U5310 ( .A1(n4766), .A2(n4768), .ZN(n4763) );
  OAI21_X1 U5311 ( .B1(n9544), .B2(n4767), .A(n7117), .ZN(n4766) );
  NAND2_X1 U5312 ( .A1(n7047), .A2(n4768), .ZN(n4764) );
  INV_X1 U5313 ( .A(n9596), .ZN(n9579) );
  NAND2_X1 U5314 ( .A1(n9179), .A2(n9621), .ZN(n9181) );
  INV_X1 U5315 ( .A(n8974), .ZN(n9186) );
  INV_X1 U5316 ( .A(n4749), .ZN(n4748) );
  AOI21_X1 U5317 ( .B1(n4749), .B2(n4747), .A(n4352), .ZN(n4746) );
  INV_X1 U5318 ( .A(n4754), .ZN(n4747) );
  INV_X1 U5319 ( .A(n4752), .ZN(n4751) );
  OAI21_X1 U5320 ( .B1(n8942), .B2(n4753), .A(n4755), .ZN(n4752) );
  NAND2_X1 U5321 ( .A1(n9032), .A2(n8940), .ZN(n4755) );
  NAND2_X1 U5322 ( .A1(n4756), .A2(n4318), .ZN(n4753) );
  NOR2_X1 U5323 ( .A1(n8942), .A2(n4757), .ZN(n4754) );
  AOI21_X1 U5324 ( .B1(n4309), .B2(n4731), .A(n4362), .ZN(n4730) );
  INV_X1 U5325 ( .A(n8674), .ZN(n9101) );
  NAND2_X1 U5326 ( .A1(n4740), .A2(n4742), .ZN(n4739) );
  INV_X1 U5327 ( .A(n8431), .ZN(n9675) );
  NAND2_X1 U5328 ( .A1(n9508), .A2(n9627), .ZN(n9702) );
  NAND2_X1 U5329 ( .A1(n5617), .A2(n5620), .ZN(n6337) );
  XNOR2_X1 U5330 ( .A(n5590), .B(n5589), .ZN(n7380) );
  XNOR2_X1 U5331 ( .A(n5157), .B(n5156), .ZN(n6332) );
  NAND2_X1 U5332 ( .A1(n5051), .A2(n5050), .ZN(n5065) );
  AND2_X1 U5333 ( .A1(n5045), .A2(n5018), .ZN(n6552) );
  AND4_X1 U5334 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n7090)
         );
  OR2_X1 U5335 ( .A1(n6863), .A2(n6802), .ZN(n5821) );
  INV_X1 U5336 ( .A(n7102), .ZN(n7596) );
  AND2_X1 U5337 ( .A1(n6597), .A2(n6596), .ZN(n7551) );
  NAND2_X1 U5338 ( .A1(n5687), .A2(n5686), .ZN(n7956) );
  INV_X1 U5339 ( .A(n7509), .ZN(n7979) );
  NAND2_X1 U5340 ( .A1(n5734), .A2(n5733), .ZN(n7980) );
  NAND2_X1 U5341 ( .A1(n6480), .A2(n4329), .ZN(n6440) );
  NAND2_X1 U5342 ( .A1(n6473), .A2(n6472), .ZN(n6841) );
  AND2_X1 U5343 ( .A1(n5953), .A2(n5962), .ZN(n7797) );
  NAND2_X1 U5344 ( .A1(n7891), .A2(n7904), .ZN(n4682) );
  INV_X1 U5345 ( .A(n7890), .ZN(n4683) );
  OR2_X1 U5346 ( .A1(n6583), .A2(n7906), .ZN(n9769) );
  INV_X1 U5347 ( .A(n7531), .ZN(n9368) );
  NAND2_X1 U5348 ( .A1(n4439), .A2(n5899), .ZN(n7294) );
  NAND2_X1 U5349 ( .A1(n6340), .A2(n7542), .ZN(n4439) );
  NAND2_X1 U5350 ( .A1(n6269), .A2(n6268), .ZN(n4636) );
  OAI21_X1 U5351 ( .B1(n4636), .B2(n4630), .A(n4634), .ZN(n4629) );
  NAND2_X1 U5352 ( .A1(n9886), .A2(n9893), .ZN(n4634) );
  NAND2_X1 U5353 ( .A1(n9884), .A2(n9841), .ZN(n4630) );
  NAND2_X1 U5354 ( .A1(n4644), .A2(n4642), .ZN(n8307) );
  NAND2_X1 U5355 ( .A1(n5588), .A2(n4643), .ZN(n4642) );
  NAND2_X1 U5356 ( .A1(n8365), .A2(n4645), .ZN(n4644) );
  INV_X1 U5357 ( .A(n5556), .ZN(n4643) );
  NOR2_X2 U5358 ( .A1(n5648), .A2(n5627), .ZN(n8495) );
  OR2_X1 U5359 ( .A1(n5479), .A2(n5478), .ZN(n8938) );
  OR2_X1 U5360 ( .A1(n5352), .A2(n5351), .ZN(n8921) );
  NAND2_X1 U5361 ( .A1(n8869), .A2(n4401), .ZN(n4511) );
  INV_X1 U5362 ( .A(n4402), .ZN(n4401) );
  OAI21_X1 U5363 ( .B1(n8870), .B2(n9479), .A(n9501), .ZN(n4402) );
  NAND2_X1 U5364 ( .A1(n4547), .A2(n4545), .ZN(n8904) );
  INV_X1 U5365 ( .A(n9244), .ZN(n9150) );
  OAI211_X1 U5366 ( .C1(n8615), .C2(n6307), .A(n5006), .B(n5005), .ZN(n6796)
         );
  OR2_X1 U5367 ( .A1(n5000), .A2(n6317), .ZN(n4955) );
  INV_X1 U5368 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5369 ( .A1(n7437), .A2(n7440), .ZN(n4427) );
  NAND2_X1 U5370 ( .A1(n4425), .A2(n4424), .ZN(n4423) );
  NOR2_X1 U5371 ( .A1(n4613), .A2(n7535), .ZN(n4424) );
  NAND2_X1 U5372 ( .A1(n7442), .A2(n7441), .ZN(n4425) );
  NAND2_X1 U5373 ( .A1(n4421), .A2(n4337), .ZN(n7454) );
  NAND2_X1 U5374 ( .A1(n4474), .A2(n4473), .ZN(n8549) );
  AOI21_X1 U5375 ( .B1(n8541), .B2(n4470), .A(n4469), .ZN(n4473) );
  NOR2_X1 U5376 ( .A1(n8663), .A2(n8766), .ZN(n4469) );
  OAI21_X1 U5377 ( .B1(n7475), .B2(n7470), .A(n7519), .ZN(n4444) );
  NAND2_X1 U5378 ( .A1(n4488), .A2(n9134), .ZN(n8566) );
  NAND2_X1 U5379 ( .A1(n4479), .A2(n8633), .ZN(n4478) );
  NAND2_X1 U5380 ( .A1(n8581), .A2(n8580), .ZN(n4479) );
  OR2_X1 U5381 ( .A1(n4313), .A2(n8645), .ZN(n8721) );
  NOR2_X1 U5382 ( .A1(n7528), .A2(n4437), .ZN(n4434) );
  INV_X1 U5383 ( .A(n7533), .ZN(n4429) );
  NAND2_X1 U5384 ( .A1(n4433), .A2(n7528), .ZN(n4432) );
  INV_X1 U5385 ( .A(n4436), .ZN(n4433) );
  NAND2_X1 U5386 ( .A1(n7685), .A2(n7993), .ZN(n4833) );
  NOR2_X1 U5387 ( .A1(n9204), .A2(n4454), .ZN(n4453) );
  INV_X1 U5388 ( .A(n4455), .ZN(n4454) );
  NOR2_X1 U5389 ( .A1(n9209), .A2(n9213), .ZN(n4455) );
  INV_X1 U5390 ( .A(n8926), .ZN(n8925) );
  AOI21_X1 U5391 ( .B1(n5590), .B2(n4780), .A(n4777), .ZN(n4776) );
  NAND2_X1 U5392 ( .A1(n4778), .A2(n6225), .ZN(n4777) );
  NOR2_X1 U5393 ( .A1(n4812), .A2(n4816), .ZN(n4811) );
  INV_X1 U5394 ( .A(n5514), .ZN(n4812) );
  OAI21_X1 U5395 ( .B1(n5530), .B2(n4816), .A(n5557), .ZN(n4815) );
  NOR2_X1 U5396 ( .A1(n4790), .A2(n4382), .ZN(n4789) );
  INV_X1 U5397 ( .A(n5423), .ZN(n4790) );
  INV_X1 U5398 ( .A(n5294), .ZN(n4801) );
  INV_X1 U5399 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5340) );
  INV_X1 U5400 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5162) );
  INV_X1 U5401 ( .A(n7336), .ZN(n4584) );
  AND2_X1 U5402 ( .A1(n6086), .A2(n5661), .ZN(n5663) );
  AND2_X1 U5403 ( .A1(n6071), .A2(n9949), .ZN(n6086) );
  AND2_X1 U5404 ( .A1(n5966), .A2(n5659), .ZN(n5986) );
  NOR2_X1 U5405 ( .A1(n5967), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5966) );
  OR2_X1 U5406 ( .A1(n5908), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5920) );
  AND2_X1 U5407 ( .A1(n8286), .A2(n6115), .ZN(n6706) );
  NOR2_X1 U5408 ( .A1(n6112), .A2(n6125), .ZN(n6280) );
  NOR2_X1 U5409 ( .A1(n4827), .A2(n7972), .ZN(n4824) );
  NAND2_X1 U5410 ( .A1(n4833), .A2(n4830), .ZN(n4829) );
  INV_X1 U5411 ( .A(n6214), .ZN(n4830) );
  OR2_X1 U5412 ( .A1(n8163), .A2(n8004), .ZN(n7487) );
  INV_X1 U5413 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9915) );
  AND2_X1 U5414 ( .A1(n4641), .A2(n6133), .ZN(n4640) );
  INV_X1 U5415 ( .A(n4857), .ZN(n4856) );
  AND2_X1 U5416 ( .A1(n5504), .A2(n5503), .ZN(n5506) );
  AOI21_X1 U5417 ( .B1(n9321), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9313), .ZN(
        n9435) );
  NAND2_X1 U5418 ( .A1(n8974), .A2(n4465), .ZN(n4464) );
  OR2_X1 U5419 ( .A1(n4464), .A2(n9179), .ZN(n4463) );
  NAND2_X1 U5420 ( .A1(n9102), .A2(n8674), .ZN(n4528) );
  NAND2_X1 U5421 ( .A1(n9377), .A2(n9150), .ZN(n4461) );
  OR2_X1 U5422 ( .A1(n9239), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U5423 ( .A1(n4313), .A2(n4522), .ZN(n4520) );
  INV_X1 U5424 ( .A(n8786), .ZN(n7043) );
  AND2_X1 U5425 ( .A1(n9071), .A2(n4452), .ZN(n9013) );
  AND2_X1 U5426 ( .A1(n4453), .A2(n9018), .ZN(n4452) );
  NAND2_X1 U5427 ( .A1(n9071), .A2(n4453), .ZN(n9027) );
  INV_X1 U5428 ( .A(n4316), .ZN(n4731) );
  INV_X1 U5429 ( .A(n8537), .ZN(n4533) );
  INV_X1 U5430 ( .A(n8663), .ZN(n4532) );
  INV_X1 U5431 ( .A(n4536), .ZN(n4534) );
  NAND2_X1 U5432 ( .A1(n7371), .A2(n7370), .ZN(n7537) );
  XNOR2_X1 U5433 ( .A(n7363), .B(n7362), .ZN(n7360) );
  NAND2_X1 U5434 ( .A1(n5491), .A2(n5490), .ZN(n5513) );
  AND2_X1 U5435 ( .A1(n5514), .A2(n5495), .ZN(n5512) );
  INV_X1 U5436 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4901) );
  AND2_X1 U5437 ( .A1(n5386), .A2(n5365), .ZN(n5385) );
  NOR2_X1 U5438 ( .A1(n5292), .A2(n4804), .ZN(n4803) );
  INV_X1 U5439 ( .A(n5289), .ZN(n4804) );
  INV_X1 U5440 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4888) );
  INV_X1 U5441 ( .A(n4806), .ZN(n4805) );
  OAI21_X1 U5442 ( .B1(n4807), .B2(n5233), .A(n5261), .ZN(n4806) );
  NAND2_X1 U5443 ( .A1(n4794), .A2(n5161), .ZN(n5205) );
  NOR2_X1 U5444 ( .A1(n5186), .A2(n4796), .ZN(n4795) );
  INV_X1 U5445 ( .A(n5087), .ZN(n4420) );
  INV_X1 U5446 ( .A(n5068), .ZN(n4419) );
  OAI21_X1 U5447 ( .B1(n4298), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4409), .ZN(
        n4971) );
  INV_X1 U5448 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4917) );
  XNOR2_X1 U5449 ( .A(n6180), .B(n5739), .ZN(n5750) );
  INV_X1 U5450 ( .A(n4600), .ZN(n4599) );
  OAI21_X1 U5451 ( .B1(n6043), .B2(n4601), .A(n7631), .ZN(n4600) );
  AOI21_X1 U5452 ( .B1(n4627), .B2(n5932), .A(n4333), .ZN(n4626) );
  XNOR2_X1 U5453 ( .A(n5739), .B(n8128), .ZN(n5782) );
  NAND2_X1 U5454 ( .A1(n4819), .A2(n7519), .ZN(n4818) );
  INV_X1 U5455 ( .A(n6594), .ZN(n6230) );
  AND4_X1 U5456 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n7338)
         );
  NAND2_X1 U5457 ( .A1(n4698), .A2(n6384), .ZN(n6485) );
  NAND2_X1 U5458 ( .A1(n4565), .A2(n6396), .ZN(n6486) );
  INV_X1 U5459 ( .A(n4566), .ZN(n4565) );
  INV_X1 U5460 ( .A(n6424), .ZN(n4720) );
  NAND2_X1 U5461 ( .A1(n4722), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4721) );
  OR2_X1 U5462 ( .A1(n6608), .A2(n6443), .ZN(n6609) );
  NAND2_X1 U5463 ( .A1(n4393), .A2(n4392), .ZN(n6431) );
  NAND2_X1 U5464 ( .A1(n6607), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5465 ( .A1(n4691), .A2(n4692), .ZN(n9759) );
  AND2_X1 U5466 ( .A1(n6833), .A2(n6832), .ZN(n9761) );
  XNOR2_X1 U5467 ( .A(n7027), .B(n6855), .ZN(n4563) );
  AND3_X1 U5468 ( .A1(n4707), .A2(n4388), .A3(n4706), .ZN(n7788) );
  NAND2_X1 U5469 ( .A1(n7763), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4560) );
  NOR2_X1 U5470 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  OR2_X1 U5471 ( .A1(n6300), .A2(n7220), .ZN(n6399) );
  AOI21_X1 U5472 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n7853), .A(n7850), .ZN(
        n7867) );
  NOR2_X1 U5473 ( .A1(n7886), .A2(n7885), .ZN(n7889) );
  INV_X1 U5474 ( .A(n7882), .ZN(n7883) );
  INV_X1 U5475 ( .A(n6156), .ZN(n7906) );
  INV_X1 U5476 ( .A(n7378), .ZN(n7926) );
  OR2_X1 U5477 ( .A1(n6146), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7378) );
  OR2_X1 U5478 ( .A1(n6061), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U5479 ( .A1(n6033), .A2(n5660), .ZN(n6059) );
  NAND2_X1 U5480 ( .A1(n5986), .A2(n9915), .ZN(n6012) );
  OR2_X1 U5481 ( .A1(n6012), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6024) );
  INV_X1 U5482 ( .A(n4853), .ZN(n4852) );
  OAI21_X1 U5483 ( .B1(n4854), .B2(n6203), .A(n6206), .ZN(n4853) );
  NAND2_X1 U5484 ( .A1(n4620), .A2(n7426), .ZN(n6998) );
  INV_X1 U5485 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U5486 ( .A1(n6816), .A2(n6195), .ZN(n6765) );
  OR2_X1 U5487 ( .A1(n5831), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5845) );
  INV_X1 U5488 ( .A(n4591), .ZN(n4590) );
  OAI21_X1 U5489 ( .B1(n4594), .B2(n6188), .A(n4592), .ZN(n4591) );
  AND2_X1 U5490 ( .A1(n7896), .A2(n7586), .ZN(n8129) );
  OR2_X1 U5491 ( .A1(n7556), .A2(n7555), .ZN(n7990) );
  NAND2_X1 U5492 ( .A1(n6032), .A2(n6031), .ZN(n7686) );
  AOI21_X1 U5493 ( .B1(n4606), .B2(n4604), .A(n4603), .ZN(n4602) );
  INV_X1 U5494 ( .A(n4606), .ZN(n4605) );
  INV_X1 U5495 ( .A(n7462), .ZN(n4603) );
  AOI21_X1 U5496 ( .B1(n4615), .B2(n4617), .A(n4613), .ZN(n4612) );
  INV_X1 U5497 ( .A(n4615), .ZN(n4614) );
  INV_X1 U5498 ( .A(n4618), .ZN(n4617) );
  NOR2_X1 U5499 ( .A1(n7069), .A2(n4837), .ZN(n4836) );
  INV_X1 U5500 ( .A(n6201), .ZN(n4837) );
  NAND2_X1 U5501 ( .A1(n7519), .A2(n6153), .ZN(n6288) );
  NOR2_X1 U5502 ( .A1(n6168), .A2(n6278), .ZN(n6292) );
  INV_X1 U5503 ( .A(n5676), .ZN(n4858) );
  INV_X1 U5504 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5982) );
  OR2_X1 U5505 ( .A1(n5935), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5936) );
  NOR2_X1 U5506 ( .A1(n5903), .A2(n5902), .ZN(n5915) );
  NAND2_X1 U5507 ( .A1(n5666), .A2(n4687), .ZN(n5785) );
  AND2_X1 U5508 ( .A1(n5588), .A2(n8367), .ZN(n4645) );
  OAI21_X1 U5509 ( .B1(n4982), .B2(n8707), .A(n4958), .ZN(n4959) );
  NOR2_X1 U5510 ( .A1(n4982), .A2(n6755), .ZN(n4947) );
  OR2_X1 U5511 ( .A1(n5498), .A2(n8415), .ZN(n5523) );
  AND2_X1 U5512 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5038) );
  AND2_X1 U5513 ( .A1(n4678), .A2(n4327), .ZN(n8422) );
  NAND2_X1 U5514 ( .A1(n7061), .A2(n7060), .ZN(n4678) );
  INV_X1 U5515 ( .A(n8908), .ZN(n8484) );
  NAND2_X1 U5516 ( .A1(n4673), .A2(n4674), .ZN(n8465) );
  OR2_X1 U5517 ( .A1(n7061), .A2(n4676), .ZN(n4673) );
  INV_X1 U5518 ( .A(n8878), .ZN(n8505) );
  OAI21_X1 U5519 ( .B1(n6619), .B2(n6630), .A(n6629), .ZN(n6628) );
  AND2_X1 U5520 ( .A1(n5333), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5521 ( .A1(n4481), .A2(n4480), .ZN(n8626) );
  NOR4_X1 U5522 ( .A1(n8964), .A2(n8981), .A3(n8996), .A4(n8655), .ZN(n8656)
         );
  NAND2_X1 U5523 ( .A1(n4723), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U5524 ( .A1(n8798), .A2(n8797), .ZN(n8796) );
  NOR2_X1 U5525 ( .A1(n9345), .A2(n6549), .ZN(n9390) );
  NAND2_X1 U5526 ( .A1(n6552), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4501) );
  AOI21_X1 U5527 ( .B1(n6555), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9405), .ZN(
        n9424) );
  AOI21_X1 U5528 ( .B1(n6560), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9329), .ZN(
        n9355) );
  NOR2_X1 U5529 ( .A1(n9325), .A2(n4377), .ZN(n9359) );
  NOR2_X1 U5530 ( .A1(n9359), .A2(n9360), .ZN(n9358) );
  NOR2_X1 U5531 ( .A1(n9358), .A2(n4498), .ZN(n8805) );
  AND2_X1 U5532 ( .A1(n6563), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4498) );
  AND2_X1 U5533 ( .A1(n4497), .A2(n4496), .ZN(n9439) );
  NAND2_X1 U5534 ( .A1(n9321), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4496) );
  INV_X1 U5535 ( .A(n4495), .ZN(n9438) );
  OR2_X1 U5536 ( .A1(n9439), .A2(n9440), .ZN(n4495) );
  NOR2_X1 U5537 ( .A1(n9452), .A2(n4500), .ZN(n9462) );
  AND2_X1 U5538 ( .A1(n9457), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4500) );
  NOR2_X1 U5539 ( .A1(n9462), .A2(n9463), .ZN(n9461) );
  XNOR2_X1 U5540 ( .A(n8834), .B(n8835), .ZN(n9481) );
  NOR2_X1 U5541 ( .A1(n9461), .A2(n4499), .ZN(n8834) );
  AND2_X1 U5542 ( .A1(n8833), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4499) );
  NOR2_X1 U5543 ( .A1(n8823), .A2(n9477), .ZN(n8824) );
  OR2_X1 U5544 ( .A1(n9493), .A2(n9494), .ZN(n9496) );
  OR2_X1 U5545 ( .A1(n9001), .A2(n4464), .ZN(n8968) );
  INV_X1 U5546 ( .A(n8903), .ZN(n4546) );
  AND2_X1 U5547 ( .A1(n4554), .A2(n4323), .ZN(n4550) );
  NAND2_X1 U5548 ( .A1(n6637), .A2(n8697), .ZN(n8908) );
  NAND2_X1 U5549 ( .A1(n4351), .A2(n9058), .ZN(n9057) );
  NOR2_X1 U5550 ( .A1(n9079), .A2(n9218), .ZN(n9071) );
  NAND2_X1 U5551 ( .A1(n9071), .A2(n9052), .ZN(n9049) );
  NAND2_X1 U5552 ( .A1(n4528), .A2(n4526), .ZN(n9065) );
  NOR2_X1 U5553 ( .A1(n8888), .A2(n4527), .ZN(n4526) );
  INV_X1 U5554 ( .A(n8744), .ZN(n4527) );
  OR2_X1 U5555 ( .A1(n5428), .A2(n8361), .ZN(n5452) );
  NAND2_X1 U5556 ( .A1(n4528), .A2(n8744), .ZN(n9086) );
  OR2_X1 U5557 ( .A1(n5391), .A2(n8350), .ZN(n5410) );
  NAND2_X1 U5558 ( .A1(n4459), .A2(n4458), .ZN(n9118) );
  NOR2_X1 U5559 ( .A1(n9121), .A2(n4460), .ZN(n4458) );
  INV_X1 U5560 ( .A(n9523), .ZN(n4459) );
  NOR2_X1 U5561 ( .A1(n9118), .A2(n9228), .ZN(n9095) );
  NAND2_X1 U5562 ( .A1(n5346), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U5563 ( .A1(n9523), .A2(n4461), .ZN(n9146) );
  NOR2_X1 U5564 ( .A1(n9523), .A2(n4460), .ZN(n9126) );
  OR2_X1 U5565 ( .A1(n5318), .A2(n5317), .ZN(n5320) );
  OR2_X1 U5566 ( .A1(n5320), .A2(n5300), .ZN(n5348) );
  NAND2_X1 U5567 ( .A1(n9510), .A2(n8664), .ZN(n9509) );
  NOR2_X1 U5568 ( .A1(n8875), .A2(n8781), .ZN(n8914) );
  OR2_X1 U5569 ( .A1(n5243), .A2(n5242), .ZN(n5270) );
  NAND2_X1 U5570 ( .A1(n7104), .A2(n8637), .ZN(n6508) );
  OR2_X1 U5571 ( .A1(n4449), .A2(n8910), .ZN(n4446) );
  NAND2_X1 U5572 ( .A1(n4450), .A2(n9700), .ZN(n4449) );
  INV_X1 U5573 ( .A(n4451), .ZN(n4450) );
  NAND2_X1 U5574 ( .A1(n4448), .A2(n4447), .ZN(n9531) );
  NOR2_X1 U5575 ( .A1(n8910), .A2(n4451), .ZN(n4447) );
  INV_X1 U5576 ( .A(n9554), .ZN(n4448) );
  NOR2_X1 U5577 ( .A1(n9554), .A2(n7119), .ZN(n7185) );
  NOR2_X1 U5578 ( .A1(n9554), .A2(n4451), .ZN(n7200) );
  NAND2_X1 U5579 ( .A1(n4760), .A2(n4764), .ZN(n4758) );
  AND2_X1 U5580 ( .A1(n5179), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5181) );
  AND2_X1 U5581 ( .A1(n5133), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5179) );
  INV_X1 U5582 ( .A(n7112), .ZN(n7174) );
  INV_X1 U5583 ( .A(n8603), .ZN(n5388) );
  INV_X1 U5584 ( .A(n9568), .ZN(n4728) );
  AOI21_X1 U5585 ( .B1(n9568), .B2(n4727), .A(n4349), .ZN(n4726) );
  INV_X1 U5586 ( .A(n6916), .ZN(n4727) );
  NOR2_X1 U5587 ( .A1(n9569), .A2(n6919), .ZN(n9570) );
  OR2_X1 U5588 ( .A1(n9588), .A2(n8393), .ZN(n9569) );
  OAI21_X1 U5589 ( .B1(n9576), .B2(n6896), .A(n6895), .ZN(n8522) );
  NAND2_X1 U5590 ( .A1(n4445), .A2(n9642), .ZN(n9588) );
  NOR2_X1 U5592 ( .A1(n6793), .A2(n6792), .ZN(n9607) );
  OR2_X1 U5593 ( .A1(n9160), .A2(n4305), .ZN(n6517) );
  OR2_X1 U5594 ( .A1(n6508), .A2(n8756), .ZN(n9160) );
  AOI21_X1 U5595 ( .B1(n9618), .B2(n6516), .A(n6515), .ZN(n6739) );
  NAND2_X1 U5596 ( .A1(n4745), .A2(n4743), .ZN(n8977) );
  NAND2_X1 U5597 ( .A1(n9035), .A2(n4326), .ZN(n4745) );
  NOR2_X1 U5598 ( .A1(n9004), .A2(n8946), .ZN(n4744) );
  OAI21_X1 U5599 ( .B1(n9063), .B2(n8933), .A(n8932), .ZN(n9048) );
  NAND2_X1 U5600 ( .A1(n9075), .A2(n8930), .ZN(n8932) );
  AND2_X1 U5601 ( .A1(n6299), .A2(n6297), .ZN(n6514) );
  NOR2_X1 U5602 ( .A1(n4343), .A2(n4770), .ZN(n4769) );
  INV_X1 U5603 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4933) );
  INV_X1 U5604 ( .A(n9298), .ZN(n4930) );
  NOR2_X1 U5605 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4929) );
  INV_X1 U5606 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4926) );
  AOI21_X1 U5607 ( .B1(n5590), .B2(n5589), .A(n4782), .ZN(n4779) );
  INV_X1 U5608 ( .A(n4813), .ZN(n5558) );
  AOI21_X1 U5609 ( .B1(n5531), .B2(n5530), .A(n4816), .ZN(n4813) );
  XNOR2_X1 U5610 ( .A(n5625), .B(n5624), .ZN(n6363) );
  XNOR2_X1 U5611 ( .A(n4907), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U5612 ( .A1(n5424), .A2(n5423), .ZN(n5440) );
  NAND2_X1 U5613 ( .A1(n5290), .A2(n5289), .ZN(n5311) );
  OAI21_X1 U5614 ( .B1(n5235), .B2(n5234), .A(n5233), .ZN(n5259) );
  AND2_X1 U5615 ( .A1(n5236), .A2(n5216), .ZN(n8831) );
  OR3_X1 U5616 ( .A1(n5167), .A2(P1_IR_REG_8__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U5617 ( .A1(n5159), .A2(n5158), .ZN(n4440) );
  NAND2_X1 U5618 ( .A1(n4793), .A2(n5109), .ZN(n5142) );
  XNOR2_X1 U5619 ( .A(n4971), .B(SI_1_), .ZN(n4970) );
  NAND2_X1 U5620 ( .A1(n8613), .A2(n4348), .ZN(n4954) );
  INV_X1 U5621 ( .A(n6660), .ZN(n5764) );
  AND2_X1 U5622 ( .A1(n4587), .A2(n4321), .ZN(n7663) );
  INV_X1 U5623 ( .A(n7729), .ZN(n7694) );
  NAND2_X1 U5624 ( .A1(n7086), .A2(n5873), .ZN(n7241) );
  INV_X1 U5625 ( .A(n8027), .ZN(n8004) );
  NAND2_X1 U5626 ( .A1(n4625), .A2(n4626), .ZN(n7305) );
  NAND2_X1 U5627 ( .A1(n4638), .A2(n6068), .ZN(n7701) );
  NAND2_X1 U5628 ( .A1(n6054), .A2(n6053), .ZN(n8159) );
  NAND2_X1 U5629 ( .A1(n6145), .A2(n8106), .ZN(n7705) );
  NAND2_X1 U5630 ( .A1(n6865), .A2(n4317), .ZN(n6983) );
  INV_X1 U5631 ( .A(n7705), .ZN(n7737) );
  NAND2_X1 U5632 ( .A1(n7326), .A2(n5977), .ZN(n7314) );
  NAND2_X1 U5633 ( .A1(n6170), .A2(n6169), .ZN(n7734) );
  NAND2_X1 U5634 ( .A1(n6078), .A2(n6077), .ZN(n7964) );
  INV_X1 U5635 ( .A(n7647), .ZN(n7745) );
  INV_X1 U5636 ( .A(n7345), .ZN(n7746) );
  OR2_X2 U5637 ( .A1(n6399), .A2(P2_U3151), .ZN(n7878) );
  OR2_X1 U5638 ( .A1(n5744), .A2(n9782), .ZN(n5762) );
  NAND2_X1 U5639 ( .A1(n6381), .A2(n6382), .ZN(n6498) );
  INV_X1 U5640 ( .A(n4690), .ZN(n6497) );
  INV_X1 U5641 ( .A(n9779), .ZN(n7915) );
  OAI22_X1 U5642 ( .A1(n6495), .A2(n6579), .B1(n6410), .B2(n6409), .ZN(n9751)
         );
  AND2_X1 U5643 ( .A1(n4690), .A2(n6382), .ZN(n9741) );
  AOI22_X1 U5644 ( .A1(n9751), .A2(n9752), .B1(n6412), .B2(n6411), .ZN(n6482)
         );
  AND2_X1 U5645 ( .A1(n4697), .A2(n4695), .ZN(n6422) );
  OR2_X1 U5646 ( .A1(n6441), .A2(n6442), .ZN(n4403) );
  NAND2_X1 U5647 ( .A1(n6841), .A2(n4394), .ZN(n9773) );
  OR2_X1 U5648 ( .A1(n6842), .A2(n6852), .ZN(n4394) );
  NOR2_X1 U5649 ( .A1(n6837), .A2(n6835), .ZN(n7011) );
  NOR2_X1 U5650 ( .A1(n7029), .A2(n4562), .ZN(n6856) );
  NOR2_X1 U5651 ( .A1(n4563), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4562) );
  AND2_X1 U5652 ( .A1(n5877), .A2(n5897), .ZN(n7028) );
  OR2_X1 U5653 ( .A1(n7158), .A2(n7142), .ZN(n4710) );
  INV_X1 U5654 ( .A(n4561), .ZN(n7762) );
  NAND2_X1 U5655 ( .A1(n4707), .A2(n4706), .ZN(n7753) );
  INV_X1 U5656 ( .A(n7913), .ZN(n9774) );
  NAND2_X1 U5657 ( .A1(n4701), .A2(n4700), .ZN(n7800) );
  NOR2_X1 U5658 ( .A1(n7801), .A2(n7802), .ZN(n7837) );
  INV_X1 U5659 ( .A(n4407), .ZN(n7819) );
  XNOR2_X1 U5660 ( .A(n7882), .B(n7852), .ZN(n7849) );
  NOR2_X1 U5661 ( .A1(n7849), .A2(n8064), .ZN(n7886) );
  NAND2_X1 U5662 ( .A1(n4849), .A2(n4848), .ZN(n8024) );
  AND2_X1 U5663 ( .A1(n4849), .A2(n4363), .ZN(n8026) );
  OAI21_X1 U5664 ( .B1(n7284), .B2(n7451), .A(n7281), .ZN(n8090) );
  OR2_X1 U5665 ( .A1(n6816), .A2(n4310), .ZN(n4842) );
  INV_X1 U5666 ( .A(n8088), .ZN(n8112) );
  OR2_X1 U5667 ( .A1(n6278), .A2(n6281), .ZN(n8106) );
  INV_X1 U5668 ( .A(n8092), .ZN(n8085) );
  INV_X1 U5669 ( .A(n8106), .ZN(n8131) );
  INV_X1 U5670 ( .A(n8080), .ZN(n8135) );
  NOR2_X1 U5671 ( .A1(n6705), .A2(n6282), .ZN(n6284) );
  AND2_X1 U5672 ( .A1(n9370), .A2(n9369), .ZN(n9373) );
  NAND2_X1 U5673 ( .A1(n4572), .A2(n4575), .ZN(n7934) );
  OR2_X1 U5674 ( .A1(n8148), .A2(n4577), .ZN(n4572) );
  NAND2_X1 U5675 ( .A1(n4574), .A2(n7512), .ZN(n7943) );
  NAND2_X1 U5676 ( .A1(n8148), .A2(n4578), .ZN(n4574) );
  NAND2_X1 U5677 ( .A1(n8148), .A2(n7510), .ZN(n7953) );
  NAND2_X1 U5678 ( .A1(n4832), .A2(n4834), .ZN(n7978) );
  INV_X1 U5679 ( .A(n4835), .ZN(n4834) );
  INV_X1 U5680 ( .A(n7686), .ZN(n8246) );
  NAND2_X1 U5681 ( .A1(n6022), .A2(n6021), .ZN(n8249) );
  AND2_X1 U5682 ( .A1(n8045), .A2(n8044), .ZN(n8248) );
  NAND2_X1 U5683 ( .A1(n4607), .A2(n4608), .ZN(n8068) );
  NAND2_X1 U5684 ( .A1(n7284), .A2(n4611), .ZN(n4607) );
  INV_X1 U5685 ( .A(n8271), .ZN(n8280) );
  NAND2_X1 U5686 ( .A1(n4620), .A2(n4618), .ZN(n7074) );
  INV_X1 U5687 ( .A(n6278), .ZN(n8285) );
  AND2_X1 U5688 ( .A1(n6301), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6359) );
  INV_X1 U5689 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U5690 ( .A1(n5690), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5692) );
  INV_X1 U5691 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5703) );
  OR2_X1 U5692 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  INV_X1 U5693 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9960) );
  INV_X1 U5694 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7103) );
  XNOR2_X1 U5695 ( .A(n6134), .B(n6133), .ZN(n7102) );
  INV_X1 U5696 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U5697 ( .A1(n5717), .A2(n5719), .ZN(n5714) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10011) );
  INV_X1 U5699 ( .A(n7896), .ZN(n7918) );
  INV_X1 U5700 ( .A(n7797), .ZN(n7805) );
  INV_X1 U5701 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U5702 ( .A(n5898), .B(n5900), .ZN(n7134) );
  INV_X1 U5703 ( .A(n7028), .ZN(n6855) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6333) );
  INV_X1 U5705 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6329) );
  XNOR2_X1 U5706 ( .A(n5860), .B(n5859), .ZN(n6854) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6325) );
  NOR3_X1 U5708 ( .A1(n5770), .A2(n4857), .A3(P2_IR_REG_5__SCAN_IN), .ZN(n5825) );
  INV_X1 U5709 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6318) );
  NOR2_X1 U5710 ( .A1(n5770), .A2(n4857), .ZN(n5804) );
  INV_X1 U5711 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6312) );
  CLKBUF_X1 U5712 ( .A(n6380), .Z(n4397) );
  AND2_X1 U5713 ( .A1(n6363), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6297) );
  OR2_X1 U5714 ( .A1(n8603), .A2(n7381), .ZN(n5565) );
  AND2_X1 U5715 ( .A1(n5641), .A2(n5570), .ZN(n8986) );
  AOI21_X1 U5716 ( .B1(n4662), .B2(n4664), .A(n4660), .ZN(n4659) );
  INV_X1 U5717 ( .A(n8481), .ZN(n4660) );
  NAND2_X1 U5718 ( .A1(n4962), .A2(n4963), .ZN(n6620) );
  NAND2_X1 U5719 ( .A1(n4670), .A2(n4668), .ZN(n7267) );
  INV_X1 U5720 ( .A(n5203), .ZN(n4669) );
  NAND2_X1 U5721 ( .A1(n8365), .A2(n8367), .ZN(n8366) );
  NOR2_X1 U5722 ( .A1(n4647), .A2(n5055), .ZN(n8387) );
  NAND2_X1 U5723 ( .A1(n4650), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5724 ( .A1(n5334), .A2(n5333), .ZN(n8401) );
  INV_X1 U5725 ( .A(n4543), .ZN(n4542) );
  NAND2_X1 U5726 ( .A1(n6332), .A2(n8608), .ZN(n4544) );
  OAI21_X1 U5727 ( .B1(n8603), .B2(n6336), .A(n5124), .ZN(n4543) );
  NAND2_X1 U5728 ( .A1(n8615), .A2(n9312), .ZN(n4920) );
  NAND2_X1 U5729 ( .A1(n8355), .A2(n4653), .ZN(n4657) );
  AND2_X1 U5730 ( .A1(n5459), .A2(n5439), .ZN(n4653) );
  NAND2_X1 U5731 ( .A1(n4661), .A2(n4665), .ZN(n8482) );
  NAND2_X1 U5732 ( .A1(n5334), .A2(n4666), .ZN(n4661) );
  INV_X1 U5733 ( .A(n8949), .ZN(n8951) );
  INV_X1 U5734 ( .A(n8596), .ZN(n8947) );
  OR2_X1 U5735 ( .A1(n5455), .A2(n5454), .ZN(n8935) );
  OR2_X1 U5736 ( .A1(n5413), .A2(n5412), .ZN(n8928) );
  OR2_X1 U5737 ( .A1(n5378), .A2(n5377), .ZN(n8922) );
  OR2_X1 U5738 ( .A1(n5136), .A2(n5135), .ZN(n8785) );
  NAND4_X1 U5739 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n8788)
         );
  NAND2_X1 U5740 ( .A1(n4996), .A2(n4995), .ZN(n8790) );
  CLKBUF_X2 U5741 ( .A(P1_U3973), .Z(n8792) );
  INV_X1 U5742 ( .A(n4506), .ZN(n9341) );
  INV_X1 U5743 ( .A(n4504), .ZN(n9393) );
  INV_X1 U5744 ( .A(n4502), .ZN(n9392) );
  INV_X1 U5745 ( .A(n4497), .ZN(n9316) );
  AND2_X1 U5746 ( .A1(n4495), .A2(n4494), .ZN(n6536) );
  NAND2_X1 U5747 ( .A1(n6565), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4494) );
  INV_X1 U5748 ( .A(n9476), .ZN(n9489) );
  NAND2_X1 U5749 ( .A1(n4510), .A2(n4509), .ZN(n4508) );
  INV_X1 U5750 ( .A(n8874), .ZN(n4509) );
  NAND2_X1 U5751 ( .A1(n9400), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4510) );
  INV_X1 U5752 ( .A(n9223), .ZN(n9083) );
  NAND2_X1 U5753 ( .A1(n9142), .A2(n8669), .ZN(n9133) );
  NAND2_X1 U5754 ( .A1(n4535), .A2(n8537), .ZN(n8662) );
  OR2_X1 U5755 ( .A1(n7196), .A2(n8646), .ZN(n4535) );
  NAND2_X1 U5756 ( .A1(n4762), .A2(n4763), .ZN(n7182) );
  OR2_X1 U5757 ( .A1(n9541), .A2(n4764), .ZN(n4762) );
  NAND2_X1 U5758 ( .A1(n9541), .A2(n9544), .ZN(n4765) );
  OR2_X1 U5759 ( .A1(n9616), .A2(n9535), .ZN(n9167) );
  OR2_X1 U5760 ( .A1(n9616), .A2(n6750), .ZN(n9153) );
  INV_X1 U5761 ( .A(n9605), .ZN(n9519) );
  INV_X1 U5762 ( .A(n9167), .ZN(n9612) );
  INV_X1 U5763 ( .A(n9160), .ZN(n9608) );
  NAND2_X1 U5764 ( .A1(n9183), .A2(n4344), .ZN(n9250) );
  OAI21_X1 U5765 ( .B1(n9035), .B2(n4748), .A(n4746), .ZN(n8997) );
  NAND2_X1 U5766 ( .A1(n9035), .A2(n4754), .ZN(n4750) );
  OAI21_X1 U5767 ( .B1(n9035), .B2(n4318), .A(n4756), .ZN(n9021) );
  NAND2_X1 U5768 ( .A1(n4732), .A2(n4735), .ZN(n9078) );
  NAND2_X1 U5769 ( .A1(n4733), .A2(n4316), .ZN(n4732) );
  NAND2_X1 U5770 ( .A1(n4734), .A2(n4311), .ZN(n9094) );
  NAND2_X1 U5771 ( .A1(n9125), .A2(n4740), .ZN(n4734) );
  AOI21_X1 U5772 ( .B1(n9125), .B2(n9124), .A(n4742), .ZN(n9114) );
  AND2_X2 U5773 ( .A1(n6575), .A2(n6740), .ZN(n9714) );
  NAND2_X2 U5774 ( .A1(n6514), .A2(n6337), .ZN(n9618) );
  INV_X1 U5775 ( .A(n4936), .ZN(n9306) );
  CLKBUF_X1 U5776 ( .A(n6540), .Z(n8880) );
  NAND2_X1 U5777 ( .A1(n4898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4897) );
  INV_X1 U5778 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7106) );
  INV_X1 U5779 ( .A(n8769), .ZN(n7104) );
  INV_X1 U5780 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7040) );
  INV_X1 U5781 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6953) );
  XNOR2_X1 U5782 ( .A(n4909), .B(n4908), .ZN(n6955) );
  INV_X1 U5783 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4908) );
  INV_X1 U5784 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6362) );
  INV_X1 U5785 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6349) );
  INV_X1 U5786 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6336) );
  INV_X1 U5787 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6331) );
  INV_X1 U5788 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U5789 ( .A1(n4515), .A2(n5068), .ZN(n5088) );
  INV_X1 U5790 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6320) );
  INV_X1 U5791 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U5792 ( .A1(n4415), .A2(n5004), .ZN(n5020) );
  NAND2_X1 U5793 ( .A1(n5002), .A2(n5001), .ZN(n4415) );
  NAND2_X1 U5794 ( .A1(n9384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4493) );
  OR2_X1 U5795 ( .A1(n6177), .A2(n6176), .ZN(P2_U3154) );
  AND2_X1 U5796 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  OAI21_X1 U5797 ( .B1(n6295), .B2(n9847), .A(n4398), .ZN(P2_U3488) );
  NOR2_X1 U5798 ( .A1(n4378), .A2(n4399), .ZN(n4398) );
  NOR2_X1 U5799 ( .A1(n9849), .A2(n6285), .ZN(n4399) );
  INV_X1 U5800 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5801 ( .A1(n5630), .A2(n4864), .ZN(n5655) );
  NAND2_X1 U5802 ( .A1(n4513), .A2(n4305), .ZN(n4512) );
  AOI21_X1 U5803 ( .B1(n4511), .B2(n9535), .A(n4508), .ZN(n4507) );
  OAI22_X1 U5804 ( .A1(n8871), .A2(n9479), .B1(n8872), .B2(n9476), .ZN(n4513)
         );
  NAND2_X1 U5805 ( .A1(n4525), .A2(n4523), .ZN(P1_U3519) );
  OR2_X1 U5806 ( .A1(n9714), .A2(n4524), .ZN(n4523) );
  NAND2_X1 U5807 ( .A1(n9250), .A2(n9714), .ZN(n4525) );
  INV_X1 U5808 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5809 ( .A1(n4516), .A2(n4517), .ZN(n4518) );
  NOR2_X1 U5810 ( .A1(n7559), .A2(n7558), .ZN(n4308) );
  NAND2_X1 U5811 ( .A1(n9306), .A2(n4935), .ZN(n4992) );
  AND2_X1 U5812 ( .A1(n4735), .A2(n4335), .ZN(n4309) );
  AND2_X1 U5813 ( .A1(n7090), .A2(n9809), .ZN(n4310) );
  OR2_X1 U5814 ( .A1(n6608), .A2(n4721), .ZN(n4718) );
  AND2_X1 U5815 ( .A1(n4360), .A2(n4739), .ZN(n4311) );
  INV_X1 U5816 ( .A(n6494), .ZN(n4699) );
  OR2_X1 U5817 ( .A1(n4491), .A2(n4770), .ZN(n4312) );
  AND3_X1 U5818 ( .A1(n8643), .A2(n8523), .A3(n8641), .ZN(n4313) );
  INV_X1 U5819 ( .A(n8893), .ZN(n9058) );
  AND2_X1 U5820 ( .A1(n5450), .A2(n5449), .ZN(n9052) );
  AND2_X1 U5821 ( .A1(n7889), .A2(n7888), .ZN(n4314) );
  NOR2_X1 U5822 ( .A1(n6383), .A2(n4699), .ZN(n6386) );
  INV_X1 U5823 ( .A(n9528), .ZN(n4529) );
  INV_X1 U5824 ( .A(n8931), .ZN(n8930) );
  INV_X1 U5825 ( .A(n5739), .ZN(n5928) );
  INV_X1 U5826 ( .A(n4596), .ZN(n6868) );
  NAND2_X1 U5827 ( .A1(n5263), .A2(n4771), .ZN(n4905) );
  OR2_X1 U5828 ( .A1(n9194), .A2(n8945), .ZN(n4315) );
  AND2_X1 U5829 ( .A1(n4311), .A2(n4738), .ZN(n4316) );
  AND2_X1 U5830 ( .A1(n5837), .A2(n5824), .ZN(n4317) );
  NOR2_X1 U5831 ( .A1(n9209), .A2(n8938), .ZN(n4318) );
  XNOR2_X1 U5832 ( .A(n4297), .B(n5054), .ZN(n4319) );
  INV_X1 U5833 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U5834 ( .A1(n8719), .A2(n9559), .ZN(n4320) );
  AND2_X1 U5835 ( .A1(n5497), .A2(n5496), .ZN(n9032) );
  NAND2_X1 U5836 ( .A1(n8605), .A2(n8604), .ZN(n9179) );
  NAND2_X1 U5837 ( .A1(n5995), .A2(n8098), .ZN(n4321) );
  INV_X1 U5838 ( .A(n8910), .ZN(n9693) );
  NAND2_X1 U5839 ( .A1(n6459), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U5840 ( .A1(n4750), .A2(n4751), .ZN(n9007) );
  XNOR2_X1 U5841 ( .A(n8207), .B(n7946), .ZN(n7933) );
  NAND2_X1 U5842 ( .A1(n5361), .A2(n5360), .ZN(n5384) );
  INV_X1 U5843 ( .A(n8954), .ZN(n4483) );
  INV_X1 U5844 ( .A(n5770), .ZN(n4687) );
  INV_X1 U5845 ( .A(n6382), .ZN(n4689) );
  INV_X1 U5846 ( .A(n4597), .ZN(n4594) );
  AND2_X1 U5847 ( .A1(n8901), .A2(n4551), .ZN(n4323) );
  NAND2_X1 U5848 ( .A1(n5344), .A2(n5343), .ZN(n9239) );
  AND2_X1 U5849 ( .A1(n4502), .A2(n4501), .ZN(n4324) );
  AND4_X1 U5850 ( .A1(n5914), .A2(n5948), .A3(n5901), .A4(n5669), .ZN(n4325)
         );
  AND2_X1 U5851 ( .A1(n4746), .A2(n4315), .ZN(n4326) );
  NAND2_X1 U5852 ( .A1(n5098), .A2(n5099), .ZN(n4327) );
  NAND2_X1 U5853 ( .A1(n7748), .A2(n6245), .ZN(n4328) );
  AND2_X1 U5854 ( .A1(n6417), .A2(n6416), .ZN(n4329) );
  INV_X1 U5855 ( .A(n7568), .ZN(n4621) );
  AND2_X1 U5856 ( .A1(n4531), .A2(n4529), .ZN(n4330) );
  AND2_X1 U5857 ( .A1(n6459), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4331) );
  AND2_X1 U5858 ( .A1(n8226), .A2(n7964), .ZN(n4332) );
  AND2_X1 U5859 ( .A1(n5934), .A2(n7744), .ZN(n4333) );
  NAND2_X1 U5860 ( .A1(n5682), .A2(n5757), .ZN(n5741) );
  INV_X1 U5861 ( .A(n9121), .ZN(n9233) );
  NAND2_X1 U5862 ( .A1(n5371), .A2(n5370), .ZN(n9121) );
  AND2_X1 U5863 ( .A1(n4580), .A2(n7711), .ZN(n4334) );
  OR2_X1 U5864 ( .A1(n9223), .A2(n8928), .ZN(n4335) );
  AND2_X1 U5865 ( .A1(n4432), .A2(n4434), .ZN(n4336) );
  AND2_X1 U5866 ( .A1(n7575), .A2(n7449), .ZN(n4337) );
  NAND2_X1 U5867 ( .A1(n9071), .A2(n4455), .ZN(n4456) );
  OR2_X1 U5868 ( .A1(n7686), .A2(n7742), .ZN(n4338) );
  AND2_X1 U5869 ( .A1(n4719), .A2(n4711), .ZN(n4339) );
  NAND2_X1 U5870 ( .A1(n8659), .A2(n8612), .ZN(n4340) );
  INV_X1 U5871 ( .A(n9629), .ZN(n6792) );
  AND3_X1 U5872 ( .A1(n4981), .A2(n4980), .A3(n4979), .ZN(n9629) );
  NAND2_X1 U5873 ( .A1(n6716), .A2(n4342), .ZN(n4652) );
  AND2_X1 U5874 ( .A1(n5886), .A2(n5873), .ZN(n4341) );
  AND2_X1 U5875 ( .A1(n4319), .A2(n5037), .ZN(n4342) );
  NAND2_X1 U5876 ( .A1(n4913), .A2(n4912), .ZN(n4343) );
  AND2_X1 U5877 ( .A1(n4867), .A2(n4724), .ZN(n4344) );
  AND2_X1 U5878 ( .A1(n4648), .A2(n8388), .ZN(n4345) );
  OR2_X1 U5879 ( .A1(n7352), .A2(n7647), .ZN(n7440) );
  INV_X1 U5880 ( .A(n7440), .ZN(n4613) );
  INV_X1 U5881 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4896) );
  OR2_X1 U5882 ( .A1(n6378), .A2(n4397), .ZN(n4346) );
  INV_X1 U5883 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U5884 ( .A1(n7664), .A2(n4321), .ZN(n4586) );
  NOR2_X1 U5885 ( .A1(n7748), .A2(n6245), .ZN(n4347) );
  AND2_X1 U5886 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4348) );
  AND2_X1 U5887 ( .A1(n6918), .A2(n9655), .ZN(n4349) );
  OR2_X1 U5888 ( .A1(n7304), .A2(n5973), .ZN(n4350) );
  NAND2_X1 U5889 ( .A1(n7582), .A2(n7532), .ZN(n7526) );
  INV_X1 U5890 ( .A(n7526), .ZN(n4438) );
  INV_X1 U5891 ( .A(n4757), .ZN(n4756) );
  NOR2_X1 U5892 ( .A1(n9045), .A2(n8939), .ZN(n4757) );
  AND2_X1 U5893 ( .A1(n8892), .A2(n8891), .ZN(n4351) );
  NOR2_X1 U5894 ( .A1(n9018), .A2(n8944), .ZN(n4352) );
  INV_X1 U5895 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5805) );
  OR2_X1 U5896 ( .A1(n9199), .A2(n8943), .ZN(n4353) );
  AND3_X1 U5897 ( .A1(n5263), .A2(n4457), .A3(n4771), .ZN(n4894) );
  NAND2_X1 U5898 ( .A1(n4893), .A2(n4896), .ZN(n4770) );
  AND2_X1 U5899 ( .A1(n7525), .A2(n4436), .ZN(n4354) );
  NAND2_X1 U5900 ( .A1(n9190), .A2(n8596), .ZN(n8902) );
  AND2_X1 U5901 ( .A1(n5316), .A2(n5315), .ZN(n9377) );
  NOR2_X1 U5902 ( .A1(n7655), .A2(n7979), .ZN(n4355) );
  AND2_X1 U5903 ( .A1(n8226), .A2(n7993), .ZN(n7501) );
  AND2_X1 U5904 ( .A1(n5337), .A2(n5336), .ZN(n4356) );
  AND2_X1 U5905 ( .A1(n5022), .A2(SI_3_), .ZN(n4357) );
  AND2_X1 U5906 ( .A1(n5090), .A2(SI_6_), .ZN(n4358) );
  AND2_X1 U5907 ( .A1(n4748), .A2(n4315), .ZN(n4359) );
  OR2_X1 U5908 ( .A1(n9233), .A2(n8923), .ZN(n4360) );
  INV_X1 U5909 ( .A(n7047), .ZN(n4767) );
  OR2_X1 U5910 ( .A1(n4905), .A2(n4890), .ZN(n4361) );
  NOR2_X1 U5911 ( .A1(n9083), .A2(n8929), .ZN(n4362) );
  NAND2_X1 U5912 ( .A1(n5520), .A2(n5519), .ZN(n9199) );
  NAND2_X1 U5913 ( .A1(n8249), .A2(n8052), .ZN(n4363) );
  AND2_X1 U5914 ( .A1(n4548), .A2(n4552), .ZN(n4364) );
  OR2_X1 U5915 ( .A1(n7190), .A2(n8783), .ZN(n4365) );
  AND2_X1 U5916 ( .A1(n8523), .A2(n8716), .ZN(n4366) );
  AND3_X2 U5917 ( .A1(n4957), .A2(n4956), .A3(n4955), .ZN(n8707) );
  INV_X1 U5918 ( .A(n8707), .ZN(n9620) );
  INV_X1 U5919 ( .A(n8876), .ZN(n9175) );
  AND2_X1 U5920 ( .A1(n5170), .A2(n5169), .ZN(n9688) );
  OR2_X1 U5921 ( .A1(n7557), .A2(n7519), .ZN(n4367) );
  NOR2_X1 U5922 ( .A1(n9760), .A2(n6471), .ZN(n4368) );
  AND2_X1 U5923 ( .A1(n6357), .A2(n6135), .ZN(n4369) );
  NOR2_X1 U5924 ( .A1(n8876), .A2(n4463), .ZN(n4370) );
  AND2_X1 U5925 ( .A1(n4632), .A2(n4635), .ZN(n4371) );
  AND2_X1 U5926 ( .A1(n8536), .A2(n8722), .ZN(n7181) );
  INV_X1 U5927 ( .A(n7181), .ZN(n4761) );
  INV_X1 U5928 ( .A(n4553), .ZN(n4552) );
  OAI21_X1 U5929 ( .B1(n8684), .B2(n8981), .A(n8902), .ZN(n4553) );
  NAND2_X1 U5930 ( .A1(n8410), .A2(n5511), .ZN(n8365) );
  AND2_X1 U5931 ( .A1(n7443), .A2(n7444), .ZN(n7574) );
  OR2_X1 U5932 ( .A1(n8179), .A2(n7668), .ZN(n7458) );
  AND2_X1 U5933 ( .A1(n5106), .A2(n4417), .ZN(n4372) );
  OR2_X1 U5934 ( .A1(n5996), .A2(n4858), .ZN(n4373) );
  INV_X1 U5935 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6133) );
  INV_X1 U5936 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5826) );
  INV_X1 U5937 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4783) );
  AND2_X1 U5938 ( .A1(n7691), .A2(n6043), .ZN(n4374) );
  NOR2_X1 U5939 ( .A1(n7305), .A2(n7304), .ZN(n4375) );
  OR2_X1 U5940 ( .A1(n9523), .A2(n9165), .ZN(n4376) );
  AND2_X1 U5941 ( .A1(n5263), .A2(n4887), .ZN(n5265) );
  BUF_X1 U5942 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9384) );
  NAND2_X1 U5943 ( .A1(n5427), .A2(n5426), .ZN(n9218) );
  INV_X1 U5944 ( .A(n9218), .ZN(n9075) );
  AND2_X1 U5945 ( .A1(n6560), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4377) );
  INV_X1 U5946 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4559) );
  INV_X1 U5947 ( .A(n7630), .ZN(n4601) );
  INV_X1 U5948 ( .A(n9190), .ZN(n4465) );
  NAND2_X1 U5949 ( .A1(n4598), .A2(n4599), .ZN(n7632) );
  NOR2_X1 U5950 ( .A1(n7928), .A2(n8180), .ZN(n4378) );
  AND2_X1 U5951 ( .A1(n4530), .A2(n4531), .ZN(n4379) );
  NOR2_X1 U5952 ( .A1(n7793), .A2(n7755), .ZN(n4380) );
  NOR2_X1 U5953 ( .A1(n7129), .A2(n7142), .ZN(n4381) );
  AND2_X1 U5954 ( .A1(n5442), .A2(n5441), .ZN(n4382) );
  AND2_X1 U5955 ( .A1(n8668), .A2(n8667), .ZN(n4383) );
  NAND2_X1 U5956 ( .A1(n6854), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4384) );
  AND2_X1 U5957 ( .A1(n4705), .A2(n4704), .ZN(n4385) );
  AND2_X1 U5958 ( .A1(n5713), .A2(n6357), .ZN(n6115) );
  AND2_X1 U5959 ( .A1(n6294), .A2(n6293), .ZN(n9886) );
  NOR2_X1 U5960 ( .A1(n6583), .A2(n6156), .ZN(n7920) );
  NAND2_X1 U5961 ( .A1(n6983), .A2(n5856), .ZN(n6984) );
  INV_X1 U5962 ( .A(n8398), .ZN(n4667) );
  INV_X1 U5963 ( .A(n7149), .ZN(n7763) );
  OAI21_X1 U5964 ( .B1(n6917), .B2(n4728), .A(n4726), .ZN(n7042) );
  NAND2_X1 U5965 ( .A1(n4765), .A2(n7047), .ZN(n7118) );
  NAND2_X1 U5966 ( .A1(n6917), .A2(n6916), .ZN(n9567) );
  XNOR2_X1 U5967 ( .A(n4897), .B(n4896), .ZN(n5615) );
  INV_X1 U5968 ( .A(n7710), .ZN(n4583) );
  AOI21_X1 U5969 ( .B1(n8522), .B2(n8716), .A(n4320), .ZN(n8517) );
  INV_X1 U5970 ( .A(n8517), .ZN(n4522) );
  NAND2_X1 U5971 ( .A1(n6865), .A2(n5824), .ZN(n6926) );
  NAND2_X1 U5972 ( .A1(n4838), .A2(n6201), .ZN(n7068) );
  NOR2_X1 U5973 ( .A1(n4446), .A2(n9554), .ZN(n9522) );
  AND2_X1 U5974 ( .A1(n7805), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4386) );
  AND2_X1 U5975 ( .A1(n4710), .A2(n4709), .ZN(n4387) );
  OR2_X1 U5976 ( .A1(n7149), .A2(n7224), .ZN(n4388) );
  NAND2_X1 U5977 ( .A1(n7805), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4703) );
  AND3_X2 U5978 ( .A1(n6704), .A2(n6284), .A3(n6283), .ZN(n9849) );
  NAND2_X1 U5979 ( .A1(n4720), .A2(n4722), .ZN(n4719) );
  AND2_X1 U5980 ( .A1(n4718), .A2(n4719), .ZN(n4389) );
  NAND2_X1 U5981 ( .A1(n9607), .A2(n9637), .ZN(n9587) );
  INV_X1 U5982 ( .A(n9587), .ZN(n4445) );
  NAND2_X1 U5983 ( .A1(n7076), .A2(n9826), .ZN(n4633) );
  AND3_X1 U5984 ( .A1(n4698), .A2(n6384), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n4390) );
  XOR2_X1 U5985 ( .A(n6459), .B(n6432), .Z(n4391) );
  INV_X1 U5986 ( .A(n4305), .ZN(n9535) );
  NAND2_X1 U5987 ( .A1(n6394), .A2(n6396), .ZN(n4564) );
  AOI22_X1 U5988 ( .A1(n6604), .A2(n6603), .B1(n6445), .B2(n6605), .ZN(n6448)
         );
  NAND2_X1 U5989 ( .A1(n6423), .A2(n6605), .ZN(n6424) );
  INV_X1 U5990 ( .A(n6605), .ZN(n4392) );
  NOR2_X1 U5991 ( .A1(n7804), .A2(n8184), .ZN(n7820) );
  NOR2_X1 U5992 ( .A1(n7871), .A2(n7870), .ZN(n7895) );
  INV_X1 U5993 ( .A(n6430), .ZN(n4393) );
  NOR2_X1 U5994 ( .A1(n7820), .A2(n7821), .ZN(n7823) );
  NOR2_X1 U5995 ( .A1(n7869), .A2(n7868), .ZN(n7871) );
  OAI21_X1 U5996 ( .B1(n6411), .B2(n9946), .A(n4405), .ZN(n9744) );
  XNOR2_X1 U5997 ( .A(n6851), .B(n6852), .ZN(n6461) );
  NAND2_X1 U5998 ( .A1(n9743), .A2(n9744), .ZN(n9742) );
  INV_X1 U5999 ( .A(n5205), .ZN(n5208) );
  NAND2_X1 U6000 ( .A1(n5159), .A2(n4795), .ZN(n4794) );
  NAND2_X2 U6001 ( .A1(n5285), .A2(n5284), .ZN(n5290) );
  AND4_X2 U6002 ( .A1(n5668), .A2(n5859), .A3(n5951), .A4(n5667), .ZN(n4873)
         );
  NOR2_X1 U6003 ( .A1(n6844), .A2(n9776), .ZN(n6845) );
  AOI21_X1 U6004 ( .B1(n7874), .B2(n7884), .A(n7873), .ZN(n7876) );
  NOR2_X1 U6005 ( .A1(n7147), .A2(n7159), .ZN(n7758) );
  NOR2_X1 U6006 ( .A1(n7144), .A2(n7143), .ZN(n7160) );
  NOR2_X1 U6007 ( .A1(n7775), .A2(n7774), .ZN(n7777) );
  NAND2_X2 U6008 ( .A1(n8437), .A2(n5418), .ZN(n8356) );
  NAND2_X1 U6009 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  INV_X1 U6010 ( .A(n7754), .ZN(n4395) );
  AOI21_X1 U6011 ( .B1(n7921), .B2(n7920), .A(n7919), .ZN(n7922) );
  XNOR2_X2 U6012 ( .A(n5795), .B(n5794), .ZN(n6427) );
  AOI21_X1 U6013 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7134), .A(n7126), .ZN(
        n7127) );
  NOR2_X1 U6014 ( .A1(n9981), .A2(n7851), .ZN(n7869) );
  NAND2_X1 U6015 ( .A1(n4556), .A2(n4555), .ZN(n6851) );
  NAND2_X1 U6016 ( .A1(n6999), .A2(n6200), .ZN(n4838) );
  OAI21_X2 U6017 ( .B1(n8051), .B2(n6213), .A(n6212), .ZN(n8037) );
  INV_X1 U6018 ( .A(n7280), .ZN(n6207) );
  AOI21_X2 U6019 ( .B1(n9057), .B2(n8897), .A(n8896), .ZN(n9024) );
  NAND2_X1 U6020 ( .A1(n5115), .A2(n5114), .ZN(n5157) );
  OAI21_X1 U6021 ( .B1(n8668), .B2(n4540), .A(n4538), .ZN(n9108) );
  NAND2_X1 U6022 ( .A1(n5290), .A2(n4803), .ZN(n4802) );
  NAND2_X1 U6023 ( .A1(n4802), .A2(n5294), .ZN(n5339) );
  NOR2_X1 U6024 ( .A1(n8982), .A2(n8981), .ZN(n8980) );
  NAND2_X4 U6025 ( .A1(n4911), .A2(n6299), .ZN(n5601) );
  NAND2_X1 U6026 ( .A1(n4657), .A2(n8323), .ZN(n8456) );
  NAND2_X1 U6027 ( .A1(n5208), .A2(n5207), .ZN(n5210) );
  INV_X1 U6028 ( .A(n4636), .ZN(n4635) );
  NAND2_X1 U6029 ( .A1(n4788), .A2(n5444), .ZN(n5464) );
  INV_X1 U6030 ( .A(n5004), .ZN(n4413) );
  NAND2_X1 U6031 ( .A1(n4414), .A2(n4412), .ZN(n4514) );
  NOR2_X4 U6032 ( .A1(n5062), .A2(n4886), .ZN(n5263) );
  OAI21_X2 U6033 ( .B1(n5290), .B2(n4799), .A(n4797), .ZN(n5357) );
  AND2_X1 U6034 ( .A1(n6851), .A2(n6852), .ZN(n4400) );
  NAND2_X1 U6035 ( .A1(n4512), .A2(n4507), .ZN(P1_U3262) );
  NAND2_X1 U6036 ( .A1(n4873), .A2(n4325), .ZN(n5670) );
  NOR2_X2 U6037 ( .A1(n7033), .A2(n7032), .ZN(n7133) );
  OAI21_X1 U6038 ( .B1(n5736), .B2(n5768), .A(n5767), .ZN(n5769) );
  NOR2_X1 U6039 ( .A1(n7165), .A2(n7136), .ZN(n7138) );
  NAND2_X1 U6040 ( .A1(n4975), .A2(n4783), .ZN(n4409) );
  NAND3_X1 U6041 ( .A1(n4517), .A2(n4917), .A3(n4516), .ZN(n4410) );
  NAND3_X1 U6042 ( .A1(n5001), .A2(n5002), .A3(n5019), .ZN(n4414) );
  NAND2_X1 U6043 ( .A1(n4515), .A2(n4418), .ZN(n4416) );
  NAND2_X1 U6044 ( .A1(n4416), .A2(n4372), .ZN(n4793) );
  OAI21_X1 U6045 ( .B1(n4515), .B2(n4420), .A(n4418), .ZN(n5107) );
  NAND3_X1 U6046 ( .A1(n4422), .A2(n7573), .A3(n7445), .ZN(n4421) );
  NAND3_X1 U6047 ( .A1(n4426), .A2(n4423), .A3(n7574), .ZN(n4422) );
  INV_X1 U6048 ( .A(n7525), .ZN(n4431) );
  AND2_X1 U6049 ( .A1(n7529), .A2(n7582), .ZN(n4435) );
  INV_X1 U6050 ( .A(n7527), .ZN(n4437) );
  NAND3_X1 U6051 ( .A1(n7435), .A2(n4442), .A3(n4441), .ZN(n7439) );
  OAI211_X1 U6052 ( .C1(n7433), .C2(n7427), .A(n7438), .B(n7426), .ZN(n4443)
         );
  NAND3_X1 U6053 ( .A1(n7476), .A2(n4367), .A3(n4444), .ZN(n7483) );
  INV_X1 U6054 ( .A(n4456), .ZN(n9041) );
  NAND2_X1 U6055 ( .A1(n4925), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4922) );
  NAND4_X1 U6056 ( .A1(n5263), .A2(n4769), .A3(n4771), .A4(n4457), .ZN(n4925)
         );
  INV_X1 U6057 ( .A(n9001), .ZN(n4462) );
  NAND2_X1 U6058 ( .A1(n4370), .A2(n4462), .ZN(n8884) );
  NOR2_X1 U6059 ( .A1(n9001), .A2(n4463), .ZN(n8955) );
  NOR2_X1 U6060 ( .A1(n9001), .A2(n9190), .ZN(n8978) );
  AOI21_X1 U6061 ( .B1(n4466), .B2(n8527), .A(n8526), .ZN(n8528) );
  NAND2_X1 U6062 ( .A1(n4467), .A2(n8524), .ZN(n4466) );
  NAND2_X1 U6063 ( .A1(n4468), .A2(n8719), .ZN(n4467) );
  NAND2_X1 U6064 ( .A1(n8718), .A2(n4366), .ZN(n4468) );
  AOI21_X1 U6065 ( .B1(n8549), .B2(n9512), .A(n8548), .ZN(n8551) );
  NAND2_X1 U6066 ( .A1(n8542), .A2(n8766), .ZN(n4474) );
  INV_X1 U6067 ( .A(n8583), .ZN(n4475) );
  INV_X1 U6068 ( .A(n8582), .ZN(n4476) );
  NAND2_X1 U6069 ( .A1(n4478), .A2(n4340), .ZN(n4477) );
  NAND3_X1 U6070 ( .A1(n4490), .A2(n4489), .A3(n8559), .ZN(n4488) );
  NAND3_X1 U6071 ( .A1(n8552), .A2(n8612), .A3(n8737), .ZN(n4490) );
  MUX2_X1 U6072 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6525), .S(n4300), .Z(n8798)
         );
  NAND2_X1 U6073 ( .A1(n4514), .A2(n5047), .ZN(n5051) );
  XNOR2_X1 U6074 ( .A(n4514), .B(n5047), .ZN(n6311) );
  AND2_X1 U6075 ( .A1(n4519), .A2(n4518), .ZN(n6683) );
  INV_X1 U6076 ( .A(n6682), .ZN(n4519) );
  NAND2_X1 U6077 ( .A1(n4521), .A2(n4520), .ZN(n7112) );
  INV_X1 U6078 ( .A(n8645), .ZN(n4521) );
  NAND2_X2 U6079 ( .A1(n4298), .A2(P1_U3086), .ZN(n9308) );
  NAND2_X2 U6080 ( .A1(n4298), .A2(P2_U3151), .ZN(n8304) );
  MUX2_X1 U6081 ( .A(n6308), .B(n6322), .S(n4975), .Z(n5021) );
  MUX2_X1 U6082 ( .A(n6310), .B(n6312), .S(n4298), .Z(n5048) );
  MUX2_X1 U6083 ( .A(n6320), .B(n6318), .S(n4298), .Z(n5066) );
  MUX2_X1 U6084 ( .A(n6323), .B(n6325), .S(n4298), .Z(n5089) );
  MUX2_X1 U6085 ( .A(n6331), .B(n6329), .S(n4298), .Z(n5111) );
  MUX2_X1 U6086 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n4298), .Z(n5108) );
  MUX2_X1 U6087 ( .A(n6336), .B(n6333), .S(n4298), .Z(n5117) );
  MUX2_X1 U6088 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n4298), .Z(n5160) );
  MUX2_X1 U6089 ( .A(n6362), .B(n6352), .S(n4298), .Z(n5231) );
  MUX2_X1 U6090 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n4298), .Z(n5260) );
  MUX2_X1 U6091 ( .A(n6349), .B(n5162), .S(n4298), .Z(n5164) );
  MUX2_X1 U6092 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n4298), .Z(n5286) );
  MUX2_X1 U6093 ( .A(n6600), .B(n5291), .S(n4298), .Z(n5309) );
  MUX2_X1 U6094 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n4298), .Z(n5335) );
  MUX2_X1 U6095 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n4298), .Z(n5362) );
  MUX2_X1 U6096 ( .A(n5340), .B(n5341), .S(n4298), .Z(n5359) );
  MUX2_X1 U6097 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n4298), .Z(n5400) );
  MUX2_X1 U6098 ( .A(n6953), .B(n10011), .S(n4298), .Z(n5422) );
  MUX2_X1 U6099 ( .A(n7040), .B(n6996), .S(n4298), .Z(n5442) );
  MUX2_X1 U6100 ( .A(n7106), .B(n7103), .S(n4298), .Z(n5446) );
  MUX2_X1 U6101 ( .A(n7217), .B(n9960), .S(n4298), .Z(n5466) );
  MUX2_X1 U6102 ( .A(n7230), .B(n7278), .S(n4298), .Z(n5493) );
  MUX2_X1 U6103 ( .A(n7288), .B(n7276), .S(n4298), .Z(n5516) );
  MUX2_X1 U6104 ( .A(n9309), .B(n8301), .S(n4298), .Z(n5534) );
  MUX2_X1 U6105 ( .A(n7381), .B(n8297), .S(n4298), .Z(n5562) );
  MUX2_X1 U6106 ( .A(n9303), .B(n8293), .S(n4298), .Z(n7367) );
  NAND2_X1 U6107 ( .A1(n8991), .A2(n4550), .ZN(n4547) );
  NAND2_X1 U6108 ( .A1(n8991), .A2(n4323), .ZN(n4548) );
  AOI21_X1 U6109 ( .B1(n8991), .B2(n8901), .A(n8900), .ZN(n8982) );
  NOR2_X4 U6110 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5736) );
  OAI21_X1 U6111 ( .B1(n6607), .B2(n4557), .A(n4558), .ZN(n6460) );
  NAND2_X1 U6112 ( .A1(n6607), .A2(n4558), .ZN(n4555) );
  AOI21_X1 U6113 ( .B1(n4558), .B2(n4557), .A(n4331), .ZN(n4556) );
  INV_X1 U6114 ( .A(n6433), .ZN(n4557) );
  AND2_X2 U6115 ( .A1(n4561), .A2(n4560), .ZN(n7773) );
  NAND2_X1 U6116 ( .A1(n4566), .A2(n6396), .ZN(n4567) );
  NAND2_X1 U6117 ( .A1(n8029), .A2(n7486), .ZN(n4568) );
  NAND2_X1 U6118 ( .A1(n4569), .A2(n7477), .ZN(n8029) );
  NAND2_X1 U6119 ( .A1(n8035), .A2(n7478), .ZN(n4569) );
  NAND4_X1 U6120 ( .A1(n5736), .A2(n4856), .A3(n4570), .A4(n5826), .ZN(n5838)
         );
  NAND2_X1 U6121 ( .A1(n8148), .A2(n4575), .ZN(n4571) );
  NAND2_X1 U6122 ( .A1(n4571), .A2(n4573), .ZN(n6257) );
  NAND2_X1 U6123 ( .A1(n7337), .A2(n4582), .ZN(n4581) );
  OAI21_X1 U6124 ( .B1(n6594), .B2(n6421), .A(n5801), .ZN(n4597) );
  NAND2_X1 U6125 ( .A1(n4596), .A2(n4595), .ZN(n7410) );
  NAND2_X1 U6126 ( .A1(n4588), .A2(n4594), .ZN(n4596) );
  INV_X1 U6127 ( .A(n4593), .ZN(n4588) );
  NAND2_X1 U6128 ( .A1(n4590), .A2(n7402), .ZN(n6946) );
  NOR2_X1 U6129 ( .A1(n4593), .A2(n4595), .ZN(n4589) );
  NAND2_X1 U6130 ( .A1(n4593), .A2(n4595), .ZN(n4592) );
  INV_X1 U6131 ( .A(n6030), .ZN(n7691) );
  NAND2_X1 U6132 ( .A1(n6030), .A2(n7630), .ZN(n4598) );
  OAI21_X2 U6133 ( .B1(n7284), .B2(n4605), .A(n4602), .ZN(n8059) );
  OR2_X1 U6134 ( .A1(n6250), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U6135 ( .A1(n7451), .A2(n7281), .ZN(n4610) );
  OAI21_X2 U6136 ( .B1(n6935), .B2(n4614), .A(n4612), .ZN(n7209) );
  NAND2_X1 U6137 ( .A1(n7290), .A2(n4627), .ZN(n4625) );
  NAND2_X2 U6138 ( .A1(n4625), .A2(n4623), .ZN(n7326) );
  AND2_X1 U6139 ( .A1(n7648), .A2(n5931), .ZN(n4627) );
  AOI21_X1 U6140 ( .B1(n7931), .B2(n4633), .A(n4636), .ZN(n6295) );
  NAND2_X1 U6141 ( .A1(n7931), .A2(n8127), .ZN(n4632) );
  OAI21_X1 U6142 ( .B1(n7931), .B2(n4631), .A(n4628), .ZN(n6296) );
  OR2_X2 U6143 ( .A1(n4636), .A2(n9886), .ZN(n4631) );
  NAND2_X2 U6144 ( .A1(n5871), .A2(n7083), .ZN(n7086) );
  NAND2_X2 U6145 ( .A1(n4637), .A2(n5726), .ZN(n5739) );
  NAND2_X1 U6146 ( .A1(n5713), .A2(n4369), .ZN(n4637) );
  NAND3_X1 U6147 ( .A1(n4638), .A2(n6068), .A3(n8016), .ZN(n7699) );
  NAND2_X1 U6148 ( .A1(n5717), .A2(n4640), .ZN(n4639) );
  OAI21_X2 U6149 ( .B1(n7984), .B2(n7501), .A(n7502), .ZN(n7971) );
  NAND2_X1 U6150 ( .A1(n6257), .A2(n6256), .ZN(n7548) );
  NAND3_X1 U6151 ( .A1(n5822), .A2(n6862), .A3(n5821), .ZN(n6865) );
  NAND2_X2 U6152 ( .A1(n7314), .A2(n5979), .ZN(n7337) );
  OAI21_X1 U6153 ( .B1(n8308), .B2(n8307), .A(n8495), .ZN(n8312) );
  INV_X1 U6154 ( .A(n4652), .ZN(n5055) );
  NAND3_X1 U6155 ( .A1(n4650), .A2(n4345), .A3(n4652), .ZN(n8386) );
  OAI21_X2 U6156 ( .B1(n8356), .B2(n4656), .A(n4654), .ZN(n8323) );
  NAND2_X1 U6157 ( .A1(n5334), .A2(n4662), .ZN(n4658) );
  NAND2_X1 U6158 ( .A1(n4658), .A2(n4659), .ZN(n8347) );
  NAND2_X1 U6159 ( .A1(n7061), .A2(n4671), .ZN(n4670) );
  OAI21_X2 U6160 ( .B1(n5296), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5342) );
  OAI21_X1 U6161 ( .B1(n7892), .B2(n9769), .A(n4680), .ZN(P2_U3200) );
  AND2_X1 U6162 ( .A1(n4684), .A2(n4681), .ZN(n4680) );
  OAI21_X1 U6163 ( .B1(n7900), .B2(n4314), .A(n7920), .ZN(n4684) );
  NAND3_X1 U6164 ( .A1(n5771), .A2(n5777), .A3(n5770), .ZN(n4685) );
  NAND2_X1 U6165 ( .A1(n6458), .A2(n4368), .ZN(n4691) );
  NAND3_X1 U6166 ( .A1(n4695), .A2(n4865), .A3(n4697), .ZN(n6423) );
  NAND3_X1 U6167 ( .A1(n4698), .A2(n4696), .A3(n6384), .ZN(n4695) );
  INV_X1 U6168 ( .A(n4705), .ZN(n7790) );
  INV_X1 U6169 ( .A(n7791), .ZN(n4704) );
  INV_X1 U6170 ( .A(n4710), .ZN(n7157) );
  INV_X1 U6171 ( .A(n7128), .ZN(n4709) );
  INV_X1 U6172 ( .A(n4322), .ZN(n4712) );
  NAND2_X1 U6173 ( .A1(n4723), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U6174 ( .A1(n4723), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6175 ( .A1(n4723), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U6176 ( .A1(n4723), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U6177 ( .A1(n4723), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6178 ( .A1(n4723), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6179 ( .A1(n4723), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6180 ( .A1(n4723), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6181 ( .A1(n4723), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6182 ( .A1(n4723), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6183 ( .A1(n4723), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6184 ( .A1(n4723), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6185 ( .A1(n4723), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6186 ( .A1(n4723), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6187 ( .A1(n4723), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6188 ( .A1(n4723), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6189 ( .A1(n4723), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6190 ( .A1(n4723), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U6191 ( .A1(n9177), .A2(n9702), .ZN(n4724) );
  XNOR2_X1 U6192 ( .A(n4725), .B(n4483), .ZN(n9177) );
  NAND2_X1 U6193 ( .A1(n8953), .A2(n8952), .ZN(n4725) );
  NAND2_X1 U6194 ( .A1(n7042), .A2(n8515), .ZN(n7045) );
  INV_X1 U6195 ( .A(n9125), .ZN(n4733) );
  NAND2_X1 U6196 ( .A1(n4729), .A2(n4730), .ZN(n9063) );
  NAND2_X1 U6197 ( .A1(n9125), .A2(n4309), .ZN(n4729) );
  AND2_X1 U6198 ( .A1(n9239), .A2(n8921), .ZN(n4742) );
  NAND2_X1 U6199 ( .A1(n9541), .A2(n4760), .ZN(n4759) );
  NAND3_X1 U6200 ( .A1(n4759), .A2(n4758), .A3(n4365), .ZN(n7194) );
  NAND2_X1 U6201 ( .A1(n4894), .A2(n4893), .ZN(n4898) );
  NAND2_X1 U6202 ( .A1(n5263), .A2(n4773), .ZN(n5296) );
  INV_X1 U6203 ( .A(n4776), .ZN(n7363) );
  NAND2_X1 U6204 ( .A1(n5361), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U6205 ( .A1(n5424), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U6206 ( .A1(n4793), .A2(n4791), .ZN(n5115) );
  INV_X1 U6207 ( .A(n5283), .ZN(n5285) );
  NAND3_X1 U6208 ( .A1(n7523), .A2(n7582), .A3(n4809), .ZN(n7525) );
  NAND2_X1 U6209 ( .A1(n5515), .A2(n5514), .ZN(n5531) );
  NAND2_X1 U6210 ( .A1(n4810), .A2(n4814), .ZN(n5560) );
  NAND2_X1 U6211 ( .A1(n5515), .A2(n4811), .ZN(n4810) );
  NAND3_X1 U6212 ( .A1(n4820), .A2(n4818), .A3(n7550), .ZN(n4817) );
  NAND3_X1 U6213 ( .A1(n7534), .A2(n7535), .A3(n7529), .ZN(n4820) );
  NAND2_X1 U6214 ( .A1(n4821), .A2(n6184), .ZN(n6956) );
  AOI21_X1 U6215 ( .B1(n8124), .B2(n4821), .A(n8123), .ZN(n8125) );
  NAND2_X1 U6216 ( .A1(n6183), .A2(n6182), .ZN(n4821) );
  NAND2_X1 U6217 ( .A1(n7991), .A2(n4824), .ZN(n4823) );
  NOR2_X1 U6218 ( .A1(n8231), .A2(n8003), .ZN(n4835) );
  NAND2_X1 U6219 ( .A1(n6816), .A2(n4841), .ZN(n4839) );
  NAND2_X1 U6220 ( .A1(n4839), .A2(n4840), .ZN(n6936) );
  AOI21_X1 U6221 ( .B1(n4841), .B2(n4310), .A(n4347), .ZN(n4840) );
  NAND2_X1 U6222 ( .A1(n4842), .A2(n4843), .ZN(n6876) );
  AND2_X1 U6223 ( .A1(n4843), .A2(n4328), .ZN(n4841) );
  OAI21_X1 U6224 ( .B1(n6195), .B2(n4310), .A(n6196), .ZN(n4844) );
  NAND2_X2 U6225 ( .A1(n4847), .A2(n4845), .ZN(n8014) );
  NAND3_X1 U6226 ( .A1(n8025), .A2(n4363), .A3(n8036), .ZN(n4846) );
  NAND2_X1 U6227 ( .A1(n8037), .A2(n4848), .ZN(n4847) );
  INV_X1 U6228 ( .A(n4849), .ZN(n8039) );
  INV_X2 U6229 ( .A(n6180), .ZN(n9783) );
  OAI211_X2 U6230 ( .C1(n4783), .C2(n7543), .A(n4346), .B(n4850), .ZN(n6180)
         );
  OAI21_X1 U6231 ( .B1(n7206), .B2(n6204), .A(n6203), .ZN(n7258) );
  NAND2_X1 U6232 ( .A1(n6204), .A2(n6203), .ZN(n4855) );
  NOR2_X2 U6233 ( .A1(n5695), .A2(n4859), .ZN(n5707) );
  NAND2_X1 U6234 ( .A1(n5765), .A2(n5764), .ZN(n6657) );
  INV_X1 U6235 ( .A(n7602), .ZN(n7604) );
  NAND2_X1 U6236 ( .A1(n4922), .A2(n4921), .ZN(n4934) );
  NOR2_X1 U6237 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4879) );
  XNOR2_X1 U6238 ( .A(n6774), .B(n8707), .ZN(n6773) );
  AOI21_X1 U6239 ( .B1(n6751), .B2(n4943), .A(n4870), .ZN(n4944) );
  NAND2_X1 U6240 ( .A1(n7537), .A2(n7536), .ZN(n7541) );
  NAND2_X1 U6241 ( .A1(n5749), .A2(n4851), .ZN(n5751) );
  NOR2_X1 U6242 ( .A1(n6143), .A2(n6144), .ZN(n7620) );
  NAND2_X1 U6243 ( .A1(n7722), .A2(n6111), .ZN(n6143) );
  XNOR2_X1 U6244 ( .A(n6130), .B(n6129), .ZN(n6301) );
  NAND2_X1 U6245 ( .A1(n5742), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5746) );
  OR2_X2 U6246 ( .A1(n5682), .A2(n5681), .ZN(n5744) );
  OR2_X1 U6247 ( .A1(n5789), .A2(n5740), .ZN(n5747) );
  NAND2_X1 U6248 ( .A1(n4952), .A2(n8613), .ZN(n5000) );
  XNOR2_X2 U6249 ( .A(n5003), .B(n4976), .ZN(n5001) );
  AOI21_X2 U6250 ( .B1(n7677), .B2(n7657), .A(n7656), .ZN(n7725) );
  AOI22_X1 U6251 ( .A1(n7194), .A2(n8646), .B1(n9688), .B2(n7193), .ZN(n8912)
         );
  INV_X1 U6252 ( .A(n5681), .ZN(n5757) );
  AND2_X2 U6253 ( .A1(n6709), .A2(n8106), .ZN(n8080) );
  AND2_X1 U6254 ( .A1(n6512), .A2(n5626), .ZN(n9621) );
  INV_X1 U6255 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4923) );
  AND2_X1 U6256 ( .A1(n5760), .A2(n5759), .ZN(n4861) );
  INV_X1 U6257 ( .A(n9308), .ZN(n9300) );
  NAND2_X1 U6258 ( .A1(n6108), .A2(n6107), .ZN(n7963) );
  AND2_X1 U6259 ( .A1(n5016), .A2(n4880), .ZN(n4862) );
  AND2_X1 U6260 ( .A1(n5256), .A2(n5255), .ZN(n4863) );
  AND3_X1 U6261 ( .A1(n5629), .A2(n8495), .A3(n5628), .ZN(n4864) );
  AND2_X1 U6262 ( .A1(n9182), .A2(n9181), .ZN(n4867) );
  OR2_X1 U6263 ( .A1(n7928), .A2(n8271), .ZN(n4868) );
  AND4_X1 U6264 ( .A1(n7585), .A2(n7584), .A3(n7583), .A4(n7582), .ZN(n4869)
         );
  AND2_X1 U6265 ( .A1(n4946), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4870) );
  AND2_X1 U6266 ( .A1(n5621), .A2(n5624), .ZN(n4871) );
  OR2_X1 U6267 ( .A1(n7543), .A2(n8293), .ZN(n4872) );
  AND2_X1 U6268 ( .A1(n6237), .A2(n6236), .ZN(n8123) );
  INV_X1 U6269 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5341) );
  AND2_X1 U6270 ( .A1(n8279), .A2(n8097), .ZN(n4874) );
  OR2_X1 U6271 ( .A1(n8279), .A2(n8097), .ZN(n4875) );
  OR2_X1 U6272 ( .A1(n9052), .A2(n8934), .ZN(n4876) );
  AND2_X1 U6273 ( .A1(n5653), .A2(n5652), .ZN(n4877) );
  AND2_X1 U6274 ( .A1(n8424), .A2(n5152), .ZN(n4878) );
  NAND2_X2 U6275 ( .A1(n6741), .A2(n9602), .ZN(n9138) );
  INV_X1 U6276 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5669) );
  INV_X1 U6277 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5667) );
  INV_X1 U6278 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5673) );
  INV_X1 U6279 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4880) );
  OAI211_X1 U6280 ( .C1(n7946), .C2(n4354), .A(n7549), .B(n4296), .ZN(n7534)
         );
  INV_X1 U6281 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U6282 ( .A1(n5757), .A2(n6405), .ZN(n5758) );
  INV_X1 U6283 ( .A(n5035), .ZN(n5036) );
  INV_X1 U6284 ( .A(n8888), .ZN(n8889) );
  NAND2_X1 U6285 ( .A1(n4306), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6286 ( .A1(n4713), .A2(n6852), .ZN(n6832) );
  INV_X1 U6287 ( .A(n7564), .ZN(n6193) );
  INV_X1 U6288 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6289 ( .A1(n9065), .A2(n8890), .ZN(n8892) );
  OR2_X1 U6290 ( .A1(n6774), .A2(n9620), .ZN(n6775) );
  INV_X1 U6291 ( .A(n7242), .ZN(n5886) );
  INV_X1 U6292 ( .A(n6852), .ZN(n6456) );
  NOR2_X1 U6293 ( .A1(n5920), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5919) );
  NOR2_X1 U6294 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5697) );
  OAI21_X1 U6295 ( .B1(n5154), .B2(n8424), .A(n5153), .ZN(n5155) );
  INV_X1 U6296 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5317) );
  INV_X1 U6297 ( .A(n5452), .ZN(n5451) );
  INV_X1 U6298 ( .A(n5348), .ZN(n5346) );
  INV_X1 U6299 ( .A(n4952), .ZN(n5120) );
  OR2_X1 U6300 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  INV_X1 U6301 ( .A(SI_25_), .ZN(n9906) );
  INV_X1 U6302 ( .A(SI_9_), .ZN(n5116) );
  INV_X1 U6303 ( .A(n7963), .ZN(n6110) );
  NOR2_X1 U6304 ( .A1(n6072), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6071) );
  AND2_X1 U6305 ( .A1(n6023), .A2(n7693), .ZN(n6033) );
  OR2_X1 U6306 ( .A1(n6059), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6061) );
  OR2_X1 U6307 ( .A1(n5956), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5967) );
  OR2_X1 U6308 ( .A1(n5889), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5908) );
  INV_X1 U6309 ( .A(n8062), .ZN(n8041) );
  INV_X1 U6310 ( .A(n8781), .ZN(n8913) );
  OR2_X1 U6311 ( .A1(n5474), .A2(n8329), .ZN(n5498) );
  NAND2_X1 U6312 ( .A1(n9186), .A2(n8951), .ZN(n8952) );
  NAND2_X1 U6313 ( .A1(n5408), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5428) );
  INV_X1 U6314 ( .A(n5270), .ZN(n5269) );
  OR2_X1 U6315 ( .A1(n9520), .A2(n8915), .ZN(n8916) );
  AND2_X1 U6316 ( .A1(n5490), .A2(n5468), .ZN(n5469) );
  INV_X1 U6317 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5366) );
  AND2_X1 U6318 ( .A1(n5844), .A2(n7089), .ZN(n5864) );
  INV_X1 U6319 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5656) );
  INV_X1 U6320 ( .A(n6927), .ZN(n5837) );
  OR2_X1 U6321 ( .A1(n6159), .A2(n6158), .ZN(n7731) );
  OAI21_X1 U6322 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7590) );
  OR2_X1 U6323 ( .A1(n5741), .A2(n6414), .ZN(n5790) );
  INV_X1 U6324 ( .A(n7980), .ZN(n8003) );
  AND2_X1 U6325 ( .A1(n6873), .A2(n7428), .ZN(n7566) );
  AND2_X1 U6326 ( .A1(n6271), .A2(n6288), .ZN(n8127) );
  INV_X1 U6327 ( .A(n6115), .ZN(n6139) );
  INV_X1 U6328 ( .A(n7956), .ZN(n7732) );
  INV_X1 U6329 ( .A(n7964), .ZN(n7993) );
  AND2_X1 U6330 ( .A1(n7448), .A2(n7447), .ZN(n7573) );
  INV_X1 U6331 ( .A(n6946), .ZN(n7560) );
  OR2_X1 U6332 ( .A1(n6112), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6114) );
  INV_X1 U6333 ( .A(n5980), .ZN(n5981) );
  AND2_X1 U6334 ( .A1(n8406), .A2(n5488), .ZN(n8324) );
  INV_X1 U6335 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7253) );
  AND2_X1 U6336 ( .A1(n5038), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5056) );
  AND2_X1 U6337 ( .A1(n5511), .A2(n5509), .ZN(n8407) );
  INV_X1 U6338 ( .A(n8506), .ZN(n8459) );
  AND2_X1 U6339 ( .A1(n5056), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5080) );
  OR2_X1 U6340 ( .A1(n9621), .A2(n8697), .ZN(n5627) );
  NAND2_X1 U6341 ( .A1(n8760), .A2(n8759), .ZN(n8761) );
  INV_X1 U6342 ( .A(n5640), .ZN(n6637) );
  OR2_X1 U6343 ( .A1(n9386), .A2(n9382), .ZN(n9476) );
  OR2_X1 U6344 ( .A1(n9386), .A2(n6637), .ZN(n9501) );
  NAND2_X1 U6345 ( .A1(n5269), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6346 ( .A1(n5181), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6347 ( .A1(n9616), .A2(n9534), .ZN(n9605) );
  AND2_X1 U6348 ( .A1(n5640), .A2(n8697), .ZN(n8878) );
  INV_X1 U6349 ( .A(n8928), .ZN(n8929) );
  NOR2_X1 U6350 ( .A1(n5188), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5212) );
  AND2_X1 U6351 ( .A1(n6292), .A2(n6160), .ZN(n7729) );
  NAND2_X1 U6352 ( .A1(n5751), .A2(n5766), .ZN(n6659) );
  INV_X1 U6353 ( .A(n7731), .ZN(n7680) );
  INV_X1 U6354 ( .A(n7707), .ZN(n7726) );
  AND2_X1 U6355 ( .A1(n6597), .A2(n6234), .ZN(n7740) );
  AND4_X1 U6356 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n7644)
         );
  AND4_X1 U6357 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n7647)
         );
  INV_X1 U6358 ( .A(n7917), .ZN(n9767) );
  INV_X1 U6359 ( .A(n7968), .ZN(n8111) );
  INV_X1 U6360 ( .A(n8118), .ZN(n8099) );
  OR2_X1 U6361 ( .A1(n9824), .A2(n8129), .ZN(n7968) );
  INV_X1 U6362 ( .A(n9824), .ZN(n9836) );
  INV_X1 U6363 ( .A(n8180), .ZN(n8192) );
  NAND2_X1 U6364 ( .A1(n6273), .A2(n6139), .ZN(n6283) );
  NAND2_X1 U6365 ( .A1(n7102), .A2(n7588), .ZN(n9824) );
  NAND2_X1 U6366 ( .A1(n7076), .A2(n9826), .ZN(n9807) );
  AND2_X1 U6367 ( .A1(n7102), .A2(n8129), .ZN(n9791) );
  NAND2_X1 U6368 ( .A1(n6300), .A2(n6359), .ZN(n6278) );
  INV_X1 U6369 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5900) );
  NOR2_X1 U6370 ( .A1(n5132), .A2(n7253), .ZN(n5133) );
  NAND2_X1 U6371 ( .A1(n5639), .A2(n8770), .ZN(n8475) );
  NOR2_X1 U6372 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  AND2_X1 U6373 ( .A1(n5600), .A2(n5599), .ZN(n8949) );
  OR2_X1 U6374 ( .A1(n5394), .A2(n5393), .ZN(n8926) );
  INV_X1 U6375 ( .A(n6342), .ZN(n9321) );
  INV_X1 U6376 ( .A(n9479), .ZN(n9497) );
  INV_X1 U6377 ( .A(n9501), .ZN(n9485) );
  INV_X1 U6378 ( .A(n9602), .ZN(n9581) );
  INV_X1 U6379 ( .A(n9153), .ZN(n9590) );
  AOI21_X1 U6380 ( .B1(n5618), .B2(n10007), .A(n6339), .ZN(n6574) );
  AND2_X1 U6381 ( .A1(n8992), .A2(n8681), .ZN(n9009) );
  AND2_X1 U6382 ( .A1(n8669), .A2(n8737), .ZN(n9143) );
  AND2_X1 U6383 ( .A1(n6739), .A2(n6519), .ZN(n6575) );
  AND2_X1 U6384 ( .A1(n5140), .A2(n5139), .ZN(n6563) );
  AND2_X1 U6385 ( .A1(n4302), .A2(P1_U3086), .ZN(n7215) );
  NAND2_X1 U6386 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  AND2_X1 U6387 ( .A1(n6142), .A2(n6141), .ZN(n7707) );
  INV_X1 U6388 ( .A(n7734), .ZN(n7341) );
  NAND2_X1 U6389 ( .A1(n6152), .A2(n6151), .ZN(n7946) );
  INV_X1 U6390 ( .A(n7338), .ZN(n8077) );
  INV_X1 U6391 ( .A(n7644), .ZN(n7743) );
  OR2_X1 U6392 ( .A1(P2_U3150), .A2(n6400), .ZN(n9779) );
  INV_X1 U6393 ( .A(n7920), .ZN(n9762) );
  OR2_X1 U6394 ( .A1(n8080), .A2(n6813), .ZN(n8088) );
  OR2_X1 U6395 ( .A1(n6709), .A2(n7968), .ZN(n8092) );
  NAND2_X1 U6396 ( .A1(n9849), .A2(n9836), .ZN(n8180) );
  NAND2_X1 U6397 ( .A1(n9849), .A2(n9807), .ZN(n8189) );
  INV_X1 U6398 ( .A(n9849), .ZN(n9847) );
  OR2_X1 U6399 ( .A1(n7551), .A2(n7377), .ZN(n9369) );
  OR2_X1 U6400 ( .A1(n9886), .A2(n9824), .ZN(n8271) );
  OR2_X1 U6401 ( .A1(n9886), .A2(n9841), .ZN(n8273) );
  INV_X2 U6402 ( .A(n9886), .ZN(n9884) );
  AND2_X1 U6403 ( .A1(n8285), .A2(n6112), .ZN(n6356) );
  INV_X1 U6404 ( .A(n6356), .ZN(n6347) );
  INV_X1 U6405 ( .A(n6478), .ZN(n8300) );
  INV_X1 U6406 ( .A(n4295), .ZN(n8419) );
  INV_X1 U6407 ( .A(n8475), .ZN(n8508) );
  INV_X1 U6408 ( .A(n8495), .ZN(n8511) );
  INV_X1 U6409 ( .A(n8945), .ZN(n8946) );
  OR2_X1 U6410 ( .A1(n5325), .A2(n5324), .ZN(n8919) );
  OR2_X1 U6411 ( .A1(n9386), .A2(n6541), .ZN(n9479) );
  NAND2_X1 U6412 ( .A1(n6514), .A2(n5633), .ZN(n9602) );
  NAND2_X1 U6413 ( .A1(n9738), .A2(n9702), .ZN(n9247) );
  AND2_X2 U6414 ( .A1(n6575), .A2(n6574), .ZN(n9738) );
  INV_X1 U6415 ( .A(n9738), .ZN(n9735) );
  NAND2_X1 U6416 ( .A1(n9714), .A2(n9702), .ZN(n9295) );
  INV_X1 U6417 ( .A(n9714), .ZN(n9712) );
  AND2_X1 U6418 ( .A1(n9311), .A2(n7232), .ZN(n6339) );
  INV_X1 U6419 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7288) );
  INV_X1 U6420 ( .A(n8708), .ZN(n8637) );
  INV_X1 U6421 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6600) );
  INV_X1 U6422 ( .A(n7878), .ZN(P2_U3893) );
  NOR2_X1 U6423 ( .A1(n6299), .A2(n6298), .ZN(P1_U3973) );
  NOR2_X2 U6424 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4977) );
  NAND2_X1 U6425 ( .A1(n4977), .A2(n4879), .ZN(n5015) );
  INV_X1 U6426 ( .A(n5015), .ZN(n4881) );
  NOR2_X1 U6427 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4885) );
  NAND4_X1 U6428 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4886)
         );
  INV_X1 U6429 ( .A(n4894), .ZN(n4891) );
  NAND2_X1 U6430 ( .A1(n4891), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4892) );
  INV_X1 U6431 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4899) );
  NAND2_X2 U6432 ( .A1(n4900), .A2(n5620), .ZN(n6299) );
  NAND2_X1 U6433 ( .A1(n5342), .A2(n4901), .ZN(n4902) );
  NAND2_X1 U6434 ( .A1(n4902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6435 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  NAND2_X1 U6436 ( .A1(n4906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U6437 ( .A1(n4905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U6438 ( .A1(n5626), .A2(n6749), .ZN(n4910) );
  NAND2_X1 U6439 ( .A1(n6509), .A2(n4910), .ZN(n4911) );
  XNOR2_X1 U6440 ( .A(n4922), .B(n4926), .ZN(n5640) );
  NAND2_X1 U6441 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4914) );
  NAND2_X1 U6442 ( .A1(n4915), .A2(n4914), .ZN(n4916) );
  NAND2_X1 U6443 ( .A1(n8613), .A2(SI_0_), .ZN(n4919) );
  XNOR2_X1 U6444 ( .A(n4919), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U6445 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4921) );
  INV_X1 U6446 ( .A(n4925), .ZN(n4928) );
  AND3_X1 U6447 ( .A1(n4933), .A2(n4923), .A3(n4926), .ZN(n4927) );
  NAND2_X1 U6448 ( .A1(n4928), .A2(n4927), .ZN(n9298) );
  NOR2_X1 U6449 ( .A1(n4930), .A2(n4929), .ZN(n4931) );
  NAND2_X1 U6450 ( .A1(n4932), .A2(n4931), .ZN(n4937) );
  NAND2_X1 U6451 ( .A1(n5594), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U6452 ( .A1(n8620), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U6453 ( .A1(n5040), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4938) );
  INV_X1 U6454 ( .A(n6749), .ZN(n4942) );
  INV_X1 U6455 ( .A(n6299), .ZN(n4946) );
  INV_X1 U6456 ( .A(n4944), .ZN(n4945) );
  NOR2_X1 U6457 ( .A1(n4947), .A2(n4945), .ZN(n6374) );
  AOI222_X1 U6458 ( .A1(n6751), .A2(n5551), .B1(n6756), .B2(n5456), .C1(n9384), 
        .C2(n4946), .ZN(n6373) );
  OAI22_X1 U6459 ( .A1(n6374), .A2(n6373), .B1(n4947), .B2(n4297), .ZN(n6621)
         );
  NAND2_X1 U6460 ( .A1(n5594), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6461 ( .A1(n8620), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6462 ( .A1(n5040), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4948) );
  NAND4_X2 U6463 ( .A1(n4951), .A2(n4950), .A3(n4949), .A4(n4948), .ZN(n6774)
         );
  NAND2_X1 U6464 ( .A1(n6774), .A2(n4943), .ZN(n4958) );
  NAND2_X1 U6465 ( .A1(n4952), .A2(n4298), .ZN(n4999) );
  INV_X1 U6466 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6314) );
  OR2_X1 U6467 ( .A1(n4999), .A2(n6314), .ZN(n4957) );
  NAND2_X1 U6468 ( .A1(n5120), .A2(n4300), .ZN(n4956) );
  AND2_X1 U6469 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6470 ( .A1(n4298), .A2(n4953), .ZN(n5754) );
  NAND2_X1 U6471 ( .A1(n5754), .A2(n4954), .ZN(n4969) );
  XNOR2_X1 U6472 ( .A(n4970), .B(n4969), .ZN(n6317) );
  XNOR2_X1 U6473 ( .A(n4959), .B(n5602), .ZN(n4961) );
  AOI22_X1 U6474 ( .A1(n6774), .A2(n5551), .B1(n9620), .B2(n5456), .ZN(n4960)
         );
  NAND2_X1 U6475 ( .A1(n4961), .A2(n4960), .ZN(n4963) );
  INV_X1 U6476 ( .A(n4963), .ZN(n6630) );
  NAND2_X1 U6477 ( .A1(n5594), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6478 ( .A1(n8620), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U6479 ( .A1(n5040), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6480 ( .A1(n8791), .A2(n5456), .ZN(n4983) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4968) );
  OR2_X1 U6482 ( .A1(n4999), .A2(n4968), .ZN(n4981) );
  NAND2_X1 U6483 ( .A1(n4970), .A2(n4969), .ZN(n4974) );
  INV_X1 U6484 ( .A(n4971), .ZN(n4972) );
  NAND2_X1 U6485 ( .A1(n4972), .A2(SI_1_), .ZN(n4973) );
  NAND2_X1 U6486 ( .A1(n4974), .A2(n4973), .ZN(n5002) );
  MUX2_X1 U6487 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4302), .Z(n5003) );
  INV_X1 U6488 ( .A(SI_2_), .ZN(n4976) );
  XNOR2_X1 U6489 ( .A(n5002), .B(n5001), .ZN(n6315) );
  OR2_X1 U6490 ( .A1(n5000), .A2(n6315), .ZN(n4980) );
  OR2_X1 U6491 ( .A1(n4977), .A2(n4899), .ZN(n4978) );
  NAND2_X1 U6492 ( .A1(n5120), .A2(n6646), .ZN(n4979) );
  AOI22_X1 U6493 ( .A1(n8791), .A2(n5551), .B1(n6792), .B2(n4943), .ZN(n4985)
         );
  NAND2_X1 U6494 ( .A1(n4984), .A2(n4985), .ZN(n4989) );
  INV_X1 U6495 ( .A(n4984), .ZN(n4987) );
  INV_X1 U6496 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6497 ( .A1(n4987), .A2(n4986), .ZN(n4988) );
  AND2_X1 U6498 ( .A1(n4989), .A2(n4988), .ZN(n6629) );
  NAND2_X1 U6499 ( .A1(n6628), .A2(n4989), .ZN(n6686) );
  INV_X1 U6500 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n4990) );
  OAI22_X1 U6501 ( .A1(n5131), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n5372), .B2(
        n4990), .ZN(n4991) );
  INV_X1 U6502 ( .A(n4991), .ZN(n4996) );
  INV_X1 U6503 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6791) );
  INV_X1 U6504 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U6505 ( .A1(n5645), .A2(n6791), .B1(n5476), .B2(n4993), .ZN(n4994)
         );
  INV_X1 U6506 ( .A(n4994), .ZN(n4995) );
  INV_X1 U6507 ( .A(n8790), .ZN(n6779) );
  OR3_X1 U6508 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        n9384), .ZN(n4997) );
  NAND2_X1 U6509 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4997), .ZN(n4998) );
  INV_X1 U6510 ( .A(n9350), .ZN(n6307) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6308) );
  OR2_X1 U6512 ( .A1(n4999), .A2(n6308), .ZN(n5006) );
  NAND2_X1 U6513 ( .A1(n5003), .A2(SI_2_), .ZN(n5004) );
  INV_X1 U6514 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6322) );
  XNOR2_X1 U6515 ( .A(n5021), .B(SI_3_), .ZN(n5019) );
  XNOR2_X1 U6516 ( .A(n5020), .B(n5019), .ZN(n6321) );
  OR2_X1 U6517 ( .A1(n5000), .A2(n6321), .ZN(n5005) );
  OAI22_X1 U6518 ( .A1(n6779), .A2(n5601), .B1(n9637), .B2(n5550), .ZN(n5030)
         );
  NAND2_X1 U6519 ( .A1(n8790), .A2(n5456), .ZN(n5008) );
  NAND2_X1 U6520 ( .A1(n6796), .A2(n5567), .ZN(n5007) );
  NAND2_X1 U6521 ( .A1(n5008), .A2(n5007), .ZN(n5009) );
  XNOR2_X1 U6522 ( .A(n5009), .B(n4297), .ZN(n5029) );
  XOR2_X1 U6523 ( .A(n5030), .B(n5029), .Z(n6687) );
  NAND2_X1 U6524 ( .A1(n6686), .A2(n6687), .ZN(n6685) );
  NOR2_X1 U6525 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5010) );
  NOR2_X1 U6526 ( .A1(n5038), .A2(n5010), .ZN(n9582) );
  NAND2_X1 U6527 ( .A1(n5594), .A2(n9582), .ZN(n5013) );
  NAND2_X1 U6528 ( .A1(n8620), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6529 ( .A1(n5040), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5011) );
  NAND4_X1 U6530 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n8789)
         );
  NAND2_X1 U6531 ( .A1(n8789), .A2(n5456), .ZN(n5026) );
  NAND2_X1 U6532 ( .A1(n5015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6533 ( .A1(n5017), .A2(n5016), .ZN(n5045) );
  OR2_X1 U6534 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  INV_X1 U6535 ( .A(n6552), .ZN(n9398) );
  OR2_X1 U6536 ( .A1(n4999), .A2(n6310), .ZN(n5024) );
  INV_X1 U6537 ( .A(n5021), .ZN(n5022) );
  XNOR2_X1 U6538 ( .A(n5048), .B(SI_4_), .ZN(n5047) );
  OR2_X1 U6539 ( .A1(n5000), .A2(n6311), .ZN(n5023) );
  OAI211_X1 U6540 ( .C1(n8615), .C2(n9398), .A(n5024), .B(n5023), .ZN(n6903)
         );
  NAND2_X1 U6541 ( .A1(n6903), .A2(n5567), .ZN(n5025) );
  NAND2_X1 U6542 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  XNOR2_X1 U6543 ( .A(n5027), .B(n4297), .ZN(n5034) );
  AND2_X1 U6544 ( .A1(n6903), .A2(n5456), .ZN(n5028) );
  AOI21_X1 U6545 ( .B1(n8789), .B2(n5551), .A(n5028), .ZN(n5035) );
  XNOR2_X1 U6546 ( .A(n5034), .B(n5035), .ZN(n6717) );
  INV_X1 U6547 ( .A(n5029), .ZN(n5032) );
  INV_X1 U6548 ( .A(n5030), .ZN(n5031) );
  NAND2_X1 U6549 ( .A1(n5032), .A2(n5031), .ZN(n6715) );
  AND2_X1 U6550 ( .A1(n6717), .A2(n6715), .ZN(n5033) );
  NAND2_X1 U6551 ( .A1(n5034), .A2(n5036), .ZN(n5037) );
  NOR2_X1 U6552 ( .A1(n5038), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U6553 ( .A1(n5056), .A2(n5039), .ZN(n8392) );
  NAND2_X1 U6554 ( .A1(n5594), .A2(n8392), .ZN(n5044) );
  NAND2_X1 U6555 ( .A1(n8620), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6556 ( .A1(n5040), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6557 ( .A1(n5045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5046) );
  XNOR2_X1 U6558 ( .A(n5046), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6555) );
  INV_X1 U6559 ( .A(n6555), .ZN(n9414) );
  INV_X1 U6560 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6561 ( .A1(n5049), .A2(SI_4_), .ZN(n5050) );
  XNOR2_X1 U6562 ( .A(n5066), .B(SI_5_), .ZN(n5064) );
  XNOR2_X1 U6563 ( .A(n5065), .B(n5064), .ZN(n6319) );
  OR2_X1 U6564 ( .A1(n5000), .A2(n6319), .ZN(n5053) );
  OR2_X1 U6565 ( .A1(n4999), .A2(n6320), .ZN(n5052) );
  OAI211_X1 U6566 ( .C1(n8615), .C2(n9414), .A(n5053), .B(n5052), .ZN(n8393)
         );
  AOI22_X1 U6567 ( .A1(n8788), .A2(n5456), .B1(n8393), .B2(n5567), .ZN(n5054)
         );
  AOI22_X1 U6568 ( .A1(n8788), .A2(n5551), .B1(n5456), .B2(n8393), .ZN(n8388)
         );
  NAND2_X1 U6569 ( .A1(n8386), .A2(n4652), .ZN(n6972) );
  NOR2_X1 U6570 ( .A1(n5056), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U6571 ( .A1(n5080), .A2(n5057), .ZN(n9564) );
  NAND2_X1 U6572 ( .A1(n5594), .A2(n9564), .ZN(n5061) );
  NAND2_X1 U6573 ( .A1(n5040), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6574 ( .A1(n8620), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5058) );
  NAND4_X1 U6575 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n8787)
         );
  NAND2_X1 U6576 ( .A1(n8787), .A2(n5456), .ZN(n5072) );
  NAND2_X1 U6577 ( .A1(n5062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5063) );
  XNOR2_X1 U6578 ( .A(n5063), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6557) );
  INV_X1 U6579 ( .A(n6557), .ZN(n9429) );
  INV_X1 U6580 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6581 ( .A1(n5067), .A2(SI_5_), .ZN(n5068) );
  XNOR2_X1 U6582 ( .A(n5089), .B(SI_6_), .ZN(n5087) );
  XNOR2_X1 U6583 ( .A(n5088), .B(n5087), .ZN(n6324) );
  OR2_X1 U6584 ( .A1(n5000), .A2(n6324), .ZN(n5070) );
  OR2_X1 U6585 ( .A1(n4999), .A2(n6323), .ZN(n5069) );
  OAI211_X1 U6586 ( .C1(n8615), .C2(n9429), .A(n5070), .B(n5069), .ZN(n6919)
         );
  NAND2_X1 U6587 ( .A1(n6919), .A2(n5567), .ZN(n5071) );
  NAND2_X1 U6588 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  XNOR2_X1 U6589 ( .A(n5073), .B(n4297), .ZN(n5076) );
  NAND2_X1 U6590 ( .A1(n8787), .A2(n5551), .ZN(n5075) );
  NAND2_X1 U6591 ( .A1(n6919), .A2(n5456), .ZN(n5074) );
  NAND2_X1 U6592 ( .A1(n5075), .A2(n5074), .ZN(n5077) );
  NAND2_X1 U6593 ( .A1(n5076), .A2(n5077), .ZN(n6973) );
  NAND2_X1 U6594 ( .A1(n6972), .A2(n6973), .ZN(n6971) );
  INV_X1 U6595 ( .A(n5076), .ZN(n5079) );
  INV_X1 U6596 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6597 ( .A1(n5079), .A2(n5078), .ZN(n6975) );
  NAND2_X1 U6598 ( .A1(n5080), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5132) );
  OAI21_X1 U6599 ( .B1(n5080), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5132), .ZN(
        n5081) );
  INV_X1 U6600 ( .A(n5081), .ZN(n7065) );
  NAND2_X1 U6601 ( .A1(n5594), .A2(n7065), .ZN(n5085) );
  NAND2_X1 U6602 ( .A1(n5040), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6603 ( .A1(n8620), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5082) );
  NAND4_X1 U6604 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n8786)
         );
  NOR2_X1 U6605 ( .A1(n5062), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6606 ( .A1(n5122), .A2(n4899), .ZN(n5086) );
  XNOR2_X1 U6607 ( .A(n5086), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6560) );
  INV_X1 U6608 ( .A(n6560), .ZN(n9335) );
  INV_X1 U6609 ( .A(n5089), .ZN(n5090) );
  XNOR2_X1 U6610 ( .A(n5108), .B(SI_7_), .ZN(n5105) );
  XNOR2_X1 U6611 ( .A(n5107), .B(n5105), .ZN(n5841) );
  INV_X1 U6612 ( .A(n5841), .ZN(n6327) );
  OR2_X1 U6613 ( .A1(n5000), .A2(n6327), .ZN(n5092) );
  INV_X1 U6614 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6328) );
  OR2_X1 U6615 ( .A1(n8603), .A2(n6328), .ZN(n5091) );
  OAI211_X1 U6616 ( .C1(n8615), .C2(n9335), .A(n5092), .B(n5091), .ZN(n6920)
         );
  OAI22_X1 U6617 ( .A1(n7043), .A2(n5601), .B1(n9662), .B2(n5550), .ZN(n5097)
         );
  NAND2_X1 U6618 ( .A1(n8786), .A2(n4943), .ZN(n5094) );
  NAND2_X1 U6619 ( .A1(n6920), .A2(n5567), .ZN(n5093) );
  NAND2_X1 U6620 ( .A1(n5094), .A2(n5093), .ZN(n5095) );
  XNOR2_X1 U6621 ( .A(n5095), .B(n4297), .ZN(n5096) );
  XOR2_X1 U6622 ( .A(n5097), .B(n5096), .Z(n7060) );
  INV_X1 U6623 ( .A(n5096), .ZN(n5099) );
  INV_X1 U6624 ( .A(n5097), .ZN(n5098) );
  NOR2_X1 U6625 ( .A1(n5133), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5100) );
  NOR2_X1 U6626 ( .A1(n5179), .A2(n5100), .ZN(n8432) );
  NAND2_X1 U6627 ( .A1(n5594), .A2(n8432), .ZN(n5104) );
  NAND2_X1 U6628 ( .A1(n5040), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6629 ( .A1(n8620), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5101) );
  NAND4_X1 U6630 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n8784)
         );
  NAND2_X1 U6631 ( .A1(n8784), .A2(n5456), .ZN(n5126) );
  INV_X1 U6632 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6633 ( .A1(n5108), .A2(SI_7_), .ZN(n5109) );
  INV_X1 U6634 ( .A(SI_8_), .ZN(n5110) );
  NAND2_X1 U6635 ( .A1(n5111), .A2(n5110), .ZN(n5114) );
  INV_X1 U6636 ( .A(n5111), .ZN(n5112) );
  NAND2_X1 U6637 ( .A1(n5112), .A2(SI_8_), .ZN(n5113) );
  NAND2_X1 U6638 ( .A1(n5114), .A2(n5113), .ZN(n5141) );
  NAND2_X1 U6639 ( .A1(n5117), .A2(n5116), .ZN(n5158) );
  INV_X1 U6640 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6641 ( .A1(n5118), .A2(SI_9_), .ZN(n5119) );
  INV_X1 U6642 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6643 ( .A1(n5122), .A2(n5121), .ZN(n5167) );
  NAND2_X1 U6644 ( .A1(n5167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  INV_X1 U6645 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6646 ( .A1(n5138), .A2(n5137), .ZN(n5140) );
  NAND2_X1 U6647 ( .A1(n5140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U6648 ( .A(n5123), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U6649 ( .A1(n5387), .A2(n8813), .ZN(n5124) );
  NAND2_X1 U6650 ( .A1(n8431), .A2(n5567), .ZN(n5125) );
  NAND2_X1 U6651 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  XNOR2_X1 U6652 ( .A(n5127), .B(n5602), .ZN(n8424) );
  AND2_X1 U6653 ( .A1(n8431), .A2(n5456), .ZN(n5128) );
  AOI21_X1 U6654 ( .B1(n8784), .B2(n5551), .A(n5128), .ZN(n5152) );
  INV_X1 U6655 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5130) );
  INV_X1 U6656 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5129) );
  OAI22_X1 U6657 ( .A1(n5645), .A2(n5130), .B1(n5372), .B2(n5129), .ZN(n5136)
         );
  AND2_X1 U6658 ( .A1(n5132), .A2(n7253), .ZN(n5134) );
  OR2_X1 U6659 ( .A1(n5134), .A2(n5133), .ZN(n9549) );
  INV_X1 U6660 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10025) );
  OAI22_X1 U6661 ( .A1(n5642), .A2(n9549), .B1(n5476), .B2(n10025), .ZN(n5135)
         );
  NAND2_X1 U6662 ( .A1(n8785), .A2(n4943), .ZN(n5146) );
  OR2_X1 U6663 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  INV_X1 U6664 ( .A(n6563), .ZN(n9364) );
  XNOR2_X1 U6665 ( .A(n5142), .B(n5141), .ZN(n5857) );
  INV_X1 U6666 ( .A(n5857), .ZN(n6330) );
  OR2_X1 U6667 ( .A1(n5000), .A2(n6330), .ZN(n5144) );
  OR2_X1 U6668 ( .A1(n4999), .A2(n6331), .ZN(n5143) );
  OAI211_X1 U6669 ( .C1(n8615), .C2(n9364), .A(n5144), .B(n5143), .ZN(n7255)
         );
  NAND2_X1 U6670 ( .A1(n7255), .A2(n5567), .ZN(n5145) );
  NAND2_X1 U6671 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  XNOR2_X1 U6672 ( .A(n5147), .B(n4297), .ZN(n8421) );
  NAND2_X1 U6673 ( .A1(n8785), .A2(n5551), .ZN(n5149) );
  NAND2_X1 U6674 ( .A1(n7255), .A2(n5456), .ZN(n5148) );
  NAND2_X1 U6675 ( .A1(n5149), .A2(n5148), .ZN(n7247) );
  NOR2_X1 U6676 ( .A1(n8421), .A2(n7247), .ZN(n5150) );
  NOR2_X1 U6677 ( .A1(n4878), .A2(n5150), .ZN(n5151) );
  INV_X1 U6678 ( .A(n5152), .ZN(n8423) );
  AOI21_X1 U6679 ( .B1(n8421), .B2(n7247), .A(n8423), .ZN(n5154) );
  NAND3_X1 U6680 ( .A1(n8421), .A2(n7247), .A3(n8423), .ZN(n5153) );
  NAND2_X1 U6681 ( .A1(n5157), .A2(n5156), .ZN(n5159) );
  XNOR2_X1 U6682 ( .A(n5160), .B(SI_10_), .ZN(n5186) );
  NAND2_X1 U6683 ( .A1(n5160), .A2(SI_10_), .ZN(n5161) );
  NAND2_X1 U6684 ( .A1(n5164), .A2(n5163), .ZN(n5209) );
  INV_X1 U6685 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6686 ( .A1(n5165), .A2(SI_11_), .ZN(n5166) );
  NAND2_X1 U6687 ( .A1(n5209), .A2(n5166), .ZN(n5206) );
  XNOR2_X1 U6688 ( .A(n5205), .B(n5206), .ZN(n6345) );
  NAND2_X1 U6689 ( .A1(n6345), .A2(n8608), .ZN(n5170) );
  OR2_X1 U6690 ( .A1(n5212), .A2(n4899), .ZN(n5168) );
  XNOR2_X1 U6691 ( .A(n5168), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6565) );
  AOI22_X1 U6692 ( .A1(n5388), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5387), .B2(
        n6565), .ZN(n5169) );
  INV_X1 U6693 ( .A(n9688), .ZN(n8473) );
  OR2_X1 U6694 ( .A1(n5181), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5171) );
  AND2_X1 U6695 ( .A1(n5243), .A2(n5171), .ZN(n8474) );
  NAND2_X1 U6696 ( .A1(n5594), .A2(n8474), .ZN(n5175) );
  NAND2_X1 U6697 ( .A1(n5040), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6698 ( .A1(n8620), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5172) );
  NAND4_X1 U6699 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n8782)
         );
  AOI22_X1 U6700 ( .A1(n8473), .A2(n5567), .B1(n5456), .B2(n8782), .ZN(n5176)
         );
  XNOR2_X1 U6701 ( .A(n5176), .B(n4297), .ZN(n8468) );
  OR2_X1 U6702 ( .A1(n9688), .A2(n5550), .ZN(n5178) );
  NAND2_X1 U6703 ( .A1(n8782), .A2(n5551), .ZN(n5177) );
  NAND2_X1 U6704 ( .A1(n5178), .A2(n5177), .ZN(n8467) );
  INV_X1 U6705 ( .A(n8467), .ZN(n5199) );
  NOR2_X1 U6706 ( .A1(n5179), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6707 ( .A1(n5181), .A2(n5180), .ZN(n7183) );
  INV_X1 U6708 ( .A(n7183), .ZN(n8340) );
  NAND2_X1 U6709 ( .A1(n5594), .A2(n8340), .ZN(n5185) );
  NAND2_X1 U6710 ( .A1(n8620), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6711 ( .A1(n5040), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5182) );
  NAND4_X1 U6712 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n8783)
         );
  NAND2_X1 U6713 ( .A1(n8783), .A2(n5551), .ZN(n5195) );
  INV_X1 U6714 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6715 ( .A1(n6340), .A2(n8608), .ZN(n5193) );
  NAND2_X1 U6716 ( .A1(n5188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6717 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5189), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5191) );
  INV_X1 U6718 ( .A(n5212), .ZN(n5190) );
  NAND2_X1 U6719 ( .A1(n5191), .A2(n5190), .ZN(n6342) );
  AOI22_X1 U6720 ( .A1(n5388), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5387), .B2(
        n9321), .ZN(n5192) );
  NAND2_X1 U6721 ( .A1(n5193), .A2(n5192), .ZN(n7190) );
  NAND2_X1 U6722 ( .A1(n7190), .A2(n5456), .ZN(n5194) );
  NAND2_X1 U6723 ( .A1(n5195), .A2(n5194), .ZN(n5200) );
  INV_X1 U6724 ( .A(n5200), .ZN(n8335) );
  NAND2_X1 U6725 ( .A1(n8783), .A2(n4943), .ZN(n5197) );
  NAND2_X1 U6726 ( .A1(n7190), .A2(n5567), .ZN(n5196) );
  NAND2_X1 U6727 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  XNOR2_X1 U6728 ( .A(n5198), .B(n4297), .ZN(n8466) );
  INV_X1 U6729 ( .A(n8466), .ZN(n8333) );
  OAI22_X1 U6730 ( .A1(n8468), .A2(n5199), .B1(n8335), .B2(n8333), .ZN(n5204)
         );
  OAI21_X1 U6731 ( .B1(n8466), .B2(n5200), .A(n8467), .ZN(n5202) );
  NOR3_X1 U6732 ( .A1(n8466), .A2(n8467), .A3(n5200), .ZN(n5201) );
  AOI21_X1 U6733 ( .B1(n8468), .B2(n5202), .A(n5201), .ZN(n5203) );
  INV_X1 U6734 ( .A(n5206), .ZN(n5207) );
  XNOR2_X1 U6735 ( .A(n5231), .B(SI_12_), .ZN(n5230) );
  XNOR2_X1 U6736 ( .A(n5235), .B(n5230), .ZN(n6351) );
  NAND2_X1 U6737 ( .A1(n6351), .A2(n8608), .ZN(n5218) );
  INV_X1 U6738 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6739 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  NAND2_X1 U6740 ( .A1(n5213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5215) );
  INV_X1 U6741 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6742 ( .A1(n5215), .A2(n5214), .ZN(n5236) );
  OR2_X1 U6743 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  AOI22_X1 U6744 ( .A1(n5388), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5387), .B2(
        n8831), .ZN(n5217) );
  XNOR2_X1 U6745 ( .A(n5243), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U6746 ( .A1(n5594), .A2(n7268), .ZN(n5222) );
  NAND2_X1 U6747 ( .A1(n8620), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6748 ( .A1(n5040), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5219) );
  NAND4_X1 U6749 ( .A1(n5222), .A2(n5221), .A3(n5220), .A4(n5219), .ZN(n8909)
         );
  INV_X1 U6750 ( .A(n8909), .ZN(n7195) );
  OAI22_X1 U6751 ( .A1(n9693), .A2(n5550), .B1(n7195), .B2(n5601), .ZN(n5226)
         );
  NAND2_X1 U6752 ( .A1(n8910), .A2(n5567), .ZN(n5224) );
  NAND2_X1 U6753 ( .A1(n8909), .A2(n4943), .ZN(n5223) );
  NAND2_X1 U6754 ( .A1(n5224), .A2(n5223), .ZN(n5225) );
  XNOR2_X1 U6755 ( .A(n5225), .B(n4297), .ZN(n5227) );
  XOR2_X1 U6756 ( .A(n5226), .B(n5227), .Z(n7266) );
  NAND2_X1 U6757 ( .A1(n7267), .A2(n7266), .ZN(n5229) );
  OR2_X1 U6758 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  INV_X1 U6759 ( .A(n5230), .ZN(n5234) );
  INV_X1 U6760 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U6761 ( .A1(n5232), .A2(SI_12_), .ZN(n5233) );
  XNOR2_X1 U6762 ( .A(n5260), .B(SI_13_), .ZN(n5257) );
  XNOR2_X1 U6763 ( .A(n5259), .B(n5257), .ZN(n6368) );
  NAND2_X1 U6764 ( .A1(n6368), .A2(n8608), .ZN(n5239) );
  NAND2_X1 U6765 ( .A1(n5236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6766 ( .A(n5237), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9457) );
  AOI22_X1 U6767 ( .A1(n5388), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5387), .B2(
        n9457), .ZN(n5238) );
  NAND2_X1 U6768 ( .A1(n5239), .A2(n5238), .ZN(n8875) );
  INV_X1 U6769 ( .A(n8875), .ZN(n9700) );
  INV_X1 U6770 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5241) );
  INV_X1 U6771 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5240) );
  OAI21_X1 U6772 ( .B1(n5243), .B2(n5241), .A(n5240), .ZN(n5244) );
  NAND2_X1 U6773 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5242) );
  NAND2_X1 U6774 ( .A1(n5244), .A2(n5270), .ZN(n9540) );
  INV_X1 U6775 ( .A(n9540), .ZN(n5245) );
  NAND2_X1 U6776 ( .A1(n5594), .A2(n5245), .ZN(n5248) );
  NAND2_X1 U6777 ( .A1(n8620), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6778 ( .A1(n5040), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5246) );
  NAND4_X1 U6779 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n8781)
         );
  OAI22_X1 U6780 ( .A1(n9700), .A2(n5550), .B1(n8913), .B2(n5601), .ZN(n5254)
         );
  NAND2_X1 U6781 ( .A1(n8875), .A2(n5567), .ZN(n5251) );
  NAND2_X1 U6782 ( .A1(n8781), .A2(n4943), .ZN(n5250) );
  NAND2_X1 U6783 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  XNOR2_X1 U6784 ( .A(n5252), .B(n4297), .ZN(n5253) );
  XOR2_X1 U6785 ( .A(n5254), .B(n5253), .Z(n8447) );
  INV_X1 U6786 ( .A(n5253), .ZN(n5256) );
  INV_X1 U6787 ( .A(n5254), .ZN(n5255) );
  AOI21_X2 U6788 ( .B1(n8448), .B2(n8447), .A(n4863), .ZN(n5279) );
  INV_X1 U6789 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6790 ( .A1(n5260), .A2(SI_13_), .ZN(n5261) );
  XNOR2_X1 U6791 ( .A(n5286), .B(SI_14_), .ZN(n5262) );
  XNOR2_X1 U6792 ( .A(n5283), .B(n5262), .ZN(n6452) );
  NAND2_X1 U6793 ( .A1(n6452), .A2(n8608), .ZN(n5268) );
  NOR2_X1 U6794 ( .A1(n5263), .A2(n4899), .ZN(n5264) );
  MUX2_X1 U6795 ( .A(n4899), .B(n5264), .S(P1_IR_REG_14__SCAN_IN), .Z(n5266)
         );
  OR2_X1 U6796 ( .A1(n5266), .A2(n5265), .ZN(n9471) );
  INV_X1 U6797 ( .A(n9471), .ZN(n8833) );
  AOI22_X1 U6798 ( .A1(n5388), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5387), .B2(
        n8833), .ZN(n5267) );
  NAND2_X1 U6799 ( .A1(n9520), .A2(n5567), .ZN(n5277) );
  INV_X1 U6800 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U6801 ( .A1(n5270), .A2(n10002), .ZN(n5271) );
  AND2_X1 U6802 ( .A1(n5318), .A2(n5271), .ZN(n9518) );
  NAND2_X1 U6803 ( .A1(n5594), .A2(n9518), .ZN(n5275) );
  NAND2_X1 U6804 ( .A1(n5040), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6805 ( .A1(n8620), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5272) );
  NAND4_X1 U6806 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n8915)
         );
  NAND2_X1 U6807 ( .A1(n8915), .A2(n4943), .ZN(n5276) );
  NAND2_X1 U6808 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  XNOR2_X1 U6809 ( .A(n5278), .B(n5602), .ZN(n5280) );
  XNOR2_X1 U6810 ( .A(n5279), .B(n5280), .ZN(n8314) );
  AOI22_X1 U6811 ( .A1(n9520), .A2(n5456), .B1(n5551), .B2(n8915), .ZN(n8315)
         );
  NAND2_X1 U6812 ( .A1(n8314), .A2(n8315), .ZN(n8313) );
  INV_X1 U6813 ( .A(n5279), .ZN(n5281) );
  NAND2_X1 U6814 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6815 ( .A1(n8313), .A2(n5282), .ZN(n8373) );
  NAND2_X1 U6816 ( .A1(n5286), .A2(SI_14_), .ZN(n5284) );
  INV_X1 U6817 ( .A(n5286), .ZN(n5288) );
  NAND2_X1 U6818 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  NOR2_X1 U6819 ( .A1(n5293), .A2(SI_15_), .ZN(n5292) );
  NAND2_X1 U6820 ( .A1(n5293), .A2(SI_15_), .ZN(n5294) );
  XNOR2_X1 U6821 ( .A(n5335), .B(SI_16_), .ZN(n5295) );
  XNOR2_X1 U6822 ( .A(n5339), .B(n5295), .ZN(n6653) );
  NAND2_X1 U6823 ( .A1(n6653), .A2(n8608), .ZN(n5299) );
  NAND2_X1 U6824 ( .A1(n5296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6825 ( .A(n5297), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8846) );
  AOI22_X1 U6826 ( .A1(n5388), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5387), .B2(
        n8846), .ZN(n5298) );
  NAND2_X1 U6827 ( .A1(n9244), .A2(n5567), .ZN(n5307) );
  INV_X1 U6828 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6829 ( .A1(n5320), .A2(n5300), .ZN(n5301) );
  AND2_X1 U6830 ( .A1(n5348), .A2(n5301), .ZN(n9147) );
  NAND2_X1 U6831 ( .A1(n5594), .A2(n9147), .ZN(n5305) );
  NAND2_X1 U6832 ( .A1(n5040), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6833 ( .A1(n8620), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5302) );
  NAND4_X1 U6834 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n8780)
         );
  NAND2_X1 U6835 ( .A1(n8780), .A2(n4943), .ZN(n5306) );
  NAND2_X1 U6836 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  XNOR2_X1 U6837 ( .A(n5308), .B(n4297), .ZN(n5330) );
  OAI22_X1 U6838 ( .A1(n9150), .A2(n5550), .B1(n8920), .B2(n5601), .ZN(n8376)
         );
  XNOR2_X1 U6839 ( .A(n5309), .B(SI_15_), .ZN(n5310) );
  XNOR2_X1 U6840 ( .A(n5311), .B(n5310), .ZN(n6477) );
  NAND2_X1 U6841 ( .A1(n6477), .A2(n8608), .ZN(n5316) );
  NOR2_X1 U6842 ( .A1(n5265), .A2(n4899), .ZN(n5312) );
  MUX2_X1 U6843 ( .A(n4899), .B(n5312), .S(P1_IR_REG_15__SCAN_IN), .Z(n5313)
         );
  INV_X1 U6844 ( .A(n5313), .ZN(n5314) );
  NAND2_X1 U6845 ( .A1(n5314), .A2(n5296), .ZN(n8835) );
  INV_X1 U6846 ( .A(n8835), .ZN(n9484) );
  AOI22_X1 U6847 ( .A1(n5388), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5387), .B2(
        n9484), .ZN(n5315) );
  NAND2_X1 U6848 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  NAND2_X1 U6849 ( .A1(n5320), .A2(n5319), .ZN(n9163) );
  INV_X1 U6850 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5321) );
  OAI22_X1 U6851 ( .A1(n5642), .A2(n9163), .B1(n5372), .B2(n5321), .ZN(n5325)
         );
  INV_X1 U6852 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5323) );
  INV_X1 U6853 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5322) );
  OAI22_X1 U6854 ( .A1(n5645), .A2(n5323), .B1(n5476), .B2(n5322), .ZN(n5324)
         );
  INV_X1 U6855 ( .A(n8919), .ZN(n8917) );
  OAI22_X1 U6856 ( .A1(n9377), .A2(n4982), .B1(n8917), .B2(n5550), .ZN(n5326)
         );
  XNOR2_X1 U6857 ( .A(n5326), .B(n4297), .ZN(n8374) );
  OR2_X1 U6858 ( .A1(n9377), .A2(n5550), .ZN(n5328) );
  NAND2_X1 U6859 ( .A1(n8919), .A2(n5551), .ZN(n5327) );
  NAND2_X1 U6860 ( .A1(n5328), .A2(n5327), .ZN(n8503) );
  AOI22_X1 U6861 ( .A1(n5330), .A2(n8376), .B1(n8374), .B2(n8503), .ZN(n5329)
         );
  NAND2_X1 U6862 ( .A1(n8373), .A2(n5329), .ZN(n5334) );
  INV_X1 U6863 ( .A(n5330), .ZN(n8377) );
  OAI21_X1 U6864 ( .B1(n8374), .B2(n8503), .A(n8376), .ZN(n5332) );
  NOR3_X1 U6865 ( .A1(n8376), .A2(n8374), .A3(n8503), .ZN(n5331) );
  AOI21_X1 U6866 ( .B1(n8377), .B2(n5332), .A(n5331), .ZN(n5333) );
  AND2_X1 U6867 ( .A1(n5335), .A2(SI_16_), .ZN(n5338) );
  INV_X1 U6868 ( .A(n5335), .ZN(n5337) );
  INV_X1 U6869 ( .A(SI_16_), .ZN(n5336) );
  XNOR2_X1 U6870 ( .A(n5359), .B(SI_17_), .ZN(n5356) );
  XNOR2_X1 U6871 ( .A(n5357), .B(n5356), .ZN(n6702) );
  NAND2_X1 U6872 ( .A1(n6702), .A2(n8608), .ZN(n5344) );
  XNOR2_X1 U6873 ( .A(n5342), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8858) );
  AOI22_X1 U6874 ( .A1(n5388), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5387), .B2(
        n8858), .ZN(n5343) );
  INV_X1 U6875 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9130) );
  INV_X1 U6876 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5345) );
  OAI22_X1 U6877 ( .A1(n5645), .A2(n9130), .B1(n5372), .B2(n5345), .ZN(n5352)
         );
  INV_X1 U6878 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6879 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6880 ( .A1(n5375), .A2(n5349), .ZN(n9129) );
  INV_X1 U6881 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5350) );
  OAI22_X1 U6882 ( .A1(n5642), .A2(n9129), .B1(n5476), .B2(n5350), .ZN(n5351)
         );
  AOI22_X1 U6883 ( .A1(n9239), .A2(n5567), .B1(n5456), .B2(n8921), .ZN(n5353)
         );
  XOR2_X1 U6884 ( .A(n4297), .B(n5353), .Z(n5355) );
  INV_X1 U6885 ( .A(n9239), .ZN(n9128) );
  INV_X1 U6886 ( .A(n8921), .ZN(n8560) );
  OAI22_X1 U6887 ( .A1(n9128), .A2(n5550), .B1(n8560), .B2(n5601), .ZN(n5354)
         );
  NAND2_X1 U6888 ( .A1(n5355), .A2(n5354), .ZN(n8399) );
  NOR2_X1 U6889 ( .A1(n5355), .A2(n5354), .ZN(n8398) );
  NAND2_X1 U6890 ( .A1(n5357), .A2(n5356), .ZN(n5361) );
  INV_X1 U6891 ( .A(SI_17_), .ZN(n5358) );
  NAND2_X1 U6892 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X1 U6893 ( .A1(n5362), .A2(SI_18_), .ZN(n5386) );
  INV_X1 U6894 ( .A(n5362), .ZN(n5364) );
  INV_X1 U6895 ( .A(SI_18_), .ZN(n5363) );
  NAND2_X1 U6896 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  XNOR2_X1 U6897 ( .A(n5384), .B(n5385), .ZN(n6761) );
  NAND2_X1 U6898 ( .A1(n6761), .A2(n8608), .ZN(n5371) );
  OR2_X1 U6899 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  AND2_X1 U6900 ( .A1(n5369), .A2(n5368), .ZN(n8865) );
  AOI22_X1 U6901 ( .A1(n5388), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5387), .B2(
        n8865), .ZN(n5370) );
  NAND2_X1 U6902 ( .A1(n9121), .A2(n5567), .ZN(n5380) );
  INV_X1 U6903 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9117) );
  INV_X1 U6904 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9235) );
  OAI22_X1 U6905 ( .A1(n5645), .A2(n9117), .B1(n5372), .B2(n9235), .ZN(n5378)
         );
  INV_X1 U6906 ( .A(n5375), .ZN(n5373) );
  NAND2_X1 U6907 ( .A1(n5373), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5391) );
  INV_X1 U6908 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6909 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  NAND2_X1 U6910 ( .A1(n5391), .A2(n5376), .ZN(n9116) );
  INV_X1 U6911 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10005) );
  OAI22_X1 U6912 ( .A1(n5642), .A2(n9116), .B1(n5476), .B2(n10005), .ZN(n5377)
         );
  NAND2_X1 U6913 ( .A1(n8922), .A2(n5456), .ZN(n5379) );
  NAND2_X1 U6914 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  XNOR2_X1 U6915 ( .A(n5381), .B(n5602), .ZN(n5383) );
  AOI22_X1 U6916 ( .A1(n9121), .A2(n5456), .B1(n5551), .B2(n8922), .ZN(n5382)
         );
  NAND2_X1 U6917 ( .A1(n5383), .A2(n5382), .ZN(n8480) );
  OR2_X1 U6918 ( .A1(n5383), .A2(n5382), .ZN(n8481) );
  XNOR2_X1 U6919 ( .A(n5400), .B(SI_19_), .ZN(n5404) );
  XNOR2_X1 U6920 ( .A(n5405), .B(n5404), .ZN(n6882) );
  NAND2_X1 U6921 ( .A1(n6882), .A2(n8608), .ZN(n5390) );
  AOI22_X1 U6922 ( .A1(n5388), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5387), .B2(
        n9535), .ZN(n5389) );
  INV_X1 U6923 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9098) );
  INV_X1 U6924 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9229) );
  OAI22_X1 U6925 ( .A1(n5645), .A2(n9098), .B1(n5372), .B2(n9229), .ZN(n5394)
         );
  INV_X1 U6926 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U6927 ( .A1(n5391), .A2(n8350), .ZN(n5392) );
  NAND2_X1 U6928 ( .A1(n5410), .A2(n5392), .ZN(n9097) );
  INV_X1 U6929 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10012) );
  OAI22_X1 U6930 ( .A1(n5642), .A2(n9097), .B1(n5476), .B2(n10012), .ZN(n5393)
         );
  OAI22_X1 U6931 ( .A1(n9096), .A2(n4982), .B1(n8925), .B2(n5550), .ZN(n5395)
         );
  XNOR2_X1 U6932 ( .A(n5395), .B(n5602), .ZN(n5399) );
  OR2_X1 U6933 ( .A1(n9096), .A2(n5550), .ZN(n5397) );
  NAND2_X1 U6934 ( .A1(n8926), .A2(n5551), .ZN(n5396) );
  AND2_X1 U6935 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NOR2_X1 U6936 ( .A1(n5399), .A2(n5398), .ZN(n8345) );
  NAND2_X1 U6937 ( .A1(n5399), .A2(n5398), .ZN(n8343) );
  OAI21_X2 U6938 ( .B1(n8347), .B2(n8345), .A(n8343), .ZN(n8438) );
  INV_X1 U6939 ( .A(n5400), .ZN(n5402) );
  INV_X1 U6940 ( .A(SI_19_), .ZN(n5401) );
  NAND2_X1 U6941 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  XNOR2_X1 U6942 ( .A(n5422), .B(SI_20_), .ZN(n5419) );
  XNOR2_X1 U6943 ( .A(n5420), .B(n5419), .ZN(n6944) );
  NAND2_X1 U6944 ( .A1(n6944), .A2(n8608), .ZN(n5407) );
  OR2_X1 U6945 ( .A1(n4999), .A2(n6953), .ZN(n5406) );
  INV_X1 U6946 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9082) );
  INV_X1 U6947 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9224) );
  OAI22_X1 U6948 ( .A1(n5645), .A2(n9082), .B1(n5372), .B2(n9224), .ZN(n5413)
         );
  INV_X1 U6949 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6950 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  NAND2_X1 U6951 ( .A1(n5428), .A2(n5411), .ZN(n9090) );
  INV_X1 U6952 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9283) );
  OAI22_X1 U6953 ( .A1(n5642), .A2(n9090), .B1(n5476), .B2(n9283), .ZN(n5412)
         );
  AOI22_X1 U6954 ( .A1(n9223), .A2(n5567), .B1(n5456), .B2(n8928), .ZN(n5414)
         );
  XOR2_X1 U6955 ( .A(n4297), .B(n5414), .Z(n5416) );
  OAI22_X1 U6956 ( .A1(n9083), .A2(n5550), .B1(n8929), .B2(n5601), .ZN(n5415)
         );
  NOR2_X1 U6957 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  AOI21_X1 U6958 ( .B1(n5416), .B2(n5415), .A(n5417), .ZN(n8439) );
  NAND2_X1 U6959 ( .A1(n8438), .A2(n8439), .ZN(n8437) );
  INV_X1 U6960 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6961 ( .A1(n5420), .A2(n5419), .ZN(n5424) );
  INV_X1 U6962 ( .A(SI_20_), .ZN(n5421) );
  NAND2_X1 U6963 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  XNOR2_X1 U6964 ( .A(n5442), .B(SI_21_), .ZN(n5425) );
  XNOR2_X1 U6965 ( .A(n5440), .B(n5425), .ZN(n6995) );
  NAND2_X1 U6966 ( .A1(n6995), .A2(n8608), .ZN(n5427) );
  OR2_X1 U6967 ( .A1(n8603), .A2(n7040), .ZN(n5426) );
  INV_X1 U6968 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U6969 ( .A1(n5428), .A2(n8361), .ZN(n5429) );
  AND2_X1 U6970 ( .A1(n5452), .A2(n5429), .ZN(n9072) );
  NAND2_X1 U6971 ( .A1(n5594), .A2(n9072), .ZN(n5433) );
  NAND2_X1 U6972 ( .A1(n5040), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6973 ( .A1(n8620), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5430) );
  NAND4_X1 U6974 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n8931)
         );
  OAI22_X1 U6975 ( .A1(n9075), .A2(n5550), .B1(n8930), .B2(n5601), .ZN(n5436)
         );
  OAI22_X1 U6976 ( .A1(n9075), .A2(n4982), .B1(n8930), .B2(n5550), .ZN(n5434)
         );
  XNOR2_X1 U6977 ( .A(n5434), .B(n4297), .ZN(n5435) );
  XOR2_X1 U6978 ( .A(n5436), .B(n5435), .Z(n8357) );
  INV_X1 U6979 ( .A(n5435), .ZN(n5438) );
  INV_X1 U6980 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6981 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  INV_X1 U6982 ( .A(SI_21_), .ZN(n5441) );
  INV_X1 U6983 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6984 ( .A1(n5443), .A2(SI_21_), .ZN(n5444) );
  INV_X1 U6985 ( .A(SI_22_), .ZN(n5445) );
  NAND2_X1 U6986 ( .A1(n5446), .A2(n5445), .ZN(n5462) );
  INV_X1 U6987 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6988 ( .A1(n5447), .A2(SI_22_), .ZN(n5448) );
  NAND2_X1 U6989 ( .A1(n5462), .A2(n5448), .ZN(n5463) );
  XNOR2_X1 U6990 ( .A(n5464), .B(n5463), .ZN(n7101) );
  NAND2_X1 U6991 ( .A1(n7101), .A2(n8608), .ZN(n5450) );
  OR2_X1 U6992 ( .A1(n4999), .A2(n7106), .ZN(n5449) );
  INV_X1 U6993 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9054) );
  INV_X1 U6994 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9214) );
  OAI22_X1 U6995 ( .A1(n5645), .A2(n9054), .B1(n5372), .B2(n9214), .ZN(n5455)
         );
  INV_X1 U6996 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U6997 ( .A1(n5452), .A2(n8458), .ZN(n5453) );
  NAND2_X1 U6998 ( .A1(n5474), .A2(n5453), .ZN(n9053) );
  INV_X1 U6999 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9275) );
  OAI22_X1 U7000 ( .A1(n5642), .A2(n9053), .B1(n5476), .B2(n9275), .ZN(n5454)
         );
  AOI22_X1 U7001 ( .A1(n9213), .A2(n5567), .B1(n5456), .B2(n8935), .ZN(n5457)
         );
  XNOR2_X1 U7002 ( .A(n5457), .B(n4297), .ZN(n5458) );
  INV_X1 U7003 ( .A(n5458), .ZN(n5459) );
  INV_X1 U7004 ( .A(n8456), .ZN(n5461) );
  OAI22_X1 U7005 ( .A1(n9052), .A2(n5550), .B1(n8934), .B2(n5601), .ZN(n8457)
         );
  NAND2_X1 U7006 ( .A1(n5461), .A2(n5460), .ZN(n8322) );
  NAND2_X1 U7007 ( .A1(n8322), .A2(n8323), .ZN(n5489) );
  INV_X1 U7008 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7217) );
  INV_X1 U7009 ( .A(SI_23_), .ZN(n5465) );
  NAND2_X1 U7010 ( .A1(n5466), .A2(n5465), .ZN(n5490) );
  INV_X1 U7011 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U7012 ( .A1(n5467), .A2(SI_23_), .ZN(n5468) );
  NAND2_X1 U7013 ( .A1(n5470), .A2(n5469), .ZN(n5491) );
  OR2_X1 U7014 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7015 ( .A1(n5491), .A2(n5471), .ZN(n7219) );
  NAND2_X1 U7016 ( .A1(n7219), .A2(n8608), .ZN(n5473) );
  OR2_X1 U7017 ( .A1(n4999), .A2(n7217), .ZN(n5472) );
  NAND2_X1 U7018 ( .A1(n9209), .A2(n5567), .ZN(n5481) );
  INV_X1 U7019 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U7020 ( .A1(n5474), .A2(n8329), .ZN(n5475) );
  NAND2_X1 U7021 ( .A1(n5498), .A2(n5475), .ZN(n8328) );
  INV_X1 U7022 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9271) );
  OAI22_X1 U7023 ( .A1(n8328), .A2(n5642), .B1(n5476), .B2(n9271), .ZN(n5479)
         );
  INV_X1 U7024 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5477) );
  INV_X1 U7025 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10024) );
  OAI22_X1 U7026 ( .A1(n5645), .A2(n5477), .B1(n5372), .B2(n10024), .ZN(n5478)
         );
  NAND2_X1 U7027 ( .A1(n8938), .A2(n4943), .ZN(n5480) );
  NAND2_X1 U7028 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  XNOR2_X1 U7029 ( .A(n5482), .B(n5602), .ZN(n5484) );
  AND2_X1 U7030 ( .A1(n8938), .A2(n5551), .ZN(n5483) );
  AOI21_X1 U7031 ( .B1(n9209), .B2(n5456), .A(n5483), .ZN(n5485) );
  NAND2_X1 U7032 ( .A1(n5484), .A2(n5485), .ZN(n8406) );
  INV_X1 U7033 ( .A(n5484), .ZN(n5487) );
  INV_X1 U7034 ( .A(n5485), .ZN(n5486) );
  NAND2_X1 U7035 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U7036 ( .A1(n5489), .A2(n8324), .ZN(n8326) );
  NAND2_X1 U7037 ( .A1(n8326), .A2(n8406), .ZN(n5510) );
  INV_X1 U7038 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7278) );
  INV_X1 U7039 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7230) );
  INV_X1 U7040 ( .A(SI_24_), .ZN(n5492) );
  NAND2_X1 U7041 ( .A1(n5493), .A2(n5492), .ZN(n5514) );
  INV_X1 U7042 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7043 ( .A1(n5494), .A2(SI_24_), .ZN(n5495) );
  XNOR2_X1 U7044 ( .A(n5513), .B(n5512), .ZN(n7229) );
  NAND2_X1 U7045 ( .A1(n7229), .A2(n8608), .ZN(n5497) );
  OR2_X1 U7046 ( .A1(n8603), .A2(n7230), .ZN(n5496) );
  INV_X1 U7047 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U7048 ( .A1(n5498), .A2(n8415), .ZN(n5499) );
  NAND2_X1 U7049 ( .A1(n5523), .A2(n5499), .ZN(n8413) );
  AOI22_X1 U7050 ( .A1(n8620), .A2(P1_REG1_REG_24__SCAN_IN), .B1(n5040), .B2(
        P1_REG0_REG_24__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U7051 ( .C1(n8413), .C2(n5642), .A(n5501), .B(n5500), .ZN(n8941)
         );
  INV_X1 U7052 ( .A(n8941), .ZN(n8940) );
  OAI22_X1 U7053 ( .A1(n9032), .A2(n4982), .B1(n8940), .B2(n5550), .ZN(n5502)
         );
  XNOR2_X1 U7054 ( .A(n5502), .B(n5602), .ZN(n5505) );
  OR2_X1 U7055 ( .A1(n9032), .A2(n5550), .ZN(n5504) );
  NAND2_X1 U7056 ( .A1(n8941), .A2(n5551), .ZN(n5503) );
  NAND2_X1 U7057 ( .A1(n5505), .A2(n5506), .ZN(n5511) );
  INV_X1 U7058 ( .A(n5505), .ZN(n5508) );
  INV_X1 U7059 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U7060 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  NAND2_X1 U7061 ( .A1(n5510), .A2(n8407), .ZN(n8410) );
  NAND2_X1 U7062 ( .A1(n5513), .A2(n5512), .ZN(n5515) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U7064 ( .A1(n5516), .A2(n9906), .ZN(n5532) );
  INV_X1 U7065 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U7066 ( .A1(n5517), .A2(SI_25_), .ZN(n5518) );
  XNOR2_X1 U7067 ( .A(n5531), .B(n5530), .ZN(n7275) );
  NAND2_X1 U7068 ( .A1(n7275), .A2(n8608), .ZN(n5520) );
  OR2_X1 U7069 ( .A1(n4999), .A2(n7288), .ZN(n5519) );
  INV_X1 U7070 ( .A(n9199), .ZN(n9018) );
  INV_X1 U7071 ( .A(n5523), .ZN(n5521) );
  NAND2_X1 U7072 ( .A1(n5521), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5541) );
  INV_X1 U7073 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7074 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  NAND2_X1 U7075 ( .A1(n5541), .A2(n5524), .ZN(n9014) );
  AOI22_X1 U7076 ( .A1(n8620), .A2(P1_REG1_REG_25__SCAN_IN), .B1(n5040), .B2(
        P1_REG0_REG_25__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7077 ( .C1(n9014), .C2(n5642), .A(n5526), .B(n5525), .ZN(n8943)
         );
  INV_X1 U7078 ( .A(n8943), .ZN(n8944) );
  OAI22_X1 U7079 ( .A1(n9018), .A2(n5550), .B1(n8944), .B2(n5601), .ZN(n5554)
         );
  NAND2_X1 U7080 ( .A1(n9199), .A2(n5567), .ZN(n5528) );
  NAND2_X1 U7081 ( .A1(n8943), .A2(n5456), .ZN(n5527) );
  NAND2_X1 U7082 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U7083 ( .A(n5529), .B(n4297), .ZN(n5555) );
  XOR2_X1 U7084 ( .A(n5554), .B(n5555), .Z(n8367) );
  INV_X1 U7085 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8301) );
  INV_X1 U7086 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9309) );
  INV_X1 U7087 ( .A(SI_26_), .ZN(n5533) );
  NAND2_X1 U7088 ( .A1(n5534), .A2(n5533), .ZN(n5559) );
  INV_X1 U7089 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7090 ( .A1(n5535), .A2(SI_26_), .ZN(n5536) );
  NAND2_X1 U7091 ( .A1(n8299), .A2(n8608), .ZN(n5538) );
  OR2_X1 U7092 ( .A1(n8603), .A2(n9309), .ZN(n5537) );
  INV_X1 U7093 ( .A(n5541), .ZN(n5539) );
  NAND2_X1 U7094 ( .A1(n5539), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5569) );
  INV_X1 U7095 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7096 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  NAND2_X1 U7097 ( .A1(n5569), .A2(n5542), .ZN(n9000) );
  OR2_X1 U7098 ( .A1(n9000), .A2(n5642), .ZN(n5547) );
  INV_X1 U7099 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U7100 ( .A1(n8620), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7101 ( .A1(n5040), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7102 ( .C1(n5645), .C2(n8999), .A(n5544), .B(n5543), .ZN(n5545)
         );
  INV_X1 U7103 ( .A(n5545), .ZN(n5546) );
  OAI22_X1 U7104 ( .A1(n9194), .A2(n4982), .B1(n8945), .B2(n5550), .ZN(n5549)
         );
  XNOR2_X1 U7105 ( .A(n5549), .B(n4297), .ZN(n5585) );
  OR2_X1 U7106 ( .A1(n9194), .A2(n5550), .ZN(n5553) );
  NAND2_X1 U7107 ( .A1(n8946), .A2(n5551), .ZN(n5552) );
  NAND2_X1 U7108 ( .A1(n5553), .A2(n5552), .ZN(n5584) );
  XNOR2_X1 U7109 ( .A(n5585), .B(n5584), .ZN(n8491) );
  NOR2_X1 U7110 ( .A1(n5555), .A2(n5554), .ZN(n8492) );
  NOR2_X1 U7111 ( .A1(n8491), .A2(n8492), .ZN(n5556) );
  NAND2_X1 U7112 ( .A1(n5560), .A2(n5559), .ZN(n5590) );
  INV_X1 U7113 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8297) );
  INV_X1 U7114 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7381) );
  INV_X1 U7115 ( .A(SI_27_), .ZN(n5561) );
  NAND2_X1 U7116 ( .A1(n5562), .A2(n5561), .ZN(n5591) );
  INV_X1 U7117 ( .A(n5562), .ZN(n5563) );
  NAND2_X1 U7118 ( .A1(n5563), .A2(SI_27_), .ZN(n5564) );
  NAND2_X1 U7119 ( .A1(n7380), .A2(n8608), .ZN(n5566) );
  NAND2_X1 U7120 ( .A1(n9190), .A2(n5567), .ZN(n5577) );
  INV_X1 U7121 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7122 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  NAND2_X1 U7123 ( .A1(n8986), .A2(n5594), .ZN(n5575) );
  INV_X1 U7124 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U7125 ( .A1(n5040), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7126 ( .A1(n8620), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5571) );
  OAI211_X1 U7127 ( .C1(n5645), .C2(n8979), .A(n5572), .B(n5571), .ZN(n5573)
         );
  INV_X1 U7128 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7129 ( .A1(n8947), .A2(n5456), .ZN(n5576) );
  NAND2_X1 U7130 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  XNOR2_X1 U7131 ( .A(n5578), .B(n5602), .ZN(n5581) );
  INV_X1 U7132 ( .A(n5581), .ZN(n5583) );
  NOR2_X1 U7133 ( .A1(n8596), .A2(n5601), .ZN(n5579) );
  AOI21_X1 U7134 ( .B1(n9190), .B2(n4943), .A(n5579), .ZN(n5580) );
  INV_X1 U7135 ( .A(n5580), .ZN(n5582) );
  AOI21_X1 U7136 ( .B1(n5583), .B2(n5582), .A(n5631), .ZN(n8305) );
  INV_X1 U7137 ( .A(n8305), .ZN(n5587) );
  NAND2_X1 U7138 ( .A1(n5585), .A2(n5584), .ZN(n8306) );
  INV_X1 U7139 ( .A(n8306), .ZN(n5586) );
  NOR2_X1 U7140 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  INV_X1 U7141 ( .A(n8307), .ZN(n5630) );
  INV_X1 U7142 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8295) );
  INV_X1 U7143 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7601) );
  MUX2_X1 U7144 ( .A(n8295), .B(n7601), .S(n8613), .Z(n6224) );
  XNOR2_X1 U7145 ( .A(n6224), .B(SI_28_), .ZN(n6221) );
  NAND2_X1 U7146 ( .A1(n7600), .A2(n8608), .ZN(n5593) );
  OR2_X1 U7147 ( .A1(n8603), .A2(n7601), .ZN(n5592) );
  XNOR2_X1 U7148 ( .A(n5641), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U7149 ( .A1(n8971), .A2(n5594), .ZN(n5600) );
  INV_X1 U7150 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7151 ( .A1(n8620), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7152 ( .A1(n5040), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7153 ( .C1(n5645), .C2(n5597), .A(n5596), .B(n5595), .ZN(n5598)
         );
  INV_X1 U7154 ( .A(n5598), .ZN(n5599) );
  OAI22_X1 U7155 ( .A1(n8974), .A2(n5550), .B1(n8949), .B2(n5601), .ZN(n5603)
         );
  XNOR2_X1 U7156 ( .A(n5603), .B(n5602), .ZN(n5605) );
  OAI22_X1 U7157 ( .A1(n8974), .A2(n4982), .B1(n8949), .B2(n5550), .ZN(n5604)
         );
  XNOR2_X1 U7158 ( .A(n5605), .B(n5604), .ZN(n5632) );
  INV_X1 U7159 ( .A(n5632), .ZN(n5629) );
  NOR2_X1 U7160 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n10030) );
  NOR4_X1 U7161 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5608) );
  NOR4_X1 U7162 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5607) );
  NOR4_X1 U7163 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5606) );
  NAND4_X1 U7164 ( .A1(n10030), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n5614)
         );
  NOR4_X1 U7165 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5612) );
  NOR4_X1 U7166 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5611) );
  NOR4_X1 U7167 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5610) );
  NOR4_X1 U7168 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5609) );
  NAND4_X1 U7169 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), .ZN(n5613)
         );
  NOR2_X1 U7170 ( .A1(n5614), .A2(n5613), .ZN(n6513) );
  NAND2_X1 U7171 ( .A1(n5615), .A2(P1_B_REG_SCAN_IN), .ZN(n5616) );
  MUX2_X1 U7172 ( .A(P1_B_REG_SCAN_IN), .B(n5616), .S(n7232), .Z(n5617) );
  INV_X1 U7173 ( .A(n6337), .ZN(n5618) );
  INV_X1 U7174 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10007) );
  INV_X1 U7175 ( .A(n5620), .ZN(n9311) );
  INV_X1 U7176 ( .A(n5615), .ZN(n5619) );
  OR2_X1 U7177 ( .A1(n5620), .A2(n5619), .ZN(n9297) );
  OAI21_X1 U7178 ( .B1(n6337), .B2(P1_D_REG_1__SCAN_IN), .A(n9297), .ZN(n6518)
         );
  INV_X1 U7179 ( .A(n6518), .ZN(n6738) );
  OAI211_X1 U7180 ( .C1(n6513), .C2(n6337), .A(n6574), .B(n6738), .ZN(n5634)
         );
  NAND2_X1 U7181 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  NAND2_X1 U7182 ( .A1(n5623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  INV_X1 U7183 ( .A(n6514), .ZN(n8514) );
  OR2_X1 U7184 ( .A1(n5634), .A2(n8514), .ZN(n5648) );
  INV_X1 U7185 ( .A(n6508), .ZN(n6512) );
  INV_X1 U7186 ( .A(n5631), .ZN(n5628) );
  NAND3_X1 U7187 ( .A1(n8307), .A2(n8495), .A3(n5632), .ZN(n5654) );
  NAND3_X1 U7188 ( .A1(n5632), .A2(n5631), .A3(n8495), .ZN(n5653) );
  OR2_X1 U7189 ( .A1(n6508), .A2(n6955), .ZN(n9534) );
  INV_X1 U7190 ( .A(n6517), .ZN(n5633) );
  INV_X1 U7191 ( .A(n9534), .ZN(n5635) );
  OAI21_X1 U7192 ( .B1(n5635), .B2(n9180), .A(n5634), .ZN(n5637) );
  INV_X1 U7193 ( .A(n6515), .ZN(n5636) );
  NAND3_X1 U7194 ( .A1(n5637), .A2(n5636), .A3(n6299), .ZN(n5638) );
  NAND2_X1 U7195 ( .A1(n5638), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5639) );
  OR2_X1 U7196 ( .A1(n6363), .A2(P1_U3086), .ZN(n8770) );
  INV_X1 U7197 ( .A(n8971), .ZN(n5650) );
  INV_X1 U7198 ( .A(n5641), .ZN(n8956) );
  INV_X1 U7199 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U7200 ( .A1(n5642), .A2(n9918), .ZN(n5647) );
  INV_X1 U7201 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U7202 ( .A1(n8620), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7203 ( .A1(n5040), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U7204 ( .C1(n5645), .C2(n8959), .A(n5644), .B(n5643), .ZN(n5646)
         );
  AOI21_X1 U7205 ( .B1(n8956), .B2(n5647), .A(n5646), .ZN(n8606) );
  OAI22_X1 U7206 ( .A1(n8596), .A2(n8908), .B1(n8606), .B2(n8505), .ZN(n8965)
         );
  NOR2_X2 U7207 ( .A1(n5648), .A2(n5626), .ZN(n8506) );
  AOI22_X1 U7208 ( .A1(n8965), .A2(n8506), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5649) );
  OAI21_X1 U7209 ( .B1(n8508), .B2(n5650), .A(n5649), .ZN(n5651) );
  AOI21_X1 U7210 ( .B1(n9186), .B2(n4295), .A(n5651), .ZN(n5652) );
  NAND3_X1 U7211 ( .A1(n5655), .A2(n5654), .A3(n4877), .ZN(P1_U3220) );
  NOR2_X1 U7212 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5798) );
  NAND2_X1 U7213 ( .A1(n5798), .A2(n5656), .ZN(n5831) );
  NAND2_X1 U7214 ( .A1(n5864), .A2(n5657), .ZN(n5889) );
  INV_X1 U7215 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7216 ( .A1(n5919), .A2(n5658), .ZN(n5956) );
  INV_X1 U7217 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5659) );
  INV_X1 U7218 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7693) );
  INV_X1 U7219 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5660) );
  INV_X1 U7220 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9949) );
  INV_X1 U7221 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5661) );
  INV_X1 U7222 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7223 ( .A1(n5663), .A2(n5662), .ZN(n6146) );
  INV_X1 U7224 ( .A(n5663), .ZN(n6102) );
  NAND2_X1 U7225 ( .A1(n6102), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7226 ( .A1(n6146), .A2(n5664), .ZN(n7949) );
  NOR2_X2 U7227 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5668) );
  INV_X2 U7228 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7229 ( .A1(n5980), .A2(n5982), .ZN(n5695) );
  NOR2_X1 U7230 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5672) );
  NAND4_X1 U7231 ( .A1(n5672), .A2(n5671), .A3(n5723), .A4(n5696), .ZN(n5675)
         );
  NAND4_X1 U7232 ( .A1(n5673), .A2(n6133), .A3(n5699), .A4(n6129), .ZN(n5674)
         );
  NAND2_X1 U7233 ( .A1(n5707), .A2(n5688), .ZN(n5690) );
  NOR2_X2 U7234 ( .A1(n5690), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7235 ( .A1(n5679), .A2(n5678), .ZN(n8287) );
  XNOR2_X2 U7236 ( .A(n5680), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7237 ( .A1(n7949), .A2(n6229), .ZN(n5687) );
  INV_X1 U7238 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7948) );
  INV_X1 U7239 ( .A(n5682), .ZN(n5756) );
  INV_X2 U7240 ( .A(n5789), .ZN(n5775) );
  NAND2_X1 U7241 ( .A1(n5775), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7242 ( .A1(n6103), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7243 ( .C1(n7948), .C2(n6594), .A(n5684), .B(n5683), .ZN(n5685)
         );
  INV_X1 U7244 ( .A(n5685), .ZN(n5686) );
  XNOR2_X2 U7245 ( .A(n5692), .B(n5691), .ZN(n6154) );
  NAND2_X4 U7246 ( .A1(n6155), .A2(n6154), .ZN(n6378) );
  NAND2_X2 U7247 ( .A1(n6378), .A2(n4298), .ZN(n5772) );
  NAND2_X1 U7248 ( .A1(n7380), .A2(n7542), .ZN(n5694) );
  NAND2_X4 U7249 ( .A1(n6378), .A2(n8613), .ZN(n7543) );
  OR2_X1 U7250 ( .A1(n7543), .A2(n8297), .ZN(n5693) );
  AND2_X2 U7251 ( .A1(n5721), .A2(n5697), .ZN(n5717) );
  NAND2_X1 U7252 ( .A1(n6130), .A2(n6129), .ZN(n5698) );
  XNOR2_X1 U7253 ( .A(n5712), .B(P2_B_REG_SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7254 ( .A1(n5705), .A2(n7277), .ZN(n5711) );
  NAND2_X1 U7255 ( .A1(n4373), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5706) );
  MUX2_X1 U7256 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5706), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5709) );
  INV_X1 U7257 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7258 ( .A1(n5709), .A2(n5708), .ZN(n8302) );
  INV_X1 U7259 ( .A(n8302), .ZN(n5710) );
  NAND2_X1 U7260 ( .A1(n5711), .A2(n5710), .ZN(n6112) );
  OR2_X2 U7261 ( .A1(n6112), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7262 ( .A1(n5712), .A2(n8302), .ZN(n6357) );
  NAND2_X1 U7263 ( .A1(n5714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5715) );
  MUX2_X1 U7264 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5715), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5716) );
  INV_X1 U7265 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7266 ( .A1(n5718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5720) );
  INV_X1 U7267 ( .A(n7586), .ZN(n6270) );
  AND2_X1 U7268 ( .A1(n7588), .A2(n6270), .ZN(n6135) );
  NAND2_X1 U7269 ( .A1(n7389), .A2(n7586), .ZN(n6258) );
  INV_X1 U7270 ( .A(n5721), .ZN(n5722) );
  NAND2_X1 U7271 ( .A1(n5722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7272 ( .A1(n6009), .A2(n5723), .ZN(n5724) );
  NAND2_X1 U7273 ( .A1(n5724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7274 ( .A1(n7918), .A2(n7586), .ZN(n6163) );
  AND2_X1 U7275 ( .A1(n6258), .A2(n6163), .ZN(n5726) );
  XNOR2_X1 U7276 ( .A(n8213), .B(n7622), .ZN(n7619) );
  XOR2_X1 U7277 ( .A(n7956), .B(n7619), .Z(n6144) );
  NAND2_X1 U7278 ( .A1(n7219), .A2(n7542), .ZN(n5728) );
  OR2_X1 U7279 ( .A1(n7543), .A2(n9960), .ZN(n5727) );
  XNOR2_X1 U7280 ( .A(n7997), .B(n5928), .ZN(n6080) );
  NAND2_X1 U7281 ( .A1(n6061), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7282 ( .A1(n6072), .A2(n5729), .ZN(n7996) );
  NAND2_X1 U7283 ( .A1(n7996), .A2(n6229), .ZN(n5734) );
  INV_X1 U7284 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U7285 ( .A1(n5775), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7286 ( .A1(n6103), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U7287 ( .C1(n7995), .C2(n6594), .A(n5731), .B(n5730), .ZN(n5732)
         );
  INV_X1 U7288 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7289 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5735) );
  MUX2_X1 U7290 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5735), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5738) );
  INV_X1 U7291 ( .A(n5736), .ZN(n5737) );
  INV_X1 U7292 ( .A(n5750), .ZN(n5749) );
  INV_X1 U7293 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5740) );
  INV_X1 U7294 ( .A(n5741), .ZN(n5742) );
  INV_X1 U7295 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7297 ( .A1(n4306), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7298 ( .A1(n5750), .A2(n6178), .ZN(n5766) );
  INV_X1 U7299 ( .A(n6659), .ZN(n5765) );
  INV_X1 U7300 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6581) );
  INV_X1 U7301 ( .A(SI_0_), .ZN(n5753) );
  INV_X1 U7302 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5752) );
  OAI21_X1 U7303 ( .B1(n8613), .B2(n5753), .A(n5752), .ZN(n5755) );
  NAND2_X1 U7304 ( .A1(n5755), .A2(n5754), .ZN(n6305) );
  MUX2_X1 U7305 ( .A(n6581), .B(n6305), .S(n6378), .Z(n8196) );
  INV_X1 U7306 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9782) );
  INV_X1 U7307 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7308 ( .A1(n5756), .A2(n5758), .ZN(n5759) );
  INV_X1 U7309 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7310 ( .A1(n5741), .A2(n6406), .ZN(n5761) );
  NAND3_X1 U7311 ( .A1(n5762), .A2(n4861), .A3(n5761), .ZN(n6353) );
  INV_X1 U7312 ( .A(n6353), .ZN(n5763) );
  AOI21_X1 U7313 ( .B1(n5928), .B2(n8196), .A(n6726), .ZN(n6660) );
  NAND2_X1 U7314 ( .A1(n6657), .A2(n5766), .ZN(n6693) );
  INV_X1 U7315 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6309) );
  OR2_X1 U7316 ( .A1(n7543), .A2(n6309), .ZN(n5774) );
  OR2_X1 U7317 ( .A1(n5772), .A2(n6315), .ZN(n5773) );
  OAI211_X1 U7318 ( .C1(n6378), .C2(n6411), .A(n5774), .B(n5773), .ZN(n8128)
         );
  NAND2_X1 U7319 ( .A1(n5775), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5781) );
  OR2_X1 U7320 ( .A1(n5744), .A2(n9792), .ZN(n5780) );
  INV_X1 U7321 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5776) );
  OR2_X1 U7322 ( .A1(n4307), .A2(n5776), .ZN(n5779) );
  INV_X1 U7323 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5777) );
  OR2_X1 U7324 ( .A1(n5741), .A2(n5777), .ZN(n5778) );
  NAND4_X2 U7325 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n6181)
         );
  XNOR2_X1 U7326 ( .A(n5782), .B(n6181), .ZN(n6694) );
  NAND2_X1 U7327 ( .A1(n6693), .A2(n6694), .ZN(n6692) );
  INV_X1 U7328 ( .A(n6181), .ZN(n6729) );
  NAND2_X1 U7329 ( .A1(n5782), .A2(n6729), .ZN(n5783) );
  NAND2_X1 U7330 ( .A1(n6692), .A2(n5783), .ZN(n6826) );
  NAND2_X1 U7331 ( .A1(n5770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5784) );
  MUX2_X1 U7332 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5784), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5786) );
  NAND2_X1 U7333 ( .A1(n5786), .A2(n5785), .ZN(n6494) );
  OR2_X1 U7334 ( .A1(n7543), .A2(n6322), .ZN(n5788) );
  OR2_X1 U7335 ( .A1(n5772), .A2(n6321), .ZN(n5787) );
  OAI211_X1 U7336 ( .C1(n6378), .C2(n6494), .A(n5788), .B(n5787), .ZN(n6240)
         );
  XNOR2_X1 U7337 ( .A(n5739), .B(n6240), .ZN(n5819) );
  NAND2_X1 U7338 ( .A1(n6103), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5793) );
  INV_X1 U7339 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6413) );
  OR2_X1 U7340 ( .A1(n6589), .A2(n6413), .ZN(n5792) );
  OR2_X1 U7341 ( .A1(n4307), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5791) );
  INV_X1 U7342 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6414) );
  XNOR2_X1 U7343 ( .A(n5819), .B(n8119), .ZN(n6827) );
  NAND2_X1 U7344 ( .A1(n5785), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  OR2_X1 U7345 ( .A1(n5772), .A2(n6311), .ZN(n5797) );
  OR2_X1 U7346 ( .A1(n7543), .A2(n6312), .ZN(n5796) );
  OAI211_X1 U7347 ( .C1(n6378), .C2(n6427), .A(n5797), .B(n5796), .ZN(n6188)
         );
  XNOR2_X1 U7348 ( .A(n5739), .B(n6188), .ZN(n5815) );
  NAND2_X1 U7349 ( .A1(n5775), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5802) );
  OR2_X1 U7350 ( .A1(n5744), .A2(n9802), .ZN(n5801) );
  INV_X1 U7351 ( .A(n5798), .ZN(n5809) );
  NAND2_X1 U7352 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5799) );
  AND2_X1 U7353 ( .A1(n5809), .A2(n5799), .ZN(n6949) );
  OR2_X1 U7354 ( .A1(n4307), .A2(n6949), .ZN(n5800) );
  INV_X1 U7355 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U7356 ( .A1(n5815), .A2(n6868), .ZN(n5818) );
  INV_X1 U7357 ( .A(n5818), .ZN(n6863) );
  OR2_X1 U7358 ( .A1(n6827), .A2(n6863), .ZN(n5803) );
  OR2_X1 U7359 ( .A1(n6826), .A2(n5803), .ZN(n5822) );
  OR2_X1 U7360 ( .A1(n5804), .A2(n5904), .ZN(n5806) );
  XNOR2_X1 U7361 ( .A(n5806), .B(n5805), .ZN(n6605) );
  OR2_X1 U7362 ( .A1(n5772), .A2(n6319), .ZN(n5808) );
  OR2_X1 U7363 ( .A1(n7543), .A2(n6318), .ZN(n5807) );
  OAI211_X1 U7364 ( .C1(n6378), .C2(n6605), .A(n5808), .B(n5807), .ZN(n9837)
         );
  XNOR2_X1 U7365 ( .A(n7622), .B(n9837), .ZN(n5823) );
  NAND2_X1 U7366 ( .A1(n6103), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7367 ( .A1(n6589), .A2(n4559), .ZN(n5813) );
  NAND2_X1 U7368 ( .A1(n5809), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5810) );
  AND2_X1 U7369 ( .A1(n5831), .A2(n5810), .ZN(n6965) );
  OR2_X1 U7370 ( .A1(n4307), .A2(n6965), .ZN(n5812) );
  INV_X1 U7371 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6443) );
  OR2_X1 U7372 ( .A1(n6594), .A2(n6443), .ZN(n5811) );
  XNOR2_X1 U7373 ( .A(n5823), .B(n7751), .ZN(n6862) );
  INV_X1 U7374 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7375 ( .A1(n5816), .A2(n4596), .ZN(n5817) );
  AND2_X1 U7376 ( .A1(n5818), .A2(n5817), .ZN(n6803) );
  INV_X1 U7377 ( .A(n5819), .ZN(n5820) );
  INV_X1 U7378 ( .A(n8119), .ZN(n7752) );
  NAND2_X1 U7379 ( .A1(n5820), .A2(n7752), .ZN(n6801) );
  AND2_X1 U7380 ( .A1(n6803), .A2(n6801), .ZN(n6802) );
  INV_X1 U7381 ( .A(n7751), .ZN(n6929) );
  NAND2_X1 U7382 ( .A1(n5823), .A2(n6929), .ZN(n5824) );
  OR2_X1 U7383 ( .A1(n5825), .A2(n5904), .ZN(n5827) );
  OR2_X1 U7384 ( .A1(n5772), .A2(n6324), .ZN(n5829) );
  OR2_X1 U7385 ( .A1(n7543), .A2(n6325), .ZN(n5828) );
  OAI211_X1 U7386 ( .C1(n6378), .C2(n6459), .A(n5829), .B(n5828), .ZN(n6815)
         );
  XNOR2_X1 U7387 ( .A(n7622), .B(n6815), .ZN(n5854) );
  NAND2_X1 U7388 ( .A1(n5775), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5836) );
  INV_X1 U7389 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5830) );
  OR2_X1 U7390 ( .A1(n5744), .A2(n5830), .ZN(n5835) );
  NAND2_X1 U7391 ( .A1(n5831), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5832) );
  AND2_X1 U7392 ( .A1(n5845), .A2(n5832), .ZN(n6934) );
  OR2_X1 U7393 ( .A1(n4307), .A2(n6934), .ZN(n5834) );
  INV_X1 U7394 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6821) );
  OR2_X1 U7395 ( .A1(n6594), .A2(n6821), .ZN(n5833) );
  XNOR2_X1 U7396 ( .A(n5854), .B(n6989), .ZN(n6927) );
  NAND2_X1 U7397 ( .A1(n5858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  INV_X1 U7398 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5839) );
  XNOR2_X1 U7399 ( .A(n5840), .B(n5839), .ZN(n6852) );
  NAND2_X1 U7400 ( .A1(n5841), .A2(n7542), .ZN(n5843) );
  INV_X1 U7401 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6326) );
  OR2_X1 U7402 ( .A1(n7543), .A2(n6326), .ZN(n5842) );
  OAI211_X1 U7403 ( .C1(n6378), .C2(n6852), .A(n5843), .B(n5842), .ZN(n6244)
         );
  XNOR2_X1 U7404 ( .A(n7622), .B(n6244), .ZN(n5851) );
  NAND2_X1 U7405 ( .A1(n6103), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5850) );
  INV_X1 U7406 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6470) );
  OR2_X1 U7407 ( .A1(n6589), .A2(n6470), .ZN(n5849) );
  INV_X1 U7408 ( .A(n5844), .ZN(n5865) );
  NAND2_X1 U7409 ( .A1(n5845), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5846) );
  AND2_X1 U7410 ( .A1(n5865), .A2(n5846), .ZN(n6994) );
  OR2_X1 U7411 ( .A1(n4307), .A2(n6994), .ZN(n5848) );
  INV_X1 U7412 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6471) );
  OR2_X1 U7413 ( .A1(n6594), .A2(n6471), .ZN(n5847) );
  NAND2_X1 U7414 ( .A1(n5851), .A2(n7090), .ZN(n7082) );
  INV_X1 U7415 ( .A(n5851), .ZN(n5852) );
  INV_X1 U7416 ( .A(n7090), .ZN(n7749) );
  NAND2_X1 U7417 ( .A1(n5852), .A2(n7749), .ZN(n5853) );
  AND2_X1 U7418 ( .A1(n7082), .A2(n5853), .ZN(n6985) );
  INV_X1 U7419 ( .A(n5854), .ZN(n5855) );
  INV_X1 U7420 ( .A(n6989), .ZN(n7750) );
  NAND2_X1 U7421 ( .A1(n5855), .A2(n7750), .ZN(n6982) );
  AND2_X1 U7422 ( .A1(n6985), .A2(n6982), .ZN(n5856) );
  NAND2_X1 U7423 ( .A1(n6984), .A2(n7082), .ZN(n5871) );
  NAND2_X1 U7424 ( .A1(n5857), .A2(n7542), .ZN(n5862) );
  NAND2_X1 U7425 ( .A1(n5874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  INV_X1 U7426 ( .A(n6854), .ZN(n9766) );
  AOI22_X1 U7427 ( .A1(n6020), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6303), .B2(
        n9766), .ZN(n5861) );
  NAND2_X1 U7428 ( .A1(n5862), .A2(n5861), .ZN(n6245) );
  XNOR2_X1 U7429 ( .A(n7622), .B(n6245), .ZN(n5872) );
  NAND2_X1 U7430 ( .A1(n6103), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5870) );
  INV_X1 U7431 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7432 ( .A1(n6589), .A2(n5863), .ZN(n5869) );
  INV_X1 U7433 ( .A(n5864), .ZN(n5880) );
  NAND2_X1 U7434 ( .A1(n5865), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5866) );
  AND2_X1 U7435 ( .A1(n5880), .A2(n5866), .ZN(n7094) );
  OR2_X1 U7436 ( .A1(n4307), .A2(n7094), .ZN(n5868) );
  INV_X1 U7437 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10006) );
  OR2_X1 U7438 ( .A1(n6594), .A2(n10006), .ZN(n5867) );
  NAND4_X1 U7439 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n7748)
         );
  XNOR2_X1 U7440 ( .A(n5872), .B(n7748), .ZN(n7083) );
  INV_X1 U7441 ( .A(n7748), .ZN(n6937) );
  NAND2_X1 U7442 ( .A1(n5872), .A2(n6937), .ZN(n5873) );
  NAND2_X1 U7443 ( .A1(n6332), .A2(n7542), .ZN(n5879) );
  NAND2_X1 U7444 ( .A1(n5875), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5877) );
  INV_X1 U7445 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U7446 ( .A1(n5876), .A2(n5901), .ZN(n5897) );
  AOI22_X1 U7447 ( .A1(n6020), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6303), .B2(
        n7028), .ZN(n5878) );
  XNOR2_X1 U7448 ( .A(n7622), .B(n9819), .ZN(n5887) );
  NAND2_X1 U7449 ( .A1(n6103), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5885) );
  INV_X1 U7450 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6836) );
  OR2_X1 U7451 ( .A1(n6589), .A2(n6836), .ZN(n5884) );
  NAND2_X1 U7452 ( .A1(n5880), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5881) );
  AND2_X1 U7453 ( .A1(n5889), .A2(n5881), .ZN(n7233) );
  OR2_X1 U7454 ( .A1(n4307), .A2(n7233), .ZN(n5883) );
  INV_X1 U7455 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6837) );
  OR2_X1 U7456 ( .A1(n6594), .A2(n6837), .ZN(n5882) );
  NAND4_X1 U7457 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n7747)
         );
  XNOR2_X1 U7458 ( .A(n5887), .B(n7747), .ZN(n7242) );
  NAND2_X1 U7459 ( .A1(n5887), .A2(n7747), .ZN(n5888) );
  NAND2_X1 U7460 ( .A1(n7239), .A2(n5888), .ZN(n7290) );
  NAND2_X1 U7461 ( .A1(n6103), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5896) );
  INV_X1 U7462 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7005) );
  OR2_X1 U7463 ( .A1(n6594), .A2(n7005), .ZN(n5895) );
  NAND2_X1 U7464 ( .A1(n5889), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5890) );
  AND2_X1 U7465 ( .A1(n5908), .A2(n5890), .ZN(n7295) );
  OR2_X1 U7466 ( .A1(n4307), .A2(n7295), .ZN(n5894) );
  INV_X1 U7467 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5892) );
  OR2_X1 U7468 ( .A1(n6589), .A2(n5892), .ZN(n5893) );
  NAND2_X1 U7469 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5898) );
  INV_X1 U7470 ( .A(n7134), .ZN(n7037) );
  AOI22_X1 U7471 ( .A1(n6020), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6303), .B2(
        n7037), .ZN(n5899) );
  XNOR2_X1 U7472 ( .A(n7622), .B(n7294), .ZN(n7291) );
  NAND2_X1 U7473 ( .A1(n6345), .A2(n7542), .ZN(n5907) );
  NAND2_X1 U7474 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  OR2_X1 U7475 ( .A1(n5915), .A2(n5904), .ZN(n5905) );
  XNOR2_X1 U7476 ( .A(n5905), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7171) );
  AOI22_X1 U7477 ( .A1(n6020), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6303), .B2(
        n7171), .ZN(n5906) );
  NAND2_X1 U7478 ( .A1(n5907), .A2(n5906), .ZN(n7352) );
  NAND2_X1 U7479 ( .A1(n6103), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5913) );
  INV_X1 U7480 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7167) );
  OR2_X1 U7481 ( .A1(n6589), .A2(n7167), .ZN(n5912) );
  NAND2_X1 U7482 ( .A1(n5908), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5909) );
  AND2_X1 U7483 ( .A1(n5920), .A2(n5909), .ZN(n7097) );
  OR2_X1 U7484 ( .A1(n4307), .A2(n7097), .ZN(n5911) );
  INV_X1 U7485 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7142) );
  OR2_X1 U7486 ( .A1(n6594), .A2(n7142), .ZN(n5910) );
  NAND2_X1 U7487 ( .A1(n7352), .A2(n7647), .ZN(n7441) );
  NAND2_X1 U7488 ( .A1(n7440), .A2(n7441), .ZN(n7570) );
  XNOR2_X1 U7489 ( .A(n7570), .B(n5928), .ZN(n7646) );
  OAI21_X1 U7490 ( .B1(n7345), .B2(n7291), .A(n7646), .ZN(n5932) );
  NAND2_X1 U7491 ( .A1(n6351), .A2(n7542), .ZN(n5918) );
  NAND2_X1 U7492 ( .A1(n5915), .A2(n5914), .ZN(n5935) );
  NAND2_X1 U7493 ( .A1(n5935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U7494 ( .A(n5916), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7149) );
  AOI22_X1 U7495 ( .A1(n6020), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6303), .B2(
        n7149), .ZN(n5917) );
  NAND2_X1 U7496 ( .A1(n5918), .A2(n5917), .ZN(n7653) );
  XNOR2_X1 U7497 ( .A(n7653), .B(n7622), .ZN(n5933) );
  NAND2_X1 U7498 ( .A1(n5775), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5925) );
  INV_X1 U7499 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7208) );
  OR2_X1 U7500 ( .A1(n5744), .A2(n7208), .ZN(n5924) );
  INV_X1 U7501 ( .A(n5919), .ZN(n5939) );
  NAND2_X1 U7502 ( .A1(n5920), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5921) );
  AND2_X1 U7503 ( .A1(n5939), .A2(n5921), .ZN(n7225) );
  OR2_X1 U7504 ( .A1(n4307), .A2(n7225), .ZN(n5923) );
  INV_X1 U7505 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7224) );
  OR2_X1 U7506 ( .A1(n6594), .A2(n7224), .ZN(n5922) );
  NAND4_X1 U7507 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n7744)
         );
  XNOR2_X1 U7508 ( .A(n5933), .B(n7744), .ZN(n7648) );
  NAND3_X1 U7509 ( .A1(n7622), .A2(n7345), .A3(n7294), .ZN(n5926) );
  OAI21_X1 U7510 ( .B1(n7622), .B2(n7745), .A(n5926), .ZN(n5930) );
  INV_X1 U7511 ( .A(n7294), .ZN(n9825) );
  NAND3_X1 U7512 ( .A1(n5928), .A2(n7345), .A3(n9825), .ZN(n5927) );
  OAI211_X1 U7513 ( .C1(n5928), .C2(n7745), .A(n7570), .B(n5927), .ZN(n5929)
         );
  OAI21_X1 U7514 ( .B1(n7570), .B2(n5930), .A(n5929), .ZN(n5931) );
  INV_X1 U7515 ( .A(n5933), .ZN(n5934) );
  NAND2_X1 U7516 ( .A1(n6368), .A2(n7542), .ZN(n5938) );
  NAND2_X1 U7517 ( .A1(n5936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7518 ( .A(n5949), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7789) );
  AOI22_X1 U7519 ( .A1(n6020), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6303), .B2(
        n7789), .ZN(n5937) );
  XNOR2_X1 U7520 ( .A(n8110), .B(n7622), .ZN(n5945) );
  NAND2_X1 U7521 ( .A1(n6103), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5944) );
  INV_X1 U7522 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7755) );
  OR2_X1 U7523 ( .A1(n6594), .A2(n7755), .ZN(n5943) );
  NAND2_X1 U7524 ( .A1(n5939), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5940) );
  AND2_X1 U7525 ( .A1(n5956), .A2(n5940), .ZN(n8105) );
  OR2_X1 U7526 ( .A1(n4307), .A2(n8105), .ZN(n5942) );
  INV_X1 U7527 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7764) );
  OR2_X1 U7528 ( .A1(n6589), .A2(n7764), .ZN(n5941) );
  NAND2_X1 U7529 ( .A1(n5945), .A2(n7644), .ZN(n7322) );
  INV_X1 U7530 ( .A(n5945), .ZN(n5946) );
  NAND2_X1 U7531 ( .A1(n5946), .A2(n7743), .ZN(n5947) );
  NAND2_X1 U7532 ( .A1(n7322), .A2(n5947), .ZN(n7304) );
  NAND2_X1 U7533 ( .A1(n6452), .A2(n7542), .ZN(n5955) );
  NAND2_X1 U7534 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7535 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7536 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7537 ( .A1(n5952), .A2(n5951), .ZN(n5962) );
  AOI22_X1 U7538 ( .A1(n6020), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6303), .B2(
        n7797), .ZN(n5954) );
  XNOR2_X1 U7539 ( .A(n8279), .B(n7622), .ZN(n5974) );
  NAND2_X1 U7540 ( .A1(n6103), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5961) );
  INV_X1 U7541 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8191) );
  OR2_X1 U7542 ( .A1(n6589), .A2(n8191), .ZN(n5960) );
  NAND2_X1 U7543 ( .A1(n5956), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5957) );
  AND2_X1 U7544 ( .A1(n5967), .A2(n5957), .ZN(n7330) );
  OR2_X1 U7545 ( .A1(n4307), .A2(n7330), .ZN(n5959) );
  INV_X1 U7546 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7792) );
  OR2_X1 U7547 ( .A1(n6594), .A2(n7792), .ZN(n5958) );
  NAND4_X1 U7548 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n8097)
         );
  XNOR2_X1 U7549 ( .A(n5974), .B(n8097), .ZN(n7323) );
  INV_X1 U7550 ( .A(n7323), .ZN(n5973) );
  NAND2_X1 U7551 ( .A1(n6477), .A2(n7542), .ZN(n5965) );
  NAND2_X1 U7552 ( .A1(n5962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7553 ( .A(n5963), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7835) );
  AOI22_X1 U7554 ( .A1(n7835), .A2(n6303), .B1(n6020), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7555 ( .A1(n5965), .A2(n5964), .ZN(n8186) );
  XNOR2_X1 U7556 ( .A(n8186), .B(n5928), .ZN(n5978) );
  NAND2_X1 U7557 ( .A1(n6103), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5972) );
  INV_X1 U7558 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8184) );
  OR2_X1 U7559 ( .A1(n6589), .A2(n8184), .ZN(n5971) );
  INV_X1 U7560 ( .A(n5966), .ZN(n5987) );
  NAND2_X1 U7561 ( .A1(n5967), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5968) );
  AND2_X1 U7562 ( .A1(n5987), .A2(n5968), .ZN(n8091) );
  OR2_X1 U7563 ( .A1(n4307), .A2(n8091), .ZN(n5970) );
  INV_X1 U7564 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7802) );
  OR2_X1 U7565 ( .A1(n6594), .A2(n7802), .ZN(n5969) );
  NAND4_X1 U7566 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n8076)
         );
  XNOR2_X1 U7567 ( .A(n5978), .B(n8076), .ZN(n7312) );
  INV_X1 U7568 ( .A(n7312), .ZN(n5976) );
  OR2_X1 U7569 ( .A1(n5973), .A2(n7322), .ZN(n7325) );
  INV_X1 U7570 ( .A(n8097), .ZN(n7317) );
  NAND2_X1 U7571 ( .A1(n5974), .A2(n7317), .ZN(n5975) );
  AND2_X1 U7572 ( .A1(n7325), .A2(n5975), .ZN(n7311) );
  AND2_X1 U7573 ( .A1(n5976), .A2(n7311), .ZN(n5977) );
  NAND2_X1 U7574 ( .A1(n5978), .A2(n8076), .ZN(n5979) );
  NAND2_X1 U7575 ( .A1(n6653), .A2(n7542), .ZN(n5985) );
  NAND2_X1 U7576 ( .A1(n5981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7577 ( .A(n5983), .B(n5982), .ZN(n7853) );
  INV_X1 U7578 ( .A(n7853), .ZN(n7843) );
  AOI22_X1 U7579 ( .A1(n6020), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6303), .B2(
        n7843), .ZN(n5984) );
  XNOR2_X1 U7580 ( .A(n8179), .B(n7622), .ZN(n5994) );
  NAND2_X1 U7581 ( .A1(n6103), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5993) );
  INV_X1 U7582 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8081) );
  OR2_X1 U7583 ( .A1(n6594), .A2(n8081), .ZN(n5992) );
  INV_X1 U7584 ( .A(n5986), .ZN(n6000) );
  NAND2_X1 U7585 ( .A1(n5987), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5988) );
  AND2_X1 U7586 ( .A1(n6000), .A2(n5988), .ZN(n8083) );
  OR2_X1 U7587 ( .A1(n4307), .A2(n8083), .ZN(n5991) );
  INV_X1 U7588 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7589 ( .A1(n6589), .A2(n5989), .ZN(n5990) );
  NAND4_X1 U7590 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n8098)
         );
  XNOR2_X1 U7591 ( .A(n5994), .B(n8098), .ZN(n7336) );
  INV_X1 U7592 ( .A(n5994), .ZN(n5995) );
  NAND2_X1 U7593 ( .A1(n6702), .A2(n7542), .ZN(n5999) );
  NAND2_X1 U7594 ( .A1(n5996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7595 ( .A(n5997), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7884) );
  AOI22_X1 U7596 ( .A1(n6020), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6303), .B2(
        n7884), .ZN(n5998) );
  XNOR2_X1 U7597 ( .A(n8261), .B(n7622), .ZN(n6006) );
  NAND2_X1 U7598 ( .A1(n6103), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6005) );
  INV_X1 U7599 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8064) );
  OR2_X1 U7600 ( .A1(n6594), .A2(n8064), .ZN(n6004) );
  NAND2_X1 U7601 ( .A1(n6000), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6001) );
  AND2_X1 U7602 ( .A1(n6012), .A2(n6001), .ZN(n7666) );
  OR2_X1 U7603 ( .A1(n4307), .A2(n7666), .ZN(n6003) );
  INV_X1 U7604 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9981) );
  OR2_X1 U7605 ( .A1(n6589), .A2(n9981), .ZN(n6002) );
  NAND2_X1 U7606 ( .A1(n6006), .A2(n7338), .ZN(n7710) );
  INV_X1 U7607 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7608 ( .A1(n6007), .A2(n8077), .ZN(n6008) );
  AND2_X1 U7609 ( .A1(n7710), .A2(n6008), .ZN(n7664) );
  NAND2_X1 U7610 ( .A1(n6761), .A2(n7542), .ZN(n6011) );
  XNOR2_X1 U7611 ( .A(n6009), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7904) );
  AOI22_X1 U7612 ( .A1(n6020), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6303), .B2(
        n7904), .ZN(n6010) );
  XNOR2_X1 U7613 ( .A(n8255), .B(n7622), .ZN(n6018) );
  NAND2_X1 U7614 ( .A1(n6012), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7615 ( .A1(n6024), .A2(n6013), .ZN(n8055) );
  NAND2_X1 U7616 ( .A1(n6229), .A2(n8055), .ZN(n6017) );
  INV_X1 U7617 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8174) );
  OR2_X1 U7618 ( .A1(n6589), .A2(n8174), .ZN(n6016) );
  INV_X1 U7619 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8254) );
  OR2_X1 U7620 ( .A1(n5744), .A2(n8254), .ZN(n6015) );
  INV_X1 U7621 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8054) );
  OR2_X1 U7622 ( .A1(n6594), .A2(n8054), .ZN(n6014) );
  NAND4_X1 U7623 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n8062)
         );
  XNOR2_X1 U7624 ( .A(n6018), .B(n8062), .ZN(n7711) );
  NAND2_X1 U7625 ( .A1(n6018), .A2(n8041), .ZN(n6019) );
  NAND2_X1 U7626 ( .A1(n7713), .A2(n6019), .ZN(n7612) );
  NAND2_X1 U7627 ( .A1(n6882), .A2(n7542), .ZN(n6022) );
  AOI22_X1 U7628 ( .A1(n6020), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7896), .B2(
        n6303), .ZN(n6021) );
  XNOR2_X1 U7629 ( .A(n8249), .B(n5928), .ZN(n6042) );
  INV_X1 U7630 ( .A(n6023), .ZN(n6034) );
  NAND2_X1 U7631 ( .A1(n6024), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7632 ( .A1(n6034), .A2(n6025), .ZN(n8047) );
  NAND2_X1 U7633 ( .A1(n8047), .A2(n6229), .ZN(n6029) );
  NAND2_X1 U7634 ( .A1(n6103), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7635 ( .A1(n6230), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7636 ( .A1(n5775), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6026) );
  NAND4_X1 U7637 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n8052)
         );
  XNOR2_X1 U7638 ( .A(n6042), .B(n8052), .ZN(n7611) );
  NOR2_X1 U7639 ( .A1(n7612), .A2(n7611), .ZN(n6030) );
  NAND2_X1 U7640 ( .A1(n6944), .A2(n7542), .ZN(n6032) );
  OR2_X1 U7641 ( .A1(n7543), .A2(n10011), .ZN(n6031) );
  XNOR2_X1 U7642 ( .A(n7686), .B(n7622), .ZN(n6039) );
  INV_X1 U7643 ( .A(n6033), .ZN(n6046) );
  NAND2_X1 U7644 ( .A1(n6034), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7645 ( .A1(n6046), .A2(n6035), .ZN(n8031) );
  NAND2_X1 U7646 ( .A1(n8031), .A2(n6229), .ZN(n6038) );
  AOI22_X1 U7647 ( .A1(n5775), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6103), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7648 ( .A1(n6230), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7649 ( .A1(n6039), .A2(n8042), .ZN(n7630) );
  INV_X1 U7650 ( .A(n6039), .ZN(n6040) );
  INV_X1 U7651 ( .A(n8042), .ZN(n7742) );
  NAND2_X1 U7652 ( .A1(n6040), .A2(n7742), .ZN(n6041) );
  NAND2_X1 U7653 ( .A1(n7630), .A2(n6041), .ZN(n7688) );
  AND2_X1 U7654 ( .A1(n6042), .A2(n8052), .ZN(n7687) );
  NOR2_X1 U7655 ( .A1(n7688), .A2(n7687), .ZN(n6043) );
  NAND2_X1 U7656 ( .A1(n6995), .A2(n7542), .ZN(n6045) );
  OR2_X1 U7657 ( .A1(n7543), .A2(n6996), .ZN(n6044) );
  XNOR2_X1 U7658 ( .A(n8163), .B(n7622), .ZN(n6051) );
  INV_X1 U7659 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7660 ( .A1(n6046), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7661 ( .A1(n6059), .A2(n6047), .ZN(n8019) );
  NAND2_X1 U7662 ( .A1(n8019), .A2(n6229), .ZN(n6049) );
  AOI22_X1 U7663 ( .A1(n5775), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6103), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U7664 ( .C1(n6594), .C2(n6050), .A(n6049), .B(n6048), .ZN(n8027)
         );
  XNOR2_X1 U7665 ( .A(n6051), .B(n8027), .ZN(n7631) );
  NAND2_X1 U7666 ( .A1(n6051), .A2(n8004), .ZN(n6052) );
  NAND2_X1 U7667 ( .A1(n7101), .A2(n7542), .ZN(n6054) );
  OR2_X1 U7668 ( .A1(n7543), .A2(n7103), .ZN(n6053) );
  XNOR2_X1 U7669 ( .A(n8159), .B(n7622), .ZN(n6056) );
  INV_X1 U7670 ( .A(n6055), .ZN(n6058) );
  INV_X1 U7671 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7672 ( .A1(n6059), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7673 ( .A1(n6061), .A2(n6060), .ZN(n8009) );
  NAND2_X1 U7674 ( .A1(n8009), .A2(n6229), .ZN(n6067) );
  INV_X1 U7675 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7676 ( .A1(n5775), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7677 ( .A1(n6103), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6062) );
  OAI211_X1 U7678 ( .C1(n6064), .C2(n6594), .A(n6063), .B(n6062), .ZN(n6065)
         );
  INV_X1 U7679 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7680 ( .A1(n6067), .A2(n6066), .ZN(n7741) );
  AND2_X2 U7681 ( .A1(n7699), .A2(n6068), .ZN(n7602) );
  OAI21_X1 U7682 ( .B1(n6080), .B2(n7980), .A(n7602), .ZN(n6082) );
  NAND2_X1 U7683 ( .A1(n7229), .A2(n7542), .ZN(n6070) );
  OR2_X1 U7684 ( .A1(n7543), .A2(n7278), .ZN(n6069) );
  XNOR2_X1 U7685 ( .A(n8226), .B(n5928), .ZN(n6079) );
  INV_X1 U7686 ( .A(n6071), .ZN(n6087) );
  NAND2_X1 U7687 ( .A1(n6072), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7688 ( .A1(n6087), .A2(n6073), .ZN(n7982) );
  NAND2_X1 U7689 ( .A1(n7982), .A2(n6229), .ZN(n6078) );
  INV_X1 U7690 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U7691 ( .A1(n5775), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7692 ( .A1(n6103), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7693 ( .C1(n7986), .C2(n6594), .A(n6075), .B(n6074), .ZN(n6076)
         );
  INV_X1 U7694 ( .A(n6076), .ZN(n6077) );
  NOR2_X1 U7695 ( .A1(n6079), .A2(n7964), .ZN(n6083) );
  AOI21_X1 U7696 ( .B1(n6079), .B2(n7964), .A(n6083), .ZN(n7675) );
  INV_X1 U7697 ( .A(n6080), .ZN(n7603) );
  NAND2_X1 U7698 ( .A1(n6082), .A2(n6081), .ZN(n7677) );
  INV_X1 U7699 ( .A(n6083), .ZN(n7657) );
  NAND2_X1 U7700 ( .A1(n7275), .A2(n7542), .ZN(n6085) );
  OR2_X1 U7701 ( .A1(n7543), .A2(n7276), .ZN(n6084) );
  XNOR2_X1 U7702 ( .A(n7655), .B(n7622), .ZN(n6094) );
  INV_X1 U7703 ( .A(n6086), .ZN(n6100) );
  NAND2_X1 U7704 ( .A1(n6087), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7705 ( .A1(n6100), .A2(n6088), .ZN(n7966) );
  NAND2_X1 U7706 ( .A1(n7966), .A2(n6229), .ZN(n6093) );
  INV_X1 U7707 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U7708 ( .A1(n6103), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7709 ( .A1(n5775), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7710 ( .C1(n7977), .C2(n6594), .A(n6090), .B(n6089), .ZN(n6091)
         );
  INV_X1 U7711 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7712 ( .A1(n6094), .A2(n7509), .ZN(n6097) );
  INV_X1 U7713 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7714 ( .A1(n6095), .A2(n7979), .ZN(n6096) );
  NAND2_X1 U7715 ( .A1(n6097), .A2(n6096), .ZN(n7656) );
  INV_X1 U7716 ( .A(n6097), .ZN(n7724) );
  NAND2_X1 U7717 ( .A1(n8299), .A2(n7542), .ZN(n6099) );
  OR2_X1 U7718 ( .A1(n7543), .A2(n8301), .ZN(n6098) );
  XNOR2_X1 U7719 ( .A(n8219), .B(n7622), .ZN(n6109) );
  NAND2_X1 U7720 ( .A1(n6100), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7721 ( .A1(n6102), .A2(n6101), .ZN(n7959) );
  NAND2_X1 U7722 ( .A1(n7959), .A2(n6229), .ZN(n6108) );
  INV_X1 U7723 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U7724 ( .A1(n5775), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7725 ( .A1(n6103), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6104) );
  OAI211_X1 U7726 ( .C1(n7958), .C2(n6594), .A(n6105), .B(n6104), .ZN(n6106)
         );
  INV_X1 U7727 ( .A(n6106), .ZN(n6107) );
  XNOR2_X1 U7728 ( .A(n6109), .B(n7963), .ZN(n7723) );
  NAND2_X1 U7729 ( .A1(n6109), .A2(n6110), .ZN(n6111) );
  NAND2_X1 U7730 ( .A1(n7277), .A2(n8302), .ZN(n6113) );
  INV_X1 U7731 ( .A(n6273), .ZN(n8286) );
  NOR2_X1 U7732 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n10031) );
  NOR4_X1 U7733 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6118) );
  NOR4_X1 U7734 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6117) );
  NOR4_X1 U7735 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6116) );
  NAND4_X1 U7736 ( .A1(n10031), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n6124)
         );
  NOR4_X1 U7737 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6122) );
  NOR4_X1 U7738 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6121) );
  NOR4_X1 U7739 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6120) );
  NOR4_X1 U7740 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6119) );
  NAND4_X1 U7741 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n6123)
         );
  NOR2_X1 U7742 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  INV_X1 U7743 ( .A(n6280), .ZN(n6126) );
  NAND2_X1 U7744 ( .A1(n6706), .A2(n6126), .ZN(n6162) );
  INV_X1 U7745 ( .A(n6162), .ZN(n6131) );
  NOR2_X1 U7746 ( .A1(n5712), .A2(n8302), .ZN(n6127) );
  NAND2_X1 U7747 ( .A1(n6128), .A2(n6127), .ZN(n6300) );
  NAND2_X1 U7748 ( .A1(n6132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  AND2_X1 U7749 ( .A1(n7535), .A2(n9824), .ZN(n6137) );
  NAND2_X1 U7750 ( .A1(n7596), .A2(n7896), .ZN(n6237) );
  INV_X1 U7751 ( .A(n6135), .ZN(n6136) );
  NAND2_X1 U7752 ( .A1(n6137), .A2(n6287), .ZN(n6161) );
  INV_X1 U7753 ( .A(n6161), .ZN(n6138) );
  NAND2_X1 U7754 ( .A1(n6290), .A2(n6138), .ZN(n6142) );
  INV_X1 U7755 ( .A(n6287), .ZN(n6140) );
  NAND2_X1 U7756 ( .A1(n6292), .A2(n6140), .ZN(n6141) );
  AOI211_X1 U7757 ( .C1(n6144), .C2(n6143), .A(n7707), .B(n7620), .ZN(n6177)
         );
  NAND2_X1 U7758 ( .A1(n6290), .A2(n8111), .ZN(n6145) );
  NAND2_X1 U7759 ( .A1(n9791), .A2(n7588), .ZN(n6281) );
  NAND2_X1 U7760 ( .A1(n8213), .A2(n7705), .ZN(n6175) );
  NAND2_X1 U7761 ( .A1(n6146), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7762 ( .A1(n7378), .A2(n6147), .ZN(n7940) );
  NAND2_X1 U7763 ( .A1(n7940), .A2(n6229), .ZN(n6152) );
  INV_X1 U7764 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U7765 ( .A1(n5775), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7766 ( .A1(n6230), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7767 ( .C1(n5744), .C2(n9996), .A(n6149), .B(n6148), .ZN(n6150)
         );
  INV_X1 U7768 ( .A(n6150), .ZN(n6151) );
  INV_X1 U7769 ( .A(n7946), .ZN(n7524) );
  INV_X1 U7770 ( .A(n6292), .ZN(n6159) );
  INV_X1 U7771 ( .A(n6163), .ZN(n6153) );
  INV_X1 U7772 ( .A(n6288), .ZN(n6710) );
  INV_X1 U7773 ( .A(n6154), .ZN(n7593) );
  NAND2_X1 U7774 ( .A1(n7593), .A2(n7906), .ZN(n6157) );
  NAND2_X1 U7775 ( .A1(n6378), .A2(n6157), .ZN(n6266) );
  NAND2_X1 U7776 ( .A1(n6710), .A2(n6266), .ZN(n6158) );
  NOR2_X1 U7777 ( .A1(n6288), .A2(n6266), .ZN(n6160) );
  AOI22_X1 U7778 ( .A1(n7963), .A2(n7729), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6172) );
  INV_X1 U7779 ( .A(n6168), .ZN(n6166) );
  NAND2_X1 U7780 ( .A1(n6161), .A2(n7968), .ZN(n6291) );
  NAND2_X1 U7781 ( .A1(n6162), .A2(n6291), .ZN(n6165) );
  NAND2_X1 U7782 ( .A1(n7519), .A2(n6163), .ZN(n6277) );
  AND3_X1 U7783 ( .A1(n6300), .A2(n6301), .A3(n6277), .ZN(n6164) );
  OAI211_X1 U7784 ( .C1(n6166), .C2(n6287), .A(n6165), .B(n6164), .ZN(n6167)
         );
  NAND2_X1 U7785 ( .A1(n6167), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6170) );
  NOR2_X1 U7786 ( .A1(n6278), .A2(n6288), .ZN(n7594) );
  NAND2_X1 U7787 ( .A1(n6168), .A2(n7594), .ZN(n6169) );
  NAND2_X1 U7788 ( .A1(n7734), .A2(n7949), .ZN(n6171) );
  OAI211_X1 U7789 ( .C1(n7524), .C2(n7731), .A(n6172), .B(n6171), .ZN(n6173)
         );
  INV_X1 U7790 ( .A(n6173), .ZN(n6174) );
  INV_X1 U7791 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7792 ( .A1(n6178), .A2(n6180), .ZN(n7390) );
  INV_X1 U7793 ( .A(n8196), .ZN(n6730) );
  NAND2_X1 U7794 ( .A1(n6353), .A2(n6730), .ZN(n6179) );
  NAND2_X1 U7795 ( .A1(n6178), .A2(n9783), .ZN(n8121) );
  NAND2_X1 U7796 ( .A1(n6728), .A2(n8121), .ZN(n6183) );
  INV_X1 U7797 ( .A(n8128), .ZN(n6698) );
  OR2_X1 U7798 ( .A1(n6181), .A2(n6698), .ZN(n7394) );
  NAND2_X1 U7799 ( .A1(n6181), .A2(n6698), .ZN(n7395) );
  NAND2_X1 U7800 ( .A1(n7394), .A2(n7395), .ZN(n6182) );
  OR2_X1 U7801 ( .A1(n6181), .A2(n8128), .ZN(n6184) );
  INV_X1 U7802 ( .A(n6240), .ZN(n9795) );
  OR2_X1 U7803 ( .A1(n8119), .A2(n9795), .ZN(n6185) );
  NAND2_X1 U7804 ( .A1(n6956), .A2(n6185), .ZN(n6187) );
  NAND2_X1 U7805 ( .A1(n8119), .A2(n9795), .ZN(n6186) );
  NAND2_X1 U7806 ( .A1(n6187), .A2(n6186), .ZN(n6945) );
  NAND2_X1 U7807 ( .A1(n6945), .A2(n6946), .ZN(n6190) );
  NAND2_X1 U7808 ( .A1(n6868), .A2(n4595), .ZN(n6189) );
  NAND2_X1 U7809 ( .A1(n6190), .A2(n6189), .ZN(n6963) );
  OR2_X1 U7810 ( .A1(n7751), .A2(n6966), .ZN(n7412) );
  NAND2_X1 U7811 ( .A1(n7751), .A2(n6966), .ZN(n7409) );
  NAND2_X1 U7812 ( .A1(n6963), .A2(n7561), .ZN(n6192) );
  OR2_X1 U7813 ( .A1(n7751), .A2(n9837), .ZN(n6191) );
  NAND2_X1 U7814 ( .A1(n6192), .A2(n6191), .ZN(n6817) );
  INV_X1 U7815 ( .A(n6817), .ZN(n6194) );
  OR2_X1 U7816 ( .A1(n6989), .A2(n6815), .ZN(n7414) );
  NAND2_X1 U7817 ( .A1(n6989), .A2(n6815), .ZN(n7413) );
  AND2_X1 U7818 ( .A1(n7414), .A2(n7413), .ZN(n7564) );
  INV_X1 U7819 ( .A(n6815), .ZN(n9805) );
  OR2_X1 U7820 ( .A1(n6989), .A2(n9805), .ZN(n6195) );
  INV_X1 U7821 ( .A(n6244), .ZN(n9809) );
  OR2_X1 U7822 ( .A1(n7090), .A2(n9809), .ZN(n6196) );
  INV_X1 U7823 ( .A(n7747), .ZN(n6878) );
  OR2_X1 U7824 ( .A1(n9819), .A2(n6878), .ZN(n6197) );
  NAND2_X1 U7825 ( .A1(n6936), .A2(n6197), .ZN(n6199) );
  NAND2_X1 U7826 ( .A1(n9819), .A2(n6878), .ZN(n6198) );
  NAND2_X1 U7827 ( .A1(n6199), .A2(n6198), .ZN(n6999) );
  NAND2_X1 U7828 ( .A1(n7294), .A2(n7746), .ZN(n6200) );
  OR2_X1 U7829 ( .A1(n7294), .A2(n7746), .ZN(n6201) );
  INV_X1 U7830 ( .A(n7570), .ZN(n7069) );
  NAND2_X1 U7831 ( .A1(n7352), .A2(n7745), .ZN(n6202) );
  AND2_X1 U7832 ( .A1(n7653), .A2(n7744), .ZN(n6204) );
  OR2_X1 U7833 ( .A1(n7653), .A2(n7744), .ZN(n6203) );
  NAND2_X1 U7834 ( .A1(n8110), .A2(n7743), .ZN(n6205) );
  OR2_X1 U7835 ( .A1(n8110), .A2(n7743), .ZN(n6206) );
  AOI21_X2 U7836 ( .B1(n6207), .B2(n4875), .A(n4874), .ZN(n8094) );
  INV_X1 U7837 ( .A(n8076), .ZN(n7329) );
  OR2_X1 U7838 ( .A1(n8186), .A2(n7329), .ZN(n7459) );
  NAND2_X1 U7839 ( .A1(n8186), .A2(n7329), .ZN(n7456) );
  NAND2_X1 U7840 ( .A1(n7459), .A2(n7456), .ZN(n8093) );
  NAND2_X1 U7841 ( .A1(n8094), .A2(n8093), .ZN(n8069) );
  INV_X1 U7842 ( .A(n8098), .ZN(n7668) );
  NAND2_X1 U7843 ( .A1(n8179), .A2(n7668), .ZN(n7462) );
  NAND2_X1 U7844 ( .A1(n7458), .A2(n7462), .ZN(n8071) );
  OR2_X1 U7845 ( .A1(n8186), .A2(n8076), .ZN(n8070) );
  AND2_X1 U7846 ( .A1(n8071), .A2(n8070), .ZN(n6208) );
  NAND2_X1 U7847 ( .A1(n8069), .A2(n6208), .ZN(n8074) );
  NAND2_X1 U7848 ( .A1(n8179), .A2(n8098), .ZN(n6209) );
  NAND2_X1 U7849 ( .A1(n8074), .A2(n6209), .ZN(n8060) );
  NAND2_X1 U7850 ( .A1(n8261), .A2(n7338), .ZN(n7461) );
  NAND2_X1 U7851 ( .A1(n7471), .A2(n7461), .ZN(n8058) );
  NAND2_X1 U7852 ( .A1(n8060), .A2(n8058), .ZN(n6211) );
  NAND2_X1 U7853 ( .A1(n8261), .A2(n8077), .ZN(n6210) );
  NAND2_X1 U7854 ( .A1(n6211), .A2(n6210), .ZN(n8051) );
  AND2_X1 U7855 ( .A1(n8255), .A2(n8062), .ZN(n6213) );
  OR2_X1 U7856 ( .A1(n8255), .A2(n8062), .ZN(n6212) );
  INV_X1 U7857 ( .A(n8052), .ZN(n7717) );
  NAND2_X1 U7858 ( .A1(n8249), .A2(n7717), .ZN(n7477) );
  OR2_X1 U7859 ( .A1(n7686), .A2(n8042), .ZN(n7486) );
  NAND2_X1 U7860 ( .A1(n7686), .A2(n8042), .ZN(n7480) );
  NAND2_X1 U7861 ( .A1(n7486), .A2(n7480), .ZN(n8025) );
  NAND2_X1 U7862 ( .A1(n8163), .A2(n8004), .ZN(n7492) );
  NAND2_X1 U7863 ( .A1(n7487), .A2(n7492), .ZN(n8017) );
  INV_X1 U7864 ( .A(n8163), .ZN(n7639) );
  XNOR2_X1 U7865 ( .A(n8159), .B(n7741), .ZN(n8005) );
  NOR2_X1 U7866 ( .A1(n7997), .A2(n7980), .ZN(n6214) );
  INV_X1 U7867 ( .A(n7997), .ZN(n8231) );
  INV_X1 U7868 ( .A(n8226), .ZN(n7685) );
  NOR2_X1 U7869 ( .A1(n8219), .A2(n7963), .ZN(n6215) );
  INV_X1 U7870 ( .A(n8219), .ZN(n7738) );
  INV_X1 U7871 ( .A(n8213), .ZN(n6216) );
  NOR2_X1 U7872 ( .A1(n6216), .A2(n7732), .ZN(n6217) );
  OAI22_X2 U7873 ( .A1(n7945), .A2(n6217), .B1(n7956), .B2(n8213), .ZN(n7936)
         );
  NAND2_X1 U7874 ( .A1(n7600), .A2(n7542), .ZN(n6219) );
  OR2_X1 U7875 ( .A1(n7543), .A2(n8295), .ZN(n6218) );
  NAND2_X2 U7876 ( .A1(n6219), .A2(n6218), .ZN(n8207) );
  NOR2_X1 U7877 ( .A1(n8207), .A2(n7946), .ZN(n6220) );
  INV_X1 U7878 ( .A(n8207), .ZN(n7528) );
  INV_X1 U7879 ( .A(SI_28_), .ZN(n6223) );
  NAND2_X1 U7880 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  INV_X1 U7881 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6226) );
  INV_X1 U7882 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9307) );
  MUX2_X1 U7883 ( .A(n6226), .B(n9307), .S(n8613), .Z(n7362) );
  NAND2_X1 U7884 ( .A1(n8602), .A2(n7542), .ZN(n6228) );
  OR2_X1 U7885 ( .A1(n7543), .A2(n6226), .ZN(n6227) );
  NAND2_X1 U7886 ( .A1(n7926), .A2(n6229), .ZN(n6597) );
  INV_X1 U7887 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U7888 ( .A1(n5775), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7889 ( .A1(n6230), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6231) );
  OAI211_X1 U7890 ( .C1(n5744), .C2(n9893), .A(n6232), .B(n6231), .ZN(n6233)
         );
  INV_X1 U7891 ( .A(n6233), .ZN(n6234) );
  OR2_X2 U7892 ( .A1(n6286), .A2(n7740), .ZN(n7582) );
  NAND2_X1 U7893 ( .A1(n6286), .A2(n7740), .ZN(n7532) );
  XNOR2_X1 U7894 ( .A(n6235), .B(n4438), .ZN(n6239) );
  NAND2_X1 U7895 ( .A1(n7389), .A2(n6270), .ZN(n6236) );
  INV_X1 U7896 ( .A(n8123), .ZN(n6238) );
  NAND2_X1 U7897 ( .A1(n6239), .A2(n6238), .ZN(n6269) );
  INV_X1 U7898 ( .A(n7386), .ZN(n6724) );
  NAND2_X1 U7899 ( .A1(n6724), .A2(n6726), .ZN(n6725) );
  NAND2_X1 U7900 ( .A1(n6725), .A2(n7390), .ZN(n8116) );
  AND2_X1 U7901 ( .A1(n7394), .A2(n7395), .ZN(n8122) );
  NAND2_X1 U7902 ( .A1(n8116), .A2(n8122), .ZN(n8117) );
  NAND2_X1 U7903 ( .A1(n8117), .A2(n7394), .ZN(n6959) );
  OR2_X1 U7904 ( .A1(n8119), .A2(n6240), .ZN(n7401) );
  NAND2_X1 U7905 ( .A1(n8119), .A2(n6240), .ZN(n7407) );
  AND2_X1 U7906 ( .A1(n7401), .A2(n7407), .ZN(n6957) );
  NAND2_X1 U7907 ( .A1(n6959), .A2(n6957), .ZN(n6241) );
  NAND2_X1 U7908 ( .A1(n6241), .A2(n7407), .ZN(n6948) );
  NAND2_X1 U7909 ( .A1(n6948), .A2(n7560), .ZN(n6242) );
  NAND2_X1 U7910 ( .A1(n6242), .A2(n7402), .ZN(n6967) );
  NAND2_X1 U7911 ( .A1(n6967), .A2(n7409), .ZN(n6243) );
  INV_X1 U7912 ( .A(n7413), .ZN(n7404) );
  OR2_X1 U7913 ( .A1(n7090), .A2(n6244), .ZN(n6873) );
  NAND2_X1 U7914 ( .A1(n7090), .A2(n6244), .ZN(n7428) );
  INV_X1 U7915 ( .A(n6245), .ZN(n9814) );
  NAND2_X1 U7916 ( .A1(n9814), .A2(n7748), .ZN(n7420) );
  AND2_X1 U7917 ( .A1(n6873), .A2(n7420), .ZN(n7427) );
  NAND2_X1 U7918 ( .A1(n6937), .A2(n6245), .ZN(n7429) );
  NAND2_X1 U7919 ( .A1(n6246), .A2(n7429), .ZN(n6935) );
  OR2_X1 U7920 ( .A1(n9819), .A2(n7747), .ZN(n7430) );
  NAND2_X1 U7921 ( .A1(n9819), .A2(n7747), .ZN(n7426) );
  NAND2_X1 U7922 ( .A1(n7430), .A2(n7426), .ZN(n7568) );
  NOR2_X1 U7923 ( .A1(n7294), .A2(n7345), .ZN(n7425) );
  NAND2_X1 U7924 ( .A1(n7294), .A2(n7345), .ZN(n7431) );
  AND2_X1 U7925 ( .A1(n7441), .A2(n7431), .ZN(n7436) );
  INV_X1 U7926 ( .A(n7744), .ZN(n6247) );
  OR2_X1 U7927 ( .A1(n7653), .A2(n6247), .ZN(n7443) );
  NAND2_X1 U7928 ( .A1(n7653), .A2(n6247), .ZN(n7444) );
  NAND2_X1 U7929 ( .A1(n7209), .A2(n7574), .ZN(n6248) );
  NAND2_X1 U7930 ( .A1(n6248), .A2(n7443), .ZN(n7260) );
  NAND2_X1 U7931 ( .A1(n8110), .A2(n7644), .ZN(n7447) );
  NAND2_X1 U7932 ( .A1(n7260), .A2(n7447), .ZN(n6249) );
  OR2_X1 U7933 ( .A1(n8110), .A2(n7644), .ZN(n7448) );
  NAND2_X1 U7934 ( .A1(n6249), .A2(n7448), .ZN(n7284) );
  NOR2_X1 U7935 ( .A1(n8279), .A2(n7317), .ZN(n7451) );
  NAND2_X1 U7936 ( .A1(n8279), .A2(n7317), .ZN(n7281) );
  INV_X1 U7937 ( .A(n7456), .ZN(n6250) );
  INV_X1 U7938 ( .A(n7461), .ZN(n6251) );
  OAI21_X2 U7939 ( .B1(n8059), .B2(n6251), .A(n7471), .ZN(n8050) );
  NOR2_X1 U7940 ( .A1(n8255), .A2(n8041), .ZN(n7559) );
  NAND2_X1 U7941 ( .A1(n8255), .A2(n8041), .ZN(n7557) );
  INV_X1 U7942 ( .A(n7492), .ZN(n6252) );
  NAND2_X1 U7943 ( .A1(n8006), .A2(n8005), .ZN(n8008) );
  INV_X1 U7944 ( .A(n7741), .ZN(n8016) );
  OR2_X1 U7945 ( .A1(n8159), .A2(n8016), .ZN(n7494) );
  NAND2_X1 U7946 ( .A1(n8008), .A2(n7494), .ZN(n7989) );
  INV_X1 U7947 ( .A(n7989), .ZN(n6254) );
  NOR2_X1 U7948 ( .A1(n7997), .A2(n8003), .ZN(n7556) );
  INV_X1 U7949 ( .A(n7556), .ZN(n6253) );
  NAND2_X1 U7950 ( .A1(n6254), .A2(n6253), .ZN(n6255) );
  NAND2_X1 U7951 ( .A1(n7997), .A2(n8003), .ZN(n7500) );
  NAND2_X1 U7952 ( .A1(n7971), .A2(n7972), .ZN(n8148) );
  OR2_X1 U7953 ( .A1(n7655), .A2(n7509), .ZN(n7510) );
  NOR2_X1 U7954 ( .A1(n8219), .A2(n6110), .ZN(n7515) );
  NAND2_X1 U7955 ( .A1(n8219), .A2(n6110), .ZN(n7512) );
  OR2_X1 U7956 ( .A1(n8213), .A2(n7732), .ZN(n7521) );
  OR2_X1 U7957 ( .A1(n8207), .A2(n7524), .ZN(n6256) );
  AOI21_X1 U7958 ( .B1(n6258), .B2(n7102), .A(n7896), .ZN(n6271) );
  INV_X1 U7959 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6262) );
  INV_X1 U7960 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6259) );
  OR2_X1 U7961 ( .A1(n6589), .A2(n6259), .ZN(n6261) );
  INV_X1 U7962 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9374) );
  OR2_X1 U7963 ( .A1(n5744), .A2(n9374), .ZN(n6260) );
  OAI211_X1 U7964 ( .C1(n6594), .C2(n6262), .A(n6261), .B(n6260), .ZN(n6263)
         );
  INV_X1 U7965 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7966 ( .A1(n6597), .A2(n6264), .ZN(n7739) );
  AND2_X1 U7967 ( .A1(n6378), .A2(P2_B_REG_SCAN_IN), .ZN(n6265) );
  NOR2_X1 U7968 ( .A1(n8118), .A2(n6265), .ZN(n7376) );
  INV_X1 U7969 ( .A(n6266), .ZN(n6267) );
  AOI22_X1 U7970 ( .A1(n7739), .A2(n7376), .B1(n7946), .B2(n8096), .ZN(n6268)
         );
  NAND2_X1 U7971 ( .A1(n6271), .A2(n6270), .ZN(n6272) );
  NAND2_X1 U7972 ( .A1(n6272), .A2(n7535), .ZN(n6274) );
  OR2_X1 U7973 ( .A1(n6273), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7974 ( .A1(n6115), .A2(n6274), .ZN(n6275) );
  INV_X1 U7975 ( .A(n6277), .ZN(n6279) );
  INV_X1 U7976 ( .A(n6281), .ZN(n6282) );
  INV_X1 U7977 ( .A(n6286), .ZN(n7928) );
  NAND2_X1 U7978 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  NAND2_X1 U7979 ( .A1(n6290), .A2(n6289), .ZN(n6294) );
  NAND2_X1 U7980 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X1 U7981 ( .A1(n6296), .A2(n4868), .ZN(P2_U3456) );
  INV_X1 U7982 ( .A(n6297), .ZN(n6298) );
  INV_X1 U7983 ( .A(n6301), .ZN(n7220) );
  NAND2_X1 U7984 ( .A1(n6301), .A2(n7519), .ZN(n6302) );
  NAND2_X1 U7985 ( .A1(n6399), .A2(n6302), .ZN(n6377) );
  OR2_X1 U7986 ( .A1(n6377), .A2(n6303), .ZN(n6304) );
  NAND2_X1 U7987 ( .A1(n6304), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U7988 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U7989 ( .A(n6305), .B(n6581), .S(P2_STATE_REG_SCAN_IN), .Z(n6306) );
  INV_X1 U7990 ( .A(n6306), .ZN(P2_U3295) );
  INV_X2 U7991 ( .A(n7215), .ZN(n7231) );
  OAI222_X1 U7992 ( .A1(n9308), .A2(n6308), .B1(n7231), .B2(n6321), .C1(
        P1_U3086), .C2(n6307), .ZN(P1_U3352) );
  NAND2_X1 U7993 ( .A1(n8613), .A2(P2_U3151), .ZN(n8294) );
  OAI222_X1 U7994 ( .A1(n8294), .A2(n6309), .B1(n8304), .B2(n6315), .C1(
        P2_U3151), .C2(n6411), .ZN(P2_U3293) );
  OAI222_X1 U7995 ( .A1(n9308), .A2(n6310), .B1(n7231), .B2(n6311), .C1(
        P1_U3086), .C2(n9398), .ZN(P1_U3351) );
  OAI222_X1 U7996 ( .A1(n8294), .A2(n6312), .B1(n8304), .B2(n6311), .C1(
        P2_U3151), .C2(n6427), .ZN(P2_U3291) );
  INV_X1 U7997 ( .A(n4300), .ZN(n6313) );
  OAI222_X1 U7998 ( .A1(n9308), .A2(n6314), .B1(n7231), .B2(n6317), .C1(
        P1_U3086), .C2(n6313), .ZN(P1_U3354) );
  INV_X1 U7999 ( .A(n6646), .ZN(n6316) );
  OAI222_X1 U8000 ( .A1(P1_U3086), .A2(n6316), .B1(n7231), .B2(n6315), .C1(
        n9308), .C2(n4968), .ZN(P1_U3353) );
  INV_X1 U8001 ( .A(n8304), .ZN(n7218) );
  OAI222_X1 U8002 ( .A1(n8294), .A2(n4783), .B1(n8304), .B2(n6317), .C1(
        P2_U3151), .C2(n4397), .ZN(P2_U3294) );
  OAI222_X1 U8003 ( .A1(n8294), .A2(n6318), .B1(n8304), .B2(n6319), .C1(
        P2_U3151), .C2(n6605), .ZN(P2_U3290) );
  OAI222_X1 U8004 ( .A1(n9308), .A2(n6320), .B1(n7231), .B2(n6319), .C1(
        P1_U3086), .C2(n9414), .ZN(P1_U3350) );
  INV_X1 U8005 ( .A(n8294), .ZN(n6478) );
  OAI222_X1 U8006 ( .A1(n8300), .A2(n6322), .B1(n8304), .B2(n6321), .C1(
        P2_U3151), .C2(n6494), .ZN(P2_U3292) );
  OAI222_X1 U8007 ( .A1(n9308), .A2(n6323), .B1(n7231), .B2(n6324), .C1(
        P1_U3086), .C2(n9429), .ZN(P1_U3349) );
  OAI222_X1 U8008 ( .A1(n8294), .A2(n6325), .B1(n8304), .B2(n6324), .C1(
        P2_U3151), .C2(n6459), .ZN(P2_U3289) );
  OAI222_X1 U8009 ( .A1(n8294), .A2(n6326), .B1(n8304), .B2(n6327), .C1(
        P2_U3151), .C2(n6852), .ZN(P2_U3288) );
  OAI222_X1 U8010 ( .A1(n9308), .A2(n6328), .B1(n7231), .B2(n6327), .C1(
        P1_U3086), .C2(n9335), .ZN(P1_U3348) );
  OAI222_X1 U8011 ( .A1(n8294), .A2(n6329), .B1(n8304), .B2(n6330), .C1(
        P2_U3151), .C2(n6854), .ZN(P2_U3287) );
  OAI222_X1 U8012 ( .A1(n9308), .A2(n6331), .B1(n7231), .B2(n6330), .C1(
        P1_U3086), .C2(n9364), .ZN(P1_U3347) );
  INV_X1 U8013 ( .A(n6332), .ZN(n6335) );
  OAI222_X1 U8014 ( .A1(n8304), .A2(n6335), .B1(n6855), .B2(P2_U3151), .C1(
        n6333), .C2(n8300), .ZN(P2_U3286) );
  INV_X1 U8015 ( .A(n8813), .ZN(n6334) );
  OAI222_X1 U8016 ( .A1(n9308), .A2(n6336), .B1(n7231), .B2(n6335), .C1(n6334), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U8017 ( .A1(n9618), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U8018 ( .B1(n9618), .B2(n6339), .A(n6338), .ZN(P1_U3439) );
  INV_X1 U8019 ( .A(n6340), .ZN(n6343) );
  INV_X1 U8020 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6341) );
  OAI222_X1 U8021 ( .A1(n8304), .A2(n6343), .B1(n7134), .B2(P2_U3151), .C1(
        n6341), .C2(n8300), .ZN(P2_U3285) );
  INV_X1 U8022 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U8023 ( .A1(n6356), .A2(n9917), .ZN(P2_U3261) );
  INV_X1 U8024 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U8025 ( .A1(n6356), .A2(n9956), .ZN(P2_U3239) );
  INV_X1 U8026 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9941) );
  NOR2_X1 U8027 ( .A1(n6356), .A2(n9941), .ZN(P2_U3249) );
  INV_X1 U8028 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U8029 ( .A1(n6356), .A2(n9890), .ZN(P2_U3237) );
  INV_X1 U8030 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6344) );
  OAI222_X1 U8031 ( .A1(n9308), .A2(n6344), .B1(n7231), .B2(n6343), .C1(n6342), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8032 ( .A(n6345), .ZN(n6348) );
  AOI22_X1 U8033 ( .A1(n7171), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6478), .ZN(n6346) );
  OAI21_X1 U8034 ( .B1(n6348), .B2(n8304), .A(n6346), .ZN(P2_U3284) );
  AND2_X1 U8035 ( .A1(n6347), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8036 ( .A1(n6347), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8037 ( .A1(n6347), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8038 ( .A1(n6347), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8039 ( .A1(n6347), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8040 ( .A1(n6347), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8041 ( .A1(n6347), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8042 ( .A1(n6347), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8043 ( .A1(n6347), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  INV_X1 U8044 ( .A(n6565), .ZN(n9444) );
  OAI222_X1 U8045 ( .A1(n9308), .A2(n6349), .B1(n7231), .B2(n6348), .C1(
        P1_U3086), .C2(n9444), .ZN(P1_U3344) );
  NAND2_X1 U8046 ( .A1(P2_U3893), .A2(n6181), .ZN(n6350) );
  OAI21_X1 U8047 ( .B1(P2_U3893), .B2(n4968), .A(n6350), .ZN(P2_U3493) );
  INV_X1 U8048 ( .A(n6351), .ZN(n6361) );
  OAI222_X1 U8049 ( .A1(n8304), .A2(n6361), .B1(n7763), .B2(P2_U3151), .C1(
        n6352), .C2(n8300), .ZN(P2_U3283) );
  INV_X1 U8050 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8051 ( .A1(P2_U3893), .A2(n6353), .ZN(n6354) );
  OAI21_X1 U8052 ( .B1(P2_U3893), .B2(n6355), .A(n6354), .ZN(P2_U3491) );
  INV_X1 U8053 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6360) );
  INV_X1 U8054 ( .A(n6357), .ZN(n6358) );
  AOI22_X1 U8055 ( .A1(n6347), .A2(n6360), .B1(n6359), .B2(n6358), .ZN(
        P2_U3376) );
  INV_X1 U8056 ( .A(n8831), .ZN(n6569) );
  OAI222_X1 U8057 ( .A1(n9308), .A2(n6362), .B1(n7231), .B2(n6361), .C1(n6569), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  AND2_X1 U8058 ( .A1(n6347), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8059 ( .A1(n6347), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8060 ( .A1(n6347), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8061 ( .A1(n6347), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8062 ( .A1(n6347), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8063 ( .A1(n6347), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8064 ( .A1(n6347), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8065 ( .A1(n6347), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8066 ( .A1(n6347), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8067 ( .A1(n6347), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8068 ( .A1(n6347), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8069 ( .A1(n6347), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8070 ( .A1(n6347), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8071 ( .A1(n6347), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8072 ( .A1(n6347), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8073 ( .A1(n6347), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8074 ( .A1(n6347), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  NAND2_X1 U8075 ( .A1(n8697), .A2(n6363), .ZN(n6364) );
  AND2_X1 U8076 ( .A1(n8615), .A2(n6364), .ZN(n6538) );
  INV_X1 U8077 ( .A(n6538), .ZN(n6365) );
  NAND2_X1 U8078 ( .A1(n8514), .A2(n8770), .ZN(n6539) );
  AND2_X1 U8079 ( .A1(n6365), .A2(n6539), .ZN(n9400) );
  NOR2_X1 U8080 ( .A1(n9400), .A2(n8792), .ZN(P1_U3085) );
  INV_X1 U8081 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8082 ( .A1(n8926), .A2(P1_U3973), .ZN(n6366) );
  OAI21_X1 U8083 ( .B1(n6883), .B2(n8792), .A(n6366), .ZN(P1_U3573) );
  INV_X1 U8084 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U8085 ( .A1(n8922), .A2(P1_U3973), .ZN(n6367) );
  OAI21_X1 U8086 ( .B1(n6762), .B2(n8792), .A(n6367), .ZN(P1_U3572) );
  INV_X1 U8087 ( .A(n6368), .ZN(n6371) );
  AOI22_X1 U8088 ( .A1(n7789), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6478), .ZN(n6369) );
  OAI21_X1 U8089 ( .B1(n6371), .B2(n8304), .A(n6369), .ZN(P2_U3282) );
  AOI22_X1 U8090 ( .A1(n9457), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9300), .ZN(n6370) );
  OAI21_X1 U8091 ( .B1(n6371), .B2(n7231), .A(n6370), .ZN(P1_U3342) );
  NAND2_X1 U8092 ( .A1(n8921), .A2(n8792), .ZN(n6372) );
  OAI21_X1 U8093 ( .B1(n5341), .B2(n8792), .A(n6372), .ZN(P1_U3571) );
  XNOR2_X1 U8094 ( .A(n6374), .B(n6373), .ZN(n6636) );
  AND2_X1 U8095 ( .A1(n6774), .A2(n8878), .ZN(n6744) );
  AOI22_X1 U8096 ( .A1(n4295), .A2(n6756), .B1(n8506), .B2(n6744), .ZN(n6376)
         );
  NOR2_X1 U8097 ( .A1(n8475), .A2(P1_U3086), .ZN(n6635) );
  INV_X1 U8098 ( .A(n6635), .ZN(n6623) );
  NAND2_X1 U8099 ( .A1(n6623), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U8100 ( .C1(n6636), .C2(n8511), .A(n6376), .B(n6375), .ZN(P1_U3232) );
  NOR2_X1 U8101 ( .A1(n6377), .A2(P2_U3151), .ZN(n6387) );
  MUX2_X1 U8102 ( .A(P2_U3893), .B(n6387), .S(n6154), .Z(n6379) );
  NAND2_X1 U8103 ( .A1(n6379), .A2(n6378), .ZN(n7917) );
  INV_X1 U8104 ( .A(n6380), .ZN(n6410) );
  OAI21_X1 U8105 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6406), .A(n6410), .ZN(n6381) );
  NAND2_X1 U8106 ( .A1(n5736), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6382) );
  INV_X1 U8107 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6499) );
  AOI21_X1 U8108 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6411), .A(n9739), .ZN(
        n6383) );
  INV_X1 U8109 ( .A(n6386), .ZN(n6384) );
  MUX2_X1 U8110 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6421), .S(n6427), .Z(n6385)
         );
  OR3_X1 U8111 ( .A1(n6386), .A2(n6385), .A3(n4390), .ZN(n6389) );
  INV_X1 U8112 ( .A(n6387), .ZN(n6388) );
  OR2_X1 U8113 ( .A1(n6388), .A2(n6154), .ZN(n6583) );
  AOI21_X1 U8114 ( .B1(n6422), .B2(n6389), .A(n9762), .ZN(n6404) );
  AND2_X1 U8115 ( .A1(n6581), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8116 ( .A1(n5736), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6391) );
  OAI21_X1 U8117 ( .B1(n6380), .B2(n6390), .A(n6391), .ZN(n6502) );
  NAND2_X1 U8118 ( .A1(n6500), .A2(n6391), .ZN(n9743) );
  INV_X1 U8119 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U8120 ( .A1(n6411), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8121 ( .A1(n9742), .A2(n6392), .ZN(n6393) );
  NAND2_X1 U8122 ( .A1(n6393), .A2(n6494), .ZN(n6396) );
  INV_X1 U8123 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9834) );
  MUX2_X1 U8124 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9834), .S(n6427), .Z(n6395)
         );
  INV_X1 U8125 ( .A(n6395), .ZN(n6397) );
  NAND3_X1 U8126 ( .A1(n6486), .A2(n6397), .A3(n6396), .ZN(n6398) );
  AOI21_X1 U8127 ( .B1(n6429), .B2(n6398), .A(n9769), .ZN(n6403) );
  INV_X1 U8128 ( .A(n6399), .ZN(n6400) );
  INV_X1 U8129 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8130 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6806) );
  OAI21_X1 U8131 ( .B1(n9779), .B2(n6401), .A(n6806), .ZN(n6402) );
  NOR3_X1 U8132 ( .A1(n6404), .A2(n6403), .A3(n6402), .ZN(n6420) );
  MUX2_X1 U8133 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6155), .Z(n6408) );
  XNOR2_X1 U8134 ( .A(n6408), .B(n4397), .ZN(n6495) );
  MUX2_X1 U8135 ( .A(n6406), .B(n6405), .S(n6156), .Z(n6407) );
  AND2_X1 U8136 ( .A1(n6407), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6579) );
  INV_X1 U8137 ( .A(n6408), .ZN(n6409) );
  MUX2_X1 U8138 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6156), .Z(n6412) );
  INV_X1 U8139 ( .A(n6411), .ZN(n9750) );
  XNOR2_X1 U8140 ( .A(n6412), .B(n9750), .ZN(n9752) );
  MUX2_X1 U8141 ( .A(n6414), .B(n6413), .S(n6156), .Z(n6415) );
  XNOR2_X1 U8142 ( .A(n6415), .B(n6494), .ZN(n6481) );
  NAND2_X1 U8143 ( .A1(n6482), .A2(n6481), .ZN(n6480) );
  NAND2_X1 U8144 ( .A1(n6415), .A2(n4699), .ZN(n6416) );
  AND2_X1 U8145 ( .A1(n6480), .A2(n6416), .ZN(n6418) );
  MUX2_X1 U8146 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6156), .Z(n6439) );
  INV_X1 U8147 ( .A(n6427), .ZN(n6442) );
  XNOR2_X1 U8148 ( .A(n6439), .B(n6442), .ZN(n6417) );
  NAND2_X1 U8149 ( .A1(P2_U3893), .A2(n6154), .ZN(n7913) );
  OAI211_X1 U8150 ( .C1(n6418), .C2(n6417), .A(n9774), .B(n6440), .ZN(n6419)
         );
  OAI211_X1 U8151 ( .C1(n7917), .C2(n6427), .A(n6420), .B(n6419), .ZN(P2_U3186) );
  OAI21_X1 U8152 ( .B1(n6423), .B2(n6605), .A(n6424), .ZN(n6608) );
  XNOR2_X1 U8153 ( .A(n6459), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6425) );
  NAND3_X1 U8154 ( .A1(n6609), .A2(n6425), .A3(n6424), .ZN(n6426) );
  AOI21_X1 U8155 ( .B1(n4389), .B2(n6426), .A(n9762), .ZN(n6438) );
  NAND2_X1 U8156 ( .A1(n6427), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8157 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  INV_X1 U8158 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6432) );
  NAND3_X1 U8159 ( .A1(n6606), .A2(n4391), .A3(n6433), .ZN(n6434) );
  AOI21_X1 U8160 ( .B1(n6460), .B2(n6434), .A(n9769), .ZN(n6437) );
  INV_X1 U8161 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U8162 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9927), .ZN(n6931) );
  INV_X1 U8163 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U8164 ( .A1(n9779), .A2(n6435), .ZN(n6436) );
  NOR4_X1 U8165 ( .A1(n6438), .A2(n6437), .A3(n6931), .A4(n6436), .ZN(n6451)
         );
  INV_X1 U8166 ( .A(n6439), .ZN(n6441) );
  MUX2_X1 U8167 ( .A(n6443), .B(n4559), .S(n6156), .Z(n6444) );
  XNOR2_X1 U8168 ( .A(n6444), .B(n6605), .ZN(n6603) );
  INV_X1 U8169 ( .A(n6444), .ZN(n6445) );
  MUX2_X1 U8170 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6156), .Z(n6446) );
  NOR2_X1 U8171 ( .A1(n6446), .A2(n6459), .ZN(n6467) );
  AOI21_X1 U8172 ( .B1(n6446), .B2(n6459), .A(n6467), .ZN(n6447) );
  NAND2_X1 U8173 ( .A1(n6448), .A2(n6447), .ZN(n6469) );
  OAI21_X1 U8174 ( .B1(n6448), .B2(n6447), .A(n6469), .ZN(n6449) );
  NAND2_X1 U8175 ( .A1(n6449), .A2(n9774), .ZN(n6450) );
  OAI211_X1 U8176 ( .C1(n7917), .C2(n6459), .A(n6451), .B(n6450), .ZN(P2_U3188) );
  INV_X1 U8177 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6453) );
  INV_X1 U8178 ( .A(n6452), .ZN(n6454) );
  OAI222_X1 U8179 ( .A1(n9308), .A2(n6453), .B1(n7231), .B2(n6454), .C1(
        P1_U3086), .C2(n9471), .ZN(P1_U3341) );
  INV_X1 U8180 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6455) );
  OAI222_X1 U8181 ( .A1(n8294), .A2(n6455), .B1(n8304), .B2(n6454), .C1(
        P2_U3151), .C2(n7805), .ZN(P2_U3281) );
  INV_X1 U8182 ( .A(n6457), .ZN(n6458) );
  OAI21_X1 U8183 ( .B1(n6458), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6833), .ZN(
        n6466) );
  AOI21_X1 U8184 ( .B1(n6470), .B2(n6461), .A(n6850), .ZN(n6462) );
  NOR2_X1 U8185 ( .A1(n9769), .A2(n6462), .ZN(n6465) );
  INV_X1 U8186 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8187 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6988) );
  OAI21_X1 U8188 ( .B1(n9779), .B2(n6463), .A(n6988), .ZN(n6464) );
  AOI211_X1 U8189 ( .C1(n6466), .C2(n7920), .A(n6465), .B(n6464), .ZN(n6476)
         );
  INV_X1 U8190 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U8191 ( .A1(n6469), .A2(n6468), .ZN(n6473) );
  MUX2_X1 U8192 ( .A(n6471), .B(n6470), .S(n6156), .Z(n6840) );
  XNOR2_X1 U8193 ( .A(n6840), .B(n6852), .ZN(n6472) );
  OAI21_X1 U8194 ( .B1(n6473), .B2(n6472), .A(n6841), .ZN(n6474) );
  NAND2_X1 U8195 ( .A1(n6474), .A2(n9774), .ZN(n6475) );
  OAI211_X1 U8196 ( .C1(n7917), .C2(n6852), .A(n6476), .B(n6475), .ZN(P2_U3189) );
  INV_X1 U8197 ( .A(n6477), .ZN(n6599) );
  AOI22_X1 U8198 ( .A1(n7835), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n6478), .ZN(n6479) );
  OAI21_X1 U8199 ( .B1(n6599), .B2(n8304), .A(n6479), .ZN(P2_U3280) );
  OAI21_X1 U8200 ( .B1(n6482), .B2(n6481), .A(n6480), .ZN(n6492) );
  INV_X1 U8201 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6484) );
  INV_X1 U8202 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6483) );
  OAI22_X1 U8203 ( .A1(n9779), .A2(n6484), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6483), .ZN(n6491) );
  AOI21_X1 U8204 ( .B1(n6414), .B2(n6485), .A(n4390), .ZN(n6489) );
  INV_X1 U8205 ( .A(n6486), .ZN(n6487) );
  AOI21_X1 U8206 ( .B1(n6413), .B2(n4564), .A(n6487), .ZN(n6488) );
  OAI22_X1 U8207 ( .A1(n9762), .A2(n6489), .B1(n6488), .B2(n9769), .ZN(n6490)
         );
  AOI211_X1 U8208 ( .C1(n9774), .C2(n6492), .A(n6491), .B(n6490), .ZN(n6493)
         );
  OAI21_X1 U8209 ( .B1(n6494), .B2(n7917), .A(n6493), .ZN(P2_U3185) );
  XNOR2_X1 U8210 ( .A(n6495), .B(n6579), .ZN(n6496) );
  INV_X1 U8211 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6727) );
  OAI22_X1 U8212 ( .A1(n7913), .A2(n6496), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6727), .ZN(n6506) );
  AOI21_X1 U8213 ( .B1(n6499), .B2(n6498), .A(n6497), .ZN(n6504) );
  INV_X1 U8214 ( .A(n6500), .ZN(n6501) );
  AOI21_X1 U8215 ( .B1(n5740), .B2(n6502), .A(n6501), .ZN(n6503) );
  OAI22_X1 U8216 ( .A1(n9762), .A2(n6504), .B1(n6503), .B2(n9769), .ZN(n6505)
         );
  AOI211_X1 U8217 ( .C1(n7915), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6506), .B(
        n6505), .ZN(n6507) );
  OAI21_X1 U8218 ( .B1(n4397), .B2(n7917), .A(n6507), .ZN(P2_U3183) );
  NAND2_X1 U8219 ( .A1(n8769), .A2(n9535), .ZN(n8630) );
  NAND2_X1 U8220 ( .A1(n8708), .A2(n8756), .ZN(n8768) );
  OR2_X1 U8221 ( .A1(n6509), .A2(n6749), .ZN(n8513) );
  NAND2_X1 U8222 ( .A1(n8513), .A2(n6508), .ZN(n6742) );
  AND2_X1 U8223 ( .A1(n6509), .A2(n5626), .ZN(n6510) );
  OR2_X1 U8224 ( .A1(n6742), .A2(n6510), .ZN(n9508) );
  NAND2_X1 U8225 ( .A1(n7104), .A2(n9535), .ZN(n8766) );
  OR2_X1 U8226 ( .A1(n8766), .A2(n8756), .ZN(n9627) );
  INV_X1 U8227 ( .A(n9702), .ZN(n9625) );
  AND2_X1 U8228 ( .A1(n6751), .A2(n6755), .ZN(n8706) );
  NOR2_X1 U8229 ( .A1(n6780), .A2(n8706), .ZN(n8638) );
  AOI21_X1 U8230 ( .B1(n9596), .B2(n9625), .A(n8638), .ZN(n6511) );
  AOI211_X1 U8231 ( .C1(n6512), .C2(n6756), .A(n6744), .B(n6511), .ZN(n6576)
         );
  NAND2_X1 U8232 ( .A1(n6514), .A2(n6513), .ZN(n6516) );
  AND2_X1 U8233 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  NAND2_X1 U8234 ( .A1(n9735), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6520) );
  OAI21_X1 U8235 ( .B1(n6576), .B2(n9735), .A(n6520), .ZN(P1_U3522) );
  NOR2_X1 U8236 ( .A1(n8831), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6521) );
  AOI21_X1 U8237 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8831), .A(n6521), .ZN(
        n6537) );
  NAND2_X1 U8238 ( .A1(n9321), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U8239 ( .B1(n9321), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6522), .ZN(
        n9317) );
  NOR2_X1 U8240 ( .A1(n8813), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6523) );
  AOI21_X1 U8241 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n8813), .A(n6523), .ZN(
        n8806) );
  INV_X1 U8242 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6524) );
  MUX2_X1 U8243 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6524), .S(n6646), .Z(n6645)
         );
  INV_X1 U8244 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6525) );
  INV_X1 U8245 ( .A(n9384), .ZN(n6526) );
  INV_X1 U8246 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U8247 ( .A1(n6526), .A2(n6746), .ZN(n8797) );
  NAND2_X1 U8248 ( .A1(n4300), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8249 ( .A1(n8796), .A2(n6527), .ZN(n6644) );
  NAND2_X1 U8250 ( .A1(n6645), .A2(n6644), .ZN(n6643) );
  NAND2_X1 U8251 ( .A1(n6646), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8252 ( .A1(n6643), .A2(n6528), .ZN(n9340) );
  OAI21_X1 U8253 ( .B1(n9350), .B2(P1_REG2_REG_3__SCAN_IN), .A(n4505), .ZN(
        n9342) );
  INV_X1 U8254 ( .A(n9342), .ZN(n6529) );
  NAND2_X1 U8255 ( .A1(n6552), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U8256 ( .B1(n6552), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6530), .ZN(
        n9394) );
  NAND2_X1 U8257 ( .A1(n6555), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6531) );
  OAI21_X1 U8258 ( .B1(n6555), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6531), .ZN(
        n9410) );
  NOR2_X1 U8259 ( .A1(n4324), .A2(n9410), .ZN(n9409) );
  AOI21_X1 U8260 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6555), .A(n9409), .ZN(
        n9420) );
  INV_X1 U8261 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6532) );
  AOI22_X1 U8262 ( .A1(n6557), .A2(n6532), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9429), .ZN(n9421) );
  NOR2_X1 U8263 ( .A1(n9420), .A2(n9421), .ZN(n9419) );
  AOI21_X1 U8264 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6557), .A(n9419), .ZN(
        n9326) );
  NAND2_X1 U8265 ( .A1(n6560), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U8266 ( .B1(n6560), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6533), .ZN(
        n9327) );
  NOR2_X1 U8267 ( .A1(n9326), .A2(n9327), .ZN(n9325) );
  NAND2_X1 U8268 ( .A1(n6563), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6534) );
  OAI21_X1 U8269 ( .B1(n6563), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6534), .ZN(
        n9360) );
  OAI21_X1 U8270 ( .B1(n8813), .B2(P1_REG2_REG_9__SCAN_IN), .A(n8804), .ZN(
        n9318) );
  NAND2_X1 U8271 ( .A1(n6565), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6535) );
  OAI21_X1 U8272 ( .B1(n6565), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6535), .ZN(
        n9440) );
  NAND2_X1 U8273 ( .A1(n6537), .A2(n6536), .ZN(n8830) );
  OAI21_X1 U8274 ( .B1(n6537), .B2(n6536), .A(n8830), .ZN(n6542) );
  NAND2_X1 U8275 ( .A1(n6539), .A2(n6538), .ZN(n9386) );
  OR2_X1 U8276 ( .A1(n5640), .A2(n8880), .ZN(n6541) );
  NAND2_X1 U8277 ( .A1(n6542), .A2(n9497), .ZN(n6573) );
  NAND2_X1 U8278 ( .A1(n9321), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U8279 ( .B1(n9321), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6543), .ZN(
        n9314) );
  NOR2_X1 U8280 ( .A1(n8813), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6544) );
  AOI21_X1 U8281 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n8813), .A(n6544), .ZN(
        n8811) );
  INV_X1 U8282 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U8283 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9717), .S(n6646), .Z(n6642)
         );
  INV_X1 U8284 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U8285 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9715), .S(n8799), .Z(n8795)
         );
  AND2_X1 U8286 ( .A1(n9384), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U8287 ( .A1(n8795), .A2(n8794), .ZN(n8793) );
  NAND2_X1 U8288 ( .A1(n4300), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8289 ( .A1(n8793), .A2(n6545), .ZN(n6641) );
  NAND2_X1 U8290 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  NAND2_X1 U8291 ( .A1(n6646), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8292 ( .A1(n6640), .A2(n6546), .ZN(n9344) );
  NAND2_X1 U8293 ( .A1(n9350), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U8294 ( .B1(n9350), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6547), .ZN(
        n9346) );
  INV_X1 U8295 ( .A(n9346), .ZN(n6548) );
  AND2_X1 U8296 ( .A1(n9344), .A2(n6548), .ZN(n9345) );
  AND2_X1 U8297 ( .A1(n9350), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6549) );
  OR2_X1 U8298 ( .A1(n6552), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8299 ( .A1(n6552), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8300 ( .A1(n6551), .A2(n6550), .ZN(n9389) );
  NOR2_X1 U8301 ( .A1(n9390), .A2(n9389), .ZN(n9388) );
  AOI21_X1 U8302 ( .B1(n6552), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9388), .ZN(
        n9406) );
  OR2_X1 U8303 ( .A1(n6555), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8304 ( .A1(n6555), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U8305 ( .A1(n6554), .A2(n6553), .ZN(n9407) );
  NOR2_X1 U8306 ( .A1(n9406), .A2(n9407), .ZN(n9405) );
  INV_X1 U8307 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6556) );
  MUX2_X1 U8308 ( .A(n6556), .B(P1_REG1_REG_6__SCAN_IN), .S(n6557), .Z(n9425)
         );
  NOR2_X1 U8309 ( .A1(n9424), .A2(n9425), .ZN(n9423) );
  AOI21_X1 U8310 ( .B1(n6557), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9423), .ZN(
        n9330) );
  OR2_X1 U8311 ( .A1(n6560), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8312 ( .A1(n6560), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8313 ( .A1(n6559), .A2(n6558), .ZN(n9331) );
  NOR2_X1 U8314 ( .A1(n9330), .A2(n9331), .ZN(n9329) );
  OR2_X1 U8315 ( .A1(n6563), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8316 ( .A1(n6563), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8317 ( .A1(n6562), .A2(n6561), .ZN(n9356) );
  NOR2_X1 U8318 ( .A1(n9355), .A2(n9356), .ZN(n9354) );
  AOI21_X1 U8319 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6563), .A(n9354), .ZN(
        n8810) );
  NAND2_X1 U8320 ( .A1(n8811), .A2(n8810), .ZN(n8809) );
  OAI21_X1 U8321 ( .B1(n8813), .B2(P1_REG1_REG_9__SCAN_IN), .A(n8809), .ZN(
        n9315) );
  NOR2_X1 U8322 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  INV_X1 U8323 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U8324 ( .A(n6564), .B(P1_REG1_REG_11__SCAN_IN), .S(n6565), .Z(n9436)
         );
  NOR2_X1 U8325 ( .A1(n9435), .A2(n9436), .ZN(n9434) );
  AOI21_X1 U8326 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6565), .A(n9434), .ZN(
        n6567) );
  INV_X1 U8327 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9732) );
  AOI22_X1 U8328 ( .A1(n8831), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9732), .B2(
        n6569), .ZN(n6566) );
  NAND2_X1 U8329 ( .A1(n6567), .A2(n6566), .ZN(n8819) );
  OAI21_X1 U8330 ( .B1(n6567), .B2(n6566), .A(n8819), .ZN(n6571) );
  INV_X1 U8331 ( .A(n8880), .ZN(n9382) );
  NAND2_X1 U8332 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7270) );
  NAND2_X1 U8333 ( .A1(n9400), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6568) );
  OAI211_X1 U8334 ( .C1(n9501), .C2(n6569), .A(n7270), .B(n6568), .ZN(n6570)
         );
  AOI21_X1 U8335 ( .B1(n6571), .B2(n9489), .A(n6570), .ZN(n6572) );
  NAND2_X1 U8336 ( .A1(n6573), .A2(n6572), .ZN(P1_U3255) );
  INV_X1 U8337 ( .A(n6574), .ZN(n6740) );
  INV_X1 U8338 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6578) );
  OR2_X1 U8339 ( .A1(n6576), .A2(n9712), .ZN(n6577) );
  OAI21_X1 U8340 ( .B1(n9714), .B2(n6578), .A(n6577), .ZN(P1_U3453) );
  INV_X1 U8341 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6587) );
  MUX2_X1 U8342 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n6156), .Z(n6580) );
  AOI21_X1 U8343 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(n6582) );
  AOI21_X1 U8344 ( .B1(n6583), .B2(n7913), .A(n6582), .ZN(n6584) );
  AOI21_X1 U8345 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6584), .ZN(
        n6586) );
  NAND2_X1 U8346 ( .A1(n9767), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6585) );
  OAI211_X1 U8347 ( .C1(n9779), .C2(n6587), .A(n6586), .B(n6585), .ZN(P2_U3182) );
  INV_X1 U8348 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6593) );
  INV_X1 U8349 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6588) );
  OR2_X1 U8350 ( .A1(n6589), .A2(n6588), .ZN(n6592) );
  INV_X1 U8351 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6590) );
  OR2_X1 U8352 ( .A1(n5744), .A2(n6590), .ZN(n6591) );
  OAI211_X1 U8353 ( .C1(n6594), .C2(n6593), .A(n6592), .B(n6591), .ZN(n6595)
         );
  INV_X1 U8354 ( .A(n6595), .ZN(n6596) );
  NAND2_X1 U8355 ( .A1(n7878), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6598) );
  OAI21_X1 U8356 ( .B1(n7551), .B2(n7878), .A(n6598), .ZN(P2_U3522) );
  OAI222_X1 U8357 ( .A1(n9308), .A2(n6600), .B1(n7231), .B2(n6599), .C1(n8835), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8358 ( .A(n8606), .ZN(n6601) );
  NAND2_X1 U8359 ( .A1(n6601), .A2(n8792), .ZN(n6602) );
  OAI21_X1 U8360 ( .B1(n6226), .B2(n8792), .A(n6602), .ZN(P1_U3583) );
  XNOR2_X1 U8361 ( .A(n6604), .B(n6603), .ZN(n6618) );
  INV_X1 U8362 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6615) );
  INV_X1 U8363 ( .A(n9769), .ZN(n9746) );
  OAI21_X1 U8364 ( .B1(n6607), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6606), .ZN(
        n6612) );
  INV_X1 U8365 ( .A(n6608), .ZN(n6610) );
  OAI21_X1 U8366 ( .B1(n6610), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6609), .ZN(
        n6611) );
  AOI22_X1 U8367 ( .A1(n9746), .A2(n6612), .B1(n7920), .B2(n6611), .ZN(n6614)
         );
  AND2_X1 U8368 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6870) );
  INV_X1 U8369 ( .A(n6870), .ZN(n6613) );
  OAI211_X1 U8370 ( .C1(n6615), .C2(n9779), .A(n6614), .B(n6613), .ZN(n6616)
         );
  AOI21_X1 U8371 ( .B1(n4392), .B2(n9767), .A(n6616), .ZN(n6617) );
  OAI21_X1 U8372 ( .B1(n7913), .B2(n6618), .A(n6617), .ZN(P2_U3187) );
  AOI21_X1 U8373 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(n6625) );
  AOI22_X1 U8374 ( .A1(n8484), .A2(n6751), .B1(n8791), .B2(n8878), .ZN(n6752)
         );
  OAI22_X1 U8375 ( .A1(n6752), .A2(n8459), .B1(n8419), .B2(n8707), .ZN(n6622)
         );
  AOI21_X1 U8376 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6623), .A(n6622), .ZN(
        n6624) );
  OAI21_X1 U8377 ( .B1(n6625), .B2(n8511), .A(n6624), .ZN(P1_U3222) );
  NAND2_X1 U8378 ( .A1(n6353), .A2(n8196), .ZN(n7382) );
  NAND2_X1 U8379 ( .A1(n7388), .A2(n7382), .ZN(n8199) );
  INV_X1 U8380 ( .A(n8199), .ZN(n6711) );
  NAND2_X1 U8381 ( .A1(n7341), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8382 ( .A1(n6695), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U8383 ( .A1(n7705), .A2(n6730), .B1(n7680), .B2(n4851), .ZN(n6626)
         );
  OAI211_X1 U8384 ( .C1(n6711), .C2(n7707), .A(n6627), .B(n6626), .ZN(P2_U3172) );
  INV_X1 U8385 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9601) );
  INV_X1 U8386 ( .A(n6628), .ZN(n6632) );
  NOR3_X1 U8387 ( .A1(n6619), .A2(n6630), .A3(n6629), .ZN(n6631) );
  OAI21_X1 U8388 ( .B1(n6632), .B2(n6631), .A(n8495), .ZN(n6634) );
  INV_X1 U8389 ( .A(n6774), .ZN(n6782) );
  OAI22_X1 U8390 ( .A1(n6782), .A2(n8908), .B1(n6779), .B2(n8505), .ZN(n9599)
         );
  AOI22_X1 U8391 ( .A1(n9599), .A2(n8506), .B1(n6792), .B2(n4295), .ZN(n6633)
         );
  OAI211_X1 U8392 ( .C1(n6635), .C2(n9601), .A(n6634), .B(n6633), .ZN(P1_U3237) );
  AOI21_X1 U8393 ( .B1(n9382), .B2(n6746), .A(n5640), .ZN(n9381) );
  MUX2_X1 U8394 ( .A(n8797), .B(n6636), .S(n8880), .Z(n6638) );
  NAND2_X1 U8395 ( .A1(n6638), .A2(n6637), .ZN(n6639) );
  OAI211_X1 U8396 ( .C1(n9384), .C2(n9381), .A(n6639), .B(P1_U3973), .ZN(n9402) );
  INV_X1 U8397 ( .A(n9402), .ZN(n6652) );
  OAI211_X1 U8398 ( .C1(n6642), .C2(n6641), .A(n9489), .B(n6640), .ZN(n6650)
         );
  OAI211_X1 U8399 ( .C1(n6645), .C2(n6644), .A(n9497), .B(n6643), .ZN(n6649)
         );
  AOI22_X1 U8400 ( .A1(n9400), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6648) );
  NAND2_X1 U8401 ( .A1(n9485), .A2(n6646), .ZN(n6647) );
  NAND4_X1 U8402 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n6651)
         );
  OR2_X1 U8403 ( .A1(n6652), .A2(n6651), .ZN(P1_U3245) );
  INV_X1 U8404 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6654) );
  INV_X1 U8405 ( .A(n6653), .ZN(n6655) );
  INV_X1 U8406 ( .A(n8846), .ZN(n8828) );
  OAI222_X1 U8407 ( .A1(n9308), .A2(n6654), .B1(n7231), .B2(n6655), .C1(
        P1_U3086), .C2(n8828), .ZN(P1_U3339) );
  INV_X1 U8408 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6656) );
  OAI222_X1 U8409 ( .A1(n8294), .A2(n6656), .B1(n8304), .B2(n6655), .C1(
        P2_U3151), .C2(n7853), .ZN(P2_U3279) );
  INV_X1 U8410 ( .A(n6657), .ZN(n6658) );
  AOI21_X1 U8411 ( .B1(n6660), .B2(n6659), .A(n6658), .ZN(n6664) );
  AOI22_X1 U8412 ( .A1(n7680), .A2(n6181), .B1(n7729), .B2(n6353), .ZN(n6661)
         );
  OAI21_X1 U8413 ( .B1(n7737), .B2(n9783), .A(n6661), .ZN(n6662) );
  AOI21_X1 U8414 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6695), .A(n6662), .ZN(
        n6663) );
  OAI21_X1 U8415 ( .B1(n6664), .B2(n7707), .A(n6663), .ZN(P2_U3162) );
  INV_X1 U8416 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9859) );
  INV_X1 U8417 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9505) );
  INV_X1 U8418 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10001) );
  INV_X1 U8419 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U8420 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10001), .B2(n6665), .ZN(n9862) );
  NOR2_X1 U8421 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6666) );
  AOI21_X1 U8422 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6666), .ZN(n9865) );
  NOR2_X1 U8423 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6667) );
  AOI21_X1 U8424 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6667), .ZN(n9868) );
  NOR2_X1 U8425 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6668) );
  AOI21_X1 U8426 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6668), .ZN(n9871) );
  NOR2_X1 U8427 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6669) );
  AOI21_X1 U8428 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6669), .ZN(n9874) );
  NOR2_X1 U8429 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6670) );
  AOI21_X1 U8430 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6670), .ZN(n9877) );
  NOR2_X1 U8431 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6671) );
  AOI21_X1 U8432 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6671), .ZN(n9880) );
  NOR2_X1 U8433 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6672) );
  AOI21_X1 U8434 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6672), .ZN(n9883) );
  NOR2_X1 U8435 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6673) );
  AOI21_X1 U8436 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6673), .ZN(n10051) );
  INV_X1 U8437 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9780) );
  INV_X1 U8438 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U8439 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .B1(n9780), .B2(n9903), .ZN(n10057) );
  NOR2_X1 U8440 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6674) );
  AOI21_X1 U8441 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6674), .ZN(n10054) );
  NOR2_X1 U8442 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6675) );
  AOI21_X1 U8443 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6675), .ZN(n10045) );
  NOR2_X1 U8444 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6676) );
  AOI21_X1 U8445 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6676), .ZN(n10048) );
  AND2_X1 U8446 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6677) );
  NOR2_X1 U8447 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6677), .ZN(n9851) );
  INV_X1 U8448 ( .A(n9851), .ZN(n9852) );
  INV_X1 U8449 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9854) );
  NAND3_X1 U8450 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U8451 ( .A1(n9854), .A2(n9853), .ZN(n9850) );
  NAND2_X1 U8452 ( .A1(n9852), .A2(n9850), .ZN(n10060) );
  NAND2_X1 U8453 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6678) );
  OAI21_X1 U8454 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n6678), .ZN(n10059) );
  NOR2_X1 U8455 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  AOI21_X1 U8456 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10058), .ZN(n10063) );
  NAND2_X1 U8457 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6679) );
  OAI21_X1 U8458 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6679), .ZN(n10062) );
  NOR2_X1 U8459 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  AOI21_X1 U8460 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10061), .ZN(n10066) );
  NOR2_X1 U8461 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6680) );
  AOI21_X1 U8462 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6680), .ZN(n10065) );
  NAND2_X1 U8463 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  OAI21_X1 U8464 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10064), .ZN(n10047) );
  NAND2_X1 U8465 ( .A1(n10048), .A2(n10047), .ZN(n10046) );
  OAI21_X1 U8466 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10046), .ZN(n10044) );
  NAND2_X1 U8467 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  OAI21_X1 U8468 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10043), .ZN(n10053) );
  NAND2_X1 U8469 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  OAI21_X1 U8470 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10052), .ZN(n10056) );
  NAND2_X1 U8471 ( .A1(n10057), .A2(n10056), .ZN(n10055) );
  OAI21_X1 U8472 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10055), .ZN(n10050) );
  NAND2_X1 U8473 ( .A1(n10051), .A2(n10050), .ZN(n10049) );
  OAI21_X1 U8474 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10049), .ZN(n9882) );
  NAND2_X1 U8475 ( .A1(n9883), .A2(n9882), .ZN(n9881) );
  OAI21_X1 U8476 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9881), .ZN(n9879) );
  NAND2_X1 U8477 ( .A1(n9880), .A2(n9879), .ZN(n9878) );
  OAI21_X1 U8478 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9878), .ZN(n9876) );
  NAND2_X1 U8479 ( .A1(n9877), .A2(n9876), .ZN(n9875) );
  OAI21_X1 U8480 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9875), .ZN(n9873) );
  NAND2_X1 U8481 ( .A1(n9874), .A2(n9873), .ZN(n9872) );
  OAI21_X1 U8482 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9872), .ZN(n9870) );
  NAND2_X1 U8483 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  OAI21_X1 U8484 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9869), .ZN(n9867) );
  NAND2_X1 U8485 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  OAI21_X1 U8486 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9866), .ZN(n9864) );
  NAND2_X1 U8487 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  OAI21_X1 U8488 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9863), .ZN(n9861) );
  NAND2_X1 U8489 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  OAI21_X1 U8490 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9860), .ZN(n6681) );
  OR2_X1 U8491 ( .A1(n9505), .A2(n6681), .ZN(n9858) );
  NAND2_X1 U8492 ( .A1(n9859), .A2(n9858), .ZN(n9855) );
  NAND2_X1 U8493 ( .A1(n9505), .A2(n6681), .ZN(n9857) );
  NAND2_X1 U8494 ( .A1(n9855), .A2(n9857), .ZN(n6684) );
  XNOR2_X1 U8495 ( .A(n6684), .B(n6683), .ZN(ADD_1068_U4) );
  OAI21_X1 U8496 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(n6690) );
  MUX2_X1 U8497 ( .A(n8475), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n6689) );
  AOI22_X1 U8498 ( .A1(n8484), .A2(n8791), .B1(n8789), .B2(n8878), .ZN(n6789)
         );
  OAI22_X1 U8499 ( .A1(n6789), .A2(n8459), .B1(n8419), .B2(n9637), .ZN(n6688)
         );
  AOI211_X1 U8500 ( .C1(n6690), .C2(n8495), .A(n6689), .B(n6688), .ZN(n6691)
         );
  INV_X1 U8501 ( .A(n6691), .ZN(P1_U3218) );
  OAI21_X1 U8502 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6700) );
  NAND2_X1 U8503 ( .A1(n6695), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6697) );
  AOI22_X1 U8504 ( .A1(n7680), .A2(n7752), .B1(n7729), .B2(n4851), .ZN(n6696)
         );
  OAI211_X1 U8505 ( .C1(n6698), .C2(n7737), .A(n6697), .B(n6696), .ZN(n6699)
         );
  AOI21_X1 U8506 ( .B1(n7726), .B2(n6700), .A(n6699), .ZN(n6701) );
  INV_X1 U8507 ( .A(n6701), .ZN(P2_U3177) );
  INV_X1 U8508 ( .A(n6702), .ZN(n6723) );
  AOI22_X1 U8509 ( .A1(n8858), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9300), .ZN(n6703) );
  OAI21_X1 U8510 ( .B1(n6723), .B2(n7231), .A(n6703), .ZN(P1_U3338) );
  INV_X1 U8511 ( .A(n6704), .ZN(n6708) );
  NOR2_X1 U8512 ( .A1(n6706), .A2(n6705), .ZN(n6707) );
  NAND2_X1 U8513 ( .A1(n6708), .A2(n6707), .ZN(n6709) );
  AOI22_X1 U8514 ( .A1(n8085), .A2(n6730), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8131), .ZN(n6714) );
  NOR2_X1 U8515 ( .A1(n6178), .A2(n8118), .ZN(n8198) );
  NOR3_X1 U8516 ( .A1(n6711), .A2(n6710), .A3(n9836), .ZN(n6712) );
  OAI21_X1 U8517 ( .B1(n8198), .B2(n6712), .A(n8135), .ZN(n6713) );
  OAI211_X1 U8518 ( .C1(n6406), .C2(n8135), .A(n6714), .B(n6713), .ZN(P2_U3233) );
  INV_X1 U8519 ( .A(n9582), .ZN(n6722) );
  AND2_X1 U8520 ( .A1(n6685), .A2(n6715), .ZN(n6718) );
  OAI211_X1 U8521 ( .C1(n6718), .C2(n6717), .A(n8495), .B(n6716), .ZN(n6721)
         );
  AOI22_X1 U8522 ( .A1(n8878), .A2(n8788), .B1(n8790), .B2(n8484), .ZN(n9577)
         );
  NAND2_X1 U8523 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9403) );
  OAI21_X1 U8524 ( .B1(n9577), .B2(n8459), .A(n9403), .ZN(n6719) );
  AOI21_X1 U8525 ( .B1(n6903), .B2(n4295), .A(n6719), .ZN(n6720) );
  OAI211_X1 U8526 ( .C1(n8508), .C2(n6722), .A(n6721), .B(n6720), .ZN(P1_U3230) );
  INV_X1 U8527 ( .A(n7884), .ZN(n7852) );
  OAI222_X1 U8528 ( .A1(n8304), .A2(n6723), .B1(n8300), .B2(n5341), .C1(
        P2_U3151), .C2(n7852), .ZN(P2_U3278) );
  NAND2_X1 U8529 ( .A1(n7389), .A2(n8129), .ZN(n8133) );
  INV_X1 U8530 ( .A(n8133), .ZN(n6812) );
  OAI21_X1 U8531 ( .B1(n6724), .B2(n6726), .A(n6725), .ZN(n9786) );
  NOR2_X1 U8532 ( .A1(n8106), .A2(n6727), .ZN(n6735) );
  OAI22_X1 U8533 ( .A1(n6728), .A2(n8123), .B1(n6729), .B2(n8118), .ZN(n6733)
         );
  NAND3_X1 U8534 ( .A1(n6724), .A2(n6730), .A3(n6238), .ZN(n6731) );
  AOI21_X1 U8535 ( .B1(n6731), .B2(n8120), .A(n5763), .ZN(n6732) );
  AOI211_X1 U8536 ( .C1(n8127), .C2(n9786), .A(n6733), .B(n6732), .ZN(n6734)
         );
  INV_X1 U8537 ( .A(n6734), .ZN(n9784) );
  AOI211_X1 U8538 ( .C1(n6812), .C2(n9786), .A(n6735), .B(n9784), .ZN(n6736)
         );
  MUX2_X1 U8539 ( .A(n6499), .B(n6736), .S(n8135), .Z(n6737) );
  OAI21_X1 U8540 ( .B1(n9783), .B2(n8092), .A(n6737), .ZN(P2_U3232) );
  NAND3_X1 U8541 ( .A1(n6740), .A2(n6739), .A3(n6738), .ZN(n6741) );
  AOI21_X1 U8542 ( .B1(n9612), .B2(n9608), .A(n9519), .ZN(n6748) );
  NOR2_X1 U8543 ( .A1(n8638), .A2(n6742), .ZN(n6743) );
  AOI211_X1 U8544 ( .C1(n9581), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6744), .B(
        n6743), .ZN(n6745) );
  MUX2_X1 U8545 ( .A(n6746), .B(n6745), .S(n9138), .Z(n6747) );
  OAI21_X1 U8546 ( .B1(n6748), .B2(n6755), .A(n6747), .ZN(P1_U3293) );
  OR2_X1 U8547 ( .A1(n6749), .A2(n4305), .ZN(n9521) );
  AND2_X1 U8548 ( .A1(n9508), .A2(n9521), .ZN(n6750) );
  NAND2_X1 U8549 ( .A1(n6751), .A2(n6756), .ZN(n6772) );
  XNOR2_X1 U8550 ( .A(n6781), .B(n6772), .ZN(n9624) );
  XNOR2_X1 U8551 ( .A(n6781), .B(n6780), .ZN(n6754) );
  INV_X1 U8552 ( .A(n6752), .ZN(n6753) );
  AOI21_X1 U8553 ( .B1(n6754), .B2(n9579), .A(n6753), .ZN(n9622) );
  MUX2_X1 U8554 ( .A(n9622), .B(n6525), .S(n9616), .Z(n6760) );
  NAND2_X1 U8555 ( .A1(n8707), .A2(n6755), .ZN(n6793) );
  INV_X1 U8556 ( .A(n6793), .ZN(n9610) );
  AOI211_X1 U8557 ( .C1(n6756), .C2(n9620), .A(n9160), .B(n9610), .ZN(n9619)
         );
  INV_X1 U8558 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U8559 ( .A1(n9605), .A2(n8707), .B1(n9602), .B2(n6757), .ZN(n6758)
         );
  AOI21_X1 U8560 ( .B1(n9619), .B2(n9612), .A(n6758), .ZN(n6759) );
  OAI211_X1 U8561 ( .C1(n9153), .C2(n9624), .A(n6760), .B(n6759), .ZN(P1_U3292) );
  INV_X1 U8562 ( .A(n6761), .ZN(n6800) );
  INV_X1 U8563 ( .A(n7904), .ZN(n7887) );
  OAI222_X1 U8564 ( .A1(n8304), .A2(n6800), .B1(n8300), .B2(n6762), .C1(
        P2_U3151), .C2(n7887), .ZN(P2_U3277) );
  OR2_X1 U8565 ( .A1(n6763), .A2(n7566), .ZN(n6764) );
  NAND2_X1 U8566 ( .A1(n6874), .A2(n6764), .ZN(n9810) );
  NOR2_X1 U8567 ( .A1(n8080), .A2(n8133), .ZN(n7930) );
  INV_X1 U8568 ( .A(n7930), .ZN(n7009) );
  INV_X1 U8569 ( .A(n8127), .ZN(n7076) );
  AOI22_X1 U8570 ( .A1(n7750), .A2(n8096), .B1(n8099), .B2(n7748), .ZN(n6768)
         );
  XNOR2_X1 U8571 ( .A(n6765), .B(n7566), .ZN(n6766) );
  NAND2_X1 U8572 ( .A1(n6766), .A2(n6238), .ZN(n6767) );
  OAI211_X1 U8573 ( .C1(n9810), .C2(n7076), .A(n6768), .B(n6767), .ZN(n9812)
         );
  NAND2_X1 U8574 ( .A1(n9812), .A2(n8135), .ZN(n6771) );
  OAI22_X1 U8575 ( .A1(n8092), .A2(n9809), .B1(n6994), .B2(n8106), .ZN(n6769)
         );
  AOI21_X1 U8576 ( .B1(n8080), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6769), .ZN(
        n6770) );
  OAI211_X1 U8577 ( .C1(n9810), .C2(n7009), .A(n6771), .B(n6770), .ZN(P2_U3226) );
  NAND2_X1 U8578 ( .A1(n6773), .A2(n6772), .ZN(n6776) );
  NAND2_X1 U8579 ( .A1(n6776), .A2(n6775), .ZN(n9593) );
  XNOR2_X1 U8580 ( .A(n8791), .B(n9629), .ZN(n9594) );
  NAND2_X1 U8581 ( .A1(n9593), .A2(n9594), .ZN(n6778) );
  INV_X1 U8582 ( .A(n8791), .ZN(n6786) );
  NAND2_X1 U8583 ( .A1(n6786), .A2(n9629), .ZN(n6777) );
  NAND2_X1 U8584 ( .A1(n6778), .A2(n6777), .ZN(n6887) );
  NAND2_X1 U8585 ( .A1(n6779), .A2(n6796), .ZN(n6894) );
  NAND2_X1 U8586 ( .A1(n8790), .A2(n9637), .ZN(n8712) );
  NAND2_X1 U8587 ( .A1(n6894), .A2(n8712), .ZN(n6886) );
  XOR2_X1 U8588 ( .A(n6887), .B(n6886), .Z(n9635) );
  INV_X1 U8589 ( .A(n6773), .ZN(n6781) );
  NAND2_X1 U8590 ( .A1(n6781), .A2(n6780), .ZN(n6784) );
  NAND2_X1 U8591 ( .A1(n6782), .A2(n9620), .ZN(n6783) );
  NAND2_X1 U8592 ( .A1(n6784), .A2(n6783), .ZN(n9595) );
  INV_X1 U8593 ( .A(n9594), .ZN(n6785) );
  NAND2_X1 U8594 ( .A1(n9595), .A2(n6785), .ZN(n6788) );
  NAND2_X1 U8595 ( .A1(n6786), .A2(n6792), .ZN(n6787) );
  XNOR2_X1 U8596 ( .A(n6893), .B(n6886), .ZN(n6790) );
  OAI21_X1 U8597 ( .B1(n6790), .B2(n9596), .A(n6789), .ZN(n9638) );
  NAND2_X1 U8598 ( .A1(n9638), .A2(n9138), .ZN(n6798) );
  OAI22_X1 U8599 ( .A1(n9138), .A2(n6791), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9602), .ZN(n6795) );
  OAI211_X1 U8600 ( .C1(n9607), .C2(n9637), .A(n9587), .B(n9608), .ZN(n9636)
         );
  NOR2_X1 U8601 ( .A1(n9636), .A2(n9167), .ZN(n6794) );
  AOI211_X1 U8602 ( .C1(n9519), .C2(n6796), .A(n6795), .B(n6794), .ZN(n6797)
         );
  OAI211_X1 U8603 ( .C1(n9635), .C2(n9153), .A(n6798), .B(n6797), .ZN(P1_U3290) );
  INV_X1 U8604 ( .A(n8865), .ZN(n9500) );
  INV_X1 U8605 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6799) );
  OAI222_X1 U8606 ( .A1(P1_U3086), .A2(n9500), .B1(n7231), .B2(n6800), .C1(
        n6799), .C2(n9308), .ZN(P1_U3337) );
  OR2_X1 U8607 ( .A1(n6826), .A2(n6827), .ZN(n6824) );
  AND2_X1 U8608 ( .A1(n6824), .A2(n6801), .ZN(n6804) );
  NAND2_X1 U8609 ( .A1(n6824), .A2(n6802), .ZN(n6861) );
  OAI21_X1 U8610 ( .B1(n6804), .B2(n6803), .A(n6861), .ZN(n6805) );
  NAND2_X1 U8611 ( .A1(n6805), .A2(n7726), .ZN(n6810) );
  INV_X1 U8612 ( .A(n6806), .ZN(n6808) );
  OAI22_X1 U8613 ( .A1(n7737), .A2(n4595), .B1(n7694), .B2(n8119), .ZN(n6807)
         );
  AOI211_X1 U8614 ( .C1(n7680), .C2(n7751), .A(n6808), .B(n6807), .ZN(n6809)
         );
  OAI211_X1 U8615 ( .C1(n6949), .C2(n7341), .A(n6810), .B(n6809), .ZN(P2_U3170) );
  XOR2_X1 U8616 ( .A(n7564), .B(n6811), .Z(n9803) );
  NOR2_X1 U8617 ( .A1(n8127), .A2(n6812), .ZN(n6813) );
  INV_X1 U8618 ( .A(n6934), .ZN(n6814) );
  AOI22_X1 U8619 ( .A1(n8085), .A2(n6815), .B1(n8131), .B2(n6814), .ZN(n6823)
         );
  NAND2_X1 U8620 ( .A1(n6817), .A2(n7564), .ZN(n6818) );
  NAND3_X1 U8621 ( .A1(n6816), .A2(n6238), .A3(n6818), .ZN(n6820) );
  AOI22_X1 U8622 ( .A1(n7749), .A2(n8099), .B1(n8096), .B2(n7751), .ZN(n6819)
         );
  AND2_X1 U8623 ( .A1(n6820), .A2(n6819), .ZN(n9804) );
  MUX2_X1 U8624 ( .A(n6821), .B(n9804), .S(n8135), .Z(n6822) );
  OAI211_X1 U8625 ( .C1(n9803), .C2(n8088), .A(n6823), .B(n6822), .ZN(P2_U3227) );
  INV_X1 U8626 ( .A(n6824), .ZN(n6825) );
  AOI211_X1 U8627 ( .C1(n6827), .C2(n6826), .A(n7707), .B(n6825), .ZN(n6831)
         );
  MUX2_X1 U8628 ( .A(n7341), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6829) );
  AOI22_X1 U8629 ( .A1(n7680), .A2(n4596), .B1(n7729), .B2(n6181), .ZN(n6828)
         );
  OAI211_X1 U8630 ( .C1(n9795), .C2(n7737), .A(n6829), .B(n6828), .ZN(n6830)
         );
  OR2_X1 U8631 ( .A1(n6831), .A2(n6830), .ZN(P2_U3158) );
  NAND2_X1 U8632 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6854), .ZN(n6834) );
  OAI21_X1 U8633 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6854), .A(n6834), .ZN(
        n9760) );
  XOR2_X1 U8634 ( .A(n6855), .B(n7010), .Z(n6835) );
  AOI21_X1 U8635 ( .B1(n6837), .B2(n6835), .A(n7011), .ZN(n6860) );
  MUX2_X1 U8636 ( .A(n6837), .B(n6836), .S(n6156), .Z(n6839) );
  AND2_X1 U8637 ( .A1(n6839), .A2(n7028), .ZN(n7020) );
  INV_X1 U8638 ( .A(n7020), .ZN(n6838) );
  OAI21_X1 U8639 ( .B1(n7028), .B2(n6839), .A(n6838), .ZN(n6846) );
  MUX2_X1 U8640 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6156), .Z(n6843) );
  NOR2_X1 U8641 ( .A1(n6843), .A2(n6854), .ZN(n6844) );
  INV_X1 U8642 ( .A(n6840), .ZN(n6842) );
  AOI21_X1 U8643 ( .B1(n6843), .B2(n6854), .A(n6844), .ZN(n9772) );
  AND2_X1 U8644 ( .A1(n9773), .A2(n9772), .ZN(n9776) );
  NOR2_X1 U8645 ( .A1(n6845), .A2(n6846), .ZN(n7019) );
  AOI21_X1 U8646 ( .B1(n6846), .B2(n6845), .A(n7019), .ZN(n6849) );
  NAND2_X1 U8647 ( .A1(n7915), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6848) );
  AND2_X1 U8648 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7234) );
  INV_X1 U8649 ( .A(n7234), .ZN(n6847) );
  OAI211_X1 U8650 ( .C1(n6849), .C2(n7913), .A(n6848), .B(n6847), .ZN(n6858)
         );
  NAND2_X1 U8651 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6854), .ZN(n6853) );
  OAI21_X1 U8652 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6854), .A(n6853), .ZN(
        n9757) );
  NOR2_X1 U8653 ( .A1(n6856), .A2(n9769), .ZN(n6857) );
  AOI211_X1 U8654 ( .C1(n9767), .C2(n7028), .A(n6858), .B(n6857), .ZN(n6859)
         );
  OAI21_X1 U8655 ( .B1(n6860), .B2(n9762), .A(n6859), .ZN(P2_U3191) );
  INV_X1 U8656 ( .A(n6861), .ZN(n6864) );
  NOR3_X1 U8657 ( .A1(n6864), .A2(n6863), .A3(n6862), .ZN(n6867) );
  INV_X1 U8658 ( .A(n6865), .ZN(n6866) );
  OAI21_X1 U8659 ( .B1(n6867), .B2(n6866), .A(n7726), .ZN(n6872) );
  OAI22_X1 U8660 ( .A1(n7737), .A2(n6966), .B1(n7694), .B2(n6868), .ZN(n6869)
         );
  AOI211_X1 U8661 ( .C1(n7680), .C2(n7750), .A(n6870), .B(n6869), .ZN(n6871)
         );
  OAI211_X1 U8662 ( .C1(n6965), .C2(n7341), .A(n6872), .B(n6871), .ZN(P2_U3167) );
  NAND2_X1 U8663 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  AND2_X1 U8664 ( .A1(n7429), .A2(n7420), .ZN(n7565) );
  XNOR2_X1 U8665 ( .A(n6875), .B(n7565), .ZN(n9815) );
  XOR2_X1 U8666 ( .A(n7565), .B(n6876), .Z(n6877) );
  OAI222_X1 U8667 ( .A1(n8120), .A2(n7090), .B1(n8118), .B2(n6878), .C1(n6877), 
        .C2(n8123), .ZN(n9817) );
  NAND2_X1 U8668 ( .A1(n9817), .A2(n8135), .ZN(n6881) );
  OAI22_X1 U8669 ( .A1(n8092), .A2(n9814), .B1(n7094), .B2(n8106), .ZN(n6879)
         );
  AOI21_X1 U8670 ( .B1(n8080), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6879), .ZN(
        n6880) );
  OAI211_X1 U8671 ( .C1(n9815), .C2(n8088), .A(n6881), .B(n6880), .ZN(P2_U3225) );
  INV_X1 U8672 ( .A(n6882), .ZN(n6884) );
  OAI222_X1 U8673 ( .A1(P2_U3151), .A2(n7918), .B1(n8304), .B2(n6884), .C1(
        n8300), .C2(n6883), .ZN(P2_U3276) );
  INV_X1 U8674 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6885) );
  OAI222_X1 U8675 ( .A1(n9308), .A2(n6885), .B1(n7231), .B2(n6884), .C1(
        P1_U3086), .C2(n4305), .ZN(P1_U3336) );
  NAND2_X1 U8676 ( .A1(n6887), .A2(n6886), .ZN(n6889) );
  NAND2_X1 U8677 ( .A1(n6779), .A2(n9637), .ZN(n6888) );
  NAND2_X1 U8678 ( .A1(n6889), .A2(n6888), .ZN(n9585) );
  INV_X1 U8679 ( .A(n8789), .ZN(n6890) );
  NAND2_X1 U8680 ( .A1(n6890), .A2(n6903), .ZN(n6895) );
  INV_X1 U8681 ( .A(n6903), .ZN(n9642) );
  NAND2_X1 U8682 ( .A1(n8789), .A2(n9642), .ZN(n8713) );
  NAND2_X1 U8683 ( .A1(n6895), .A2(n8713), .ZN(n9586) );
  NAND2_X1 U8684 ( .A1(n9585), .A2(n9586), .ZN(n6892) );
  NAND2_X1 U8685 ( .A1(n6890), .A2(n9642), .ZN(n6891) );
  NAND2_X1 U8686 ( .A1(n6892), .A2(n6891), .ZN(n6915) );
  INV_X1 U8687 ( .A(n8788), .ZN(n6977) );
  NAND2_X1 U8688 ( .A1(n6977), .A2(n8393), .ZN(n9559) );
  INV_X1 U8689 ( .A(n8393), .ZN(n9649) );
  NAND2_X1 U8690 ( .A1(n8788), .A2(n9649), .ZN(n8716) );
  NAND2_X1 U8691 ( .A1(n9559), .A2(n8716), .ZN(n8636) );
  XNOR2_X1 U8692 ( .A(n6915), .B(n8636), .ZN(n9647) );
  INV_X1 U8693 ( .A(n9647), .ZN(n6909) );
  INV_X1 U8694 ( .A(n8636), .ZN(n6897) );
  INV_X1 U8695 ( .A(n8713), .ZN(n6896) );
  NAND2_X1 U8696 ( .A1(n8522), .A2(n6897), .ZN(n9560) );
  OAI21_X1 U8697 ( .B1(n6897), .B2(n8522), .A(n9560), .ZN(n6898) );
  NAND2_X1 U8698 ( .A1(n6898), .A2(n9579), .ZN(n6902) );
  NAND2_X1 U8699 ( .A1(n8789), .A2(n8484), .ZN(n6900) );
  NAND2_X1 U8700 ( .A1(n8787), .A2(n8878), .ZN(n6899) );
  NAND2_X1 U8701 ( .A1(n6900), .A2(n6899), .ZN(n8391) );
  INV_X1 U8702 ( .A(n8391), .ZN(n6901) );
  NAND2_X1 U8703 ( .A1(n6902), .A2(n6901), .ZN(n9652) );
  AOI21_X1 U8704 ( .B1(n9588), .B2(n8393), .A(n9160), .ZN(n6904) );
  NAND2_X1 U8705 ( .A1(n6904), .A2(n9569), .ZN(n9648) );
  AOI22_X1 U8706 ( .A1(n9616), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8392), .B2(
        n9581), .ZN(n6906) );
  NAND2_X1 U8707 ( .A1(n9519), .A2(n8393), .ZN(n6905) );
  OAI211_X1 U8708 ( .C1(n9648), .C2(n9167), .A(n6906), .B(n6905), .ZN(n6907)
         );
  AOI21_X1 U8709 ( .B1(n9652), .B2(n9138), .A(n6907), .ZN(n6908) );
  OAI21_X1 U8710 ( .B1(n6909), .B2(n9153), .A(n6908), .ZN(P1_U3288) );
  INV_X1 U8711 ( .A(n8787), .ZN(n6918) );
  NAND2_X1 U8712 ( .A1(n6918), .A2(n6919), .ZN(n8719) );
  NAND2_X1 U8713 ( .A1(n8787), .A2(n9655), .ZN(n8523) );
  NAND2_X1 U8714 ( .A1(n4522), .A2(n8523), .ZN(n7048) );
  NAND2_X1 U8715 ( .A1(n7043), .A2(n6920), .ZN(n9542) );
  NAND2_X1 U8716 ( .A1(n8786), .A2(n9662), .ZN(n7110) );
  NAND2_X1 U8717 ( .A1(n9542), .A2(n7110), .ZN(n8515) );
  XNOR2_X1 U8718 ( .A(n7048), .B(n8515), .ZN(n6910) );
  NAND2_X1 U8719 ( .A1(n6910), .A2(n9579), .ZN(n6914) );
  NAND2_X1 U8720 ( .A1(n8787), .A2(n8484), .ZN(n6912) );
  NAND2_X1 U8721 ( .A1(n8785), .A2(n8878), .ZN(n6911) );
  NAND2_X1 U8722 ( .A1(n6912), .A2(n6911), .ZN(n7062) );
  INV_X1 U8723 ( .A(n7062), .ZN(n6913) );
  NAND2_X1 U8724 ( .A1(n6914), .A2(n6913), .ZN(n9665) );
  INV_X1 U8725 ( .A(n9665), .ZN(n6925) );
  NAND2_X1 U8726 ( .A1(n6915), .A2(n8636), .ZN(n6917) );
  NAND2_X1 U8727 ( .A1(n6977), .A2(n9649), .ZN(n6916) );
  NAND2_X1 U8728 ( .A1(n8719), .A2(n8523), .ZN(n9568) );
  XNOR2_X1 U8729 ( .A(n7042), .B(n8515), .ZN(n9660) );
  NAND2_X1 U8730 ( .A1(n9570), .A2(n9662), .ZN(n9553) );
  OAI211_X1 U8731 ( .C1(n9570), .C2(n9662), .A(n9608), .B(n9553), .ZN(n9661)
         );
  AOI22_X1 U8732 ( .A1(n9616), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7065), .B2(
        n9581), .ZN(n6922) );
  NAND2_X1 U8733 ( .A1(n9519), .A2(n6920), .ZN(n6921) );
  OAI211_X1 U8734 ( .C1(n9661), .C2(n9167), .A(n6922), .B(n6921), .ZN(n6923)
         );
  AOI21_X1 U8735 ( .B1(n9660), .B2(n9590), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8736 ( .B1(n6925), .B2(n9616), .A(n6924), .ZN(P1_U3286) );
  AOI21_X1 U8737 ( .B1(n6926), .B2(n6927), .A(n7707), .ZN(n6928) );
  NAND2_X1 U8738 ( .A1(n6928), .A2(n6983), .ZN(n6933) );
  OAI22_X1 U8739 ( .A1(n7737), .A2(n9805), .B1(n7694), .B2(n6929), .ZN(n6930)
         );
  AOI211_X1 U8740 ( .C1(n7680), .C2(n7749), .A(n6931), .B(n6930), .ZN(n6932)
         );
  OAI211_X1 U8741 ( .C1(n6934), .C2(n7341), .A(n6933), .B(n6932), .ZN(P2_U3179) );
  XNOR2_X1 U8742 ( .A(n6935), .B(n7568), .ZN(n9820) );
  XNOR2_X1 U8743 ( .A(n6936), .B(n7568), .ZN(n6939) );
  OAI22_X1 U8744 ( .A1(n6937), .A2(n8120), .B1(n7345), .B2(n8118), .ZN(n6938)
         );
  AOI21_X1 U8745 ( .B1(n6939), .B2(n6238), .A(n6938), .ZN(n6940) );
  OAI21_X1 U8746 ( .B1(n9820), .B2(n7076), .A(n6940), .ZN(n9822) );
  NAND2_X1 U8747 ( .A1(n9822), .A2(n8135), .ZN(n6943) );
  INV_X1 U8748 ( .A(n9819), .ZN(n7235) );
  OAI22_X1 U8749 ( .A1(n8135), .A2(n6837), .B1(n7233), .B2(n8106), .ZN(n6941)
         );
  AOI21_X1 U8750 ( .B1(n8085), .B2(n7235), .A(n6941), .ZN(n6942) );
  OAI211_X1 U8751 ( .C1(n9820), .C2(n7009), .A(n6943), .B(n6942), .ZN(P2_U3224) );
  INV_X1 U8752 ( .A(n6944), .ZN(n6954) );
  OAI222_X1 U8753 ( .A1(n8304), .A2(n6954), .B1(P2_U3151), .B2(n7586), .C1(
        n10011), .C2(n8300), .ZN(P2_U3275) );
  XNOR2_X1 U8754 ( .A(n6945), .B(n6946), .ZN(n6947) );
  AOI222_X1 U8755 ( .A1(n6238), .A2(n6947), .B1(n7752), .B2(n8096), .C1(n7751), 
        .C2(n8099), .ZN(n9799) );
  XNOR2_X1 U8756 ( .A(n6948), .B(n7560), .ZN(n9801) );
  OAI22_X1 U8757 ( .A1(n8092), .A2(n4595), .B1(n6949), .B2(n8106), .ZN(n6951)
         );
  NOR2_X1 U8758 ( .A1(n8135), .A2(n6421), .ZN(n6950) );
  AOI211_X1 U8759 ( .C1(n9801), .C2(n8112), .A(n6951), .B(n6950), .ZN(n6952)
         );
  OAI21_X1 U8760 ( .B1(n8080), .B2(n9799), .A(n6952), .ZN(P2_U3229) );
  OAI222_X1 U8761 ( .A1(P1_U3086), .A2(n6955), .B1(n7231), .B2(n6954), .C1(
        n6953), .C2(n9308), .ZN(P1_U3335) );
  INV_X1 U8762 ( .A(n6957), .ZN(n7562) );
  XNOR2_X1 U8763 ( .A(n6956), .B(n7562), .ZN(n6958) );
  AOI222_X1 U8764 ( .A1(n6238), .A2(n6958), .B1(n6181), .B2(n8096), .C1(n4596), 
        .C2(n8099), .ZN(n9794) );
  OAI22_X1 U8765 ( .A1(n8092), .A2(n9795), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8106), .ZN(n6961) );
  XNOR2_X1 U8766 ( .A(n6959), .B(n7562), .ZN(n9793) );
  NOR2_X1 U8767 ( .A1(n8088), .A2(n9793), .ZN(n6960) );
  AOI211_X1 U8768 ( .C1(n8080), .C2(P2_REG2_REG_3__SCAN_IN), .A(n6961), .B(
        n6960), .ZN(n6962) );
  OAI21_X1 U8769 ( .B1(n8080), .B2(n9794), .A(n6962), .ZN(P2_U3230) );
  XNOR2_X1 U8770 ( .A(n7561), .B(n6963), .ZN(n6964) );
  AOI222_X1 U8771 ( .A1(n6238), .A2(n6964), .B1(n7750), .B2(n8099), .C1(n4596), 
        .C2(n8096), .ZN(n9839) );
  OAI22_X1 U8772 ( .A1(n8092), .A2(n6966), .B1(n6965), .B2(n8106), .ZN(n6969)
         );
  XNOR2_X1 U8773 ( .A(n6967), .B(n7561), .ZN(n9840) );
  NOR2_X1 U8774 ( .A1(n9840), .A2(n8088), .ZN(n6968) );
  AOI211_X1 U8775 ( .C1(n8080), .C2(P2_REG2_REG_5__SCAN_IN), .A(n6969), .B(
        n6968), .ZN(n6970) );
  OAI21_X1 U8776 ( .B1(n8080), .B2(n9839), .A(n6970), .ZN(P2_U3228) );
  INV_X1 U8777 ( .A(n6971), .ZN(n6976) );
  AOI21_X1 U8778 ( .B1(n6973), .B2(n6975), .A(n6972), .ZN(n6974) );
  AOI21_X1 U8779 ( .B1(n6976), .B2(n6975), .A(n6974), .ZN(n6981) );
  OAI22_X1 U8780 ( .A1(n6977), .A2(n8908), .B1(n7043), .B2(n8505), .ZN(n9562)
         );
  AOI22_X1 U8781 ( .A1(n9562), .A2(n8506), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6978) );
  OAI21_X1 U8782 ( .B1(n9655), .B2(n8419), .A(n6978), .ZN(n6979) );
  AOI21_X1 U8783 ( .B1(n9564), .B2(n8475), .A(n6979), .ZN(n6980) );
  OAI21_X1 U8784 ( .B1(n6981), .B2(n8511), .A(n6980), .ZN(P1_U3239) );
  AND2_X1 U8785 ( .A1(n6983), .A2(n6982), .ZN(n6986) );
  OAI21_X1 U8786 ( .B1(n6986), .B2(n6985), .A(n6984), .ZN(n6987) );
  NAND2_X1 U8787 ( .A1(n6987), .A2(n7726), .ZN(n6993) );
  INV_X1 U8788 ( .A(n6988), .ZN(n6991) );
  OAI22_X1 U8789 ( .A1(n7737), .A2(n9809), .B1(n7694), .B2(n6989), .ZN(n6990)
         );
  AOI211_X1 U8790 ( .C1(n7680), .C2(n7748), .A(n6991), .B(n6990), .ZN(n6992)
         );
  OAI211_X1 U8791 ( .C1(n6994), .C2(n7341), .A(n6993), .B(n6992), .ZN(P2_U3153) );
  INV_X1 U8792 ( .A(n6995), .ZN(n7041) );
  OAI222_X1 U8793 ( .A1(n8304), .A2(n7041), .B1(P2_U3151), .B2(n7588), .C1(
        n6996), .C2(n8300), .ZN(P2_U3274) );
  INV_X1 U8794 ( .A(n7431), .ZN(n6997) );
  OR2_X1 U8795 ( .A1(n7425), .A2(n6997), .ZN(n7569) );
  XNOR2_X1 U8796 ( .A(n6998), .B(n7569), .ZN(n7001) );
  INV_X1 U8797 ( .A(n7001), .ZN(n9827) );
  INV_X1 U8798 ( .A(n7569), .ZN(n7000) );
  XNOR2_X1 U8799 ( .A(n6999), .B(n7000), .ZN(n7004) );
  NAND2_X1 U8800 ( .A1(n7001), .A2(n8127), .ZN(n7003) );
  AOI22_X1 U8801 ( .A1(n7745), .A2(n8099), .B1(n8096), .B2(n7747), .ZN(n7002)
         );
  OAI211_X1 U8802 ( .C1(n7004), .C2(n8123), .A(n7003), .B(n7002), .ZN(n9829)
         );
  NAND2_X1 U8803 ( .A1(n9829), .A2(n8135), .ZN(n7008) );
  OAI22_X1 U8804 ( .A1(n8135), .A2(n7005), .B1(n7295), .B2(n8106), .ZN(n7006)
         );
  AOI21_X1 U8805 ( .B1(n8085), .B2(n7294), .A(n7006), .ZN(n7007) );
  OAI211_X1 U8806 ( .C1(n9827), .C2(n7009), .A(n7008), .B(n7007), .ZN(P2_U3223) );
  NOR2_X1 U8807 ( .A1(n7028), .A2(n7010), .ZN(n7012) );
  NOR2_X1 U8808 ( .A1(n7012), .A2(n7011), .ZN(n7015) );
  NAND2_X1 U8809 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7134), .ZN(n7013) );
  OAI21_X1 U8810 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7134), .A(n7013), .ZN(
        n7014) );
  NOR2_X1 U8811 ( .A1(n7015), .A2(n7014), .ZN(n7126) );
  AOI21_X1 U8812 ( .B1(n7015), .B2(n7014), .A(n7126), .ZN(n7039) );
  INV_X1 U8813 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7026) );
  INV_X1 U8814 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7016) );
  NOR2_X1 U8815 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7016), .ZN(n7293) );
  INV_X1 U8816 ( .A(n7293), .ZN(n7025) );
  MUX2_X1 U8817 ( .A(n7005), .B(n5892), .S(n6156), .Z(n7018) );
  AND2_X1 U8818 ( .A1(n7018), .A2(n7037), .ZN(n7144) );
  INV_X1 U8819 ( .A(n7144), .ZN(n7017) );
  OAI21_X1 U8820 ( .B1(n7037), .B2(n7018), .A(n7017), .ZN(n7022) );
  NOR2_X1 U8821 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  NOR2_X1 U8822 ( .A1(n7021), .A2(n7022), .ZN(n7143) );
  AOI21_X1 U8823 ( .B1(n7022), .B2(n7021), .A(n7143), .ZN(n7023) );
  OR2_X1 U8824 ( .A1(n7913), .A2(n7023), .ZN(n7024) );
  OAI211_X1 U8825 ( .C1(n9779), .C2(n7026), .A(n7025), .B(n7024), .ZN(n7036)
         );
  NOR2_X1 U8826 ( .A1(n7028), .A2(n7027), .ZN(n7030) );
  NAND2_X1 U8827 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7134), .ZN(n7031) );
  OAI21_X1 U8828 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7134), .A(n7031), .ZN(
        n7032) );
  AOI21_X1 U8829 ( .B1(n7033), .B2(n7032), .A(n7133), .ZN(n7034) );
  NOR2_X1 U8830 ( .A1(n7034), .A2(n9769), .ZN(n7035) );
  AOI211_X1 U8831 ( .C1(n9767), .C2(n7037), .A(n7036), .B(n7035), .ZN(n7038)
         );
  OAI21_X1 U8832 ( .B1(n7039), .B2(n9762), .A(n7038), .ZN(P2_U3192) );
  OAI222_X1 U8833 ( .A1(P1_U3086), .A2(n8637), .B1(n7231), .B2(n7041), .C1(
        n7040), .C2(n9308), .ZN(P1_U3334) );
  NAND2_X1 U8834 ( .A1(n7043), .A2(n9662), .ZN(n7044) );
  NAND2_X1 U8835 ( .A1(n7045), .A2(n7044), .ZN(n9541) );
  INV_X1 U8836 ( .A(n8785), .ZN(n7046) );
  NAND2_X1 U8837 ( .A1(n7046), .A2(n7255), .ZN(n8518) );
  INV_X1 U8838 ( .A(n7255), .ZN(n9668) );
  NAND2_X1 U8839 ( .A1(n8785), .A2(n9668), .ZN(n7109) );
  NAND2_X1 U8840 ( .A1(n8518), .A2(n7109), .ZN(n9544) );
  NAND2_X1 U8841 ( .A1(n7046), .A2(n9668), .ZN(n7047) );
  INV_X1 U8842 ( .A(n8784), .ZN(n7116) );
  NAND2_X1 U8843 ( .A1(n7116), .A2(n8431), .ZN(n8534) );
  NAND2_X1 U8844 ( .A1(n8784), .A2(n9675), .ZN(n8641) );
  NAND2_X1 U8845 ( .A1(n8534), .A2(n8641), .ZN(n7117) );
  XNOR2_X1 U8846 ( .A(n7118), .B(n7117), .ZN(n9673) );
  INV_X1 U8847 ( .A(n9673), .ZN(n7059) );
  OR2_X1 U8848 ( .A1(n7048), .A2(n8515), .ZN(n9543) );
  NAND2_X1 U8849 ( .A1(n9542), .A2(n8518), .ZN(n7107) );
  INV_X1 U8850 ( .A(n7107), .ZN(n8527) );
  NAND2_X1 U8851 ( .A1(n9543), .A2(n8527), .ZN(n7049) );
  NAND2_X1 U8852 ( .A1(n7049), .A2(n7109), .ZN(n7050) );
  XNOR2_X1 U8853 ( .A(n7050), .B(n7117), .ZN(n7051) );
  NAND2_X1 U8854 ( .A1(n7051), .A2(n9579), .ZN(n7052) );
  NAND2_X1 U8855 ( .A1(n8785), .A2(n8484), .ZN(n8428) );
  NAND2_X1 U8856 ( .A1(n7052), .A2(n8428), .ZN(n9678) );
  OR2_X1 U8857 ( .A1(n9553), .A2(n7255), .ZN(n9554) );
  XNOR2_X1 U8858 ( .A(n9554), .B(n9675), .ZN(n7054) );
  NAND2_X1 U8859 ( .A1(n8783), .A2(n8878), .ZN(n8429) );
  INV_X1 U8860 ( .A(n8429), .ZN(n7053) );
  AOI21_X1 U8861 ( .B1(n7054), .B2(n9608), .A(n7053), .ZN(n9674) );
  AOI22_X1 U8862 ( .A1(n9616), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8432), .B2(
        n9581), .ZN(n7056) );
  NAND2_X1 U8863 ( .A1(n9519), .A2(n8431), .ZN(n7055) );
  OAI211_X1 U8864 ( .C1(n9674), .C2(n9167), .A(n7056), .B(n7055), .ZN(n7057)
         );
  AOI21_X1 U8865 ( .B1(n9678), .B2(n9138), .A(n7057), .ZN(n7058) );
  OAI21_X1 U8866 ( .B1(n7059), .B2(n9153), .A(n7058), .ZN(P1_U3284) );
  XOR2_X1 U8867 ( .A(n7061), .B(n7060), .Z(n7067) );
  AOI22_X1 U8868 ( .A1(n8506), .A2(n7062), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7063) );
  OAI21_X1 U8869 ( .B1(n8419), .B2(n9662), .A(n7063), .ZN(n7064) );
  AOI21_X1 U8870 ( .B1(n7065), .B2(n8475), .A(n7064), .ZN(n7066) );
  OAI21_X1 U8871 ( .B1(n7067), .B2(n8511), .A(n7066), .ZN(P1_U3213) );
  NAND2_X1 U8872 ( .A1(n7068), .A2(n7069), .ZN(n7070) );
  NAND3_X1 U8873 ( .A1(n7071), .A2(n6238), .A3(n7070), .ZN(n7073) );
  AOI22_X1 U8874 ( .A1(n7746), .A2(n8096), .B1(n8099), .B2(n7744), .ZN(n7072)
         );
  NAND2_X1 U8875 ( .A1(n7073), .A2(n7072), .ZN(n7095) );
  MUX2_X1 U8876 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n7095), .S(n9884), .Z(n7078)
         );
  NAND2_X1 U8877 ( .A1(n7074), .A2(n7431), .ZN(n7075) );
  XNOR2_X1 U8878 ( .A(n7075), .B(n7570), .ZN(n7100) );
  INV_X1 U8879 ( .A(n9791), .ZN(n9826) );
  INV_X1 U8880 ( .A(n9807), .ZN(n9841) );
  INV_X1 U8881 ( .A(n7352), .ZN(n7079) );
  OAI22_X1 U8882 ( .A1(n7100), .A2(n8273), .B1(n7079), .B2(n8271), .ZN(n7077)
         );
  OR2_X1 U8883 ( .A1(n7078), .A2(n7077), .ZN(P2_U3423) );
  MUX2_X1 U8884 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7095), .S(n9849), .Z(n7081)
         );
  OAI22_X1 U8885 ( .A1(n7100), .A2(n8189), .B1(n7079), .B2(n8180), .ZN(n7080)
         );
  OR2_X1 U8886 ( .A1(n7081), .A2(n7080), .ZN(P2_U3470) );
  INV_X1 U8887 ( .A(n6984), .ZN(n7085) );
  INV_X1 U8888 ( .A(n7082), .ZN(n7084) );
  NOR3_X1 U8889 ( .A1(n7085), .A2(n7084), .A3(n7083), .ZN(n7088) );
  INV_X1 U8890 ( .A(n7086), .ZN(n7087) );
  OAI21_X1 U8891 ( .B1(n7088), .B2(n7087), .A(n7726), .ZN(n7093) );
  NOR2_X1 U8892 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7089), .ZN(n9765) );
  OAI22_X1 U8893 ( .A1(n7737), .A2(n9814), .B1(n7694), .B2(n7090), .ZN(n7091)
         );
  AOI211_X1 U8894 ( .C1(n7680), .C2(n7747), .A(n9765), .B(n7091), .ZN(n7092)
         );
  OAI211_X1 U8895 ( .C1(n7094), .C2(n7341), .A(n7093), .B(n7092), .ZN(P2_U3161) );
  MUX2_X1 U8896 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7095), .S(n8135), .Z(n7096)
         );
  INV_X1 U8897 ( .A(n7096), .ZN(n7099) );
  INV_X1 U8898 ( .A(n7097), .ZN(n7353) );
  AOI22_X1 U8899 ( .A1(n8085), .A2(n7352), .B1(n8131), .B2(n7353), .ZN(n7098)
         );
  OAI211_X1 U8900 ( .C1(n7100), .C2(n8088), .A(n7099), .B(n7098), .ZN(P2_U3222) );
  INV_X1 U8901 ( .A(n7101), .ZN(n7105) );
  OAI222_X1 U8902 ( .A1(n8294), .A2(n7103), .B1(n8304), .B2(n7105), .C1(n7102), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U8903 ( .A1(n9308), .A2(n7106), .B1(n7231), .B2(n7105), .C1(
        P1_U3086), .C2(n7104), .ZN(P1_U3333) );
  NAND2_X1 U8904 ( .A1(n9688), .A2(n8782), .ZN(n8537) );
  INV_X1 U8905 ( .A(n8782), .ZN(n7193) );
  NAND2_X1 U8906 ( .A1(n8473), .A2(n7193), .ZN(n8540) );
  NAND2_X1 U8907 ( .A1(n8537), .A2(n8540), .ZN(n8646) );
  AND2_X1 U8908 ( .A1(n8641), .A2(n7109), .ZN(n8525) );
  NAND2_X1 U8909 ( .A1(n7107), .A2(n8525), .ZN(n7108) );
  NAND2_X1 U8910 ( .A1(n7108), .A2(n8534), .ZN(n8645) );
  AND2_X1 U8911 ( .A1(n7110), .A2(n7109), .ZN(n8643) );
  INV_X1 U8912 ( .A(n8783), .ZN(n7111) );
  NAND2_X1 U8913 ( .A1(n7111), .A2(n7190), .ZN(n8536) );
  INV_X1 U8914 ( .A(n7190), .ZN(n9682) );
  NAND2_X1 U8915 ( .A1(n8783), .A2(n9682), .ZN(n8722) );
  NAND2_X1 U8916 ( .A1(n7112), .A2(n7181), .ZN(n7176) );
  NAND2_X1 U8917 ( .A1(n7176), .A2(n8536), .ZN(n7196) );
  XOR2_X1 U8918 ( .A(n8646), .B(n7196), .Z(n7115) );
  NAND2_X1 U8919 ( .A1(n8783), .A2(n8484), .ZN(n7114) );
  NAND2_X1 U8920 ( .A1(n8909), .A2(n8878), .ZN(n7113) );
  NAND2_X1 U8921 ( .A1(n7114), .A2(n7113), .ZN(n8472) );
  AOI21_X1 U8922 ( .B1(n7115), .B2(n9579), .A(n8472), .ZN(n9687) );
  XNOR2_X1 U8923 ( .A(n7194), .B(n8646), .ZN(n9690) );
  NAND2_X1 U8924 ( .A1(n9690), .A2(n9590), .ZN(n7125) );
  OR2_X1 U8925 ( .A1(n7190), .A2(n8431), .ZN(n7119) );
  OAI21_X1 U8926 ( .B1(n7185), .B2(n9688), .A(n9608), .ZN(n7120) );
  OR2_X1 U8927 ( .A1(n7120), .A2(n7200), .ZN(n9686) );
  INV_X1 U8928 ( .A(n9686), .ZN(n7123) );
  AOI22_X1 U8929 ( .A1(n9616), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8474), .B2(
        n9581), .ZN(n7121) );
  OAI21_X1 U8930 ( .B1(n9605), .B2(n9688), .A(n7121), .ZN(n7122) );
  AOI21_X1 U8931 ( .B1(n7123), .B2(n9612), .A(n7122), .ZN(n7124) );
  OAI211_X1 U8932 ( .C1(n9616), .C2(n9687), .A(n7125), .B(n7124), .ZN(P1_U3282) );
  NOR2_X1 U8933 ( .A1(n7171), .A2(n7127), .ZN(n7128) );
  XNOR2_X1 U8934 ( .A(n7127), .B(n7171), .ZN(n7158) );
  AOI22_X1 U8935 ( .A1(n7149), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7224), .B2(
        n7763), .ZN(n7129) );
  AOI21_X1 U8936 ( .B1(n4387), .B2(n7129), .A(n7753), .ZN(n7156) );
  INV_X1 U8937 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7132) );
  INV_X1 U8938 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7130) );
  NOR2_X1 U8939 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7130), .ZN(n7640) );
  INV_X1 U8940 ( .A(n7640), .ZN(n7131) );
  OAI21_X1 U8941 ( .B1(n9779), .B2(n7132), .A(n7131), .ZN(n7141) );
  NOR2_X1 U8942 ( .A1(n7171), .A2(n7135), .ZN(n7136) );
  XNOR2_X1 U8943 ( .A(n7135), .B(n7171), .ZN(n7166) );
  NOR2_X1 U8944 ( .A1(n7167), .A2(n7166), .ZN(n7165) );
  XNOR2_X1 U8945 ( .A(n7763), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7137) );
  AOI21_X1 U8946 ( .B1(n7138), .B2(n7137), .A(n7762), .ZN(n7139) );
  NOR2_X1 U8947 ( .A1(n7139), .A2(n9769), .ZN(n7140) );
  AOI211_X1 U8948 ( .C1(n9767), .C2(n7149), .A(n7141), .B(n7140), .ZN(n7155)
         );
  MUX2_X1 U8949 ( .A(n7142), .B(n7167), .S(n6156), .Z(n7146) );
  AND2_X1 U8950 ( .A1(n7146), .A2(n7171), .ZN(n7147) );
  INV_X1 U8951 ( .A(n7147), .ZN(n7145) );
  OAI21_X1 U8952 ( .B1(n7171), .B2(n7146), .A(n7145), .ZN(n7161) );
  NOR2_X1 U8953 ( .A1(n7160), .A2(n7161), .ZN(n7159) );
  MUX2_X1 U8954 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6156), .Z(n7148) );
  AND2_X1 U8955 ( .A1(n7148), .A2(n7763), .ZN(n7756) );
  INV_X1 U8956 ( .A(n7756), .ZN(n7151) );
  INV_X1 U8957 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7212) );
  MUX2_X1 U8958 ( .A(n7224), .B(n7212), .S(n6156), .Z(n7150) );
  NAND2_X1 U8959 ( .A1(n7150), .A2(n7149), .ZN(n7757) );
  NAND2_X1 U8960 ( .A1(n7151), .A2(n7757), .ZN(n7152) );
  XNOR2_X1 U8961 ( .A(n7758), .B(n7152), .ZN(n7153) );
  NAND2_X1 U8962 ( .A1(n7153), .A2(n9774), .ZN(n7154) );
  OAI211_X1 U8963 ( .C1(n7156), .C2(n9762), .A(n7155), .B(n7154), .ZN(P2_U3194) );
  AOI21_X1 U8964 ( .B1(n7142), .B2(n7158), .A(n7157), .ZN(n7173) );
  AOI21_X1 U8965 ( .B1(n7161), .B2(n7160), .A(n7159), .ZN(n7164) );
  NAND2_X1 U8966 ( .A1(n7915), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7163) );
  AND2_X1 U8967 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7351) );
  INV_X1 U8968 ( .A(n7351), .ZN(n7162) );
  OAI211_X1 U8969 ( .C1(n7164), .C2(n7913), .A(n7163), .B(n7162), .ZN(n7170)
         );
  AOI21_X1 U8970 ( .B1(n7167), .B2(n7166), .A(n7165), .ZN(n7168) );
  NOR2_X1 U8971 ( .A1(n7168), .A2(n9769), .ZN(n7169) );
  AOI211_X1 U8972 ( .C1(n9767), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7172)
         );
  OAI21_X1 U8973 ( .B1(n7173), .B2(n9762), .A(n7172), .ZN(P2_U3193) );
  NAND2_X1 U8974 ( .A1(n7174), .A2(n4761), .ZN(n7175) );
  NAND2_X1 U8975 ( .A1(n7176), .A2(n7175), .ZN(n7180) );
  NAND2_X1 U8976 ( .A1(n8784), .A2(n8484), .ZN(n7178) );
  NAND2_X1 U8977 ( .A1(n8782), .A2(n8878), .ZN(n7177) );
  AND2_X1 U8978 ( .A1(n7178), .A2(n7177), .ZN(n8338) );
  INV_X1 U8979 ( .A(n8338), .ZN(n7179) );
  AOI21_X1 U8980 ( .B1(n7180), .B2(n9579), .A(n7179), .ZN(n9681) );
  XNOR2_X1 U8981 ( .A(n7182), .B(n7181), .ZN(n9684) );
  NAND2_X1 U8982 ( .A1(n9684), .A2(n9590), .ZN(n7192) );
  INV_X1 U8983 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7184) );
  OAI22_X1 U8984 ( .A1(n9138), .A2(n7184), .B1(n7183), .B2(n9602), .ZN(n7189)
         );
  INV_X1 U8985 ( .A(n7185), .ZN(n7187) );
  OAI21_X1 U8986 ( .B1(n9554), .B2(n8431), .A(n7190), .ZN(n7186) );
  NAND3_X1 U8987 ( .A1(n7187), .A2(n9608), .A3(n7186), .ZN(n9680) );
  NOR2_X1 U8988 ( .A1(n9680), .A2(n9167), .ZN(n7188) );
  AOI211_X1 U8989 ( .C1(n9519), .C2(n7190), .A(n7189), .B(n7188), .ZN(n7191)
         );
  OAI211_X1 U8990 ( .C1(n9616), .C2(n9681), .A(n7192), .B(n7191), .ZN(P1_U3283) );
  NAND2_X1 U8991 ( .A1(n8910), .A2(n7195), .ZN(n8728) );
  AND2_X2 U8992 ( .A1(n8663), .A2(n8728), .ZN(n8911) );
  XNOR2_X1 U8993 ( .A(n8912), .B(n8911), .ZN(n9696) );
  INV_X1 U8994 ( .A(n9696), .ZN(n7205) );
  XNOR2_X1 U8995 ( .A(n8662), .B(n8911), .ZN(n7199) );
  NAND2_X1 U8996 ( .A1(n8782), .A2(n8484), .ZN(n7198) );
  NAND2_X1 U8997 ( .A1(n8781), .A2(n8878), .ZN(n7197) );
  AND2_X1 U8998 ( .A1(n7198), .A2(n7197), .ZN(n7271) );
  OAI21_X1 U8999 ( .B1(n7199), .B2(n9596), .A(n7271), .ZN(n9695) );
  OAI211_X1 U9000 ( .C1(n7200), .C2(n9693), .A(n9608), .B(n9531), .ZN(n9692)
         );
  AOI22_X1 U9001 ( .A1(n9616), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7268), .B2(
        n9581), .ZN(n7202) );
  NAND2_X1 U9002 ( .A1(n8910), .A2(n9519), .ZN(n7201) );
  OAI211_X1 U9003 ( .C1(n9692), .C2(n9167), .A(n7202), .B(n7201), .ZN(n7203)
         );
  AOI21_X1 U9004 ( .B1(n9695), .B2(n9138), .A(n7203), .ZN(n7204) );
  OAI21_X1 U9005 ( .B1(n7205), .B2(n9153), .A(n7204), .ZN(P1_U3281) );
  XNOR2_X1 U9006 ( .A(n7206), .B(n7574), .ZN(n7207) );
  AOI222_X1 U9007 ( .A1(n6238), .A2(n7207), .B1(n7745), .B2(n8096), .C1(n7743), 
        .C2(n8099), .ZN(n7223) );
  MUX2_X1 U9008 ( .A(n7208), .B(n7223), .S(n9884), .Z(n7211) );
  INV_X1 U9009 ( .A(n7574), .ZN(n7446) );
  XNOR2_X1 U9010 ( .A(n7209), .B(n7446), .ZN(n7222) );
  INV_X1 U9011 ( .A(n8273), .ZN(n8281) );
  AOI22_X1 U9012 ( .A1(n7222), .A2(n8281), .B1(n8280), .B2(n7653), .ZN(n7210)
         );
  NAND2_X1 U9013 ( .A1(n7211), .A2(n7210), .ZN(P2_U3426) );
  MUX2_X1 U9014 ( .A(n7212), .B(n7223), .S(n9849), .Z(n7214) );
  INV_X1 U9015 ( .A(n8189), .ZN(n8193) );
  AOI22_X1 U9016 ( .A1(n7222), .A2(n8193), .B1(n8192), .B2(n7653), .ZN(n7213)
         );
  NAND2_X1 U9017 ( .A1(n7214), .A2(n7213), .ZN(P2_U3471) );
  NAND2_X1 U9018 ( .A1(n7219), .A2(n7215), .ZN(n7216) );
  OAI211_X1 U9019 ( .C1(n7217), .C2(n9308), .A(n7216), .B(n8770), .ZN(P1_U3332) );
  NAND2_X1 U9020 ( .A1(n7219), .A2(n7218), .ZN(n7221) );
  NAND2_X1 U9021 ( .A1(n7220), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7598) );
  OAI211_X1 U9022 ( .C1(n9960), .C2(n8294), .A(n7221), .B(n7598), .ZN(P2_U3272) );
  INV_X1 U9023 ( .A(n7222), .ZN(n7228) );
  MUX2_X1 U9024 ( .A(n7224), .B(n7223), .S(n8135), .Z(n7227) );
  INV_X1 U9025 ( .A(n7225), .ZN(n7641) );
  AOI22_X1 U9026 ( .A1(n8085), .A2(n7653), .B1(n8131), .B2(n7641), .ZN(n7226)
         );
  OAI211_X1 U9027 ( .C1(n7228), .C2(n8088), .A(n7227), .B(n7226), .ZN(P2_U3221) );
  INV_X1 U9028 ( .A(n7229), .ZN(n7279) );
  OAI222_X1 U9029 ( .A1(P1_U3086), .A2(n7232), .B1(n7231), .B2(n7279), .C1(
        n7230), .C2(n9308), .ZN(P1_U3331) );
  INV_X1 U9030 ( .A(n7233), .ZN(n7245) );
  AOI21_X1 U9031 ( .B1(n7680), .B2(n7746), .A(n7234), .ZN(n7238) );
  NAND2_X1 U9032 ( .A1(n7705), .A2(n7235), .ZN(n7237) );
  NAND2_X1 U9033 ( .A1(n7729), .A2(n7748), .ZN(n7236) );
  NAND3_X1 U9034 ( .A1(n7238), .A2(n7237), .A3(n7236), .ZN(n7244) );
  INV_X1 U9035 ( .A(n7239), .ZN(n7240) );
  AOI211_X1 U9036 ( .C1(n7242), .C2(n7241), .A(n7707), .B(n7240), .ZN(n7243)
         );
  AOI211_X1 U9037 ( .C1(n7245), .C2(n7734), .A(n7244), .B(n7243), .ZN(n7246)
         );
  INV_X1 U9038 ( .A(n7246), .ZN(P2_U3171) );
  XOR2_X1 U9039 ( .A(n8421), .B(n8422), .Z(n7249) );
  INV_X1 U9040 ( .A(n7247), .ZN(n7248) );
  NAND2_X1 U9041 ( .A1(n7249), .A2(n7248), .ZN(n8420) );
  OAI21_X1 U9042 ( .B1(n7249), .B2(n7248), .A(n8420), .ZN(n7250) );
  NAND2_X1 U9043 ( .A1(n7250), .A2(n8495), .ZN(n7257) );
  NAND2_X1 U9044 ( .A1(n8786), .A2(n8484), .ZN(n7252) );
  NAND2_X1 U9045 ( .A1(n8784), .A2(n8878), .ZN(n7251) );
  AND2_X1 U9046 ( .A1(n7252), .A2(n7251), .ZN(n9546) );
  OAI22_X1 U9047 ( .A1(n8459), .A2(n9546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7253), .ZN(n7254) );
  AOI21_X1 U9048 ( .B1(n7255), .B2(n4295), .A(n7254), .ZN(n7256) );
  OAI211_X1 U9049 ( .C1(n8508), .C2(n9549), .A(n7257), .B(n7256), .ZN(P1_U3221) );
  XOR2_X1 U9050 ( .A(n7258), .B(n7573), .Z(n7259) );
  AOI222_X1 U9051 ( .A1(n6238), .A2(n7259), .B1(n7744), .B2(n8096), .C1(n8097), 
        .C2(n8099), .ZN(n8107) );
  MUX2_X1 U9052 ( .A(n7764), .B(n8107), .S(n9849), .Z(n7262) );
  XOR2_X1 U9053 ( .A(n7260), .B(n7573), .Z(n8113) );
  AOI22_X1 U9054 ( .A1(n8113), .A2(n8193), .B1(n8192), .B2(n8110), .ZN(n7261)
         );
  NAND2_X1 U9055 ( .A1(n7262), .A2(n7261), .ZN(P2_U3472) );
  INV_X1 U9056 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7263) );
  MUX2_X1 U9057 ( .A(n7263), .B(n8107), .S(n9884), .Z(n7265) );
  AOI22_X1 U9058 ( .A1(n8113), .A2(n8281), .B1(n8280), .B2(n8110), .ZN(n7264)
         );
  NAND2_X1 U9059 ( .A1(n7265), .A2(n7264), .ZN(P2_U3429) );
  XOR2_X1 U9060 ( .A(n7267), .B(n7266), .Z(n7274) );
  NAND2_X1 U9061 ( .A1(n8475), .A2(n7268), .ZN(n7269) );
  OAI211_X1 U9062 ( .C1(n8459), .C2(n7271), .A(n7270), .B(n7269), .ZN(n7272)
         );
  AOI21_X1 U9063 ( .B1(n8910), .B2(n4295), .A(n7272), .ZN(n7273) );
  OAI21_X1 U9064 ( .B1(n7274), .B2(n8511), .A(n7273), .ZN(P1_U3224) );
  INV_X1 U9065 ( .A(n7275), .ZN(n7289) );
  OAI222_X1 U9066 ( .A1(n8304), .A2(n7289), .B1(P2_U3151), .B2(n7277), .C1(
        n7276), .C2(n8300), .ZN(P2_U3270) );
  OAI222_X1 U9067 ( .A1(n8304), .A2(n7279), .B1(P2_U3151), .B2(n5712), .C1(
        n7278), .C2(n8300), .ZN(P2_U3271) );
  INV_X1 U9068 ( .A(n7281), .ZN(n7450) );
  OR2_X1 U9069 ( .A1(n7451), .A2(n7450), .ZN(n7283) );
  INV_X1 U9070 ( .A(n7283), .ZN(n7575) );
  XNOR2_X1 U9071 ( .A(n7280), .B(n7575), .ZN(n7282) );
  OAI222_X1 U9072 ( .A1(n8118), .A2(n7329), .B1(n8120), .B2(n7644), .C1(n8123), 
        .C2(n7282), .ZN(n8190) );
  AOI21_X1 U9073 ( .B1(n8111), .B2(n8279), .A(n8190), .ZN(n7287) );
  XNOR2_X1 U9074 ( .A(n7284), .B(n7283), .ZN(n8282) );
  OAI22_X1 U9075 ( .A1(n8135), .A2(n7792), .B1(n7330), .B2(n8106), .ZN(n7285)
         );
  AOI21_X1 U9076 ( .B1(n8282), .B2(n8112), .A(n7285), .ZN(n7286) );
  OAI21_X1 U9077 ( .B1(n7287), .B2(n8080), .A(n7286), .ZN(P2_U3219) );
  OAI222_X1 U9078 ( .A1(P1_U3086), .A2(n5615), .B1(n7231), .B2(n7289), .C1(
        n7288), .C2(n9308), .ZN(P1_U3330) );
  XNOR2_X1 U9079 ( .A(n7290), .B(n7345), .ZN(n7292) );
  NAND2_X1 U9080 ( .A1(n7292), .A2(n7291), .ZN(n7348) );
  OAI21_X1 U9081 ( .B1(n7292), .B2(n7291), .A(n7348), .ZN(n7302) );
  AOI21_X1 U9082 ( .B1(n7680), .B2(n7745), .A(n7293), .ZN(n7300) );
  NAND2_X1 U9083 ( .A1(n7705), .A2(n7294), .ZN(n7299) );
  INV_X1 U9084 ( .A(n7295), .ZN(n7296) );
  NAND2_X1 U9085 ( .A1(n7734), .A2(n7296), .ZN(n7298) );
  NAND2_X1 U9086 ( .A1(n7729), .A2(n7747), .ZN(n7297) );
  NAND4_X1 U9087 ( .A1(n7300), .A2(n7299), .A3(n7298), .A4(n7297), .ZN(n7301)
         );
  AOI21_X1 U9088 ( .B1(n7302), .B2(n7726), .A(n7301), .ZN(n7303) );
  INV_X1 U9089 ( .A(n7303), .ZN(P2_U3157) );
  AOI21_X1 U9090 ( .B1(n7305), .B2(n7304), .A(n4375), .ZN(n7310) );
  NAND2_X1 U9091 ( .A1(n7729), .A2(n7744), .ZN(n7306) );
  NAND2_X1 U9092 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7766) );
  OAI211_X1 U9093 ( .C1(n7317), .C2(n7731), .A(n7306), .B(n7766), .ZN(n7308)
         );
  NOR2_X1 U9094 ( .A1(n7341), .A2(n8105), .ZN(n7307) );
  AOI211_X1 U9095 ( .C1(n8110), .C2(n7705), .A(n7308), .B(n7307), .ZN(n7309)
         );
  OAI21_X1 U9096 ( .B1(n7310), .B2(n7707), .A(n7309), .ZN(P2_U3174) );
  INV_X1 U9097 ( .A(n8186), .ZN(n8272) );
  NAND2_X1 U9098 ( .A1(n7326), .A2(n7311), .ZN(n7313) );
  AOI21_X1 U9099 ( .B1(n7313), .B2(n7312), .A(n7707), .ZN(n7315) );
  NAND2_X1 U9100 ( .A1(n7315), .A2(n7314), .ZN(n7321) );
  INV_X1 U9101 ( .A(n8091), .ZN(n7319) );
  AND2_X1 U9102 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7811) );
  AOI21_X1 U9103 ( .B1(n7680), .B2(n8098), .A(n7811), .ZN(n7316) );
  OAI21_X1 U9104 ( .B1(n7317), .B2(n7694), .A(n7316), .ZN(n7318) );
  AOI21_X1 U9105 ( .B1(n7319), .B2(n7734), .A(n7318), .ZN(n7320) );
  OAI211_X1 U9106 ( .C1(n8272), .C2(n7737), .A(n7321), .B(n7320), .ZN(P2_U3181) );
  INV_X1 U9107 ( .A(n8279), .ZN(n7335) );
  INV_X1 U9108 ( .A(n7322), .ZN(n7324) );
  NOR3_X1 U9109 ( .A1(n4375), .A2(n7324), .A3(n7323), .ZN(n7328) );
  NAND2_X1 U9110 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
  OAI21_X1 U9111 ( .B1(n7328), .B2(n7327), .A(n7726), .ZN(n7334) );
  NAND2_X1 U9112 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7785) );
  OAI21_X1 U9113 ( .B1(n7731), .B2(n7329), .A(n7785), .ZN(n7332) );
  NOR2_X1 U9114 ( .A1(n7341), .A2(n7330), .ZN(n7331) );
  AOI211_X1 U9115 ( .C1(n7729), .C2(n7743), .A(n7332), .B(n7331), .ZN(n7333)
         );
  OAI211_X1 U9116 ( .C1(n7335), .C2(n7737), .A(n7334), .B(n7333), .ZN(P2_U3155) );
  XNOR2_X1 U9117 ( .A(n7337), .B(n7336), .ZN(n7344) );
  NAND2_X1 U9118 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7831) );
  OAI21_X1 U9119 ( .B1(n7731), .B2(n7338), .A(n7831), .ZN(n7339) );
  AOI21_X1 U9120 ( .B1(n7729), .B2(n8076), .A(n7339), .ZN(n7340) );
  OAI21_X1 U9121 ( .B1(n8083), .B2(n7341), .A(n7340), .ZN(n7342) );
  AOI21_X1 U9122 ( .B1(n8179), .B2(n7705), .A(n7342), .ZN(n7343) );
  OAI21_X1 U9123 ( .B1(n7344), .B2(n7707), .A(n7343), .ZN(P2_U3166) );
  INV_X1 U9124 ( .A(n7290), .ZN(n7346) );
  NAND2_X1 U9125 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  NAND3_X1 U9126 ( .A1(n7348), .A2(n7646), .A3(n7347), .ZN(n7645) );
  INV_X1 U9127 ( .A(n7645), .ZN(n7350) );
  AOI21_X1 U9128 ( .B1(n7348), .B2(n7347), .A(n7646), .ZN(n7349) );
  NOR3_X1 U9129 ( .A1(n7350), .A2(n7349), .A3(n7707), .ZN(n7359) );
  AOI21_X1 U9130 ( .B1(n7680), .B2(n7744), .A(n7351), .ZN(n7357) );
  NAND2_X1 U9131 ( .A1(n7705), .A2(n7352), .ZN(n7356) );
  NAND2_X1 U9132 ( .A1(n7734), .A2(n7353), .ZN(n7355) );
  NAND2_X1 U9133 ( .A1(n7729), .A2(n7746), .ZN(n7354) );
  NAND4_X1 U9134 ( .A1(n7357), .A2(n7356), .A3(n7355), .A4(n7354), .ZN(n7358)
         );
  OR2_X1 U9135 ( .A1(n7359), .A2(n7358), .ZN(P2_U3176) );
  INV_X1 U9136 ( .A(n7360), .ZN(n7361) );
  NAND2_X1 U9137 ( .A1(n7361), .A2(SI_29_), .ZN(n7365) );
  NAND2_X1 U9138 ( .A1(n7365), .A2(n7364), .ZN(n7373) );
  INV_X1 U9139 ( .A(n7373), .ZN(n7371) );
  INV_X1 U9140 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8293) );
  INV_X1 U9141 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9303) );
  INV_X1 U9142 ( .A(SI_30_), .ZN(n7366) );
  NAND2_X1 U9143 ( .A1(n7367), .A2(n7366), .ZN(n7536) );
  INV_X1 U9144 ( .A(n7367), .ZN(n7368) );
  NAND2_X1 U9145 ( .A1(n7368), .A2(SI_30_), .ZN(n7369) );
  NAND2_X1 U9146 ( .A1(n7536), .A2(n7369), .ZN(n7372) );
  INV_X1 U9147 ( .A(n7372), .ZN(n7370) );
  NAND2_X1 U9148 ( .A1(n7373), .A2(n7372), .ZN(n7374) );
  NAND2_X1 U9149 ( .A1(n7537), .A2(n7374), .ZN(n8609) );
  INV_X1 U9150 ( .A(n7376), .ZN(n7377) );
  OAI22_X1 U9151 ( .A1(n8080), .A2(n9369), .B1(n7378), .B2(n8106), .ZN(n7924)
         );
  AOI21_X1 U9152 ( .B1(n8080), .B2(P2_REG2_REG_30__SCAN_IN), .A(n7924), .ZN(
        n7379) );
  OAI21_X1 U9153 ( .B1(n9368), .B2(n8092), .A(n7379), .ZN(P2_U3203) );
  INV_X1 U9154 ( .A(n7380), .ZN(n8298) );
  OAI222_X1 U9155 ( .A1(n9308), .A2(n7381), .B1(P1_U3086), .B2(n8880), .C1(
        n8298), .C2(n7231), .ZN(P1_U3328) );
  NAND2_X1 U9156 ( .A1(n7382), .A2(n7596), .ZN(n7385) );
  NAND2_X1 U9157 ( .A1(n7382), .A2(n7389), .ZN(n7383) );
  NAND3_X1 U9158 ( .A1(n7390), .A2(n7535), .A3(n7383), .ZN(n7384) );
  OAI21_X1 U9159 ( .B1(n7386), .B2(n7385), .A(n7384), .ZN(n7387) );
  OAI21_X1 U9160 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7393) );
  MUX2_X1 U9161 ( .A(n7391), .B(n7390), .S(n7519), .Z(n7392) );
  NAND3_X1 U9162 ( .A1(n7393), .A2(n8122), .A3(n7392), .ZN(n7400) );
  NAND2_X1 U9163 ( .A1(n7407), .A2(n7394), .ZN(n7397) );
  NAND2_X1 U9164 ( .A1(n7401), .A2(n7395), .ZN(n7396) );
  MUX2_X1 U9165 ( .A(n7397), .B(n7396), .S(n7519), .Z(n7398) );
  INV_X1 U9166 ( .A(n7398), .ZN(n7399) );
  NAND2_X1 U9167 ( .A1(n7400), .A2(n7399), .ZN(n7408) );
  NAND3_X1 U9168 ( .A1(n7408), .A2(n7560), .A3(n7401), .ZN(n7403) );
  NAND3_X1 U9169 ( .A1(n7403), .A2(n7402), .A3(n7412), .ZN(n7406) );
  AND2_X1 U9170 ( .A1(n7414), .A2(n7409), .ZN(n7405) );
  AOI21_X1 U9171 ( .B1(n7406), .B2(n7405), .A(n7404), .ZN(n7419) );
  NAND3_X1 U9172 ( .A1(n7408), .A2(n7560), .A3(n7407), .ZN(n7411) );
  NAND3_X1 U9173 ( .A1(n7411), .A2(n7410), .A3(n7409), .ZN(n7417) );
  AND2_X1 U9174 ( .A1(n7413), .A2(n7412), .ZN(n7416) );
  INV_X1 U9175 ( .A(n7414), .ZN(n7415) );
  AOI21_X1 U9176 ( .B1(n7417), .B2(n7416), .A(n7415), .ZN(n7418) );
  MUX2_X1 U9177 ( .A(n7419), .B(n7418), .S(n7519), .Z(n7424) );
  NAND2_X1 U9178 ( .A1(n7426), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U9179 ( .A1(n7430), .A2(n7429), .ZN(n7421) );
  MUX2_X1 U9180 ( .A(n7422), .B(n7421), .S(n7535), .Z(n7433) );
  INV_X1 U9181 ( .A(n7433), .ZN(n7423) );
  NAND3_X1 U9182 ( .A1(n7424), .A2(n7566), .A3(n7423), .ZN(n7435) );
  INV_X1 U9183 ( .A(n7425), .ZN(n7438) );
  AND2_X1 U9184 ( .A1(n7429), .A2(n7428), .ZN(n7432) );
  OAI211_X1 U9185 ( .C1(n7433), .C2(n7432), .A(n7431), .B(n7430), .ZN(n7434)
         );
  NAND2_X1 U9186 ( .A1(n7439), .A2(n7436), .ZN(n7437) );
  NAND2_X1 U9187 ( .A1(n7439), .A2(n7438), .ZN(n7442) );
  MUX2_X1 U9188 ( .A(n7444), .B(n7443), .S(n7519), .Z(n7445) );
  MUX2_X1 U9189 ( .A(n7448), .B(n7447), .S(n7519), .Z(n7449) );
  MUX2_X1 U9190 ( .A(n7451), .B(n7450), .S(n7535), .Z(n7452) );
  INV_X1 U9191 ( .A(n7452), .ZN(n7453) );
  NAND2_X1 U9192 ( .A1(n7454), .A2(n7453), .ZN(n7455) );
  INV_X1 U9193 ( .A(n8093), .ZN(n8089) );
  NAND2_X1 U9194 ( .A1(n7455), .A2(n8089), .ZN(n7460) );
  NAND3_X1 U9195 ( .A1(n7460), .A2(n7456), .A3(n7462), .ZN(n7457) );
  NAND3_X1 U9196 ( .A1(n7457), .A2(n7535), .A3(n7458), .ZN(n7468) );
  INV_X1 U9197 ( .A(n8058), .ZN(n8061) );
  NAND4_X1 U9198 ( .A1(n7460), .A2(n8061), .A3(n7459), .A4(n7458), .ZN(n7466)
         );
  NAND2_X1 U9199 ( .A1(n7557), .A2(n7461), .ZN(n7464) );
  NAND2_X1 U9200 ( .A1(n7462), .A2(n7519), .ZN(n7463) );
  AOI22_X1 U9201 ( .A1(n7464), .A2(n7519), .B1(n8061), .B2(n7463), .ZN(n7465)
         );
  NAND2_X1 U9202 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  INV_X1 U9203 ( .A(n7559), .ZN(n7469) );
  NAND2_X1 U9204 ( .A1(n7469), .A2(n7478), .ZN(n7470) );
  INV_X1 U9205 ( .A(n7471), .ZN(n7472) );
  NOR2_X1 U9206 ( .A1(n7559), .A2(n7472), .ZN(n7474) );
  INV_X1 U9207 ( .A(n7477), .ZN(n7473) );
  AOI21_X1 U9208 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7476) );
  NAND3_X1 U9209 ( .A1(n7483), .A2(n7477), .A3(n7480), .ZN(n7485) );
  INV_X1 U9210 ( .A(n7478), .ZN(n7479) );
  NOR2_X1 U9211 ( .A1(n8025), .A2(n7479), .ZN(n7482) );
  NAND2_X1 U9212 ( .A1(n7492), .A2(n7480), .ZN(n7481) );
  AOI21_X1 U9213 ( .B1(n7483), .B2(n7482), .A(n7481), .ZN(n7484) );
  MUX2_X1 U9214 ( .A(n7485), .B(n7484), .S(n7535), .Z(n7490) );
  INV_X1 U9215 ( .A(n7487), .ZN(n7489) );
  AND2_X1 U9216 ( .A1(n7487), .A2(n7486), .ZN(n7488) );
  OAI22_X1 U9217 ( .A1(n7490), .A2(n7489), .B1(n7488), .B2(n7535), .ZN(n7491)
         );
  OAI211_X1 U9218 ( .C1(n7492), .C2(n7535), .A(n7491), .B(n8005), .ZN(n7499)
         );
  INV_X1 U9219 ( .A(n7501), .ZN(n7504) );
  NAND2_X1 U9220 ( .A1(n8159), .A2(n8016), .ZN(n7493) );
  AND2_X1 U9221 ( .A1(n7500), .A2(n7493), .ZN(n7497) );
  INV_X1 U9222 ( .A(n7494), .ZN(n7495) );
  NOR2_X1 U9223 ( .A1(n7556), .A2(n7495), .ZN(n7496) );
  MUX2_X1 U9224 ( .A(n7497), .B(n7496), .S(n7519), .Z(n7498) );
  NAND3_X1 U9225 ( .A1(n7499), .A2(n7985), .A3(n7498), .ZN(n7508) );
  INV_X1 U9226 ( .A(n7500), .ZN(n7555) );
  OAI21_X1 U9227 ( .B1(n7501), .B2(n7555), .A(n7502), .ZN(n7506) );
  NAND2_X1 U9228 ( .A1(n7502), .A2(n6253), .ZN(n7503) );
  NAND2_X1 U9229 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  MUX2_X1 U9230 ( .A(n7506), .B(n7505), .S(n7535), .Z(n7507) );
  NAND3_X1 U9231 ( .A1(n7508), .A2(n7972), .A3(n7507), .ZN(n7514) );
  NAND2_X1 U9232 ( .A1(n7655), .A2(n7509), .ZN(n7511) );
  MUX2_X1 U9233 ( .A(n7511), .B(n7510), .S(n7519), .Z(n7513) );
  INV_X1 U9234 ( .A(n7512), .ZN(n7516) );
  AOI21_X1 U9235 ( .B1(n7514), .B2(n7513), .A(n7954), .ZN(n7518) );
  MUX2_X1 U9236 ( .A(n7516), .B(n7515), .S(n7519), .Z(n7517) );
  OR3_X1 U9237 ( .A1(n7518), .A2(n7944), .A3(n7517), .ZN(n7523) );
  NAND2_X1 U9238 ( .A1(n8213), .A2(n7732), .ZN(n7520) );
  MUX2_X1 U9239 ( .A(n7521), .B(n7520), .S(n7519), .Z(n7522) );
  MUX2_X1 U9240 ( .A(n7524), .B(n7528), .S(n7535), .Z(n7527) );
  AND2_X1 U9241 ( .A1(n9368), .A2(n7739), .ZN(n7581) );
  INV_X1 U9242 ( .A(n7581), .ZN(n7529) );
  INV_X1 U9243 ( .A(n7739), .ZN(n7530) );
  NAND2_X1 U9244 ( .A1(n7531), .A2(n7530), .ZN(n7533) );
  INV_X1 U9245 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8289) );
  INV_X1 U9246 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7538) );
  MUX2_X1 U9247 ( .A(n8289), .B(n7538), .S(n8613), .Z(n7539) );
  XNOR2_X1 U9248 ( .A(n7539), .B(SI_31_), .ZN(n7540) );
  XNOR2_X1 U9249 ( .A(n7541), .B(n7540), .ZN(n8614) );
  NAND2_X1 U9250 ( .A1(n8614), .A2(n7542), .ZN(n7545) );
  OR2_X1 U9251 ( .A1(n7543), .A2(n8289), .ZN(n7544) );
  OR2_X1 U9252 ( .A1(n8203), .A2(n7551), .ZN(n7550) );
  NAND2_X1 U9253 ( .A1(n8203), .A2(n7551), .ZN(n7583) );
  NAND2_X1 U9254 ( .A1(n7546), .A2(n7586), .ZN(n7591) );
  INV_X1 U9255 ( .A(n7582), .ZN(n7547) );
  OAI22_X1 U9256 ( .A1(n7548), .A2(n7547), .B1(n9368), .B2(n8203), .ZN(n7553)
         );
  NAND2_X1 U9257 ( .A1(n7550), .A2(n7549), .ZN(n7554) );
  OAI21_X1 U9258 ( .B1(n7581), .B2(n7551), .A(n8203), .ZN(n7552) );
  OAI21_X1 U9259 ( .B1(n7553), .B2(n7554), .A(n7552), .ZN(n7589) );
  INV_X1 U9260 ( .A(n7554), .ZN(n7585) );
  INV_X1 U9261 ( .A(n7933), .ZN(n7935) );
  INV_X1 U9262 ( .A(n8005), .ZN(n8000) );
  INV_X1 U9263 ( .A(n8025), .ZN(n8030) );
  INV_X1 U9264 ( .A(n7557), .ZN(n7558) );
  NAND3_X1 U9265 ( .A1(n6724), .A2(n7560), .A3(n8122), .ZN(n7563) );
  NOR4_X1 U9266 ( .A1(n7563), .A2(n7562), .A3(n7561), .A4(n8199), .ZN(n7567)
         );
  NAND4_X1 U9267 ( .A1(n7567), .A2(n7566), .A3(n7565), .A4(n7564), .ZN(n7571)
         );
  NOR4_X1 U9268 ( .A1(n7571), .A2(n7570), .A3(n7569), .A4(n7568), .ZN(n7572)
         );
  NAND4_X1 U9269 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n7576)
         );
  NOR4_X1 U9270 ( .A1(n8058), .A2(n8071), .A3(n8093), .A4(n7576), .ZN(n7577)
         );
  NAND4_X1 U9271 ( .A1(n8030), .A2(n8036), .A3(n4308), .A4(n7577), .ZN(n7578)
         );
  NOR4_X1 U9272 ( .A1(n7990), .A2(n8000), .A3(n8017), .A4(n7578), .ZN(n7579)
         );
  NAND4_X1 U9273 ( .A1(n7952), .A2(n7985), .A3(n7579), .A4(n7972), .ZN(n7580)
         );
  NOR4_X1 U9274 ( .A1(n7581), .A2(n7944), .A3(n7935), .A4(n7580), .ZN(n7584)
         );
  NAND2_X1 U9275 ( .A1(n7591), .A2(n7590), .ZN(n7592) );
  XNOR2_X1 U9276 ( .A(n7592), .B(n7918), .ZN(n7599) );
  NAND3_X1 U9277 ( .A1(n7594), .A2(n7593), .A3(n6156), .ZN(n7595) );
  OAI211_X1 U9278 ( .C1(n7596), .C2(n7598), .A(n7595), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7597) );
  OAI21_X1 U9279 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(P2_U3296) );
  INV_X1 U9280 ( .A(n7600), .ZN(n8296) );
  OAI222_X1 U9281 ( .A1(n9308), .A2(n7601), .B1(n7231), .B2(n8296), .C1(n5640), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U9282 ( .A1(n7604), .A2(n7603), .ZN(n7673) );
  OAI21_X1 U9283 ( .B1(n7604), .B2(n7603), .A(n7673), .ZN(n7605) );
  NOR2_X1 U9284 ( .A1(n7605), .A2(n7980), .ZN(n7676) );
  AOI21_X1 U9285 ( .B1(n7980), .B2(n7605), .A(n7676), .ZN(n7610) );
  AOI22_X1 U9286 ( .A1(n7729), .A2(n7741), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7607) );
  NAND2_X1 U9287 ( .A1(n7734), .A2(n7996), .ZN(n7606) );
  OAI211_X1 U9288 ( .C1(n7993), .C2(n7731), .A(n7607), .B(n7606), .ZN(n7608)
         );
  AOI21_X1 U9289 ( .B1(n7997), .B2(n7705), .A(n7608), .ZN(n7609) );
  OAI21_X1 U9290 ( .B1(n7610), .B2(n7707), .A(n7609), .ZN(P2_U3156) );
  INV_X1 U9291 ( .A(n8249), .ZN(n7618) );
  AOI21_X1 U9292 ( .B1(n7612), .B2(n7611), .A(n7707), .ZN(n7613) );
  NAND2_X1 U9293 ( .A1(n7613), .A2(n7691), .ZN(n7617) );
  NAND2_X1 U9294 ( .A1(n7729), .A2(n8062), .ZN(n7614) );
  NAND2_X1 U9295 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7911) );
  OAI211_X1 U9296 ( .C1(n8042), .C2(n7731), .A(n7614), .B(n7911), .ZN(n7615)
         );
  AOI21_X1 U9297 ( .B1(n8047), .B2(n7734), .A(n7615), .ZN(n7616) );
  OAI211_X1 U9298 ( .C1(n7618), .C2(n7737), .A(n7617), .B(n7616), .ZN(P2_U3159) );
  INV_X1 U9299 ( .A(n7619), .ZN(n7621) );
  AOI21_X1 U9300 ( .B1(n7621), .B2(n7956), .A(n7620), .ZN(n7624) );
  XOR2_X1 U9301 ( .A(n7622), .B(n7933), .Z(n7623) );
  XNOR2_X1 U9302 ( .A(n7624), .B(n7623), .ZN(n7629) );
  AOI22_X1 U9303 ( .A1(n7956), .A2(n7729), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7626) );
  NAND2_X1 U9304 ( .A1(n7940), .A2(n7734), .ZN(n7625) );
  OAI211_X1 U9305 ( .C1(n7740), .C2(n7731), .A(n7626), .B(n7625), .ZN(n7627)
         );
  AOI21_X1 U9306 ( .B1(n8207), .B2(n7705), .A(n7627), .ZN(n7628) );
  OAI21_X1 U9307 ( .B1(n7629), .B2(n7707), .A(n7628), .ZN(P2_U3160) );
  NOR3_X1 U9308 ( .A1(n4374), .A2(n4601), .A3(n7631), .ZN(n7634) );
  INV_X1 U9309 ( .A(n7632), .ZN(n7633) );
  OAI21_X1 U9310 ( .B1(n7634), .B2(n7633), .A(n7726), .ZN(n7638) );
  AOI22_X1 U9311 ( .A1(n7729), .A2(n7742), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7635) );
  OAI21_X1 U9312 ( .B1(n8016), .B2(n7731), .A(n7635), .ZN(n7636) );
  AOI21_X1 U9313 ( .B1(n8019), .B2(n7734), .A(n7636), .ZN(n7637) );
  OAI211_X1 U9314 ( .C1(n7639), .C2(n7737), .A(n7638), .B(n7637), .ZN(P2_U3163) );
  AOI21_X1 U9315 ( .B1(n7729), .B2(n7745), .A(n7640), .ZN(n7643) );
  NAND2_X1 U9316 ( .A1(n7734), .A2(n7641), .ZN(n7642) );
  OAI211_X1 U9317 ( .C1(n7644), .C2(n7731), .A(n7643), .B(n7642), .ZN(n7652)
         );
  OAI21_X1 U9318 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7649) );
  XNOR2_X1 U9319 ( .A(n7649), .B(n7648), .ZN(n7650) );
  NOR2_X1 U9320 ( .A1(n7650), .A2(n7707), .ZN(n7651) );
  AOI211_X1 U9321 ( .C1(n7653), .C2(n7705), .A(n7652), .B(n7651), .ZN(n7654)
         );
  INV_X1 U9322 ( .A(n7654), .ZN(P2_U3164) );
  INV_X1 U9323 ( .A(n7655), .ZN(n8152) );
  AND3_X1 U9324 ( .A1(n7677), .A2(n7657), .A3(n7656), .ZN(n7658) );
  OAI21_X1 U9325 ( .B1(n7725), .B2(n7658), .A(n7726), .ZN(n7662) );
  AOI22_X1 U9326 ( .A1(n7963), .A2(n7680), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7659) );
  OAI21_X1 U9327 ( .B1(n7993), .B2(n7694), .A(n7659), .ZN(n7660) );
  AOI21_X1 U9328 ( .B1(n7966), .B2(n7734), .A(n7660), .ZN(n7661) );
  OAI211_X1 U9329 ( .C1(n8152), .C2(n7737), .A(n7662), .B(n7661), .ZN(P2_U3165) );
  INV_X1 U9330 ( .A(n8261), .ZN(n7672) );
  OAI21_X1 U9331 ( .B1(n7664), .B2(n7663), .A(n7709), .ZN(n7665) );
  NAND2_X1 U9332 ( .A1(n7665), .A2(n7726), .ZN(n7671) );
  INV_X1 U9333 ( .A(n7666), .ZN(n8065) );
  AND2_X1 U9334 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7859) );
  AOI21_X1 U9335 ( .B1(n7680), .B2(n8062), .A(n7859), .ZN(n7667) );
  OAI21_X1 U9336 ( .B1(n7668), .B2(n7694), .A(n7667), .ZN(n7669) );
  AOI21_X1 U9337 ( .B1(n8065), .B2(n7734), .A(n7669), .ZN(n7670) );
  OAI211_X1 U9338 ( .C1(n7672), .C2(n7737), .A(n7671), .B(n7670), .ZN(P2_U3168) );
  INV_X1 U9339 ( .A(n7673), .ZN(n7674) );
  NOR3_X1 U9340 ( .A1(n7676), .A2(n7675), .A3(n7674), .ZN(n7679) );
  INV_X1 U9341 ( .A(n7677), .ZN(n7678) );
  OAI21_X1 U9342 ( .B1(n7679), .B2(n7678), .A(n7726), .ZN(n7684) );
  AOI22_X1 U9343 ( .A1(n7979), .A2(n7680), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7681) );
  OAI21_X1 U9344 ( .B1(n8003), .B2(n7694), .A(n7681), .ZN(n7682) );
  AOI21_X1 U9345 ( .B1(n7982), .B2(n7734), .A(n7682), .ZN(n7683) );
  OAI211_X1 U9346 ( .C1(n7685), .C2(n7737), .A(n7684), .B(n7683), .ZN(P2_U3169) );
  INV_X1 U9347 ( .A(n7687), .ZN(n7690) );
  INV_X1 U9348 ( .A(n7688), .ZN(n7689) );
  AOI21_X1 U9349 ( .B1(n7691), .B2(n7690), .A(n7689), .ZN(n7692) );
  OAI21_X1 U9350 ( .B1(n4374), .B2(n7692), .A(n7726), .ZN(n7698) );
  OAI22_X1 U9351 ( .A1(n7731), .A2(n8004), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7693), .ZN(n7696) );
  NOR2_X1 U9352 ( .A1(n7694), .A2(n7717), .ZN(n7695) );
  AOI211_X1 U9353 ( .C1(n8031), .C2(n7734), .A(n7696), .B(n7695), .ZN(n7697)
         );
  OAI211_X1 U9354 ( .C1(n8246), .C2(n7737), .A(n7698), .B(n7697), .ZN(P2_U3173) );
  INV_X1 U9355 ( .A(n7699), .ZN(n7700) );
  AOI21_X1 U9356 ( .B1(n7741), .B2(n7701), .A(n7700), .ZN(n7708) );
  AOI22_X1 U9357 ( .A1(n7729), .A2(n8027), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7703) );
  NAND2_X1 U9358 ( .A1(n7734), .A2(n8009), .ZN(n7702) );
  OAI211_X1 U9359 ( .C1(n8003), .C2(n7731), .A(n7703), .B(n7702), .ZN(n7704)
         );
  AOI21_X1 U9360 ( .B1(n8159), .B2(n7705), .A(n7704), .ZN(n7706) );
  OAI21_X1 U9361 ( .B1(n7708), .B2(n7707), .A(n7706), .ZN(P2_U3175) );
  INV_X1 U9362 ( .A(n8255), .ZN(n7721) );
  INV_X1 U9363 ( .A(n7709), .ZN(n7712) );
  NOR3_X1 U9364 ( .A1(n7712), .A2(n4583), .A3(n7711), .ZN(n7715) );
  INV_X1 U9365 ( .A(n7713), .ZN(n7714) );
  OAI21_X1 U9366 ( .B1(n7715), .B2(n7714), .A(n7726), .ZN(n7720) );
  NAND2_X1 U9367 ( .A1(n7729), .A2(n8077), .ZN(n7716) );
  NAND2_X1 U9368 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7880) );
  OAI211_X1 U9369 ( .C1(n7717), .C2(n7731), .A(n7716), .B(n7880), .ZN(n7718)
         );
  AOI21_X1 U9370 ( .B1(n8055), .B2(n7734), .A(n7718), .ZN(n7719) );
  OAI211_X1 U9371 ( .C1(n7721), .C2(n7737), .A(n7720), .B(n7719), .ZN(P2_U3178) );
  INV_X1 U9372 ( .A(n7722), .ZN(n7728) );
  NOR3_X1 U9373 ( .A1(n7725), .A2(n7724), .A3(n7723), .ZN(n7727) );
  OAI21_X1 U9374 ( .B1(n7728), .B2(n7727), .A(n7726), .ZN(n7736) );
  AOI22_X1 U9375 ( .A1(n7979), .A2(n7729), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7730) );
  OAI21_X1 U9376 ( .B1(n7732), .B2(n7731), .A(n7730), .ZN(n7733) );
  AOI21_X1 U9377 ( .B1(n7959), .B2(n7734), .A(n7733), .ZN(n7735) );
  OAI211_X1 U9378 ( .C1(n7738), .C2(n7737), .A(n7736), .B(n7735), .ZN(P2_U3180) );
  MUX2_X1 U9379 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n7739), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U9380 ( .A(n7740), .ZN(n7937) );
  MUX2_X1 U9381 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n7937), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9382 ( .A(n7946), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7878), .Z(
        P2_U3519) );
  MUX2_X1 U9383 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n7956), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9384 ( .A(n7963), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7878), .Z(
        P2_U3517) );
  MUX2_X1 U9385 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n7979), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9386 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n7964), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9387 ( .A(n7980), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7878), .Z(
        P2_U3514) );
  MUX2_X1 U9388 ( .A(n7741), .B(P2_DATAO_REG_22__SCAN_IN), .S(n7878), .Z(
        P2_U3513) );
  MUX2_X1 U9389 ( .A(n8027), .B(P2_DATAO_REG_21__SCAN_IN), .S(n7878), .Z(
        P2_U3512) );
  MUX2_X1 U9390 ( .A(n7742), .B(P2_DATAO_REG_20__SCAN_IN), .S(n7878), .Z(
        P2_U3511) );
  MUX2_X1 U9391 ( .A(n8052), .B(P2_DATAO_REG_19__SCAN_IN), .S(n7878), .Z(
        P2_U3510) );
  MUX2_X1 U9392 ( .A(n8062), .B(P2_DATAO_REG_18__SCAN_IN), .S(n7878), .Z(
        P2_U3509) );
  MUX2_X1 U9393 ( .A(n8077), .B(P2_DATAO_REG_17__SCAN_IN), .S(n7878), .Z(
        P2_U3508) );
  MUX2_X1 U9394 ( .A(n8098), .B(P2_DATAO_REG_16__SCAN_IN), .S(n7878), .Z(
        P2_U3507) );
  MUX2_X1 U9395 ( .A(n8076), .B(P2_DATAO_REG_15__SCAN_IN), .S(n7878), .Z(
        P2_U3506) );
  MUX2_X1 U9396 ( .A(n8097), .B(P2_DATAO_REG_14__SCAN_IN), .S(n7878), .Z(
        P2_U3505) );
  MUX2_X1 U9397 ( .A(n7743), .B(P2_DATAO_REG_13__SCAN_IN), .S(n7878), .Z(
        P2_U3504) );
  MUX2_X1 U9398 ( .A(n7744), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7878), .Z(
        P2_U3503) );
  MUX2_X1 U9399 ( .A(n7745), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7878), .Z(
        P2_U3502) );
  MUX2_X1 U9400 ( .A(n7746), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7878), .Z(
        P2_U3501) );
  MUX2_X1 U9401 ( .A(n7747), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7878), .Z(
        P2_U3500) );
  MUX2_X1 U9402 ( .A(n7748), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7878), .Z(
        P2_U3499) );
  MUX2_X1 U9403 ( .A(n7749), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7878), .Z(
        P2_U3498) );
  MUX2_X1 U9404 ( .A(n7750), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7878), .Z(
        P2_U3497) );
  MUX2_X1 U9405 ( .A(n7751), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7878), .Z(
        P2_U3496) );
  MUX2_X1 U9406 ( .A(n4596), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7878), .Z(
        P2_U3495) );
  MUX2_X1 U9407 ( .A(n7752), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7878), .Z(
        P2_U3494) );
  MUX2_X1 U9408 ( .A(n4851), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7878), .Z(
        P2_U3492) );
  XNOR2_X1 U9409 ( .A(n7788), .B(n7789), .ZN(n7754) );
  AOI21_X1 U9410 ( .B1(n7755), .B2(n7754), .A(n7790), .ZN(n7772) );
  AOI21_X1 U9411 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7760) );
  MUX2_X1 U9412 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6156), .Z(n7778) );
  XNOR2_X1 U9413 ( .A(n7778), .B(n7789), .ZN(n7759) );
  NAND2_X1 U9414 ( .A1(n7760), .A2(n7759), .ZN(n7780) );
  OAI21_X1 U9415 ( .B1(n7760), .B2(n7759), .A(n7780), .ZN(n7761) );
  NAND2_X1 U9416 ( .A1(n7761), .A2(n9774), .ZN(n7771) );
  AOI21_X1 U9417 ( .B1(n7765), .B2(n7764), .A(n7774), .ZN(n7768) );
  NAND2_X1 U9418 ( .A1(n7915), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7767) );
  OAI211_X1 U9419 ( .C1(n9769), .C2(n7768), .A(n7767), .B(n7766), .ZN(n7769)
         );
  AOI21_X1 U9420 ( .B1(n7789), .B2(n9767), .A(n7769), .ZN(n7770) );
  OAI211_X1 U9421 ( .C1(n7772), .C2(n9762), .A(n7771), .B(n7770), .ZN(P2_U3195) );
  NOR2_X1 U9422 ( .A1(n7789), .A2(n7773), .ZN(n7775) );
  XNOR2_X1 U9423 ( .A(n7797), .B(n8191), .ZN(n7776) );
  NOR2_X1 U9424 ( .A1(n7777), .A2(n7776), .ZN(n7803) );
  AOI21_X1 U9425 ( .B1(n7777), .B2(n7776), .A(n7803), .ZN(n7799) );
  INV_X1 U9426 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7787) );
  MUX2_X1 U9427 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6156), .Z(n7806) );
  XNOR2_X1 U9428 ( .A(n7806), .B(n7797), .ZN(n7783) );
  INV_X1 U9429 ( .A(n7778), .ZN(n7779) );
  NAND2_X1 U9430 ( .A1(n7789), .A2(n7779), .ZN(n7781) );
  NAND2_X1 U9431 ( .A1(n7781), .A2(n7780), .ZN(n7782) );
  NAND2_X1 U9432 ( .A1(n7783), .A2(n7782), .ZN(n7807) );
  OAI21_X1 U9433 ( .B1(n7783), .B2(n7782), .A(n7807), .ZN(n7784) );
  NAND2_X1 U9434 ( .A1(n9774), .A2(n7784), .ZN(n7786) );
  OAI211_X1 U9435 ( .C1(n9779), .C2(n7787), .A(n7786), .B(n7785), .ZN(n7796)
         );
  NOR2_X1 U9436 ( .A1(n7789), .A2(n7788), .ZN(n7791) );
  AOI22_X1 U9437 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7797), .B1(n7805), .B2(
        n7792), .ZN(n7793) );
  AOI21_X1 U9438 ( .B1(n4385), .B2(n7793), .A(n7800), .ZN(n7794) );
  NOR2_X1 U9439 ( .A1(n7794), .A2(n9762), .ZN(n7795) );
  AOI211_X1 U9440 ( .C1(n9767), .C2(n7797), .A(n7796), .B(n7795), .ZN(n7798)
         );
  OAI21_X1 U9441 ( .B1(n7799), .B2(n9769), .A(n7798), .ZN(P2_U3196) );
  XNOR2_X1 U9442 ( .A(n7834), .B(n7835), .ZN(n7801) );
  AOI21_X1 U9443 ( .B1(n7802), .B2(n7801), .A(n7837), .ZN(n7818) );
  AOI21_X1 U9444 ( .B1(n7804), .B2(n8184), .A(n7820), .ZN(n7815) );
  NAND2_X1 U9445 ( .A1(n7915), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7814) );
  MUX2_X1 U9446 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6156), .Z(n7824) );
  XNOR2_X1 U9447 ( .A(n7835), .B(n7824), .ZN(n7810) );
  OR2_X1 U9448 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  NAND2_X1 U9449 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U9450 ( .A1(n7810), .A2(n7809), .ZN(n7826) );
  OAI21_X1 U9451 ( .B1(n7810), .B2(n7809), .A(n7826), .ZN(n7812) );
  AOI21_X1 U9452 ( .B1(n9774), .B2(n7812), .A(n7811), .ZN(n7813) );
  OAI211_X1 U9453 ( .C1(n9769), .C2(n7815), .A(n7814), .B(n7813), .ZN(n7816)
         );
  AOI21_X1 U9454 ( .B1(n7835), .B2(n9767), .A(n7816), .ZN(n7817) );
  OAI21_X1 U9455 ( .B1(n7818), .B2(n9762), .A(n7817), .ZN(P2_U3197) );
  NOR2_X1 U9456 ( .A1(n7835), .A2(n7819), .ZN(n7821) );
  XNOR2_X1 U9457 ( .A(n7853), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7822) );
  NOR2_X1 U9458 ( .A1(n7823), .A2(n7822), .ZN(n7850) );
  AOI21_X1 U9459 ( .B1(n7823), .B2(n7822), .A(n7850), .ZN(n7845) );
  INV_X1 U9460 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7833) );
  MUX2_X1 U9461 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6156), .Z(n7854) );
  XNOR2_X1 U9462 ( .A(n7854), .B(n7843), .ZN(n7829) );
  INV_X1 U9463 ( .A(n7824), .ZN(n7825) );
  NAND2_X1 U9464 ( .A1(n7835), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U9465 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  NAND2_X1 U9466 ( .A1(n7829), .A2(n7828), .ZN(n7855) );
  OAI21_X1 U9467 ( .B1(n7829), .B2(n7828), .A(n7855), .ZN(n7830) );
  NAND2_X1 U9468 ( .A1(n9774), .A2(n7830), .ZN(n7832) );
  OAI211_X1 U9469 ( .C1(n9779), .C2(n7833), .A(n7832), .B(n7831), .ZN(n7842)
         );
  NOR2_X1 U9470 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NAND2_X1 U9471 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7853), .ZN(n7846) );
  OAI21_X1 U9472 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n7853), .A(n7846), .ZN(
        n7838) );
  NOR2_X1 U9473 ( .A1(n7839), .A2(n7838), .ZN(n7848) );
  AOI21_X1 U9474 ( .B1(n7839), .B2(n7838), .A(n7848), .ZN(n7840) );
  NOR2_X1 U9475 ( .A1(n7840), .A2(n9762), .ZN(n7841) );
  AOI211_X1 U9476 ( .C1(n9767), .C2(n7843), .A(n7842), .B(n7841), .ZN(n7844)
         );
  OAI21_X1 U9477 ( .B1(n7845), .B2(n9769), .A(n7844), .ZN(P2_U3198) );
  INV_X1 U9478 ( .A(n7846), .ZN(n7847) );
  AOI21_X1 U9479 ( .B1(n8064), .B2(n7849), .A(n7886), .ZN(n7866) );
  XNOR2_X1 U9480 ( .A(n7884), .B(n7867), .ZN(n7851) );
  AOI21_X1 U9481 ( .B1(n7851), .B2(n9981), .A(n7869), .ZN(n7863) );
  NAND2_X1 U9482 ( .A1(n7915), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7862) );
  MUX2_X1 U9483 ( .A(n8064), .B(n9981), .S(n6156), .Z(n7874) );
  XNOR2_X1 U9484 ( .A(n7874), .B(n7852), .ZN(n7858) );
  OR2_X1 U9485 ( .A1(n7854), .A2(n7853), .ZN(n7856) );
  NAND2_X1 U9486 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND2_X1 U9487 ( .A1(n7858), .A2(n7857), .ZN(n7872) );
  OAI21_X1 U9488 ( .B1(n7858), .B2(n7857), .A(n7872), .ZN(n7860) );
  AOI21_X1 U9489 ( .B1(n9774), .B2(n7860), .A(n7859), .ZN(n7861) );
  OAI211_X1 U9490 ( .C1(n9769), .C2(n7863), .A(n7862), .B(n7861), .ZN(n7864)
         );
  AOI21_X1 U9491 ( .B1(n7884), .B2(n9767), .A(n7864), .ZN(n7865) );
  OAI21_X1 U9492 ( .B1(n7866), .B2(n9762), .A(n7865), .ZN(P2_U3199) );
  NOR2_X1 U9493 ( .A1(n7884), .A2(n7867), .ZN(n7868) );
  NAND2_X1 U9494 ( .A1(n7887), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7893) );
  OAI21_X1 U9495 ( .B1(n7887), .B2(P2_REG1_REG_18__SCAN_IN), .A(n7893), .ZN(
        n7870) );
  AOI21_X1 U9496 ( .B1(n7871), .B2(n7870), .A(n7895), .ZN(n7892) );
  INV_X1 U9497 ( .A(n7872), .ZN(n7873) );
  MUX2_X1 U9498 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6156), .Z(n7875) );
  NOR2_X1 U9499 ( .A1(n7876), .A2(n7875), .ZN(n7902) );
  INV_X1 U9500 ( .A(n7902), .ZN(n7877) );
  NAND2_X1 U9501 ( .A1(n7876), .A2(n7875), .ZN(n7903) );
  NAND2_X1 U9502 ( .A1(n7877), .A2(n7903), .ZN(n7879) );
  OAI21_X1 U9503 ( .B1(n7878), .B2(n7879), .A(n7917), .ZN(n7891) );
  NAND3_X1 U9504 ( .A1(n9774), .A2(n7887), .A3(n7879), .ZN(n7881) );
  OAI211_X1 U9505 ( .C1(n9779), .C2(n9859), .A(n7881), .B(n7880), .ZN(n7890)
         );
  NOR2_X1 U9506 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U9507 ( .A1(n7887), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7898) );
  OAI21_X1 U9508 ( .B1(n7887), .B2(P2_REG2_REG_18__SCAN_IN), .A(n7898), .ZN(
        n7888) );
  NOR2_X1 U9509 ( .A1(n7889), .A2(n7888), .ZN(n7900) );
  INV_X1 U9510 ( .A(n7893), .ZN(n7894) );
  NOR2_X1 U9511 ( .A1(n7895), .A2(n7894), .ZN(n7897) );
  XNOR2_X1 U9512 ( .A(n7896), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7908) );
  XNOR2_X1 U9513 ( .A(n7897), .B(n7908), .ZN(n7923) );
  INV_X1 U9514 ( .A(n7898), .ZN(n7899) );
  NOR2_X1 U9515 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  XNOR2_X1 U9516 ( .A(n7918), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n7905) );
  XNOR2_X1 U9517 ( .A(n7901), .B(n7905), .ZN(n7921) );
  AOI21_X1 U9518 ( .B1(n7904), .B2(n7903), .A(n7902), .ZN(n7910) );
  INV_X1 U9519 ( .A(n7905), .ZN(n7907) );
  MUX2_X1 U9520 ( .A(n7908), .B(n7907), .S(n7906), .Z(n7909) );
  XNOR2_X1 U9521 ( .A(n7910), .B(n7909), .ZN(n7912) );
  OAI21_X1 U9522 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7914) );
  AOI21_X1 U9523 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n7915), .A(n7914), .ZN(
        n7916) );
  OAI21_X1 U9524 ( .B1(n7918), .B2(n7917), .A(n7916), .ZN(n7919) );
  OAI21_X1 U9525 ( .B1(n7923), .B2(n9769), .A(n7922), .ZN(P2_U3201) );
  INV_X1 U9526 ( .A(n8203), .ZN(n8138) );
  AOI21_X1 U9527 ( .B1(n8080), .B2(P2_REG2_REG_31__SCAN_IN), .A(n7924), .ZN(
        n7925) );
  OAI21_X1 U9528 ( .B1(n8138), .B2(n8092), .A(n7925), .ZN(P2_U3202) );
  AOI22_X1 U9529 ( .A1(n7926), .A2(n8131), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8080), .ZN(n7927) );
  OAI21_X1 U9530 ( .B1(n7928), .B2(n8092), .A(n7927), .ZN(n7929) );
  AOI21_X1 U9531 ( .B1(n7931), .B2(n7930), .A(n7929), .ZN(n7932) );
  OAI21_X1 U9532 ( .B1(n4371), .B2(n8080), .A(n7932), .ZN(P2_U3204) );
  XNOR2_X1 U9533 ( .A(n7934), .B(n7933), .ZN(n8210) );
  XNOR2_X1 U9534 ( .A(n7936), .B(n7935), .ZN(n7938) );
  AOI222_X1 U9535 ( .A1(n6238), .A2(n7938), .B1(n7937), .B2(n8099), .C1(n7956), 
        .C2(n8096), .ZN(n8206) );
  INV_X1 U9536 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7939) );
  MUX2_X1 U9537 ( .A(n8206), .B(n7939), .S(n8080), .Z(n7942) );
  AOI22_X1 U9538 ( .A1(n8207), .A2(n8085), .B1(n8131), .B2(n7940), .ZN(n7941)
         );
  OAI211_X1 U9539 ( .C1(n8210), .C2(n8088), .A(n7942), .B(n7941), .ZN(P2_U3205) );
  XNOR2_X1 U9540 ( .A(n7943), .B(n7944), .ZN(n8216) );
  XOR2_X1 U9541 ( .A(n7945), .B(n7944), .Z(n7947) );
  AOI222_X1 U9542 ( .A1(n6238), .A2(n7947), .B1(n7946), .B2(n8099), .C1(n7963), 
        .C2(n8096), .ZN(n8211) );
  MUX2_X1 U9543 ( .A(n8211), .B(n7948), .S(n8080), .Z(n7951) );
  AOI22_X1 U9544 ( .A1(n8213), .A2(n8085), .B1(n8131), .B2(n7949), .ZN(n7950)
         );
  OAI211_X1 U9545 ( .C1(n8216), .C2(n8088), .A(n7951), .B(n7950), .ZN(P2_U3206) );
  XNOR2_X1 U9546 ( .A(n7953), .B(n7952), .ZN(n8222) );
  XNOR2_X1 U9547 ( .A(n7955), .B(n7954), .ZN(n7957) );
  AOI222_X1 U9548 ( .A1(n6238), .A2(n7957), .B1(n7956), .B2(n8099), .C1(n7979), 
        .C2(n8096), .ZN(n8217) );
  MUX2_X1 U9549 ( .A(n8217), .B(n7958), .S(n8080), .Z(n7961) );
  AOI22_X1 U9550 ( .A1(n8219), .A2(n8085), .B1(n8131), .B2(n7959), .ZN(n7960)
         );
  OAI211_X1 U9551 ( .C1(n8222), .C2(n8088), .A(n7961), .B(n7960), .ZN(P2_U3207) );
  XNOR2_X1 U9552 ( .A(n7962), .B(n7972), .ZN(n7965) );
  AOI222_X1 U9553 ( .A1(n6238), .A2(n7965), .B1(n7964), .B2(n8096), .C1(n7963), 
        .C2(n8099), .ZN(n8151) );
  INV_X1 U9554 ( .A(n8151), .ZN(n7970) );
  INV_X1 U9555 ( .A(n7966), .ZN(n7967) );
  OAI22_X1 U9556 ( .A1(n8152), .A2(n7968), .B1(n7967), .B2(n8106), .ZN(n7969)
         );
  OAI21_X1 U9557 ( .B1(n7970), .B2(n7969), .A(n8135), .ZN(n7976) );
  INV_X1 U9558 ( .A(n7971), .ZN(n7974) );
  INV_X1 U9559 ( .A(n7972), .ZN(n7973) );
  NAND2_X1 U9560 ( .A1(n7974), .A2(n7973), .ZN(n8149) );
  NAND3_X1 U9561 ( .A1(n8149), .A2(n8112), .A3(n8148), .ZN(n7975) );
  OAI211_X1 U9562 ( .C1(n8135), .C2(n7977), .A(n7976), .B(n7975), .ZN(P2_U3208) );
  XNOR2_X1 U9563 ( .A(n7978), .B(n7985), .ZN(n7981) );
  AOI222_X1 U9564 ( .A1(n6238), .A2(n7981), .B1(n7980), .B2(n8096), .C1(n7979), 
        .C2(n8099), .ZN(n8224) );
  AOI22_X1 U9565 ( .A1(n8226), .A2(n8111), .B1(n8131), .B2(n7982), .ZN(n7983)
         );
  AOI21_X1 U9566 ( .B1(n8224), .B2(n7983), .A(n8080), .ZN(n7988) );
  XOR2_X1 U9567 ( .A(n7985), .B(n7984), .Z(n8229) );
  OAI22_X1 U9568 ( .A1(n8229), .A2(n8088), .B1(n7986), .B2(n8135), .ZN(n7987)
         );
  OR2_X1 U9569 ( .A1(n7988), .A2(n7987), .ZN(P2_U3209) );
  XOR2_X1 U9570 ( .A(n7989), .B(n7990), .Z(n8232) );
  XOR2_X1 U9571 ( .A(n7991), .B(n7990), .Z(n7992) );
  OAI222_X1 U9572 ( .A1(n8120), .A2(n8016), .B1(n8118), .B2(n7993), .C1(n8123), 
        .C2(n7992), .ZN(n8230) );
  INV_X1 U9573 ( .A(n8230), .ZN(n7994) );
  MUX2_X1 U9574 ( .A(n7995), .B(n7994), .S(n8135), .Z(n7999) );
  AOI22_X1 U9575 ( .A1(n7997), .A2(n8085), .B1(n8131), .B2(n7996), .ZN(n7998)
         );
  OAI211_X1 U9576 ( .C1(n8232), .C2(n8088), .A(n7999), .B(n7998), .ZN(P2_U3210) );
  XNOR2_X1 U9577 ( .A(n8001), .B(n8000), .ZN(n8002) );
  OAI222_X1 U9578 ( .A1(n8120), .A2(n8004), .B1(n8118), .B2(n8003), .C1(n8002), 
        .C2(n8123), .ZN(n8158) );
  OR2_X1 U9579 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  NAND2_X1 U9580 ( .A1(n8008), .A2(n8007), .ZN(n8238) );
  AOI22_X1 U9581 ( .A1(n8080), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8131), .B2(
        n8009), .ZN(n8011) );
  NAND2_X1 U9582 ( .A1(n8159), .A2(n8085), .ZN(n8010) );
  OAI211_X1 U9583 ( .C1(n8238), .C2(n8088), .A(n8011), .B(n8010), .ZN(n8012)
         );
  AOI21_X1 U9584 ( .B1(n8158), .B2(n8135), .A(n8012), .ZN(n8013) );
  INV_X1 U9585 ( .A(n8013), .ZN(P2_U3211) );
  XOR2_X1 U9586 ( .A(n8014), .B(n8017), .Z(n8015) );
  OAI222_X1 U9587 ( .A1(n8120), .A2(n8042), .B1(n8118), .B2(n8016), .C1(n8123), 
        .C2(n8015), .ZN(n8162) );
  XNOR2_X1 U9588 ( .A(n8018), .B(n8017), .ZN(n8242) );
  AOI22_X1 U9589 ( .A1(n8080), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8131), .B2(
        n8019), .ZN(n8021) );
  NAND2_X1 U9590 ( .A1(n8163), .A2(n8085), .ZN(n8020) );
  OAI211_X1 U9591 ( .C1(n8242), .C2(n8088), .A(n8021), .B(n8020), .ZN(n8022)
         );
  AOI21_X1 U9592 ( .B1(n8162), .B2(n8135), .A(n8022), .ZN(n8023) );
  INV_X1 U9593 ( .A(n8023), .ZN(P2_U3212) );
  OAI21_X1 U9594 ( .B1(n8026), .B2(n8025), .A(n8024), .ZN(n8028) );
  AOI222_X1 U9595 ( .A1(n6238), .A2(n8028), .B1(n8027), .B2(n8099), .C1(n8052), 
        .C2(n8096), .ZN(n8166) );
  XNOR2_X1 U9596 ( .A(n8029), .B(n8030), .ZN(n8168) );
  AOI22_X1 U9597 ( .A1(n8080), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8131), .B2(
        n8031), .ZN(n8032) );
  OAI21_X1 U9598 ( .B1(n8246), .B2(n8092), .A(n8032), .ZN(n8033) );
  AOI21_X1 U9599 ( .B1(n8168), .B2(n8112), .A(n8033), .ZN(n8034) );
  OAI21_X1 U9600 ( .B1(n8166), .B2(n8080), .A(n8034), .ZN(P2_U3213) );
  XOR2_X1 U9601 ( .A(n8035), .B(n8036), .Z(n8252) );
  NAND2_X1 U9602 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U9603 ( .A1(n8038), .A2(n6238), .ZN(n8040) );
  OR2_X1 U9604 ( .A1(n8040), .A2(n8039), .ZN(n8045) );
  OAI22_X1 U9605 ( .A1(n8042), .A2(n8118), .B1(n8041), .B2(n8120), .ZN(n8043)
         );
  INV_X1 U9606 ( .A(n8043), .ZN(n8044) );
  INV_X1 U9607 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8046) );
  MUX2_X1 U9608 ( .A(n8248), .B(n8046), .S(n8080), .Z(n8049) );
  AOI22_X1 U9609 ( .A1(n8249), .A2(n8085), .B1(n8131), .B2(n8047), .ZN(n8048)
         );
  OAI211_X1 U9610 ( .C1(n8252), .C2(n8088), .A(n8049), .B(n8048), .ZN(P2_U3214) );
  XNOR2_X1 U9611 ( .A(n8050), .B(n4308), .ZN(n8258) );
  XNOR2_X1 U9612 ( .A(n8051), .B(n4308), .ZN(n8053) );
  AOI222_X1 U9613 ( .A1(n6238), .A2(n8053), .B1(n8077), .B2(n8096), .C1(n8052), 
        .C2(n8099), .ZN(n8253) );
  MUX2_X1 U9614 ( .A(n8054), .B(n8253), .S(n8135), .Z(n8057) );
  AOI22_X1 U9615 ( .A1(n8255), .A2(n8085), .B1(n8131), .B2(n8055), .ZN(n8056)
         );
  OAI211_X1 U9616 ( .C1(n8258), .C2(n8088), .A(n8057), .B(n8056), .ZN(P2_U3215) );
  XNOR2_X1 U9617 ( .A(n8059), .B(n8058), .ZN(n8264) );
  XNOR2_X1 U9618 ( .A(n8060), .B(n8061), .ZN(n8063) );
  AOI222_X1 U9619 ( .A1(n6238), .A2(n8063), .B1(n8062), .B2(n8099), .C1(n8098), 
        .C2(n8096), .ZN(n8259) );
  MUX2_X1 U9620 ( .A(n8064), .B(n8259), .S(n8135), .Z(n8067) );
  AOI22_X1 U9621 ( .A1(n8261), .A2(n8085), .B1(n8131), .B2(n8065), .ZN(n8066)
         );
  OAI211_X1 U9622 ( .C1(n8264), .C2(n8088), .A(n8067), .B(n8066), .ZN(P2_U3216) );
  XOR2_X1 U9623 ( .A(n8071), .B(n8068), .Z(n8267) );
  NAND2_X1 U9624 ( .A1(n8069), .A2(n8070), .ZN(n8073) );
  INV_X1 U9625 ( .A(n8071), .ZN(n8072) );
  NAND2_X1 U9626 ( .A1(n8073), .A2(n8072), .ZN(n8075) );
  NAND3_X1 U9627 ( .A1(n8075), .A2(n6238), .A3(n8074), .ZN(n8079) );
  AOI22_X1 U9628 ( .A1(n8077), .A2(n8099), .B1(n8096), .B2(n8076), .ZN(n8078)
         );
  NAND2_X1 U9629 ( .A1(n8079), .A2(n8078), .ZN(n8265) );
  INV_X1 U9630 ( .A(n8265), .ZN(n8082) );
  MUX2_X1 U9631 ( .A(n8082), .B(n8081), .S(n8080), .Z(n8087) );
  INV_X1 U9632 ( .A(n8083), .ZN(n8084) );
  AOI22_X1 U9633 ( .A1(n8179), .A2(n8085), .B1(n8131), .B2(n8084), .ZN(n8086)
         );
  OAI211_X1 U9634 ( .C1(n8267), .C2(n8088), .A(n8087), .B(n8086), .ZN(P2_U3217) );
  XNOR2_X1 U9635 ( .A(n8090), .B(n8089), .ZN(n8183) );
  OAI22_X1 U9636 ( .A1(n8272), .A2(n8092), .B1(n8091), .B2(n8106), .ZN(n8103)
         );
  OAI21_X1 U9637 ( .B1(n8094), .B2(n8093), .A(n8069), .ZN(n8095) );
  NAND2_X1 U9638 ( .A1(n8095), .A2(n6238), .ZN(n8101) );
  AOI22_X1 U9639 ( .A1(n8099), .A2(n8098), .B1(n8097), .B2(n8096), .ZN(n8100)
         );
  NAND2_X1 U9640 ( .A1(n8101), .A2(n8100), .ZN(n8270) );
  MUX2_X1 U9641 ( .A(n8270), .B(P2_REG2_REG_15__SCAN_IN), .S(n8080), .Z(n8102)
         );
  AOI211_X1 U9642 ( .C1(n8183), .C2(n8112), .A(n8103), .B(n8102), .ZN(n8104)
         );
  INV_X1 U9643 ( .A(n8104), .ZN(P2_U3218) );
  NOR2_X1 U9644 ( .A1(n8106), .A2(n8105), .ZN(n8109) );
  INV_X1 U9645 ( .A(n8107), .ZN(n8108) );
  AOI211_X1 U9646 ( .C1(n8111), .C2(n8110), .A(n8109), .B(n8108), .ZN(n8115)
         );
  AOI22_X1 U9647 ( .A1(n8113), .A2(n8112), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8080), .ZN(n8114) );
  OAI21_X1 U9648 ( .B1(n8115), .B2(n8080), .A(n8114), .ZN(P2_U3220) );
  OAI21_X1 U9649 ( .B1(n8116), .B2(n8122), .A(n8117), .ZN(n9790) );
  INV_X1 U9650 ( .A(n9790), .ZN(n8134) );
  OAI22_X1 U9651 ( .A1(n6178), .A2(n8120), .B1(n8119), .B2(n8118), .ZN(n8126)
         );
  NAND3_X1 U9652 ( .A1(n6728), .A2(n8122), .A3(n8121), .ZN(n8124) );
  AOI211_X1 U9653 ( .C1(n8127), .C2(n9790), .A(n8126), .B(n8125), .ZN(n9787)
         );
  AND2_X1 U9654 ( .A1(n8128), .A2(n9836), .ZN(n9789) );
  INV_X1 U9655 ( .A(n8129), .ZN(n8130) );
  AOI22_X1 U9656 ( .A1(n8131), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n9789), .B2(
        n8130), .ZN(n8132) );
  OAI211_X1 U9657 ( .C1(n8134), .C2(n8133), .A(n9787), .B(n8132), .ZN(n8136)
         );
  MUX2_X1 U9658 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8136), .S(n8135), .Z(
        P2_U3231) );
  MUX2_X1 U9659 ( .A(n9369), .B(n6588), .S(n9847), .Z(n8137) );
  OAI21_X1 U9660 ( .B1(n8138), .B2(n8180), .A(n8137), .ZN(P2_U3490) );
  INV_X1 U9661 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8139) );
  MUX2_X1 U9662 ( .A(n8139), .B(n8206), .S(n9849), .Z(n8141) );
  NAND2_X1 U9663 ( .A1(n8207), .A2(n8192), .ZN(n8140) );
  OAI211_X1 U9664 ( .C1(n8210), .C2(n8189), .A(n8141), .B(n8140), .ZN(P2_U3487) );
  INV_X1 U9665 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8142) );
  MUX2_X1 U9666 ( .A(n8142), .B(n8211), .S(n9849), .Z(n8144) );
  NAND2_X1 U9667 ( .A1(n8213), .A2(n8192), .ZN(n8143) );
  OAI211_X1 U9668 ( .C1(n8216), .C2(n8189), .A(n8144), .B(n8143), .ZN(P2_U3486) );
  INV_X1 U9669 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8145) );
  MUX2_X1 U9670 ( .A(n8145), .B(n8217), .S(n9849), .Z(n8147) );
  NAND2_X1 U9671 ( .A1(n8219), .A2(n8192), .ZN(n8146) );
  OAI211_X1 U9672 ( .C1(n8222), .C2(n8189), .A(n8147), .B(n8146), .ZN(P2_U3485) );
  NAND3_X1 U9673 ( .A1(n8149), .A2(n8148), .A3(n9807), .ZN(n8150) );
  OAI211_X1 U9674 ( .C1(n8152), .C2(n9824), .A(n8151), .B(n8150), .ZN(n8223)
         );
  MUX2_X1 U9675 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8223), .S(n9849), .Z(
        P2_U3484) );
  INV_X1 U9676 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8153) );
  MUX2_X1 U9677 ( .A(n8153), .B(n8224), .S(n9849), .Z(n8155) );
  NAND2_X1 U9678 ( .A1(n8226), .A2(n8192), .ZN(n8154) );
  OAI211_X1 U9679 ( .C1(n8189), .C2(n8229), .A(n8155), .B(n8154), .ZN(P2_U3483) );
  MUX2_X1 U9680 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8230), .S(n9849), .Z(n8157)
         );
  OAI22_X1 U9681 ( .A1(n8232), .A2(n8189), .B1(n8231), .B2(n8180), .ZN(n8156)
         );
  OR2_X1 U9682 ( .A1(n8157), .A2(n8156), .ZN(P2_U3482) );
  INV_X1 U9683 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8160) );
  AOI21_X1 U9684 ( .B1(n9836), .B2(n8159), .A(n8158), .ZN(n8235) );
  MUX2_X1 U9685 ( .A(n8160), .B(n8235), .S(n9849), .Z(n8161) );
  OAI21_X1 U9686 ( .B1(n8189), .B2(n8238), .A(n8161), .ZN(P2_U3481) );
  INV_X1 U9687 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8164) );
  AOI21_X1 U9688 ( .B1(n9836), .B2(n8163), .A(n8162), .ZN(n8239) );
  MUX2_X1 U9689 ( .A(n8164), .B(n8239), .S(n9849), .Z(n8165) );
  OAI21_X1 U9690 ( .B1(n8189), .B2(n8242), .A(n8165), .ZN(P2_U3480) );
  INV_X1 U9691 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8169) );
  INV_X1 U9692 ( .A(n8166), .ZN(n8167) );
  AOI21_X1 U9693 ( .B1(n8168), .B2(n9807), .A(n8167), .ZN(n8243) );
  MUX2_X1 U9694 ( .A(n8169), .B(n8243), .S(n9849), .Z(n8170) );
  OAI21_X1 U9695 ( .B1(n8246), .B2(n8180), .A(n8170), .ZN(P2_U3479) );
  INV_X1 U9696 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8171) );
  MUX2_X1 U9697 ( .A(n8248), .B(n8171), .S(n9847), .Z(n8173) );
  NAND2_X1 U9698 ( .A1(n8249), .A2(n8192), .ZN(n8172) );
  OAI211_X1 U9699 ( .C1(n8189), .C2(n8252), .A(n8173), .B(n8172), .ZN(P2_U3478) );
  MUX2_X1 U9700 ( .A(n8174), .B(n8253), .S(n9849), .Z(n8176) );
  NAND2_X1 U9701 ( .A1(n8255), .A2(n8192), .ZN(n8175) );
  OAI211_X1 U9702 ( .C1(n8258), .C2(n8189), .A(n8176), .B(n8175), .ZN(P2_U3477) );
  MUX2_X1 U9703 ( .A(n9981), .B(n8259), .S(n9849), .Z(n8178) );
  NAND2_X1 U9704 ( .A1(n8261), .A2(n8192), .ZN(n8177) );
  OAI211_X1 U9705 ( .C1(n8189), .C2(n8264), .A(n8178), .B(n8177), .ZN(P2_U3476) );
  MUX2_X1 U9706 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8265), .S(n9849), .Z(n8182)
         );
  INV_X1 U9707 ( .A(n8179), .ZN(n8266) );
  OAI22_X1 U9708 ( .A1(n8267), .A2(n8189), .B1(n8266), .B2(n8180), .ZN(n8181)
         );
  OR2_X1 U9709 ( .A1(n8182), .A2(n8181), .ZN(P2_U3475) );
  INV_X1 U9710 ( .A(n8183), .ZN(n8274) );
  INV_X1 U9711 ( .A(n8270), .ZN(n8185) );
  MUX2_X1 U9712 ( .A(n8185), .B(n8184), .S(n9847), .Z(n8188) );
  NAND2_X1 U9713 ( .A1(n8186), .A2(n8192), .ZN(n8187) );
  OAI211_X1 U9714 ( .C1(n8189), .C2(n8274), .A(n8188), .B(n8187), .ZN(P2_U3474) );
  INV_X1 U9715 ( .A(n8190), .ZN(n8277) );
  MUX2_X1 U9716 ( .A(n8191), .B(n8277), .S(n9849), .Z(n8195) );
  AOI22_X1 U9717 ( .A1(n8282), .A2(n8193), .B1(n8192), .B2(n8279), .ZN(n8194)
         );
  NAND2_X1 U9718 ( .A1(n8195), .A2(n8194), .ZN(P2_U3473) );
  NOR2_X1 U9719 ( .A1(n8196), .A2(n9824), .ZN(n8197) );
  NOR2_X1 U9720 ( .A1(n8198), .A2(n8197), .ZN(n8201) );
  OAI21_X1 U9721 ( .B1(n6238), .B2(n9807), .A(n8199), .ZN(n8200) );
  AND2_X1 U9722 ( .A1(n8201), .A2(n8200), .ZN(n9781) );
  INV_X1 U9723 ( .A(n9781), .ZN(n8202) );
  MUX2_X1 U9724 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8202), .S(n9849), .Z(
        P2_U3459) );
  NAND2_X1 U9725 ( .A1(n8203), .A2(n8280), .ZN(n8205) );
  NAND2_X1 U9726 ( .A1(n9886), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U9727 ( .C1(n9886), .C2(n9369), .A(n8205), .B(n8204), .ZN(P2_U3458) );
  MUX2_X1 U9728 ( .A(n9996), .B(n8206), .S(n9884), .Z(n8209) );
  NAND2_X1 U9729 ( .A1(n8207), .A2(n8280), .ZN(n8208) );
  OAI211_X1 U9730 ( .C1(n8210), .C2(n8273), .A(n8209), .B(n8208), .ZN(P2_U3455) );
  INV_X1 U9731 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8212) );
  MUX2_X1 U9732 ( .A(n8212), .B(n8211), .S(n9884), .Z(n8215) );
  NAND2_X1 U9733 ( .A1(n8213), .A2(n8280), .ZN(n8214) );
  OAI211_X1 U9734 ( .C1(n8216), .C2(n8273), .A(n8215), .B(n8214), .ZN(P2_U3454) );
  INV_X1 U9735 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U9736 ( .A(n8218), .B(n8217), .S(n9884), .Z(n8221) );
  NAND2_X1 U9737 ( .A1(n8219), .A2(n8280), .ZN(n8220) );
  OAI211_X1 U9738 ( .C1(n8222), .C2(n8273), .A(n8221), .B(n8220), .ZN(P2_U3453) );
  MUX2_X1 U9739 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8223), .S(n9884), .Z(
        P2_U3452) );
  INV_X1 U9740 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8225) );
  MUX2_X1 U9741 ( .A(n8225), .B(n8224), .S(n9884), .Z(n8228) );
  NAND2_X1 U9742 ( .A1(n8226), .A2(n8280), .ZN(n8227) );
  OAI211_X1 U9743 ( .C1(n8229), .C2(n8273), .A(n8228), .B(n8227), .ZN(P2_U3451) );
  MUX2_X1 U9744 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8230), .S(n9884), .Z(n8234)
         );
  OAI22_X1 U9745 ( .A1(n8232), .A2(n8273), .B1(n8231), .B2(n8271), .ZN(n8233)
         );
  OR2_X1 U9746 ( .A1(n8234), .A2(n8233), .ZN(P2_U3450) );
  INV_X1 U9747 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8236) );
  MUX2_X1 U9748 ( .A(n8236), .B(n8235), .S(n9884), .Z(n8237) );
  OAI21_X1 U9749 ( .B1(n8238), .B2(n8273), .A(n8237), .ZN(P2_U3449) );
  INV_X1 U9750 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8240) );
  MUX2_X1 U9751 ( .A(n8240), .B(n8239), .S(n9884), .Z(n8241) );
  OAI21_X1 U9752 ( .B1(n8242), .B2(n8273), .A(n8241), .ZN(P2_U3448) );
  INV_X1 U9753 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8244) );
  MUX2_X1 U9754 ( .A(n8244), .B(n8243), .S(n9884), .Z(n8245) );
  OAI21_X1 U9755 ( .B1(n8246), .B2(n8271), .A(n8245), .ZN(P2_U3447) );
  INV_X1 U9756 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8247) );
  MUX2_X1 U9757 ( .A(n8248), .B(n8247), .S(n9886), .Z(n8251) );
  NAND2_X1 U9758 ( .A1(n8249), .A2(n8280), .ZN(n8250) );
  OAI211_X1 U9759 ( .C1(n8252), .C2(n8273), .A(n8251), .B(n8250), .ZN(P2_U3446) );
  MUX2_X1 U9760 ( .A(n8254), .B(n8253), .S(n9884), .Z(n8257) );
  NAND2_X1 U9761 ( .A1(n8255), .A2(n8280), .ZN(n8256) );
  OAI211_X1 U9762 ( .C1(n8258), .C2(n8273), .A(n8257), .B(n8256), .ZN(P2_U3444) );
  INV_X1 U9763 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8260) );
  MUX2_X1 U9764 ( .A(n8260), .B(n8259), .S(n9884), .Z(n8263) );
  NAND2_X1 U9765 ( .A1(n8261), .A2(n8280), .ZN(n8262) );
  OAI211_X1 U9766 ( .C1(n8264), .C2(n8273), .A(n8263), .B(n8262), .ZN(P2_U3441) );
  MUX2_X1 U9767 ( .A(n8265), .B(P2_REG0_REG_16__SCAN_IN), .S(n9886), .Z(n8269)
         );
  OAI22_X1 U9768 ( .A1(n8267), .A2(n8273), .B1(n8266), .B2(n8271), .ZN(n8268)
         );
  OR2_X1 U9769 ( .A1(n8269), .A2(n8268), .ZN(P2_U3438) );
  MUX2_X1 U9770 ( .A(n8270), .B(P2_REG0_REG_15__SCAN_IN), .S(n9886), .Z(n8276)
         );
  OAI22_X1 U9771 ( .A1(n8274), .A2(n8273), .B1(n8272), .B2(n8271), .ZN(n8275)
         );
  OR2_X1 U9772 ( .A1(n8276), .A2(n8275), .ZN(P2_U3435) );
  INV_X1 U9773 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8278) );
  MUX2_X1 U9774 ( .A(n8278), .B(n8277), .S(n9884), .Z(n8284) );
  AOI22_X1 U9775 ( .A1(n8282), .A2(n8281), .B1(n8280), .B2(n8279), .ZN(n8283)
         );
  NAND2_X1 U9776 ( .A1(n8284), .A2(n8283), .ZN(P2_U3432) );
  MUX2_X1 U9777 ( .A(P2_D_REG_1__SCAN_IN), .B(n8286), .S(n8285), .Z(P2_U3377)
         );
  INV_X1 U9778 ( .A(n8614), .ZN(n9302) );
  INV_X1 U9779 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8288) );
  NAND3_X1 U9780 ( .A1(n8288), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8290) );
  OAI22_X1 U9781 ( .A1(n8287), .A2(n8290), .B1(n8289), .B2(n8300), .ZN(n8291)
         );
  INV_X1 U9782 ( .A(n8291), .ZN(n8292) );
  OAI21_X1 U9783 ( .B1(n9302), .B2(n8304), .A(n8292), .ZN(P2_U3264) );
  INV_X1 U9784 ( .A(n8609), .ZN(n9304) );
  OAI222_X1 U9785 ( .A1(n8294), .A2(n8293), .B1(n8304), .B2(n9304), .C1(
        P2_U3151), .C2(n5756), .ZN(P2_U3265) );
  INV_X1 U9786 ( .A(n8602), .ZN(n9305) );
  OAI222_X1 U9787 ( .A1(n8304), .A2(n9305), .B1(n8294), .B2(n6226), .C1(
        P2_U3151), .C2(n5757), .ZN(P2_U3266) );
  OAI222_X1 U9788 ( .A1(n8304), .A2(n8296), .B1(n6154), .B2(P2_U3151), .C1(
        n8295), .C2(n8300), .ZN(P2_U3267) );
  OAI222_X1 U9789 ( .A1(n8304), .A2(n8298), .B1(n6156), .B2(P2_U3151), .C1(
        n8297), .C2(n8300), .ZN(P2_U3268) );
  INV_X1 U9790 ( .A(n8299), .ZN(n9310) );
  OAI222_X1 U9791 ( .A1(n8304), .A2(n9310), .B1(P2_U3151), .B2(n8302), .C1(
        n8301), .C2(n8300), .ZN(P2_U3269) );
  AOI21_X1 U9792 ( .B1(n8494), .B2(n8306), .A(n8305), .ZN(n8308) );
  AOI22_X1 U9793 ( .A1(n8986), .A2(n8475), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8311) );
  NAND2_X1 U9794 ( .A1(n9190), .A2(n4295), .ZN(n8310) );
  OAI22_X1 U9795 ( .A1(n8949), .A2(n8505), .B1(n8945), .B2(n8908), .ZN(n8983)
         );
  NAND2_X1 U9796 ( .A1(n8983), .A2(n8506), .ZN(n8309) );
  NAND4_X1 U9797 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(
        P1_U3214) );
  INV_X1 U9798 ( .A(n9520), .ZN(n9706) );
  OAI21_X1 U9799 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8316) );
  NAND2_X1 U9800 ( .A1(n8316), .A2(n8495), .ZN(n8321) );
  NAND2_X1 U9801 ( .A1(n8919), .A2(n8878), .ZN(n8318) );
  NAND2_X1 U9802 ( .A1(n8781), .A2(n8484), .ZN(n8317) );
  AND2_X1 U9803 ( .A1(n8318), .A2(n8317), .ZN(n9515) );
  OAI22_X1 U9804 ( .A1(n8459), .A2(n9515), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10002), .ZN(n8319) );
  AOI21_X1 U9805 ( .B1(n9518), .B2(n8475), .A(n8319), .ZN(n8320) );
  OAI211_X1 U9806 ( .C1(n9706), .C2(n8419), .A(n8321), .B(n8320), .ZN(P1_U3215) );
  INV_X1 U9807 ( .A(n9209), .ZN(n9045) );
  INV_X1 U9808 ( .A(n8322), .ZN(n8455) );
  INV_X1 U9809 ( .A(n8323), .ZN(n8325) );
  NOR3_X1 U9810 ( .A1(n8455), .A2(n8325), .A3(n8324), .ZN(n8327) );
  INV_X1 U9811 ( .A(n8326), .ZN(n8409) );
  OAI21_X1 U9812 ( .B1(n8327), .B2(n8409), .A(n8495), .ZN(n8332) );
  INV_X1 U9813 ( .A(n8328), .ZN(n9042) );
  AOI22_X1 U9814 ( .A1(n8941), .A2(n8878), .B1(n8484), .B2(n8935), .ZN(n9039)
         );
  OAI22_X1 U9815 ( .A1(n9039), .A2(n8459), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8329), .ZN(n8330) );
  AOI21_X1 U9816 ( .B1(n9042), .B2(n8475), .A(n8330), .ZN(n8331) );
  OAI211_X1 U9817 ( .C1(n9045), .C2(n8419), .A(n8332), .B(n8331), .ZN(P1_U3216) );
  XNOR2_X1 U9818 ( .A(n8465), .B(n8333), .ZN(n8334) );
  NAND2_X1 U9819 ( .A1(n8334), .A2(n8335), .ZN(n8464) );
  OAI21_X1 U9820 ( .B1(n8335), .B2(n8334), .A(n8464), .ZN(n8336) );
  NAND2_X1 U9821 ( .A1(n8336), .A2(n8495), .ZN(n8342) );
  INV_X1 U9822 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8337) );
  OAI22_X1 U9823 ( .A1(n8459), .A2(n8338), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8337), .ZN(n8339) );
  AOI21_X1 U9824 ( .B1(n8340), .B2(n8475), .A(n8339), .ZN(n8341) );
  OAI211_X1 U9825 ( .C1(n9682), .C2(n8419), .A(n8342), .B(n8341), .ZN(P1_U3217) );
  INV_X1 U9826 ( .A(n8343), .ZN(n8344) );
  NOR2_X1 U9827 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  XNOR2_X1 U9828 ( .A(n8347), .B(n8346), .ZN(n8354) );
  NAND2_X1 U9829 ( .A1(n8922), .A2(n8484), .ZN(n8349) );
  NAND2_X1 U9830 ( .A1(n8928), .A2(n8878), .ZN(n8348) );
  NAND2_X1 U9831 ( .A1(n8349), .A2(n8348), .ZN(n9103) );
  NOR2_X1 U9832 ( .A1(n8350), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8874) );
  AOI21_X1 U9833 ( .B1(n8506), .B2(n9103), .A(n8874), .ZN(n8351) );
  OAI21_X1 U9834 ( .B1(n8508), .B2(n9097), .A(n8351), .ZN(n8352) );
  AOI21_X1 U9835 ( .B1(n9228), .B2(n4295), .A(n8352), .ZN(n8353) );
  OAI21_X1 U9836 ( .B1(n8354), .B2(n8511), .A(n8353), .ZN(P1_U3219) );
  OAI21_X1 U9837 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8358) );
  NAND2_X1 U9838 ( .A1(n8358), .A2(n8495), .ZN(n8364) );
  NAND2_X1 U9839 ( .A1(n8935), .A2(n8878), .ZN(n8360) );
  NAND2_X1 U9840 ( .A1(n8928), .A2(n8484), .ZN(n8359) );
  AND2_X1 U9841 ( .A1(n8360), .A2(n8359), .ZN(n9069) );
  OAI22_X1 U9842 ( .A1(n8459), .A2(n9069), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8361), .ZN(n8362) );
  AOI21_X1 U9843 ( .B1(n9072), .B2(n8475), .A(n8362), .ZN(n8363) );
  OAI211_X1 U9844 ( .C1(n9075), .C2(n8419), .A(n8364), .B(n8363), .ZN(P1_U3223) );
  OAI21_X1 U9845 ( .B1(n8367), .B2(n8365), .A(n8366), .ZN(n8371) );
  NAND2_X1 U9846 ( .A1(n9199), .A2(n4295), .ZN(n8369) );
  OAI22_X1 U9847 ( .A1(n8945), .A2(n8505), .B1(n8940), .B2(n8908), .ZN(n9010)
         );
  AOI22_X1 U9848 ( .A1(n9010), .A2(n8506), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8368) );
  OAI211_X1 U9849 ( .C1(n8508), .C2(n9014), .A(n8369), .B(n8368), .ZN(n8370)
         );
  AOI21_X1 U9850 ( .B1(n8371), .B2(n8495), .A(n8370), .ZN(n8372) );
  INV_X1 U9851 ( .A(n8372), .ZN(P1_U3225) );
  INV_X1 U9852 ( .A(n8374), .ZN(n8375) );
  XOR2_X1 U9853 ( .A(n8373), .B(n8374), .Z(n8504) );
  NOR2_X1 U9854 ( .A1(n8504), .A2(n8503), .ZN(n8502) );
  AOI21_X1 U9855 ( .B1(n8375), .B2(n8373), .A(n8502), .ZN(n8379) );
  XNOR2_X1 U9856 ( .A(n8377), .B(n8376), .ZN(n8378) );
  XNOR2_X1 U9857 ( .A(n8379), .B(n8378), .ZN(n8385) );
  NAND2_X1 U9858 ( .A1(n8921), .A2(n8878), .ZN(n8381) );
  NAND2_X1 U9859 ( .A1(n8919), .A2(n8484), .ZN(n8380) );
  AND2_X1 U9860 ( .A1(n8381), .A2(n8380), .ZN(n9144) );
  NAND2_X1 U9861 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U9862 ( .A1(n8475), .A2(n9147), .ZN(n8382) );
  OAI211_X1 U9863 ( .C1(n8459), .C2(n9144), .A(n8827), .B(n8382), .ZN(n8383)
         );
  AOI21_X1 U9864 ( .B1(n9244), .B2(n4295), .A(n8383), .ZN(n8384) );
  OAI21_X1 U9865 ( .B1(n8385), .B2(n8511), .A(n8384), .ZN(P1_U3226) );
  OAI21_X1 U9866 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8389) );
  NAND2_X1 U9867 ( .A1(n8389), .A2(n8495), .ZN(n8397) );
  NAND2_X1 U9868 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9416) );
  INV_X1 U9869 ( .A(n9416), .ZN(n8390) );
  AOI21_X1 U9870 ( .B1(n8506), .B2(n8391), .A(n8390), .ZN(n8396) );
  NAND2_X1 U9871 ( .A1(n8475), .A2(n8392), .ZN(n8395) );
  NAND2_X1 U9872 ( .A1(n4295), .A2(n8393), .ZN(n8394) );
  NAND4_X1 U9873 ( .A1(n8397), .A2(n8396), .A3(n8395), .A4(n8394), .ZN(
        P1_U3227) );
  NAND2_X1 U9874 ( .A1(n4667), .A2(n8399), .ZN(n8400) );
  XNOR2_X1 U9875 ( .A(n8401), .B(n8400), .ZN(n8405) );
  INV_X1 U9876 ( .A(n8922), .ZN(n8923) );
  OAI22_X1 U9877 ( .A1(n8920), .A2(n8908), .B1(n8923), .B2(n8505), .ZN(n9135)
         );
  NAND2_X1 U9878 ( .A1(n9135), .A2(n8506), .ZN(n8402) );
  NAND2_X1 U9879 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8851) );
  OAI211_X1 U9880 ( .C1(n8508), .C2(n9129), .A(n8402), .B(n8851), .ZN(n8403)
         );
  AOI21_X1 U9881 ( .B1(n9239), .B2(n4295), .A(n8403), .ZN(n8404) );
  OAI21_X1 U9882 ( .B1(n8405), .B2(n8511), .A(n8404), .ZN(P1_U3228) );
  INV_X1 U9883 ( .A(n8406), .ZN(n8408) );
  NOR3_X1 U9884 ( .A1(n8409), .A2(n8408), .A3(n8407), .ZN(n8412) );
  INV_X1 U9885 ( .A(n8410), .ZN(n8411) );
  OAI21_X1 U9886 ( .B1(n8412), .B2(n8411), .A(n8495), .ZN(n8418) );
  INV_X1 U9887 ( .A(n8413), .ZN(n9029) );
  AND2_X1 U9888 ( .A1(n8938), .A2(n8484), .ZN(n8414) );
  AOI21_X1 U9889 ( .B1(n8943), .B2(n8878), .A(n8414), .ZN(n9025) );
  OAI22_X1 U9890 ( .A1(n9025), .A2(n8459), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8415), .ZN(n8416) );
  AOI21_X1 U9891 ( .B1(n9029), .B2(n8475), .A(n8416), .ZN(n8417) );
  OAI211_X1 U9892 ( .C1(n9032), .C2(n8419), .A(n8418), .B(n8417), .ZN(P1_U3229) );
  OAI21_X1 U9893 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8426) );
  XNOR2_X1 U9894 ( .A(n8424), .B(n8423), .ZN(n8425) );
  XNOR2_X1 U9895 ( .A(n8426), .B(n8425), .ZN(n8427) );
  NAND2_X1 U9896 ( .A1(n8427), .A2(n8495), .ZN(n8436) );
  NAND2_X1 U9897 ( .A1(n8429), .A2(n8428), .ZN(n8430) );
  AND2_X1 U9898 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8808) );
  AOI21_X1 U9899 ( .B1(n8506), .B2(n8430), .A(n8808), .ZN(n8435) );
  NAND2_X1 U9900 ( .A1(n4295), .A2(n8431), .ZN(n8434) );
  NAND2_X1 U9901 ( .A1(n8475), .A2(n8432), .ZN(n8433) );
  NAND4_X1 U9902 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(
        P1_U3231) );
  OAI21_X1 U9903 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8445) );
  NAND2_X1 U9904 ( .A1(n9223), .A2(n4295), .ZN(n8443) );
  NAND2_X1 U9905 ( .A1(n8931), .A2(n8878), .ZN(n8441) );
  NAND2_X1 U9906 ( .A1(n8926), .A2(n8484), .ZN(n8440) );
  NAND2_X1 U9907 ( .A1(n8441), .A2(n8440), .ZN(n9087) );
  AOI22_X1 U9908 ( .A1(n8506), .A2(n9087), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8442) );
  OAI211_X1 U9909 ( .C1(n8508), .C2(n9090), .A(n8443), .B(n8442), .ZN(n8444)
         );
  AOI21_X1 U9910 ( .B1(n8445), .B2(n8495), .A(n8444), .ZN(n8446) );
  INV_X1 U9911 ( .A(n8446), .ZN(P1_U3233) );
  XOR2_X1 U9912 ( .A(n8448), .B(n8447), .Z(n8454) );
  NAND2_X1 U9913 ( .A1(n8909), .A2(n8484), .ZN(n8450) );
  NAND2_X1 U9914 ( .A1(n8915), .A2(n8878), .ZN(n8449) );
  NAND2_X1 U9915 ( .A1(n8450), .A2(n8449), .ZN(n9529) );
  AOI22_X1 U9916 ( .A1(n8506), .A2(n9529), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8451) );
  OAI21_X1 U9917 ( .B1(n8508), .B2(n9540), .A(n8451), .ZN(n8452) );
  AOI21_X1 U9918 ( .B1(n8875), .B2(n4295), .A(n8452), .ZN(n8453) );
  OAI21_X1 U9919 ( .B1(n8454), .B2(n8511), .A(n8453), .ZN(P1_U3234) );
  AOI21_X1 U9920 ( .B1(n8457), .B2(n8456), .A(n8455), .ZN(n8463) );
  NOR2_X1 U9921 ( .A1(n8508), .A2(n9053), .ZN(n8461) );
  AOI22_X1 U9922 ( .A1(n8938), .A2(n8878), .B1(n8931), .B2(n8484), .ZN(n9059)
         );
  OAI22_X1 U9923 ( .A1(n9059), .A2(n8459), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8458), .ZN(n8460) );
  AOI211_X1 U9924 ( .C1(n9213), .C2(n4295), .A(n8461), .B(n8460), .ZN(n8462)
         );
  OAI21_X1 U9925 ( .B1(n8463), .B2(n8511), .A(n8462), .ZN(P1_U3235) );
  OAI21_X1 U9926 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8470) );
  XNOR2_X1 U9927 ( .A(n8468), .B(n8467), .ZN(n8469) );
  XNOR2_X1 U9928 ( .A(n8470), .B(n8469), .ZN(n8471) );
  NAND2_X1 U9929 ( .A1(n8471), .A2(n8495), .ZN(n8479) );
  AOI22_X1 U9930 ( .A1(n8506), .A2(n8472), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8478) );
  NAND2_X1 U9931 ( .A1(n8473), .A2(n4295), .ZN(n8477) );
  NAND2_X1 U9932 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  NAND4_X1 U9933 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(
        P1_U3236) );
  NAND2_X1 U9934 ( .A1(n8481), .A2(n8480), .ZN(n8483) );
  XOR2_X1 U9935 ( .A(n8483), .B(n8482), .Z(n8490) );
  NAND2_X1 U9936 ( .A1(n8926), .A2(n8878), .ZN(n8486) );
  NAND2_X1 U9937 ( .A1(n8921), .A2(n8484), .ZN(n8485) );
  NAND2_X1 U9938 ( .A1(n8486), .A2(n8485), .ZN(n9111) );
  AOI22_X1 U9939 ( .A1(n8506), .A2(n9111), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8487) );
  OAI21_X1 U9940 ( .B1(n8508), .B2(n9116), .A(n8487), .ZN(n8488) );
  AOI21_X1 U9941 ( .B1(n9121), .B2(n4295), .A(n8488), .ZN(n8489) );
  OAI21_X1 U9942 ( .B1(n8490), .B2(n8511), .A(n8489), .ZN(P1_U3238) );
  INV_X1 U9943 ( .A(n8366), .ZN(n8493) );
  OAI21_X1 U9944 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n8496) );
  NAND3_X1 U9945 ( .A1(n8496), .A2(n8495), .A3(n8494), .ZN(n8501) );
  OAI22_X1 U9946 ( .A1(n8596), .A2(n8505), .B1(n8944), .B2(n8908), .ZN(n8994)
         );
  AOI22_X1 U9947 ( .A1(n8994), .A2(n8506), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8497) );
  OAI21_X1 U9948 ( .B1(n8508), .B2(n9000), .A(n8497), .ZN(n8498) );
  AOI21_X1 U9949 ( .B1(n9004), .B2(n4295), .A(n8498), .ZN(n8500) );
  NAND2_X1 U9950 ( .A1(n8501), .A2(n8500), .ZN(P1_U3240) );
  AOI21_X1 U9951 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(n8512) );
  INV_X1 U9952 ( .A(n8915), .ZN(n8543) );
  OAI22_X1 U9953 ( .A1(n8543), .A2(n8908), .B1(n8920), .B2(n8505), .ZN(n9158)
         );
  AOI22_X1 U9954 ( .A1(n9158), .A2(n8506), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8507) );
  OAI21_X1 U9955 ( .B1(n8508), .B2(n9163), .A(n8507), .ZN(n8509) );
  AOI21_X1 U9956 ( .B1(n9165), .B2(n4295), .A(n8509), .ZN(n8510) );
  OAI21_X1 U9957 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(P1_U3241) );
  NOR4_X1 U9958 ( .A1(n8514), .A2(n5640), .A3(n8880), .A4(n8513), .ZN(n8777)
         );
  OAI21_X1 U9959 ( .B1(n8770), .B2(n8769), .A(P1_B_REG_SCAN_IN), .ZN(n8776) );
  NAND2_X1 U9960 ( .A1(n8974), .A2(n8951), .ZN(n8689) );
  INV_X1 U9961 ( .A(n8766), .ZN(n8612) );
  OR2_X1 U9962 ( .A1(n9004), .A2(n8945), .ZN(n8632) );
  AND4_X1 U9963 ( .A1(n8689), .A2(n8612), .A3(n8658), .A4(n8632), .ZN(n8601)
         );
  OR2_X1 U9964 ( .A1(n9218), .A2(n8930), .ZN(n8676) );
  OR2_X1 U9965 ( .A1(n9223), .A2(n8929), .ZN(n9064) );
  AND2_X1 U9966 ( .A1(n8676), .A2(n9064), .ZN(n8890) );
  INV_X1 U9967 ( .A(n8523), .ZN(n8516) );
  INV_X1 U9968 ( .A(n8515), .ZN(n8524) );
  OAI21_X1 U9969 ( .B1(n8517), .B2(n8516), .A(n8524), .ZN(n8520) );
  INV_X1 U9970 ( .A(n8518), .ZN(n8519) );
  AOI21_X1 U9971 ( .B1(n8520), .B2(n8643), .A(n8519), .ZN(n8529) );
  INV_X1 U9972 ( .A(n9559), .ZN(n8521) );
  OR2_X1 U9973 ( .A1(n8522), .A2(n8521), .ZN(n8718) );
  INV_X1 U9974 ( .A(n8525), .ZN(n8526) );
  MUX2_X1 U9975 ( .A(n8529), .B(n8528), .S(n8766), .Z(n8535) );
  INV_X1 U9976 ( .A(n8535), .ZN(n8530) );
  NAND2_X1 U9977 ( .A1(n8530), .A2(n8534), .ZN(n8531) );
  NAND2_X1 U9978 ( .A1(n8540), .A2(n8536), .ZN(n8724) );
  AOI21_X1 U9979 ( .B1(n8531), .B2(n8722), .A(n8724), .ZN(n8532) );
  NAND2_X1 U9980 ( .A1(n8663), .A2(n8537), .ZN(n8725) );
  OAI21_X1 U9981 ( .B1(n8532), .B2(n8725), .A(n8728), .ZN(n8542) );
  INV_X1 U9982 ( .A(n8641), .ZN(n8533) );
  AOI21_X1 U9983 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8539) );
  INV_X1 U9984 ( .A(n8536), .ZN(n8538) );
  OAI211_X1 U9985 ( .C1(n8539), .C2(n8538), .A(n8537), .B(n8722), .ZN(n8541)
         );
  OR2_X1 U9986 ( .A1(n8875), .A2(n8913), .ZN(n8729) );
  NAND2_X1 U9987 ( .A1(n8549), .A2(n8729), .ZN(n8546) );
  NAND2_X1 U9988 ( .A1(n9520), .A2(n8543), .ZN(n8550) );
  INV_X1 U9989 ( .A(n9511), .ZN(n8545) );
  NAND2_X1 U9990 ( .A1(n8875), .A2(n8913), .ZN(n9512) );
  INV_X1 U9991 ( .A(n9512), .ZN(n8544) );
  NOR2_X1 U9992 ( .A1(n8545), .A2(n8544), .ZN(n8664) );
  NAND2_X1 U9993 ( .A1(n8546), .A2(n8664), .ZN(n8547) );
  OR2_X2 U9994 ( .A1(n9244), .A2(n8920), .ZN(n8669) );
  OR2_X1 U9995 ( .A1(n9165), .A2(n8917), .ZN(n8649) );
  AND2_X1 U9996 ( .A1(n8669), .A2(n8649), .ZN(n8733) );
  NAND3_X1 U9997 ( .A1(n8547), .A2(n8733), .A3(n9155), .ZN(n8553) );
  NAND2_X1 U9998 ( .A1(n9511), .A2(n8729), .ZN(n8548) );
  NAND2_X1 U9999 ( .A1(n9165), .A2(n8917), .ZN(n8667) );
  NAND2_X1 U10000 ( .A1(n8667), .A2(n8550), .ZN(n8732) );
  OAI21_X1 U10001 ( .B1(n8551), .B2(n8732), .A(n8669), .ZN(n8552) );
  NAND2_X1 U10002 ( .A1(n9244), .A2(n8920), .ZN(n8737) );
  INV_X1 U10003 ( .A(n8667), .ZN(n8554) );
  NAND2_X1 U10004 ( .A1(n8669), .A2(n8554), .ZN(n8555) );
  OAI211_X1 U10005 ( .C1(n9165), .C2(n8766), .A(n8555), .B(n8737), .ZN(n8558)
         );
  NAND2_X1 U10006 ( .A1(n8737), .A2(n8919), .ZN(n8556) );
  NAND2_X1 U10007 ( .A1(n8556), .A2(n8612), .ZN(n8557) );
  NAND2_X1 U10008 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NAND2_X1 U10009 ( .A1(n9239), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U10010 ( .A1(n9109), .A2(n8562), .ZN(n9124) );
  INV_X1 U10011 ( .A(n9124), .ZN(n9134) );
  OR2_X1 U10012 ( .A1(n9228), .A2(n8925), .ZN(n8634) );
  NAND2_X1 U10013 ( .A1(n9064), .A2(n8634), .ZN(n8561) );
  NAND2_X1 U10014 ( .A1(n8561), .A2(n8612), .ZN(n8572) );
  OR2_X1 U10015 ( .A1(n9121), .A2(n8923), .ZN(n8635) );
  NAND2_X1 U10016 ( .A1(n8634), .A2(n8635), .ZN(n8738) );
  NAND2_X1 U10017 ( .A1(n9121), .A2(n8923), .ZN(n8672) );
  AND2_X1 U10018 ( .A1(n8672), .A2(n8562), .ZN(n8563) );
  NOR2_X1 U10019 ( .A1(n8738), .A2(n8563), .ZN(n8742) );
  AND2_X1 U10020 ( .A1(n9223), .A2(n8929), .ZN(n8888) );
  OR2_X1 U10021 ( .A1(n8742), .A2(n8888), .ZN(n8571) );
  NAND2_X1 U10022 ( .A1(n9228), .A2(n8925), .ZN(n8744) );
  NAND2_X1 U10023 ( .A1(n8744), .A2(n8766), .ZN(n8567) );
  NAND3_X1 U10024 ( .A1(n8635), .A2(n8612), .A3(n9109), .ZN(n8564) );
  OAI21_X1 U10025 ( .B1(n8571), .B2(n8567), .A(n8564), .ZN(n8565) );
  NAND3_X1 U10026 ( .A1(n8566), .A2(n8572), .A3(n8565), .ZN(n8575) );
  INV_X1 U10027 ( .A(n8567), .ZN(n8568) );
  NAND2_X1 U10028 ( .A1(n8568), .A2(n8738), .ZN(n8570) );
  AND2_X1 U10029 ( .A1(n8744), .A2(n8672), .ZN(n8569) );
  OAI22_X1 U10030 ( .A1(n8571), .A2(n8570), .B1(n8569), .B2(n8766), .ZN(n8573)
         );
  NAND2_X1 U10031 ( .A1(n9218), .A2(n8930), .ZN(n8891) );
  NAND2_X1 U10032 ( .A1(n8891), .A2(n8889), .ZN(n8677) );
  AOI22_X1 U10033 ( .A1(n8573), .A2(n8572), .B1(n8612), .B2(n8677), .ZN(n8574)
         );
  OAI211_X1 U10034 ( .C1(n8612), .C2(n8890), .A(n8575), .B(n8574), .ZN(n8577)
         );
  MUX2_X1 U10035 ( .A(n8891), .B(n8676), .S(n8612), .Z(n8576) );
  NAND2_X1 U10036 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U10037 ( .A1(n9213), .A2(n8934), .ZN(n8579) );
  NAND2_X1 U10038 ( .A1(n9036), .A2(n8579), .ZN(n8893) );
  NAND2_X1 U10039 ( .A1(n8578), .A2(n9058), .ZN(n8581) );
  INV_X1 U10040 ( .A(n8938), .ZN(n8939) );
  NAND2_X1 U10041 ( .A1(n9209), .A2(n8939), .ZN(n8895) );
  NAND2_X1 U10042 ( .A1(n8895), .A2(n8579), .ZN(n8679) );
  NAND2_X1 U10043 ( .A1(n8679), .A2(n8766), .ZN(n8580) );
  OR2_X1 U10044 ( .A1(n9209), .A2(n8939), .ZN(n8633) );
  NAND2_X1 U10045 ( .A1(n8633), .A2(n9036), .ZN(n8659) );
  NAND2_X1 U10046 ( .A1(n9204), .A2(n8940), .ZN(n8680) );
  OAI21_X1 U10047 ( .B1(n8766), .B2(n8895), .A(n9023), .ZN(n8582) );
  MUX2_X1 U10048 ( .A(n8680), .B(n8898), .S(n8612), .Z(n8583) );
  INV_X1 U10049 ( .A(n8595), .ZN(n8584) );
  INV_X1 U10050 ( .A(n8992), .ZN(n8899) );
  NAND2_X1 U10051 ( .A1(n9004), .A2(n8945), .ZN(n8684) );
  NAND2_X1 U10052 ( .A1(n9199), .A2(n8944), .ZN(n8681) );
  OAI211_X1 U10053 ( .C1(n8584), .C2(n8899), .A(n8684), .B(n8681), .ZN(n8600)
         );
  NAND2_X1 U10054 ( .A1(n8596), .A2(n8612), .ZN(n8589) );
  INV_X1 U10055 ( .A(n8589), .ZN(n8585) );
  AOI22_X1 U10056 ( .A1(n9190), .A2(n8585), .B1(n8949), .B2(n8612), .ZN(n8594)
         );
  NAND2_X1 U10057 ( .A1(n8947), .A2(n8766), .ZN(n8587) );
  OAI22_X1 U10058 ( .A1(n9190), .A2(n8587), .B1(n8949), .B2(n8612), .ZN(n8586)
         );
  NAND2_X1 U10059 ( .A1(n8974), .A2(n8586), .ZN(n8593) );
  INV_X1 U10060 ( .A(n8587), .ZN(n8588) );
  AND2_X1 U10061 ( .A1(n8588), .A2(n8951), .ZN(n8591) );
  OAI21_X1 U10062 ( .B1(n8951), .B2(n8589), .A(n9190), .ZN(n8590) );
  OAI21_X1 U10063 ( .B1(n8591), .B2(n9190), .A(n8590), .ZN(n8592) );
  OAI211_X1 U10064 ( .C1(n8974), .C2(n8594), .A(n8593), .B(n8592), .ZN(n8599)
         );
  NAND2_X1 U10065 ( .A1(n8632), .A2(n8992), .ZN(n8675) );
  AOI21_X1 U10066 ( .B1(n8595), .B2(n8681), .A(n8675), .ZN(n8598) );
  NAND2_X1 U10067 ( .A1(n9186), .A2(n8949), .ZN(n8903) );
  NAND4_X1 U10068 ( .A1(n8903), .A2(n8902), .A3(n8766), .A4(n8684), .ZN(n8597)
         );
  NAND2_X1 U10069 ( .A1(n8602), .A2(n8608), .ZN(n8605) );
  OR2_X1 U10070 ( .A1(n8603), .A2(n9307), .ZN(n8604) );
  OR2_X1 U10071 ( .A1(n9179), .A2(n8606), .ZN(n8690) );
  NAND2_X1 U10072 ( .A1(n9179), .A2(n8606), .ZN(n8691) );
  NAND2_X1 U10073 ( .A1(n8690), .A2(n8691), .ZN(n8954) );
  MUX2_X1 U10074 ( .A(n8691), .B(n8690), .S(n8766), .Z(n8607) );
  NAND2_X1 U10075 ( .A1(n8609), .A2(n8608), .ZN(n8611) );
  OR2_X1 U10076 ( .A1(n4999), .A2(n9303), .ZN(n8610) );
  MUX2_X1 U10077 ( .A(n8625), .B(n8612), .S(n8876), .Z(n8624) );
  MUX2_X1 U10078 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8614), .S(n4302), .Z(
        n8616) );
  NAND2_X1 U10079 ( .A1(n5040), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10080 ( .A1(n8620), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8617) );
  NAND3_X1 U10081 ( .A1(n8619), .A2(n8618), .A3(n8617), .ZN(n8778) );
  NAND2_X1 U10082 ( .A1(n9172), .A2(n8778), .ZN(n8773) );
  NAND2_X1 U10083 ( .A1(n8620), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10084 ( .A1(n5040), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8621) );
  AND3_X1 U10085 ( .A1(n8623), .A2(n8622), .A3(n8621), .ZN(n8905) );
  INV_X1 U10086 ( .A(n8905), .ZN(n8779) );
  NAND2_X1 U10087 ( .A1(n8779), .A2(n8778), .ZN(n8696) );
  NAND3_X1 U10088 ( .A1(n8624), .A2(n8773), .A3(n8696), .ZN(n8629) );
  NAND3_X1 U10089 ( .A1(n8626), .A2(n8627), .A3(n8779), .ZN(n8628) );
  INV_X1 U10090 ( .A(n8778), .ZN(n8881) );
  NAND3_X1 U10091 ( .A1(n8629), .A2(n8628), .A3(n8767), .ZN(n8765) );
  INV_X1 U10092 ( .A(n8630), .ZN(n8631) );
  AOI22_X1 U10093 ( .A1(n8765), .A2(n8631), .B1(n9535), .B2(n8637), .ZN(n8704)
         );
  OAI21_X1 U10094 ( .B1(n8905), .B2(n8876), .A(n8767), .ZN(n8705) );
  INV_X1 U10095 ( .A(n8773), .ZN(n8753) );
  NAND2_X1 U10096 ( .A1(n8876), .A2(n8905), .ZN(n8692) );
  NAND2_X1 U10097 ( .A1(n8689), .A2(n8903), .ZN(n8964) );
  NAND2_X1 U10098 ( .A1(n8632), .A2(n8684), .ZN(n8996) );
  NAND2_X1 U10099 ( .A1(n8633), .A2(n8895), .ZN(n9037) );
  XNOR2_X1 U10100 ( .A(n9223), .B(n8929), .ZN(n9085) );
  NAND2_X1 U10101 ( .A1(n8676), .A2(n8891), .ZN(n9066) );
  NAND2_X1 U10102 ( .A1(n8635), .A2(n8672), .ZN(n9113) );
  NOR2_X1 U10103 ( .A1(n9568), .A2(n8636), .ZN(n8640) );
  NOR2_X1 U10104 ( .A1(n9586), .A2(n6886), .ZN(n8639) );
  AND4_X1 U10105 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n8644)
         );
  NOR2_X1 U10106 ( .A1(n9594), .A2(n6773), .ZN(n8642) );
  NAND4_X1 U10107 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n8647)
         );
  NOR4_X1 U10108 ( .A1(n8647), .A2(n8646), .A3(n4761), .A4(n8645), .ZN(n8648)
         );
  NAND2_X1 U10109 ( .A1(n8729), .A2(n9512), .ZN(n9528) );
  NAND4_X1 U10110 ( .A1(n8648), .A2(n9511), .A3(n4529), .A4(n8911), .ZN(n8650)
         );
  NOR2_X1 U10111 ( .A1(n8650), .A2(n9156), .ZN(n8651) );
  NAND3_X1 U10112 ( .A1(n9134), .A2(n9143), .A3(n8651), .ZN(n8652) );
  NOR4_X1 U10113 ( .A1(n9037), .A2(n8893), .A3(n9085), .A4(n8653), .ZN(n8654)
         );
  NAND3_X1 U10114 ( .A1(n9009), .A2(n9023), .A3(n8654), .ZN(n8655) );
  NAND2_X1 U10115 ( .A1(n8692), .A2(n8656), .ZN(n8657) );
  NOR4_X2 U10116 ( .A1(n8705), .A2(n8753), .A3(n8954), .A4(n8657), .ZN(n8703)
         );
  INV_X1 U10117 ( .A(n8658), .ZN(n8687) );
  INV_X1 U10118 ( .A(n8890), .ZN(n8661) );
  NAND2_X1 U10119 ( .A1(n8659), .A2(n8895), .ZN(n8660) );
  NAND2_X1 U10120 ( .A1(n8898), .A2(n8660), .ZN(n8683) );
  NOR4_X1 U10121 ( .A1(n8687), .A2(n8675), .A3(n8661), .A4(n8683), .ZN(n8748)
         );
  INV_X1 U10122 ( .A(n9155), .ZN(n8665) );
  NOR2_X1 U10123 ( .A1(n9156), .A2(n8665), .ZN(n8666) );
  NAND2_X1 U10124 ( .A1(n9509), .A2(n8666), .ZN(n8668) );
  INV_X1 U10125 ( .A(n9109), .ZN(n8670) );
  NOR2_X1 U10126 ( .A1(n9113), .A2(n8670), .ZN(n8671) );
  NAND2_X1 U10127 ( .A1(n9108), .A2(n8671), .ZN(n8673) );
  NAND2_X1 U10128 ( .A1(n8673), .A2(n8672), .ZN(n9102) );
  INV_X1 U10129 ( .A(n8675), .ZN(n8686) );
  AND2_X1 U10130 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  NOR2_X1 U10131 ( .A1(n8679), .A2(n8678), .ZN(n8682) );
  OAI211_X1 U10132 ( .C1(n8683), .C2(n8682), .A(n8681), .B(n8680), .ZN(n8685)
         );
  INV_X1 U10133 ( .A(n8684), .ZN(n8900) );
  AOI21_X1 U10134 ( .B1(n8686), .B2(n8685), .A(n8900), .ZN(n8688) );
  OAI211_X1 U10135 ( .C1(n8688), .C2(n8687), .A(n8903), .B(n8902), .ZN(n8746)
         );
  AOI21_X1 U10136 ( .B1(n8748), .B2(n9086), .A(n8746), .ZN(n8694) );
  NAND2_X1 U10137 ( .A1(n8690), .A2(n8689), .ZN(n8751) );
  NAND2_X1 U10138 ( .A1(n8692), .A2(n8691), .ZN(n8749) );
  AOI21_X1 U10139 ( .B1(n8881), .B2(n8876), .A(n8749), .ZN(n8693) );
  OAI21_X1 U10140 ( .B1(n8694), .B2(n8751), .A(n8693), .ZN(n8695) );
  OAI21_X1 U10141 ( .B1(n8696), .B2(n8876), .A(n8695), .ZN(n8700) );
  INV_X1 U10142 ( .A(n8697), .ZN(n8699) );
  INV_X1 U10143 ( .A(n8767), .ZN(n8698) );
  AOI211_X1 U10144 ( .C1(n8773), .C2(n8700), .A(n8699), .B(n8698), .ZN(n8701)
         );
  OAI21_X1 U10145 ( .B1(n8701), .B2(n8703), .A(n4305), .ZN(n8702) );
  OAI211_X1 U10146 ( .C1(n8704), .C2(n8703), .A(n8756), .B(n8702), .ZN(n8764)
         );
  INV_X1 U10147 ( .A(n8705), .ZN(n8755) );
  INV_X1 U10148 ( .A(n8706), .ZN(n8711) );
  NAND2_X1 U10149 ( .A1(n8791), .A2(n9629), .ZN(n8710) );
  NAND2_X1 U10150 ( .A1(n6774), .A2(n8707), .ZN(n8709) );
  NAND4_X1 U10151 ( .A1(n8711), .A2(n8710), .A3(n8709), .A4(n8708), .ZN(n8715)
         );
  NAND2_X1 U10152 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NOR2_X1 U10153 ( .A1(n8715), .A2(n8714), .ZN(n8717) );
  OAI21_X1 U10154 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8720) );
  NAND3_X1 U10155 ( .A1(n8720), .A2(n4521), .A3(n8719), .ZN(n8723) );
  NAND3_X1 U10156 ( .A1(n8723), .A2(n8722), .A3(n8721), .ZN(n8727) );
  INV_X1 U10157 ( .A(n8724), .ZN(n8726) );
  AOI21_X1 U10158 ( .B1(n8727), .B2(n8726), .A(n8725), .ZN(n8731) );
  NAND2_X1 U10159 ( .A1(n9512), .A2(n8728), .ZN(n8730) );
  OAI211_X1 U10160 ( .C1(n8731), .C2(n8730), .A(n9155), .B(n8729), .ZN(n8736)
         );
  INV_X1 U10161 ( .A(n8732), .ZN(n8735) );
  INV_X1 U10162 ( .A(n8733), .ZN(n8734) );
  AOI21_X1 U10163 ( .B1(n8736), .B2(n8735), .A(n8734), .ZN(n8741) );
  INV_X1 U10164 ( .A(n8737), .ZN(n8740) );
  INV_X1 U10165 ( .A(n8738), .ZN(n8739) );
  OAI211_X1 U10166 ( .C1(n8741), .C2(n8740), .A(n8739), .B(n9109), .ZN(n8745)
         );
  INV_X1 U10167 ( .A(n8742), .ZN(n8743) );
  NAND3_X1 U10168 ( .A1(n8745), .A2(n8744), .A3(n8743), .ZN(n8747) );
  AOI21_X1 U10169 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8752) );
  INV_X1 U10170 ( .A(n8749), .ZN(n8750) );
  OAI21_X1 U10171 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8754) );
  AOI21_X1 U10172 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(n8758) );
  NOR3_X1 U10173 ( .A1(n8758), .A2(n8756), .A3(n4305), .ZN(n8762) );
  INV_X1 U10174 ( .A(n5626), .ZN(n8757) );
  INV_X1 U10175 ( .A(n8770), .ZN(n8759) );
  NAND2_X1 U10176 ( .A1(n8764), .A2(n8763), .ZN(n8775) );
  OAI21_X1 U10177 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(n8772) );
  NOR3_X1 U10178 ( .A1(n8770), .A2(n8769), .A3(n8768), .ZN(n8771) );
  OAI211_X1 U10179 ( .C1(n8773), .C2(n4305), .A(n8772), .B(n8771), .ZN(n8774)
         );
  OAI211_X1 U10180 ( .C1(n8777), .C2(n8776), .A(n8775), .B(n8774), .ZN(
        P1_U3242) );
  MUX2_X1 U10181 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n8778), .S(n8792), .Z(
        P1_U3585) );
  MUX2_X1 U10182 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8779), .S(n8792), .Z(
        P1_U3584) );
  MUX2_X1 U10183 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8951), .S(n8792), .Z(
        P1_U3582) );
  MUX2_X1 U10184 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8947), .S(n8792), .Z(
        P1_U3581) );
  MUX2_X1 U10185 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8946), .S(n8792), .Z(
        P1_U3580) );
  MUX2_X1 U10186 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8943), .S(n8792), .Z(
        P1_U3579) );
  MUX2_X1 U10187 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8941), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8938), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10189 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8935), .S(n8792), .Z(
        P1_U3576) );
  MUX2_X1 U10190 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n8931), .S(n8792), .Z(
        P1_U3575) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n8928), .S(n8792), .Z(
        P1_U3574) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8780), .S(n8792), .Z(
        P1_U3570) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8919), .S(n8792), .Z(
        P1_U3569) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8915), .S(n8792), .Z(
        P1_U3568) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8781), .S(n8792), .Z(
        P1_U3567) );
  MUX2_X1 U10196 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8909), .S(n8792), .Z(
        P1_U3566) );
  MUX2_X1 U10197 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8782), .S(n8792), .Z(
        P1_U3565) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8783), .S(n8792), .Z(
        P1_U3564) );
  MUX2_X1 U10199 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8784), .S(n8792), .Z(
        P1_U3563) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8785), .S(n8792), .Z(
        P1_U3562) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8786), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8787), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8788), .S(n8792), .Z(
        P1_U3559) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8789), .S(n8792), .Z(
        P1_U3558) );
  MUX2_X1 U10205 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8790), .S(n8792), .Z(
        P1_U3557) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8791), .S(n8792), .Z(
        P1_U3556) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6774), .S(n8792), .Z(
        P1_U3555) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6751), .S(n8792), .Z(
        P1_U3554) );
  OAI211_X1 U10209 ( .C1(n8795), .C2(n8794), .A(n9489), .B(n8793), .ZN(n8803)
         );
  OAI211_X1 U10210 ( .C1(n8798), .C2(n8797), .A(n9497), .B(n8796), .ZN(n8802)
         );
  AOI22_X1 U10211 ( .A1(n9400), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8801) );
  NAND2_X1 U10212 ( .A1(n9485), .A2(n4300), .ZN(n8800) );
  NAND4_X1 U10213 ( .A1(n8803), .A2(n8802), .A3(n8801), .A4(n8800), .ZN(
        P1_U3244) );
  OAI21_X1 U10214 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n8807) );
  NAND2_X1 U10215 ( .A1(n8807), .A2(n9497), .ZN(n8817) );
  AOI21_X1 U10216 ( .B1(n9400), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8808), .ZN(
        n8816) );
  OAI21_X1 U10217 ( .B1(n8811), .B2(n8810), .A(n8809), .ZN(n8812) );
  NAND2_X1 U10218 ( .A1(n8812), .A2(n9489), .ZN(n8815) );
  NAND2_X1 U10219 ( .A1(n9485), .A2(n8813), .ZN(n8814) );
  NAND4_X1 U10220 ( .A1(n8817), .A2(n8816), .A3(n8815), .A4(n8814), .ZN(
        P1_U3252) );
  INV_X1 U10221 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9245) );
  AOI22_X1 U10222 ( .A1(n8846), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9245), .B2(
        n8828), .ZN(n8825) );
  INV_X1 U10223 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8818) );
  MUX2_X1 U10224 ( .A(n8818), .B(P1_REG1_REG_13__SCAN_IN), .S(n9457), .Z(n9450) );
  OAI21_X1 U10225 ( .B1(n8831), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8819), .ZN(
        n9451) );
  NOR2_X1 U10226 ( .A1(n9450), .A2(n9451), .ZN(n9449) );
  AOI21_X1 U10227 ( .B1(n9457), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9449), .ZN(
        n9467) );
  INV_X1 U10228 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U10229 ( .A1(n8833), .A2(n9736), .ZN(n8821) );
  NAND2_X1 U10230 ( .A1(n9471), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8820) );
  AND2_X1 U10231 ( .A1(n8821), .A2(n8820), .ZN(n9466) );
  NOR2_X1 U10232 ( .A1(n9467), .A2(n9466), .ZN(n9465) );
  NOR2_X1 U10233 ( .A1(n8822), .A2(n8835), .ZN(n8823) );
  XNOR2_X1 U10234 ( .A(n8835), .B(n8822), .ZN(n9478) );
  NOR2_X1 U10235 ( .A1(n5321), .A2(n9478), .ZN(n9477) );
  NAND2_X1 U10236 ( .A1(n8825), .A2(n8824), .ZN(n8845) );
  OAI21_X1 U10237 ( .B1(n8825), .B2(n8824), .A(n8845), .ZN(n8842) );
  NAND2_X1 U10238 ( .A1(n9400), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8826) );
  OAI211_X1 U10239 ( .C1(n9501), .C2(n8828), .A(n8827), .B(n8826), .ZN(n8841)
         );
  NAND2_X1 U10240 ( .A1(n9457), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8829) );
  OAI21_X1 U10241 ( .B1(n9457), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8829), .ZN(
        n9453) );
  OAI21_X1 U10242 ( .B1(n8831), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8830), .ZN(
        n9454) );
  NOR2_X1 U10243 ( .A1(n9453), .A2(n9454), .ZN(n9452) );
  NAND2_X1 U10244 ( .A1(n8833), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8832) );
  OAI21_X1 U10245 ( .B1(n8833), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8832), .ZN(
        n9463) );
  NOR2_X1 U10246 ( .A1(n8834), .A2(n8835), .ZN(n8836) );
  NOR2_X1 U10247 ( .A1(n5323), .A2(n9481), .ZN(n9480) );
  NOR2_X1 U10248 ( .A1(n8836), .A2(n9480), .ZN(n8839) );
  NAND2_X1 U10249 ( .A1(n8846), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8837) );
  OAI21_X1 U10250 ( .B1(n8846), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8837), .ZN(
        n8838) );
  NOR2_X1 U10251 ( .A1(n8839), .A2(n8838), .ZN(n8844) );
  AOI211_X1 U10252 ( .C1(n8839), .C2(n8838), .A(n8844), .B(n9479), .ZN(n8840)
         );
  AOI211_X1 U10253 ( .C1(n9489), .C2(n8842), .A(n8841), .B(n8840), .ZN(n8843)
         );
  INV_X1 U10254 ( .A(n8843), .ZN(P1_U3259) );
  AOI21_X1 U10255 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8846), .A(n8844), .ZN(
        n8856) );
  XNOR2_X1 U10256 ( .A(n8858), .B(n9130), .ZN(n8857) );
  XOR2_X1 U10257 ( .A(n8856), .B(n8857), .Z(n8855) );
  OAI21_X1 U10258 ( .B1(n8846), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8845), .ZN(
        n8849) );
  OR2_X1 U10259 ( .A1(n8858), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U10260 ( .A1(n8858), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8847) );
  AND2_X1 U10261 ( .A1(n8863), .A2(n8847), .ZN(n8848) );
  NAND2_X1 U10262 ( .A1(n8849), .A2(n8848), .ZN(n8864) );
  OAI21_X1 U10263 ( .B1(n8849), .B2(n8848), .A(n8864), .ZN(n8850) );
  NAND2_X1 U10264 ( .A1(n8850), .A2(n9489), .ZN(n8854) );
  INV_X1 U10265 ( .A(n9400), .ZN(n9506) );
  OAI21_X1 U10266 ( .B1(n9506), .B2(n10001), .A(n8851), .ZN(n8852) );
  AOI21_X1 U10267 ( .B1(n8858), .B2(n9485), .A(n8852), .ZN(n8853) );
  OAI211_X1 U10268 ( .C1(n8855), .C2(n9479), .A(n8854), .B(n8853), .ZN(
        P1_U3260) );
  NAND2_X1 U10269 ( .A1(n8865), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8861) );
  OAI21_X1 U10270 ( .B1(n8865), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8861), .ZN(
        n9493) );
  NAND2_X1 U10271 ( .A1(n8857), .A2(n8856), .ZN(n8860) );
  OR2_X1 U10272 ( .A1(n8858), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U10273 ( .A1(n8860), .A2(n8859), .ZN(n9494) );
  NAND2_X1 U10274 ( .A1(n9496), .A2(n8861), .ZN(n8862) );
  XNOR2_X1 U10275 ( .A(n8862), .B(n9098), .ZN(n8870) );
  AND2_X1 U10276 ( .A1(n8864), .A2(n8863), .ZN(n9492) );
  NAND2_X1 U10277 ( .A1(n8865), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8867) );
  OAI21_X1 U10278 ( .B1(n8865), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8867), .ZN(
        n8866) );
  INV_X1 U10279 ( .A(n8866), .ZN(n9491) );
  NAND2_X1 U10280 ( .A1(n9492), .A2(n9491), .ZN(n9490) );
  NAND2_X1 U10281 ( .A1(n9490), .A2(n8867), .ZN(n8868) );
  XNOR2_X1 U10282 ( .A(n8868), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U10283 ( .A1(n8872), .A2(n9489), .ZN(n8869) );
  INV_X1 U10284 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U10285 ( .A1(n9095), .A2(n9083), .ZN(n9079) );
  NAND2_X1 U10286 ( .A1(n9013), .A2(n9194), .ZN(n9001) );
  XNOR2_X1 U10287 ( .A(n9172), .B(n8884), .ZN(n8877) );
  NAND2_X1 U10288 ( .A1(n8877), .A2(n9608), .ZN(n9171) );
  INV_X1 U10289 ( .A(P1_B_REG_SCAN_IN), .ZN(n8879) );
  OAI21_X1 U10290 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8906) );
  OR2_X1 U10291 ( .A1(n8881), .A2(n8906), .ZN(n9173) );
  NOR2_X1 U10292 ( .A1(n9173), .A2(n9616), .ZN(n8886) );
  NOR2_X1 U10293 ( .A1(n9172), .A2(n9605), .ZN(n8882) );
  AOI211_X1 U10294 ( .C1(n9616), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8886), .B(
        n8882), .ZN(n8883) );
  OAI21_X1 U10295 ( .B1(n9171), .B2(n9167), .A(n8883), .ZN(P1_U3263) );
  OAI211_X1 U10296 ( .C1(n8955), .C2(n9175), .A(n9608), .B(n8884), .ZN(n9174)
         );
  NOR2_X1 U10297 ( .A1(n9175), .A2(n9605), .ZN(n8885) );
  AOI211_X1 U10298 ( .C1(n9616), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8886), .B(
        n8885), .ZN(n8887) );
  OAI21_X1 U10299 ( .B1(n9167), .B2(n9174), .A(n8887), .ZN(P1_U3264) );
  INV_X1 U10300 ( .A(n9036), .ZN(n8894) );
  NOR2_X1 U10301 ( .A1(n9037), .A2(n8894), .ZN(n8897) );
  INV_X1 U10302 ( .A(n8895), .ZN(n8896) );
  NAND2_X1 U10303 ( .A1(n9024), .A2(n9023), .ZN(n9022) );
  NAND2_X1 U10304 ( .A1(n9022), .A2(n8898), .ZN(n9008) );
  NAND2_X1 U10305 ( .A1(n9008), .A2(n9009), .ZN(n8991) );
  NOR2_X1 U10306 ( .A1(n8996), .A2(n8899), .ZN(n8901) );
  XNOR2_X1 U10307 ( .A(n8904), .B(n8954), .ZN(n8907) );
  OAI222_X1 U10308 ( .A1(n8908), .A2(n8949), .B1(n8907), .B2(n9596), .C1(n8906), .C2(n8905), .ZN(n9176) );
  OAI22_X1 U10309 ( .A1(n8912), .A2(n8911), .B1(n8910), .B2(n8909), .ZN(n9527)
         );
  AOI21_X1 U10310 ( .B1(n9527), .B2(n9528), .A(n8914), .ZN(n9507) );
  AOI21_X1 U10311 ( .B1(n9377), .B2(n8917), .A(n9154), .ZN(n8918) );
  AOI21_X1 U10312 ( .B1(n9165), .B2(n8919), .A(n8918), .ZN(n9141) );
  OAI22_X1 U10313 ( .A1(n9141), .A2(n9143), .B1(n9150), .B2(n8920), .ZN(n9125)
         );
  NOR2_X1 U10314 ( .A1(n9121), .A2(n8922), .ZN(n8924) );
  NOR2_X1 U10315 ( .A1(n9096), .A2(n8925), .ZN(n8927) );
  NOR2_X1 U10316 ( .A1(n9075), .A2(n8930), .ZN(n8933) );
  NOR2_X1 U10317 ( .A1(n9032), .A2(n8940), .ZN(n8942) );
  NOR2_X1 U10318 ( .A1(n9190), .A2(n8947), .ZN(n8948) );
  NAND2_X1 U10319 ( .A1(n8974), .A2(n8949), .ZN(n8950) );
  NAND2_X1 U10320 ( .A1(n8963), .A2(n8950), .ZN(n8953) );
  NAND2_X1 U10321 ( .A1(n9177), .A2(n9590), .ZN(n8962) );
  AOI211_X1 U10322 ( .C1(n9179), .C2(n8968), .A(n9160), .B(n8955), .ZN(n9178)
         );
  NAND2_X1 U10323 ( .A1(n9179), .A2(n9519), .ZN(n8958) );
  NAND3_X1 U10324 ( .A1(n8956), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n9581), .ZN(
        n8957) );
  OAI211_X1 U10325 ( .C1(n9138), .C2(n8959), .A(n8958), .B(n8957), .ZN(n8960)
         );
  AOI21_X1 U10326 ( .B1(n9178), .B2(n9612), .A(n8960), .ZN(n8961) );
  OAI211_X1 U10327 ( .C1(n9183), .C2(n9616), .A(n8962), .B(n8961), .ZN(
        P1_U3356) );
  XNOR2_X1 U10328 ( .A(n8963), .B(n8964), .ZN(n9254) );
  XOR2_X1 U10329 ( .A(n8964), .B(n4364), .Z(n8967) );
  INV_X1 U10330 ( .A(n8965), .ZN(n8966) );
  OAI21_X1 U10331 ( .B1(n8967), .B2(n9596), .A(n8966), .ZN(n9184) );
  INV_X1 U10332 ( .A(n8978), .ZN(n8970) );
  INV_X1 U10333 ( .A(n8968), .ZN(n8969) );
  AOI211_X1 U10334 ( .C1(n9186), .C2(n8970), .A(n9160), .B(n8969), .ZN(n9185)
         );
  NAND2_X1 U10335 ( .A1(n9185), .A2(n9612), .ZN(n8973) );
  AOI22_X1 U10336 ( .A1(n8971), .A2(n9581), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9616), .ZN(n8972) );
  OAI211_X1 U10337 ( .C1(n8974), .C2(n9605), .A(n8973), .B(n8972), .ZN(n8975)
         );
  AOI21_X1 U10338 ( .B1(n9184), .B2(n9138), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10339 ( .B1(n9254), .B2(n9153), .A(n8976), .ZN(P1_U3265) );
  XOR2_X1 U10340 ( .A(n8977), .B(n8981), .Z(n9257) );
  AOI211_X1 U10341 ( .C1(n9190), .C2(n9001), .A(n9160), .B(n8978), .ZN(n9189)
         );
  OAI22_X1 U10342 ( .A1(n4465), .A2(n9605), .B1(n9138), .B2(n8979), .ZN(n8989)
         );
  AOI21_X1 U10343 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8985) );
  INV_X1 U10344 ( .A(n8983), .ZN(n8984) );
  OAI21_X1 U10345 ( .B1(n8985), .B2(n9596), .A(n8984), .ZN(n9188) );
  AOI21_X1 U10346 ( .B1(n8986), .B2(n9581), .A(n9188), .ZN(n8987) );
  NOR2_X1 U10347 ( .A1(n8987), .A2(n9616), .ZN(n8988) );
  AOI211_X1 U10348 ( .C1(n9189), .C2(n9612), .A(n8989), .B(n8988), .ZN(n8990)
         );
  OAI21_X1 U10349 ( .B1(n9257), .B2(n9153), .A(n8990), .ZN(P1_U3266) );
  NAND2_X1 U10350 ( .A1(n8991), .A2(n8992), .ZN(n8993) );
  XNOR2_X1 U10351 ( .A(n8993), .B(n8996), .ZN(n8995) );
  AOI21_X1 U10352 ( .B1(n8995), .B2(n9579), .A(n8994), .ZN(n9193) );
  XNOR2_X1 U10353 ( .A(n8997), .B(n8996), .ZN(n9261) );
  INV_X1 U10354 ( .A(n9261), .ZN(n8998) );
  NAND2_X1 U10355 ( .A1(n8998), .A2(n9590), .ZN(n9006) );
  OAI22_X1 U10356 ( .A1(n9000), .A2(n9602), .B1(n9138), .B2(n8999), .ZN(n9003)
         );
  OAI211_X1 U10357 ( .C1(n9013), .C2(n9194), .A(n9001), .B(n9608), .ZN(n9192)
         );
  NOR2_X1 U10358 ( .A1(n9192), .A2(n9167), .ZN(n9002) );
  AOI211_X1 U10359 ( .C1(n9519), .C2(n9004), .A(n9003), .B(n9002), .ZN(n9005)
         );
  OAI211_X1 U10360 ( .C1(n9616), .C2(n9193), .A(n9006), .B(n9005), .ZN(
        P1_U3267) );
  XNOR2_X1 U10361 ( .A(n9007), .B(n9009), .ZN(n9265) );
  OAI211_X1 U10362 ( .C1(n9009), .C2(n9008), .A(n8991), .B(n9579), .ZN(n9012)
         );
  INV_X1 U10363 ( .A(n9010), .ZN(n9011) );
  NAND2_X1 U10364 ( .A1(n9012), .A2(n9011), .ZN(n9197) );
  AOI211_X1 U10365 ( .C1(n9199), .C2(n9027), .A(n9160), .B(n9013), .ZN(n9198)
         );
  NAND2_X1 U10366 ( .A1(n9198), .A2(n9612), .ZN(n9017) );
  INV_X1 U10367 ( .A(n9014), .ZN(n9015) );
  AOI22_X1 U10368 ( .A1(n9015), .A2(n9581), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9616), .ZN(n9016) );
  OAI211_X1 U10369 ( .C1(n9018), .C2(n9605), .A(n9017), .B(n9016), .ZN(n9019)
         );
  AOI21_X1 U10370 ( .B1(n9197), .B2(n9138), .A(n9019), .ZN(n9020) );
  OAI21_X1 U10371 ( .B1(n9265), .B2(n9153), .A(n9020), .ZN(P1_U3268) );
  XOR2_X1 U10372 ( .A(n9023), .B(n9021), .Z(n9269) );
  OAI211_X1 U10373 ( .C1(n9024), .C2(n9023), .A(n9022), .B(n9579), .ZN(n9026)
         );
  NAND2_X1 U10374 ( .A1(n9026), .A2(n9025), .ZN(n9202) );
  INV_X1 U10375 ( .A(n9027), .ZN(n9028) );
  AOI211_X1 U10376 ( .C1(n9204), .C2(n4456), .A(n9160), .B(n9028), .ZN(n9203)
         );
  NAND2_X1 U10377 ( .A1(n9203), .A2(n9612), .ZN(n9031) );
  AOI22_X1 U10378 ( .A1(n9616), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9029), .B2(
        n9581), .ZN(n9030) );
  OAI211_X1 U10379 ( .C1(n9032), .C2(n9605), .A(n9031), .B(n9030), .ZN(n9033)
         );
  AOI21_X1 U10380 ( .B1(n9138), .B2(n9202), .A(n9033), .ZN(n9034) );
  OAI21_X1 U10381 ( .B1(n9269), .B2(n9153), .A(n9034), .ZN(P1_U3269) );
  XOR2_X1 U10382 ( .A(n9035), .B(n9037), .Z(n9273) );
  NAND2_X1 U10383 ( .A1(n9057), .A2(n9036), .ZN(n9038) );
  XOR2_X1 U10384 ( .A(n9038), .B(n9037), .Z(n9040) );
  OAI21_X1 U10385 ( .B1(n9040), .B2(n9596), .A(n9039), .ZN(n9207) );
  AOI211_X1 U10386 ( .C1(n9209), .C2(n9049), .A(n9160), .B(n9041), .ZN(n9208)
         );
  NAND2_X1 U10387 ( .A1(n9208), .A2(n9612), .ZN(n9044) );
  AOI22_X1 U10388 ( .A1(n9616), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9042), .B2(
        n9581), .ZN(n9043) );
  OAI211_X1 U10389 ( .C1(n9045), .C2(n9605), .A(n9044), .B(n9043), .ZN(n9046)
         );
  AOI21_X1 U10390 ( .B1(n9207), .B2(n9138), .A(n9046), .ZN(n9047) );
  OAI21_X1 U10391 ( .B1(n9273), .B2(n9153), .A(n9047), .ZN(P1_U3270) );
  XNOR2_X1 U10392 ( .A(n9048), .B(n9058), .ZN(n9277) );
  INV_X1 U10393 ( .A(n9071), .ZN(n9051) );
  INV_X1 U10394 ( .A(n9049), .ZN(n9050) );
  AOI211_X1 U10395 ( .C1(n9213), .C2(n9051), .A(n9160), .B(n9050), .ZN(n9212)
         );
  NOR2_X1 U10396 ( .A1(n9052), .A2(n9605), .ZN(n9056) );
  OAI22_X1 U10397 ( .A1(n9138), .A2(n9054), .B1(n9053), .B2(n9602), .ZN(n9055)
         );
  AOI211_X1 U10398 ( .C1(n9212), .C2(n9612), .A(n9056), .B(n9055), .ZN(n9062)
         );
  OAI211_X1 U10399 ( .C1(n4351), .C2(n9058), .A(n9579), .B(n9057), .ZN(n9060)
         );
  NAND2_X1 U10400 ( .A1(n9060), .A2(n9059), .ZN(n9211) );
  NAND2_X1 U10401 ( .A1(n9211), .A2(n9138), .ZN(n9061) );
  OAI211_X1 U10402 ( .C1(n9277), .C2(n9153), .A(n9062), .B(n9061), .ZN(
        P1_U3271) );
  XNOR2_X1 U10403 ( .A(n9063), .B(n9066), .ZN(n9281) );
  NAND2_X1 U10404 ( .A1(n9065), .A2(n9064), .ZN(n9067) );
  XNOR2_X1 U10405 ( .A(n9067), .B(n9066), .ZN(n9068) );
  NAND2_X1 U10406 ( .A1(n9068), .A2(n9579), .ZN(n9070) );
  NAND2_X1 U10407 ( .A1(n9070), .A2(n9069), .ZN(n9216) );
  AOI211_X1 U10408 ( .C1(n9218), .C2(n9079), .A(n9160), .B(n9071), .ZN(n9217)
         );
  NAND2_X1 U10409 ( .A1(n9217), .A2(n9612), .ZN(n9074) );
  AOI22_X1 U10410 ( .A1(n9616), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9072), .B2(
        n9581), .ZN(n9073) );
  OAI211_X1 U10411 ( .C1(n9075), .C2(n9605), .A(n9074), .B(n9073), .ZN(n9076)
         );
  AOI21_X1 U10412 ( .B1(n9216), .B2(n9138), .A(n9076), .ZN(n9077) );
  OAI21_X1 U10413 ( .B1(n9281), .B2(n9153), .A(n9077), .ZN(P1_U3272) );
  XOR2_X1 U10414 ( .A(n9085), .B(n9078), .Z(n9285) );
  INV_X1 U10415 ( .A(n9095), .ZN(n9081) );
  INV_X1 U10416 ( .A(n9079), .ZN(n9080) );
  AOI211_X1 U10417 ( .C1(n9223), .C2(n9081), .A(n9160), .B(n9080), .ZN(n9222)
         );
  OAI22_X1 U10418 ( .A1(n9083), .A2(n9605), .B1(n9082), .B2(n9138), .ZN(n9084)
         );
  AOI21_X1 U10419 ( .B1(n9222), .B2(n9612), .A(n9084), .ZN(n9093) );
  XNOR2_X1 U10420 ( .A(n9086), .B(n9085), .ZN(n9089) );
  INV_X1 U10421 ( .A(n9087), .ZN(n9088) );
  OAI21_X1 U10422 ( .B1(n9089), .B2(n9596), .A(n9088), .ZN(n9221) );
  NOR2_X1 U10423 ( .A1(n9602), .A2(n9090), .ZN(n9091) );
  OAI21_X1 U10424 ( .B1(n9221), .B2(n9091), .A(n9138), .ZN(n9092) );
  OAI211_X1 U10425 ( .C1(n9285), .C2(n9153), .A(n9093), .B(n9092), .ZN(
        P1_U3273) );
  XNOR2_X1 U10426 ( .A(n9094), .B(n9101), .ZN(n9288) );
  AOI211_X1 U10427 ( .C1(n9228), .C2(n9118), .A(n9160), .B(n9095), .ZN(n9227)
         );
  NOR2_X1 U10428 ( .A1(n9096), .A2(n9605), .ZN(n9100) );
  OAI22_X1 U10429 ( .A1(n9138), .A2(n9098), .B1(n9097), .B2(n9602), .ZN(n9099)
         );
  AOI211_X1 U10430 ( .C1(n9227), .C2(n9612), .A(n9100), .B(n9099), .ZN(n9107)
         );
  XNOR2_X1 U10431 ( .A(n9102), .B(n9101), .ZN(n9105) );
  INV_X1 U10432 ( .A(n9103), .ZN(n9104) );
  OAI21_X1 U10433 ( .B1(n9105), .B2(n9596), .A(n9104), .ZN(n9226) );
  NAND2_X1 U10434 ( .A1(n9226), .A2(n9138), .ZN(n9106) );
  OAI211_X1 U10435 ( .C1(n9288), .C2(n9153), .A(n9107), .B(n9106), .ZN(
        P1_U3274) );
  NAND2_X1 U10436 ( .A1(n9108), .A2(n9109), .ZN(n9110) );
  XNOR2_X1 U10437 ( .A(n9110), .B(n9113), .ZN(n9112) );
  AOI21_X1 U10438 ( .B1(n9112), .B2(n9579), .A(n9111), .ZN(n9232) );
  XOR2_X1 U10439 ( .A(n9114), .B(n9113), .Z(n9291) );
  INV_X1 U10440 ( .A(n9291), .ZN(n9115) );
  NAND2_X1 U10441 ( .A1(n9115), .A2(n9590), .ZN(n9123) );
  OAI22_X1 U10442 ( .A1(n9138), .A2(n9117), .B1(n9116), .B2(n9602), .ZN(n9120)
         );
  OAI211_X1 U10443 ( .C1(n9126), .C2(n9233), .A(n9608), .B(n9118), .ZN(n9231)
         );
  NOR2_X1 U10444 ( .A1(n9231), .A2(n9167), .ZN(n9119) );
  AOI211_X1 U10445 ( .C1(n9519), .C2(n9121), .A(n9120), .B(n9119), .ZN(n9122)
         );
  OAI211_X1 U10446 ( .C1(n9616), .C2(n9232), .A(n9123), .B(n9122), .ZN(
        P1_U3275) );
  XNOR2_X1 U10447 ( .A(n9125), .B(n9124), .ZN(n9241) );
  INV_X1 U10448 ( .A(n9146), .ZN(n9127) );
  AOI211_X1 U10449 ( .C1(n9239), .C2(n9127), .A(n9160), .B(n9126), .ZN(n9238)
         );
  NOR2_X1 U10450 ( .A1(n9128), .A2(n9605), .ZN(n9132) );
  OAI22_X1 U10451 ( .A1(n9138), .A2(n9130), .B1(n9129), .B2(n9602), .ZN(n9131)
         );
  AOI211_X1 U10452 ( .C1(n9238), .C2(n9612), .A(n9132), .B(n9131), .ZN(n9140)
         );
  OAI211_X1 U10453 ( .C1(n9134), .C2(n9133), .A(n9108), .B(n9579), .ZN(n9137)
         );
  INV_X1 U10454 ( .A(n9135), .ZN(n9136) );
  NAND2_X1 U10455 ( .A1(n9137), .A2(n9136), .ZN(n9237) );
  NAND2_X1 U10456 ( .A1(n9237), .A2(n9138), .ZN(n9139) );
  OAI211_X1 U10457 ( .C1(n9241), .C2(n9153), .A(n9140), .B(n9139), .ZN(
        P1_U3276) );
  XNOR2_X1 U10458 ( .A(n9141), .B(n9143), .ZN(n9296) );
  OAI211_X1 U10459 ( .C1(n4383), .C2(n9143), .A(n9142), .B(n9579), .ZN(n9145)
         );
  NAND2_X1 U10460 ( .A1(n9145), .A2(n9144), .ZN(n9242) );
  AOI211_X1 U10461 ( .C1(n9244), .C2(n4376), .A(n9160), .B(n9146), .ZN(n9243)
         );
  NAND2_X1 U10462 ( .A1(n9243), .A2(n9612), .ZN(n9149) );
  AOI22_X1 U10463 ( .A1(n9616), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9147), .B2(
        n9581), .ZN(n9148) );
  OAI211_X1 U10464 ( .C1(n9150), .C2(n9605), .A(n9149), .B(n9148), .ZN(n9151)
         );
  AOI21_X1 U10465 ( .B1(n9242), .B2(n9138), .A(n9151), .ZN(n9152) );
  OAI21_X1 U10466 ( .B1(n9296), .B2(n9153), .A(n9152), .ZN(P1_U3277) );
  XNOR2_X1 U10467 ( .A(n9154), .B(n9156), .ZN(n9379) );
  NAND2_X1 U10468 ( .A1(n9509), .A2(n9155), .ZN(n9157) );
  XNOR2_X1 U10469 ( .A(n9157), .B(n9156), .ZN(n9159) );
  AOI21_X1 U10470 ( .B1(n9159), .B2(n9579), .A(n9158), .ZN(n9376) );
  NOR2_X1 U10471 ( .A1(n9376), .A2(n9616), .ZN(n9169) );
  AOI21_X1 U10472 ( .B1(n9523), .B2(n9165), .A(n9160), .ZN(n9161) );
  NAND2_X1 U10473 ( .A1(n4376), .A2(n9161), .ZN(n9375) );
  NAND2_X1 U10474 ( .A1(n9616), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9162) );
  OAI21_X1 U10475 ( .B1(n9602), .B2(n9163), .A(n9162), .ZN(n9164) );
  AOI21_X1 U10476 ( .B1(n9165), .B2(n9519), .A(n9164), .ZN(n9166) );
  OAI21_X1 U10477 ( .B1(n9375), .B2(n9167), .A(n9166), .ZN(n9168) );
  AOI211_X1 U10478 ( .C1(n9379), .C2(n9590), .A(n9169), .B(n9168), .ZN(n9170)
         );
  INV_X1 U10479 ( .A(n9170), .ZN(P1_U3278) );
  OAI211_X1 U10480 ( .C1(n9172), .C2(n9180), .A(n9171), .B(n9173), .ZN(n9248)
         );
  MUX2_X1 U10481 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9248), .S(n9738), .Z(
        P1_U3553) );
  OAI211_X1 U10482 ( .C1(n9175), .C2(n9180), .A(n9174), .B(n9173), .ZN(n9249)
         );
  MUX2_X1 U10483 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9249), .S(n9738), .Z(
        P1_U3552) );
  INV_X1 U10484 ( .A(n9176), .ZN(n9183) );
  INV_X1 U10485 ( .A(n9178), .ZN(n9182) );
  INV_X1 U10486 ( .A(n9621), .ZN(n9180) );
  MUX2_X1 U10487 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9250), .S(n9738), .Z(
        P1_U3551) );
  INV_X1 U10488 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10016) );
  AOI211_X1 U10489 ( .C1(n9621), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9251)
         );
  MUX2_X1 U10490 ( .A(n10016), .B(n9251), .S(n9738), .Z(n9187) );
  OAI21_X1 U10491 ( .B1(n9254), .B2(n9247), .A(n9187), .ZN(P1_U3550) );
  INV_X1 U10492 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9997) );
  AOI211_X1 U10493 ( .C1(n9621), .C2(n9190), .A(n9189), .B(n9188), .ZN(n9255)
         );
  MUX2_X1 U10494 ( .A(n9997), .B(n9255), .S(n9738), .Z(n9191) );
  OAI21_X1 U10495 ( .B1(n9257), .B2(n9247), .A(n9191), .ZN(P1_U3549) );
  OAI211_X1 U10496 ( .C1(n9194), .C2(n9180), .A(n9193), .B(n9192), .ZN(n9258)
         );
  MUX2_X1 U10497 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9258), .S(n9738), .Z(n9195) );
  INV_X1 U10498 ( .A(n9195), .ZN(n9196) );
  OAI21_X1 U10499 ( .B1(n9261), .B2(n9247), .A(n9196), .ZN(P1_U3548) );
  INV_X1 U10500 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9200) );
  AOI211_X1 U10501 ( .C1(n9621), .C2(n9199), .A(n9198), .B(n9197), .ZN(n9262)
         );
  MUX2_X1 U10502 ( .A(n9200), .B(n9262), .S(n9738), .Z(n9201) );
  OAI21_X1 U10503 ( .B1(n9265), .B2(n9247), .A(n9201), .ZN(P1_U3547) );
  INV_X1 U10504 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9205) );
  AOI211_X1 U10505 ( .C1(n9621), .C2(n9204), .A(n9203), .B(n9202), .ZN(n9266)
         );
  MUX2_X1 U10506 ( .A(n9205), .B(n9266), .S(n9738), .Z(n9206) );
  OAI21_X1 U10507 ( .B1(n9269), .B2(n9247), .A(n9206), .ZN(P1_U3546) );
  AOI211_X1 U10508 ( .C1(n9621), .C2(n9209), .A(n9208), .B(n9207), .ZN(n9270)
         );
  MUX2_X1 U10509 ( .A(n10024), .B(n9270), .S(n9738), .Z(n9210) );
  OAI21_X1 U10510 ( .B1(n9273), .B2(n9247), .A(n9210), .ZN(P1_U3545) );
  AOI211_X1 U10511 ( .C1(n9621), .C2(n9213), .A(n9212), .B(n9211), .ZN(n9274)
         );
  MUX2_X1 U10512 ( .A(n9214), .B(n9274), .S(n9738), .Z(n9215) );
  OAI21_X1 U10513 ( .B1(n9277), .B2(n9247), .A(n9215), .ZN(P1_U3544) );
  INV_X1 U10514 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9219) );
  AOI211_X1 U10515 ( .C1(n9621), .C2(n9218), .A(n9217), .B(n9216), .ZN(n9278)
         );
  MUX2_X1 U10516 ( .A(n9219), .B(n9278), .S(n9738), .Z(n9220) );
  OAI21_X1 U10517 ( .B1(n9281), .B2(n9247), .A(n9220), .ZN(P1_U3543) );
  AOI211_X1 U10518 ( .C1(n9621), .C2(n9223), .A(n9222), .B(n9221), .ZN(n9282)
         );
  MUX2_X1 U10519 ( .A(n9224), .B(n9282), .S(n9738), .Z(n9225) );
  OAI21_X1 U10520 ( .B1(n9285), .B2(n9247), .A(n9225), .ZN(P1_U3542) );
  AOI211_X1 U10521 ( .C1(n9621), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9286)
         );
  MUX2_X1 U10522 ( .A(n9229), .B(n9286), .S(n9738), .Z(n9230) );
  OAI21_X1 U10523 ( .B1(n9288), .B2(n9247), .A(n9230), .ZN(P1_U3541) );
  OAI211_X1 U10524 ( .C1(n9233), .C2(n9180), .A(n9232), .B(n9231), .ZN(n9234)
         );
  INV_X1 U10525 ( .A(n9234), .ZN(n9289) );
  MUX2_X1 U10526 ( .A(n9235), .B(n9289), .S(n9738), .Z(n9236) );
  OAI21_X1 U10527 ( .B1(n9291), .B2(n9247), .A(n9236), .ZN(P1_U3540) );
  AOI211_X1 U10528 ( .C1(n9621), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9240)
         );
  OAI21_X1 U10529 ( .B1(n9241), .B2(n9625), .A(n9240), .ZN(n9292) );
  MUX2_X1 U10530 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9292), .S(n9738), .Z(
        P1_U3539) );
  AOI211_X1 U10531 ( .C1(n9621), .C2(n9244), .A(n9243), .B(n9242), .ZN(n9293)
         );
  MUX2_X1 U10532 ( .A(n9245), .B(n9293), .S(n9738), .Z(n9246) );
  OAI21_X1 U10533 ( .B1(n9296), .B2(n9247), .A(n9246), .ZN(P1_U3538) );
  MUX2_X1 U10534 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9248), .S(n9714), .Z(
        P1_U3521) );
  MUX2_X1 U10535 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9249), .S(n9714), .Z(
        P1_U3520) );
  INV_X1 U10536 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9252) );
  MUX2_X1 U10537 ( .A(n9252), .B(n9251), .S(n9714), .Z(n9253) );
  OAI21_X1 U10538 ( .B1(n9254), .B2(n9295), .A(n9253), .ZN(P1_U3518) );
  INV_X1 U10539 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9888) );
  MUX2_X1 U10540 ( .A(n9888), .B(n9255), .S(n9714), .Z(n9256) );
  OAI21_X1 U10541 ( .B1(n9257), .B2(n9295), .A(n9256), .ZN(P1_U3517) );
  MUX2_X1 U10542 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9258), .S(n9714), .Z(n9259) );
  INV_X1 U10543 ( .A(n9259), .ZN(n9260) );
  OAI21_X1 U10544 ( .B1(n9261), .B2(n9295), .A(n9260), .ZN(P1_U3516) );
  INV_X1 U10545 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9263) );
  MUX2_X1 U10546 ( .A(n9263), .B(n9262), .S(n9714), .Z(n9264) );
  OAI21_X1 U10547 ( .B1(n9265), .B2(n9295), .A(n9264), .ZN(P1_U3515) );
  INV_X1 U10548 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9267) );
  MUX2_X1 U10549 ( .A(n9267), .B(n9266), .S(n9714), .Z(n9268) );
  OAI21_X1 U10550 ( .B1(n9269), .B2(n9295), .A(n9268), .ZN(P1_U3514) );
  MUX2_X1 U10551 ( .A(n9271), .B(n9270), .S(n9714), .Z(n9272) );
  OAI21_X1 U10552 ( .B1(n9273), .B2(n9295), .A(n9272), .ZN(P1_U3513) );
  MUX2_X1 U10553 ( .A(n9275), .B(n9274), .S(n9714), .Z(n9276) );
  OAI21_X1 U10554 ( .B1(n9277), .B2(n9295), .A(n9276), .ZN(P1_U3512) );
  INV_X1 U10555 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9279) );
  MUX2_X1 U10556 ( .A(n9279), .B(n9278), .S(n9714), .Z(n9280) );
  OAI21_X1 U10557 ( .B1(n9281), .B2(n9295), .A(n9280), .ZN(P1_U3511) );
  MUX2_X1 U10558 ( .A(n9283), .B(n9282), .S(n9714), .Z(n9284) );
  OAI21_X1 U10559 ( .B1(n9285), .B2(n9295), .A(n9284), .ZN(P1_U3510) );
  MUX2_X1 U10560 ( .A(n10012), .B(n9286), .S(n9714), .Z(n9287) );
  OAI21_X1 U10561 ( .B1(n9288), .B2(n9295), .A(n9287), .ZN(P1_U3509) );
  MUX2_X1 U10562 ( .A(n10005), .B(n9289), .S(n9714), .Z(n9290) );
  OAI21_X1 U10563 ( .B1(n9291), .B2(n9295), .A(n9290), .ZN(P1_U3507) );
  MUX2_X1 U10564 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9292), .S(n9714), .Z(
        P1_U3504) );
  INV_X1 U10565 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U10566 ( .A(n10003), .B(n9293), .S(n9714), .Z(n9294) );
  OAI21_X1 U10567 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(P1_U3501) );
  MUX2_X1 U10568 ( .A(n9297), .B(P1_D_REG_1__SCAN_IN), .S(n9618), .Z(P1_U3440)
         );
  NOR3_X1 U10569 ( .A1(n9298), .A2(n4899), .A3(P1_U3086), .ZN(n9299) );
  AOI21_X1 U10570 ( .B1(n9300), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9299), .ZN(
        n9301) );
  OAI21_X1 U10571 ( .B1(n9302), .B2(n7231), .A(n9301), .ZN(P1_U3324) );
  OAI222_X1 U10572 ( .A1(P1_U3086), .A2(n4937), .B1(n7231), .B2(n9304), .C1(
        n9303), .C2(n9308), .ZN(P1_U3325) );
  OAI222_X1 U10573 ( .A1(n9308), .A2(n9307), .B1(P1_U3086), .B2(n9306), .C1(
        n9305), .C2(n7231), .ZN(P1_U3326) );
  OAI222_X1 U10574 ( .A1(P1_U3086), .A2(n9311), .B1(n7231), .B2(n9310), .C1(
        n9309), .C2(n9308), .ZN(P1_U3329) );
  MUX2_X1 U10575 ( .A(n9312), .B(n9384), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10576 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9324) );
  AOI211_X1 U10577 ( .C1(n9315), .C2(n9314), .A(n9313), .B(n9476), .ZN(n9320)
         );
  AOI211_X1 U10578 ( .C1(n9318), .C2(n9317), .A(n9316), .B(n9479), .ZN(n9319)
         );
  AOI211_X1 U10579 ( .C1(n9485), .C2(n9321), .A(n9320), .B(n9319), .ZN(n9323)
         );
  NAND2_X1 U10580 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9322) );
  OAI211_X1 U10581 ( .C1(n9506), .C2(n9324), .A(n9323), .B(n9322), .ZN(
        P1_U3253) );
  INV_X1 U10582 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9339) );
  AOI21_X1 U10583 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9328) );
  NAND2_X1 U10584 ( .A1(n9497), .A2(n9328), .ZN(n9334) );
  AOI21_X1 U10585 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9332) );
  NAND2_X1 U10586 ( .A1(n9489), .A2(n9332), .ZN(n9333) );
  OAI211_X1 U10587 ( .C1(n9501), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9336)
         );
  INV_X1 U10588 ( .A(n9336), .ZN(n9338) );
  NAND2_X1 U10589 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9337) );
  OAI211_X1 U10590 ( .C1(n9506), .C2(n9339), .A(n9338), .B(n9337), .ZN(
        P1_U3250) );
  INV_X1 U10591 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9353) );
  INV_X1 U10592 ( .A(n9340), .ZN(n9343) );
  AOI211_X1 U10593 ( .C1(n9343), .C2(n9342), .A(n9341), .B(n9479), .ZN(n9349)
         );
  INV_X1 U10594 ( .A(n9344), .ZN(n9347) );
  AOI211_X1 U10595 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9476), .ZN(n9348)
         );
  AOI211_X1 U10596 ( .C1(n9485), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9352)
         );
  NAND2_X1 U10597 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9351) );
  OAI211_X1 U10598 ( .C1(n9353), .C2(n9506), .A(n9352), .B(n9351), .ZN(
        P1_U3246) );
  AOI21_X1 U10599 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(n9357) );
  NAND2_X1 U10600 ( .A1(n9489), .A2(n9357), .ZN(n9363) );
  AOI21_X1 U10601 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9361) );
  NAND2_X1 U10602 ( .A1(n9497), .A2(n9361), .ZN(n9362) );
  OAI211_X1 U10603 ( .C1(n9501), .C2(n9364), .A(n9363), .B(n9362), .ZN(n9365)
         );
  INV_X1 U10604 ( .A(n9365), .ZN(n9367) );
  NAND2_X1 U10605 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9366) );
  OAI211_X1 U10606 ( .C1(n9506), .C2(n9903), .A(n9367), .B(n9366), .ZN(
        P1_U3251) );
  OR2_X1 U10607 ( .A1(n9368), .A2(n9824), .ZN(n9370) );
  INV_X1 U10608 ( .A(n9373), .ZN(n9371) );
  OAI22_X1 U10609 ( .A1(n9847), .A2(n9371), .B1(P2_REG1_REG_30__SCAN_IN), .B2(
        n9849), .ZN(n9372) );
  INV_X1 U10610 ( .A(n9372), .ZN(P2_U3489) );
  AOI22_X1 U10611 ( .A1(n9886), .A2(n9374), .B1(n9373), .B2(n9884), .ZN(
        P2_U3457) );
  OAI211_X1 U10612 ( .C1(n9377), .C2(n9180), .A(n9376), .B(n9375), .ZN(n9378)
         );
  AOI21_X1 U10613 ( .B1(n9379), .B2(n9702), .A(n9378), .ZN(n9380) );
  AOI22_X1 U10614 ( .A1(n9738), .A2(n9380), .B1(n5321), .B2(n9735), .ZN(
        P1_U3537) );
  AOI22_X1 U10615 ( .A1(n9714), .A2(n9380), .B1(n5322), .B2(n9712), .ZN(
        P1_U3498) );
  XNOR2_X1 U10616 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U10617 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9382), .A(n9381), .ZN(
        n9383) );
  XOR2_X1 U10618 ( .A(n9384), .B(n9383), .Z(n9387) );
  AOI22_X1 U10619 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9400), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9385) );
  OAI21_X1 U10620 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(P1_U3243) );
  AOI21_X1 U10621 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9391) );
  NAND2_X1 U10622 ( .A1(n9489), .A2(n9391), .ZN(n9397) );
  AOI21_X1 U10623 ( .B1(n9394), .B2(n9393), .A(n9392), .ZN(n9395) );
  NAND2_X1 U10624 ( .A1(n9497), .A2(n9395), .ZN(n9396) );
  OAI211_X1 U10625 ( .C1(n9501), .C2(n9398), .A(n9397), .B(n9396), .ZN(n9399)
         );
  INV_X1 U10626 ( .A(n9399), .ZN(n9404) );
  NAND2_X1 U10627 ( .A1(n9400), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9401) );
  NAND4_X1 U10628 ( .A1(n9404), .A2(n9403), .A3(n9402), .A4(n9401), .ZN(
        P1_U3247) );
  INV_X1 U10629 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9418) );
  AOI21_X1 U10630 ( .B1(n9407), .B2(n9406), .A(n9405), .ZN(n9408) );
  NAND2_X1 U10631 ( .A1(n9489), .A2(n9408), .ZN(n9413) );
  AOI21_X1 U10632 ( .B1(n9410), .B2(n4324), .A(n9409), .ZN(n9411) );
  NAND2_X1 U10633 ( .A1(n9497), .A2(n9411), .ZN(n9412) );
  OAI211_X1 U10634 ( .C1(n9501), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9415)
         );
  INV_X1 U10635 ( .A(n9415), .ZN(n9417) );
  OAI211_X1 U10636 ( .C1(n9506), .C2(n9418), .A(n9417), .B(n9416), .ZN(
        P1_U3248) );
  INV_X1 U10637 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9433) );
  AOI21_X1 U10638 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9422) );
  NAND2_X1 U10639 ( .A1(n9497), .A2(n9422), .ZN(n9428) );
  AOI21_X1 U10640 ( .B1(n9425), .B2(n9424), .A(n9423), .ZN(n9426) );
  NAND2_X1 U10641 ( .A1(n9489), .A2(n9426), .ZN(n9427) );
  OAI211_X1 U10642 ( .C1(n9501), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9430)
         );
  INV_X1 U10643 ( .A(n9430), .ZN(n9432) );
  NAND2_X1 U10644 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9431) );
  OAI211_X1 U10645 ( .C1(n9506), .C2(n9433), .A(n9432), .B(n9431), .ZN(
        P1_U3249) );
  INV_X1 U10646 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9448) );
  AOI21_X1 U10647 ( .B1(n9436), .B2(n9435), .A(n9434), .ZN(n9437) );
  NAND2_X1 U10648 ( .A1(n9489), .A2(n9437), .ZN(n9443) );
  AOI21_X1 U10649 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9441) );
  NAND2_X1 U10650 ( .A1(n9497), .A2(n9441), .ZN(n9442) );
  OAI211_X1 U10651 ( .C1(n9501), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9445)
         );
  INV_X1 U10652 ( .A(n9445), .ZN(n9447) );
  NAND2_X1 U10653 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9446) );
  OAI211_X1 U10654 ( .C1(n9506), .C2(n9448), .A(n9447), .B(n9446), .ZN(
        P1_U3254) );
  INV_X1 U10655 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9460) );
  AOI211_X1 U10656 ( .C1(n9451), .C2(n9450), .A(n9449), .B(n9476), .ZN(n9456)
         );
  AOI211_X1 U10657 ( .C1(n9454), .C2(n9453), .A(n9452), .B(n9479), .ZN(n9455)
         );
  AOI211_X1 U10658 ( .C1(n9485), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9459)
         );
  NAND2_X1 U10659 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9458) );
  OAI211_X1 U10660 ( .C1(n9506), .C2(n9460), .A(n9459), .B(n9458), .ZN(
        P1_U3256) );
  INV_X1 U10661 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9475) );
  AOI21_X1 U10662 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  NAND2_X1 U10663 ( .A1(n9497), .A2(n9464), .ZN(n9470) );
  AOI21_X1 U10664 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(n9468) );
  NAND2_X1 U10665 ( .A1(n9489), .A2(n9468), .ZN(n9469) );
  OAI211_X1 U10666 ( .C1(n9501), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9472)
         );
  INV_X1 U10667 ( .A(n9472), .ZN(n9474) );
  NAND2_X1 U10668 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9473) );
  OAI211_X1 U10669 ( .C1(n9506), .C2(n9475), .A(n9474), .B(n9473), .ZN(
        P1_U3257) );
  INV_X1 U10670 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9488) );
  AOI211_X1 U10671 ( .C1(n9478), .C2(n5321), .A(n9477), .B(n9476), .ZN(n9483)
         );
  AOI211_X1 U10672 ( .C1(n9481), .C2(n5323), .A(n9480), .B(n9479), .ZN(n9482)
         );
  AOI211_X1 U10673 ( .C1(n9485), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9487)
         );
  NAND2_X1 U10674 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9486) );
  OAI211_X1 U10675 ( .C1(n9506), .C2(n9488), .A(n9487), .B(n9486), .ZN(
        P1_U3258) );
  OAI211_X1 U10676 ( .C1(n9492), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9499)
         );
  NAND2_X1 U10677 ( .A1(n9494), .A2(n9493), .ZN(n9495) );
  NAND3_X1 U10678 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(n9498) );
  OAI211_X1 U10679 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9502)
         );
  INV_X1 U10680 ( .A(n9502), .ZN(n9504) );
  NAND2_X1 U10681 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9503) );
  OAI211_X1 U10682 ( .C1(n9506), .C2(n9505), .A(n9504), .B(n9503), .ZN(
        P1_U3261) );
  XNOR2_X1 U10683 ( .A(n9507), .B(n9511), .ZN(n9710) );
  INV_X1 U10684 ( .A(n9508), .ZN(n9600) );
  INV_X1 U10685 ( .A(n9509), .ZN(n9514) );
  AOI21_X1 U10686 ( .B1(n9510), .B2(n9512), .A(n9511), .ZN(n9513) );
  NOR3_X1 U10687 ( .A1(n9514), .A2(n9513), .A3(n9596), .ZN(n9517) );
  INV_X1 U10688 ( .A(n9515), .ZN(n9516) );
  AOI211_X1 U10689 ( .C1(n9710), .C2(n9600), .A(n9517), .B(n9516), .ZN(n9707)
         );
  AOI222_X1 U10690 ( .A1(n9520), .A2(n9519), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n9616), .C1(n9581), .C2(n9518), .ZN(n9526) );
  NOR2_X1 U10691 ( .A1(n9616), .A2(n9521), .ZN(n9613) );
  INV_X1 U10692 ( .A(n9522), .ZN(n9532) );
  OAI211_X1 U10693 ( .C1(n9522), .C2(n9706), .A(n9608), .B(n9523), .ZN(n9705)
         );
  INV_X1 U10694 ( .A(n9705), .ZN(n9524) );
  AOI22_X1 U10695 ( .A1(n9710), .A2(n9613), .B1(n9612), .B2(n9524), .ZN(n9525)
         );
  OAI211_X1 U10696 ( .C1(n9616), .C2(n9707), .A(n9526), .B(n9525), .ZN(
        P1_U3279) );
  XNOR2_X1 U10697 ( .A(n9527), .B(n9528), .ZN(n9703) );
  AOI22_X1 U10698 ( .A1(n9703), .A2(n9590), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9616), .ZN(n9539) );
  OAI21_X1 U10699 ( .B1(n4379), .B2(n4529), .A(n9510), .ZN(n9530) );
  AOI21_X1 U10700 ( .B1(n9530), .B2(n9579), .A(n9529), .ZN(n9699) );
  INV_X1 U10701 ( .A(n9699), .ZN(n9537) );
  INV_X1 U10702 ( .A(n9531), .ZN(n9533) );
  OAI211_X1 U10703 ( .C1(n9533), .C2(n9700), .A(n9608), .B(n9532), .ZN(n9698)
         );
  OAI22_X1 U10704 ( .A1(n9698), .A2(n9535), .B1(n9700), .B2(n9534), .ZN(n9536)
         );
  OAI21_X1 U10705 ( .B1(n9537), .B2(n9536), .A(n9138), .ZN(n9538) );
  OAI211_X1 U10706 ( .C1(n9540), .C2(n9602), .A(n9539), .B(n9538), .ZN(
        P1_U3280) );
  XNOR2_X1 U10707 ( .A(n9541), .B(n9544), .ZN(n9672) );
  NAND2_X1 U10708 ( .A1(n9543), .A2(n9542), .ZN(n9545) );
  XNOR2_X1 U10709 ( .A(n9545), .B(n9544), .ZN(n9547) );
  OAI21_X1 U10710 ( .B1(n9547), .B2(n9596), .A(n9546), .ZN(n9548) );
  AOI21_X1 U10711 ( .B1(n9600), .B2(n9672), .A(n9548), .ZN(n9669) );
  NOR2_X1 U10712 ( .A1(n9602), .A2(n9549), .ZN(n9550) );
  AOI21_X1 U10713 ( .B1(n9616), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9550), .ZN(
        n9551) );
  OAI21_X1 U10714 ( .B1(n9605), .B2(n9668), .A(n9551), .ZN(n9552) );
  INV_X1 U10715 ( .A(n9552), .ZN(n9558) );
  INV_X1 U10716 ( .A(n9553), .ZN(n9555) );
  OAI211_X1 U10717 ( .C1(n9555), .C2(n9668), .A(n9608), .B(n9554), .ZN(n9667)
         );
  INV_X1 U10718 ( .A(n9667), .ZN(n9556) );
  AOI22_X1 U10719 ( .A1(n9672), .A2(n9613), .B1(n9612), .B2(n9556), .ZN(n9557)
         );
  OAI211_X1 U10720 ( .C1(n9616), .C2(n9669), .A(n9558), .B(n9557), .ZN(
        P1_U3285) );
  NAND2_X1 U10721 ( .A1(n9560), .A2(n9559), .ZN(n9561) );
  XOR2_X1 U10722 ( .A(n9568), .B(n9561), .Z(n9563) );
  AOI21_X1 U10723 ( .B1(n9563), .B2(n9579), .A(n9562), .ZN(n9656) );
  AOI22_X1 U10724 ( .A1(n9616), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9564), .B2(
        n9581), .ZN(n9565) );
  OAI21_X1 U10725 ( .B1(n9605), .B2(n9655), .A(n9565), .ZN(n9566) );
  INV_X1 U10726 ( .A(n9566), .ZN(n9575) );
  XNOR2_X1 U10727 ( .A(n9567), .B(n9568), .ZN(n9659) );
  INV_X1 U10728 ( .A(n9569), .ZN(n9572) );
  INV_X1 U10729 ( .A(n9570), .ZN(n9571) );
  OAI211_X1 U10730 ( .C1(n9655), .C2(n9572), .A(n9571), .B(n9608), .ZN(n9654)
         );
  INV_X1 U10731 ( .A(n9654), .ZN(n9573) );
  AOI22_X1 U10732 ( .A1(n9659), .A2(n9590), .B1(n9612), .B2(n9573), .ZN(n9574)
         );
  OAI211_X1 U10733 ( .C1(n9616), .C2(n9656), .A(n9575), .B(n9574), .ZN(
        P1_U3287) );
  XNOR2_X1 U10734 ( .A(n9576), .B(n9586), .ZN(n9580) );
  INV_X1 U10735 ( .A(n9577), .ZN(n9578) );
  AOI21_X1 U10736 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(n9643) );
  AOI22_X1 U10737 ( .A1(n9616), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9582), .B2(
        n9581), .ZN(n9583) );
  OAI21_X1 U10738 ( .B1(n9605), .B2(n9642), .A(n9583), .ZN(n9584) );
  INV_X1 U10739 ( .A(n9584), .ZN(n9592) );
  XNOR2_X1 U10740 ( .A(n9585), .B(n9586), .ZN(n9646) );
  OAI211_X1 U10741 ( .C1(n4445), .C2(n9642), .A(n9608), .B(n9588), .ZN(n9641)
         );
  INV_X1 U10742 ( .A(n9641), .ZN(n9589) );
  AOI22_X1 U10743 ( .A1(n9646), .A2(n9590), .B1(n9612), .B2(n9589), .ZN(n9591)
         );
  OAI211_X1 U10744 ( .C1(n9616), .C2(n9643), .A(n9592), .B(n9591), .ZN(
        P1_U3289) );
  XNOR2_X1 U10745 ( .A(n9593), .B(n9594), .ZN(n9633) );
  XNOR2_X1 U10746 ( .A(n9595), .B(n9594), .ZN(n9597) );
  NOR2_X1 U10747 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  AOI211_X1 U10748 ( .C1(n9633), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9630)
         );
  NOR2_X1 U10749 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  AOI21_X1 U10750 ( .B1(n9616), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9603), .ZN(
        n9604) );
  OAI21_X1 U10751 ( .B1(n9605), .B2(n9629), .A(n9604), .ZN(n9606) );
  INV_X1 U10752 ( .A(n9606), .ZN(n9615) );
  INV_X1 U10753 ( .A(n9607), .ZN(n9609) );
  OAI211_X1 U10754 ( .C1(n9629), .C2(n9610), .A(n9609), .B(n9608), .ZN(n9628)
         );
  INV_X1 U10755 ( .A(n9628), .ZN(n9611) );
  AOI22_X1 U10756 ( .A1(n9633), .A2(n9613), .B1(n9612), .B2(n9611), .ZN(n9614)
         );
  OAI211_X1 U10757 ( .C1(n9616), .C2(n9630), .A(n9615), .B(n9614), .ZN(
        P1_U3291) );
  AND2_X1 U10758 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9618), .ZN(P1_U3294) );
  AND2_X1 U10759 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9618), .ZN(P1_U3295) );
  AND2_X1 U10760 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9618), .ZN(P1_U3296) );
  AND2_X1 U10761 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9618), .ZN(P1_U3297) );
  AND2_X1 U10762 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9618), .ZN(P1_U3298) );
  AND2_X1 U10763 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9618), .ZN(P1_U3299) );
  AND2_X1 U10764 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9618), .ZN(P1_U3300) );
  AND2_X1 U10765 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9618), .ZN(P1_U3301) );
  AND2_X1 U10766 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9618), .ZN(P1_U3302) );
  AND2_X1 U10767 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9618), .ZN(P1_U3303) );
  AND2_X1 U10768 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9618), .ZN(P1_U3304) );
  AND2_X1 U10769 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9618), .ZN(P1_U3305) );
  INV_X1 U10770 ( .A(n9618), .ZN(n9617) );
  INV_X1 U10771 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10004) );
  NOR2_X1 U10772 ( .A1(n9617), .A2(n10004), .ZN(P1_U3306) );
  AND2_X1 U10773 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9618), .ZN(P1_U3307) );
  AND2_X1 U10774 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9618), .ZN(P1_U3308) );
  AND2_X1 U10775 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9618), .ZN(P1_U3309) );
  AND2_X1 U10776 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9618), .ZN(P1_U3310) );
  AND2_X1 U10777 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9618), .ZN(P1_U3311) );
  AND2_X1 U10778 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9618), .ZN(P1_U3312) );
  INV_X1 U10779 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U10780 ( .A1(n9617), .A2(n9944), .ZN(P1_U3313) );
  AND2_X1 U10781 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9618), .ZN(P1_U3314) );
  AND2_X1 U10782 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9618), .ZN(P1_U3315) );
  AND2_X1 U10783 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9618), .ZN(P1_U3316) );
  AND2_X1 U10784 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9618), .ZN(P1_U3317) );
  AND2_X1 U10785 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9618), .ZN(P1_U3318) );
  AND2_X1 U10786 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9618), .ZN(P1_U3319) );
  AND2_X1 U10787 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9618), .ZN(P1_U3320) );
  INV_X1 U10788 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U10789 ( .A1(n9617), .A2(n9905), .ZN(P1_U3321) );
  AND2_X1 U10790 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9618), .ZN(P1_U3322) );
  AND2_X1 U10791 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9618), .ZN(P1_U3323) );
  AOI21_X1 U10792 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9623) );
  OAI211_X1 U10793 ( .C1(n9625), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9626)
         );
  INV_X1 U10794 ( .A(n9626), .ZN(n9716) );
  INV_X1 U10795 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U10796 ( .A1(n9714), .A2(n9716), .B1(n9947), .B2(n9712), .ZN(
        P1_U3456) );
  INV_X1 U10797 ( .A(n9627), .ZN(n9711) );
  OAI21_X1 U10798 ( .B1(n9629), .B2(n9180), .A(n9628), .ZN(n9632) );
  INV_X1 U10799 ( .A(n9630), .ZN(n9631) );
  AOI211_X1 U10800 ( .C1(n9711), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9718)
         );
  INV_X1 U10801 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9634) );
  AOI22_X1 U10802 ( .A1(n9714), .A2(n9718), .B1(n9634), .B2(n9712), .ZN(
        P1_U3459) );
  INV_X1 U10803 ( .A(n9635), .ZN(n9640) );
  OAI21_X1 U10804 ( .B1(n9637), .B2(n9180), .A(n9636), .ZN(n9639) );
  AOI211_X1 U10805 ( .C1(n9702), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9719)
         );
  AOI22_X1 U10806 ( .A1(n9714), .A2(n9719), .B1(n4993), .B2(n9712), .ZN(
        P1_U3462) );
  OAI21_X1 U10807 ( .B1(n9642), .B2(n9180), .A(n9641), .ZN(n9645) );
  INV_X1 U10808 ( .A(n9643), .ZN(n9644) );
  AOI211_X1 U10809 ( .C1(n9702), .C2(n9646), .A(n9645), .B(n9644), .ZN(n9721)
         );
  INV_X1 U10810 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U10811 ( .A1(n9714), .A2(n9721), .B1(n9972), .B2(n9712), .ZN(
        P1_U3465) );
  AND2_X1 U10812 ( .A1(n9647), .A2(n9702), .ZN(n9651) );
  OAI21_X1 U10813 ( .B1(n9649), .B2(n9180), .A(n9648), .ZN(n9650) );
  NOR3_X1 U10814 ( .A1(n9652), .A2(n9651), .A3(n9650), .ZN(n9723) );
  INV_X1 U10815 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9653) );
  AOI22_X1 U10816 ( .A1(n9714), .A2(n9723), .B1(n9653), .B2(n9712), .ZN(
        P1_U3468) );
  OAI21_X1 U10817 ( .B1(n9655), .B2(n9180), .A(n9654), .ZN(n9658) );
  INV_X1 U10818 ( .A(n9656), .ZN(n9657) );
  AOI211_X1 U10819 ( .C1(n9702), .C2(n9659), .A(n9658), .B(n9657), .ZN(n9724)
         );
  INV_X1 U10820 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U10821 ( .A1(n9714), .A2(n9724), .B1(n9943), .B2(n9712), .ZN(
        P1_U3471) );
  AND2_X1 U10822 ( .A1(n9660), .A2(n9702), .ZN(n9664) );
  OAI21_X1 U10823 ( .B1(n9662), .B2(n9180), .A(n9661), .ZN(n9663) );
  NOR3_X1 U10824 ( .A1(n9665), .A2(n9664), .A3(n9663), .ZN(n9726) );
  INV_X1 U10825 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U10826 ( .A1(n9714), .A2(n9726), .B1(n9666), .B2(n9712), .ZN(
        P1_U3474) );
  OAI21_X1 U10827 ( .B1(n9668), .B2(n9180), .A(n9667), .ZN(n9671) );
  INV_X1 U10828 ( .A(n9669), .ZN(n9670) );
  AOI211_X1 U10829 ( .C1(n9711), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9727)
         );
  AOI22_X1 U10830 ( .A1(n9714), .A2(n9727), .B1(n10025), .B2(n9712), .ZN(
        P1_U3477) );
  AND2_X1 U10831 ( .A1(n9673), .A2(n9702), .ZN(n9677) );
  OAI21_X1 U10832 ( .B1(n9675), .B2(n9180), .A(n9674), .ZN(n9676) );
  NOR3_X1 U10833 ( .A1(n9678), .A2(n9677), .A3(n9676), .ZN(n9728) );
  INV_X1 U10834 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U10835 ( .A1(n9714), .A2(n9728), .B1(n9679), .B2(n9712), .ZN(
        P1_U3480) );
  OAI211_X1 U10836 ( .C1(n9682), .C2(n9180), .A(n9681), .B(n9680), .ZN(n9683)
         );
  AOI21_X1 U10837 ( .B1(n9684), .B2(n9702), .A(n9683), .ZN(n9730) );
  INV_X1 U10838 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9685) );
  AOI22_X1 U10839 ( .A1(n9714), .A2(n9730), .B1(n9685), .B2(n9712), .ZN(
        P1_U3483) );
  OAI211_X1 U10840 ( .C1(n9688), .C2(n9180), .A(n9687), .B(n9686), .ZN(n9689)
         );
  AOI21_X1 U10841 ( .B1(n9690), .B2(n9702), .A(n9689), .ZN(n9731) );
  INV_X1 U10842 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9691) );
  AOI22_X1 U10843 ( .A1(n9714), .A2(n9731), .B1(n9691), .B2(n9712), .ZN(
        P1_U3486) );
  OAI21_X1 U10844 ( .B1(n9693), .B2(n9180), .A(n9692), .ZN(n9694) );
  AOI211_X1 U10845 ( .C1(n9696), .C2(n9702), .A(n9695), .B(n9694), .ZN(n9733)
         );
  INV_X1 U10846 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9697) );
  AOI22_X1 U10847 ( .A1(n9714), .A2(n9733), .B1(n9697), .B2(n9712), .ZN(
        P1_U3489) );
  OAI211_X1 U10848 ( .C1(n9700), .C2(n9180), .A(n9699), .B(n9698), .ZN(n9701)
         );
  AOI21_X1 U10849 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9734) );
  INV_X1 U10850 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U10851 ( .A1(n9714), .A2(n9734), .B1(n9704), .B2(n9712), .ZN(
        P1_U3492) );
  OAI21_X1 U10852 ( .B1(n9706), .B2(n9180), .A(n9705), .ZN(n9709) );
  INV_X1 U10853 ( .A(n9707), .ZN(n9708) );
  AOI211_X1 U10854 ( .C1(n9711), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9737)
         );
  INV_X1 U10855 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U10856 ( .A1(n9714), .A2(n9737), .B1(n9713), .B2(n9712), .ZN(
        P1_U3495) );
  AOI22_X1 U10857 ( .A1(n9738), .A2(n9716), .B1(n9715), .B2(n9735), .ZN(
        P1_U3523) );
  AOI22_X1 U10858 ( .A1(n9738), .A2(n9718), .B1(n9717), .B2(n9735), .ZN(
        P1_U3524) );
  AOI22_X1 U10859 ( .A1(n9738), .A2(n9719), .B1(n4990), .B2(n9735), .ZN(
        P1_U3525) );
  INV_X1 U10860 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10861 ( .A1(n9738), .A2(n9721), .B1(n9720), .B2(n9735), .ZN(
        P1_U3526) );
  INV_X1 U10862 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9722) );
  AOI22_X1 U10863 ( .A1(n9738), .A2(n9723), .B1(n9722), .B2(n9735), .ZN(
        P1_U3527) );
  AOI22_X1 U10864 ( .A1(n9738), .A2(n9724), .B1(n6556), .B2(n9735), .ZN(
        P1_U3528) );
  INV_X1 U10865 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10866 ( .A1(n9738), .A2(n9726), .B1(n9725), .B2(n9735), .ZN(
        P1_U3529) );
  AOI22_X1 U10867 ( .A1(n9738), .A2(n9727), .B1(n5129), .B2(n9735), .ZN(
        P1_U3530) );
  INV_X1 U10868 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U10869 ( .A1(n9738), .A2(n9728), .B1(n9958), .B2(n9735), .ZN(
        P1_U3531) );
  INV_X1 U10870 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U10871 ( .A1(n9738), .A2(n9730), .B1(n9729), .B2(n9735), .ZN(
        P1_U3532) );
  AOI22_X1 U10872 ( .A1(n9738), .A2(n9731), .B1(n6564), .B2(n9735), .ZN(
        P1_U3533) );
  AOI22_X1 U10873 ( .A1(n9738), .A2(n9733), .B1(n9732), .B2(n9735), .ZN(
        P1_U3534) );
  AOI22_X1 U10874 ( .A1(n9738), .A2(n9734), .B1(n8818), .B2(n9735), .ZN(
        P1_U3535) );
  AOI22_X1 U10875 ( .A1(n9738), .A2(n9737), .B1(n9736), .B2(n9735), .ZN(
        P1_U3536) );
  INV_X1 U10876 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9901) );
  AOI21_X1 U10877 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9748) );
  OAI21_X1 U10878 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(n9745) );
  AOI22_X1 U10879 ( .A1(n9746), .A2(n9745), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n9747) );
  OAI21_X1 U10880 ( .B1(n9748), .B2(n9762), .A(n9747), .ZN(n9749) );
  AOI21_X1 U10881 ( .B1(n9750), .B2(n9767), .A(n9749), .ZN(n9755) );
  XOR2_X1 U10882 ( .A(n9752), .B(n9751), .Z(n9753) );
  NAND2_X1 U10883 ( .A1(n9774), .A2(n9753), .ZN(n9754) );
  OAI211_X1 U10884 ( .C1(n9901), .C2(n9779), .A(n9755), .B(n9754), .ZN(
        P2_U3184) );
  AOI21_X1 U10885 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9770) );
  AOI21_X1 U10886 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(n9763) );
  NOR2_X1 U10887 ( .A1(n9763), .A2(n9762), .ZN(n9764) );
  AOI211_X1 U10888 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9768)
         );
  OAI21_X1 U10889 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(n9771) );
  INV_X1 U10890 ( .A(n9771), .ZN(n9778) );
  NOR2_X1 U10891 ( .A1(n9773), .A2(n9772), .ZN(n9775) );
  OAI21_X1 U10892 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9777) );
  OAI211_X1 U10893 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9777), .ZN(
        P2_U3190) );
  AOI22_X1 U10894 ( .A1(n9886), .A2(n9782), .B1(n9781), .B2(n9884), .ZN(
        P2_U3390) );
  NOR2_X1 U10895 ( .A1(n9783), .A2(n9824), .ZN(n9785) );
  AOI211_X1 U10896 ( .C1(n9791), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9831)
         );
  AOI22_X1 U10897 ( .A1(n9886), .A2(n5743), .B1(n9831), .B2(n9884), .ZN(
        P2_U3393) );
  INV_X1 U10898 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9792) );
  INV_X1 U10899 ( .A(n9787), .ZN(n9788) );
  AOI211_X1 U10900 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9832)
         );
  AOI22_X1 U10901 ( .A1(n9886), .A2(n9792), .B1(n9832), .B2(n9884), .ZN(
        P2_U3396) );
  INV_X1 U10902 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9798) );
  INV_X1 U10903 ( .A(n9793), .ZN(n9797) );
  OAI21_X1 U10904 ( .B1(n9795), .B2(n9824), .A(n9794), .ZN(n9796) );
  AOI21_X1 U10905 ( .B1(n9797), .B2(n9807), .A(n9796), .ZN(n9833) );
  AOI22_X1 U10906 ( .A1(n9886), .A2(n9798), .B1(n9833), .B2(n9884), .ZN(
        P2_U3399) );
  INV_X1 U10907 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9802) );
  OAI21_X1 U10908 ( .B1(n4595), .B2(n9824), .A(n9799), .ZN(n9800) );
  AOI21_X1 U10909 ( .B1(n9801), .B2(n9807), .A(n9800), .ZN(n9835) );
  AOI22_X1 U10910 ( .A1(n9886), .A2(n9802), .B1(n9835), .B2(n9884), .ZN(
        P2_U3402) );
  INV_X1 U10911 ( .A(n9803), .ZN(n9808) );
  OAI21_X1 U10912 ( .B1(n9805), .B2(n9824), .A(n9804), .ZN(n9806) );
  AOI21_X1 U10913 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9843) );
  AOI22_X1 U10914 ( .A1(n9886), .A2(n5830), .B1(n9843), .B2(n9884), .ZN(
        P2_U3408) );
  INV_X1 U10915 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9813) );
  OAI22_X1 U10916 ( .A1(n9810), .A2(n9826), .B1(n9809), .B2(n9824), .ZN(n9811)
         );
  NOR2_X1 U10917 ( .A1(n9812), .A2(n9811), .ZN(n9844) );
  AOI22_X1 U10918 ( .A1(n9886), .A2(n9813), .B1(n9844), .B2(n9884), .ZN(
        P2_U3411) );
  INV_X1 U10919 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9818) );
  OAI22_X1 U10920 ( .A1(n9815), .A2(n9841), .B1(n9814), .B2(n9824), .ZN(n9816)
         );
  NOR2_X1 U10921 ( .A1(n9817), .A2(n9816), .ZN(n9845) );
  AOI22_X1 U10922 ( .A1(n9886), .A2(n9818), .B1(n9845), .B2(n9884), .ZN(
        P2_U3414) );
  INV_X1 U10923 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9823) );
  OAI22_X1 U10924 ( .A1(n9820), .A2(n9826), .B1(n9819), .B2(n9824), .ZN(n9821)
         );
  NOR2_X1 U10925 ( .A1(n9822), .A2(n9821), .ZN(n9846) );
  AOI22_X1 U10926 ( .A1(n9886), .A2(n9823), .B1(n9846), .B2(n9884), .ZN(
        P2_U3417) );
  INV_X1 U10927 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9830) );
  OAI22_X1 U10928 ( .A1(n9827), .A2(n9826), .B1(n9825), .B2(n9824), .ZN(n9828)
         );
  NOR2_X1 U10929 ( .A1(n9829), .A2(n9828), .ZN(n9848) );
  AOI22_X1 U10930 ( .A1(n9886), .A2(n9830), .B1(n9848), .B2(n9884), .ZN(
        P2_U3420) );
  AOI22_X1 U10931 ( .A1(n9849), .A2(n9831), .B1(n5740), .B2(n9847), .ZN(
        P2_U3460) );
  AOI22_X1 U10932 ( .A1(n9849), .A2(n9832), .B1(n9946), .B2(n9847), .ZN(
        P2_U3461) );
  AOI22_X1 U10933 ( .A1(n9849), .A2(n9833), .B1(n6413), .B2(n9847), .ZN(
        P2_U3462) );
  AOI22_X1 U10934 ( .A1(n9849), .A2(n9835), .B1(n9834), .B2(n9847), .ZN(
        P2_U3463) );
  NAND2_X1 U10935 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  OAI211_X1 U10936 ( .C1(n9841), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9885)
         );
  OAI22_X1 U10937 ( .A1(n9847), .A2(n9885), .B1(P2_REG1_REG_5__SCAN_IN), .B2(
        n9849), .ZN(n9842) );
  INV_X1 U10938 ( .A(n9842), .ZN(P2_U3464) );
  AOI22_X1 U10939 ( .A1(n9849), .A2(n9843), .B1(n6432), .B2(n9847), .ZN(
        P2_U3465) );
  AOI22_X1 U10940 ( .A1(n9849), .A2(n9844), .B1(n6470), .B2(n9847), .ZN(
        P2_U3466) );
  AOI22_X1 U10941 ( .A1(n9849), .A2(n9845), .B1(n5863), .B2(n9847), .ZN(
        P2_U3467) );
  AOI22_X1 U10942 ( .A1(n9849), .A2(n9846), .B1(n6836), .B2(n9847), .ZN(
        P2_U3468) );
  AOI22_X1 U10943 ( .A1(n9849), .A2(n9848), .B1(n5892), .B2(n9847), .ZN(
        P2_U3469) );
  OAI222_X1 U10944 ( .A1(n9854), .A2(n9853), .B1(n9854), .B2(n9852), .C1(n9851), .C2(n9850), .ZN(ADD_1068_U5) );
  XOR2_X1 U10945 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U10946 ( .A(n9857), .ZN(n9856) );
  OAI222_X1 U10947 ( .A1(n9859), .A2(n9858), .B1(n9859), .B2(n9857), .C1(n9856), .C2(n9855), .ZN(ADD_1068_U55) );
  OAI21_X1 U10948 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(ADD_1068_U56) );
  OAI21_X1 U10949 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(ADD_1068_U57) );
  OAI21_X1 U10950 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(ADD_1068_U58) );
  OAI21_X1 U10951 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(ADD_1068_U59) );
  OAI21_X1 U10952 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(ADD_1068_U60) );
  OAI21_X1 U10953 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(ADD_1068_U61) );
  OAI21_X1 U10954 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(ADD_1068_U62) );
  OAI21_X1 U10955 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(ADD_1068_U63) );
  AOI22_X1 U10956 ( .A1(n9886), .A2(P2_REG0_REG_5__SCAN_IN), .B1(n9885), .B2(
        n9884), .ZN(n10042) );
  AOI22_X1 U10957 ( .A1(n9888), .A2(keyinput37), .B1(n9997), .B2(keyinput3), 
        .ZN(n9887) );
  OAI221_X1 U10958 ( .B1(n9888), .B2(keyinput37), .C1(n9997), .C2(keyinput3), 
        .A(n9887), .ZN(n9899) );
  AOI22_X1 U10959 ( .A1(n9890), .A2(keyinput63), .B1(keyinput23), .B2(n9996), 
        .ZN(n9889) );
  OAI221_X1 U10960 ( .B1(n9890), .B2(keyinput63), .C1(n9996), .C2(keyinput23), 
        .A(n9889), .ZN(n9898) );
  INV_X1 U10961 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10962 ( .A1(n9893), .A2(keyinput60), .B1(n9892), .B2(keyinput22), 
        .ZN(n9891) );
  OAI221_X1 U10963 ( .B1(n9893), .B2(keyinput60), .C1(n9892), .C2(keyinput22), 
        .A(n9891), .ZN(n9897) );
  XOR2_X1 U10964 ( .A(n4993), .B(keyinput52), .Z(n9895) );
  XNOR2_X1 U10965 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput30), .ZN(n9894) );
  NAND2_X1 U10966 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NOR4_X1 U10967 ( .A1(n9899), .A2(n9898), .A3(n9897), .A4(n9896), .ZN(n9939)
         );
  AOI22_X1 U10968 ( .A1(n8979), .A2(keyinput48), .B1(keyinput11), .B2(n9901), 
        .ZN(n9900) );
  OAI221_X1 U10969 ( .B1(n8979), .B2(keyinput48), .C1(n9901), .C2(keyinput11), 
        .A(n9900), .ZN(n9912) );
  AOI22_X1 U10970 ( .A1(n9903), .A2(keyinput15), .B1(n5321), .B2(keyinput50), 
        .ZN(n9902) );
  OAI221_X1 U10971 ( .B1(n9903), .B2(keyinput15), .C1(n5321), .C2(keyinput50), 
        .A(n9902), .ZN(n9911) );
  AOI22_X1 U10972 ( .A1(n9906), .A2(keyinput13), .B1(n9905), .B2(keyinput41), 
        .ZN(n9904) );
  OAI221_X1 U10973 ( .B1(n9906), .B2(keyinput13), .C1(n9905), .C2(keyinput41), 
        .A(n9904), .ZN(n9910) );
  XOR2_X1 U10974 ( .A(n7005), .B(keyinput12), .Z(n9908) );
  XNOR2_X1 U10975 ( .A(SI_2_), .B(keyinput6), .ZN(n9907) );
  NAND2_X1 U10976 ( .A1(n9908), .A2(n9907), .ZN(n9909) );
  NOR4_X1 U10977 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9938)
         );
  AOI22_X1 U10978 ( .A1(n10012), .A2(keyinput8), .B1(keyinput7), .B2(n10001), 
        .ZN(n9913) );
  OAI221_X1 U10979 ( .B1(n10012), .B2(keyinput8), .C1(n10001), .C2(keyinput7), 
        .A(n9913), .ZN(n9924) );
  AOI22_X1 U10980 ( .A1(n9915), .A2(keyinput53), .B1(keyinput55), .B2(n6413), 
        .ZN(n9914) );
  OAI221_X1 U10981 ( .B1(n9915), .B2(keyinput53), .C1(n6413), .C2(keyinput55), 
        .A(n9914), .ZN(n9923) );
  AOI22_X1 U10982 ( .A1(n9918), .A2(keyinput35), .B1(keyinput20), .B2(n9917), 
        .ZN(n9916) );
  OAI221_X1 U10983 ( .B1(n9918), .B2(keyinput35), .C1(n9917), .C2(keyinput20), 
        .A(n9916), .ZN(n9922) );
  XNOR2_X1 U10984 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput34), .ZN(n9920) );
  XNOR2_X1 U10985 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput58), .ZN(n9919)
         );
  NAND2_X1 U10986 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  NOR4_X1 U10987 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(n9937)
         );
  AOI22_X1 U10988 ( .A1(n10006), .A2(keyinput14), .B1(n10025), .B2(keyinput5), 
        .ZN(n9925) );
  OAI221_X1 U10989 ( .B1(n10006), .B2(keyinput14), .C1(n10025), .C2(keyinput5), 
        .A(n9925), .ZN(n9935) );
  AOI22_X1 U10990 ( .A1(n9927), .A2(keyinput32), .B1(n10002), .B2(keyinput10), 
        .ZN(n9926) );
  OAI221_X1 U10991 ( .B1(n9927), .B2(keyinput32), .C1(n10002), .C2(keyinput10), 
        .A(n9926), .ZN(n9934) );
  INV_X1 U10992 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9928) );
  XOR2_X1 U10993 ( .A(n9928), .B(keyinput62), .Z(n9932) );
  XNOR2_X1 U10994 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput31), .ZN(n9931) );
  XNOR2_X1 U10995 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput17), .ZN(n9930) );
  XNOR2_X1 U10996 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput42), .ZN(n9929) );
  NAND4_X1 U10997 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9933)
         );
  NOR3_X1 U10998 ( .A1(n9935), .A2(n9934), .A3(n9933), .ZN(n9936) );
  NAND4_X1 U10999 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(n9995)
         );
  AOI22_X1 U11000 ( .A1(n9941), .A2(keyinput28), .B1(n5350), .B2(keyinput57), 
        .ZN(n9940) );
  OAI221_X1 U11001 ( .B1(n9941), .B2(keyinput28), .C1(n5350), .C2(keyinput57), 
        .A(n9940), .ZN(n9953) );
  AOI22_X1 U11002 ( .A1(n9944), .A2(keyinput2), .B1(keyinput26), .B2(n9943), 
        .ZN(n9942) );
  OAI221_X1 U11003 ( .B1(n9944), .B2(keyinput2), .C1(n9943), .C2(keyinput26), 
        .A(n9942), .ZN(n9952) );
  AOI22_X1 U11004 ( .A1(n9947), .A2(keyinput27), .B1(keyinput21), .B2(n9946), 
        .ZN(n9945) );
  OAI221_X1 U11005 ( .B1(n9947), .B2(keyinput27), .C1(n9946), .C2(keyinput21), 
        .A(n9945), .ZN(n9951) );
  AOI22_X1 U11006 ( .A1(n5323), .A2(keyinput0), .B1(keyinput45), .B2(n9949), 
        .ZN(n9948) );
  OAI221_X1 U11007 ( .B1(n5323), .B2(keyinput0), .C1(n9949), .C2(keyinput45), 
        .A(n9948), .ZN(n9950) );
  NOR4_X1 U11008 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9993)
         );
  INV_X1 U11009 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11010 ( .A1(n9956), .A2(keyinput40), .B1(keyinput18), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11011 ( .B1(n9956), .B2(keyinput40), .C1(n9955), .C2(keyinput18), 
        .A(n9954), .ZN(n9967) );
  AOI22_X1 U11012 ( .A1(n6421), .A2(keyinput24), .B1(n9958), .B2(keyinput49), 
        .ZN(n9957) );
  OAI221_X1 U11013 ( .B1(n6421), .B2(keyinput24), .C1(n9958), .C2(keyinput49), 
        .A(n9957), .ZN(n9966) );
  INV_X1 U11014 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U11015 ( .A1(n9961), .A2(keyinput29), .B1(n9960), .B2(keyinput19), 
        .ZN(n9959) );
  OAI221_X1 U11016 ( .B1(n9961), .B2(keyinput29), .C1(n9960), .C2(keyinput19), 
        .A(n9959), .ZN(n9965) );
  XNOR2_X1 U11017 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput1), .ZN(n9963) );
  XNOR2_X1 U11018 ( .A(P1_REG1_REG_28__SCAN_IN), .B(keyinput59), .ZN(n9962) );
  NAND2_X1 U11019 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  NOR4_X1 U11020 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n9992)
         );
  AOI22_X1 U11021 ( .A1(n10011), .A2(keyinput61), .B1(keyinput16), .B2(n6226), 
        .ZN(n9968) );
  OAI221_X1 U11022 ( .B1(n10011), .B2(keyinput61), .C1(n6226), .C2(keyinput16), 
        .A(n9968), .ZN(n9978) );
  INV_X1 U11023 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10010) );
  INV_X1 U11024 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11025 ( .A1(n10010), .A2(keyinput33), .B1(n9970), .B2(keyinput44), 
        .ZN(n9969) );
  OAI221_X1 U11026 ( .B1(n10010), .B2(keyinput33), .C1(n9970), .C2(keyinput44), 
        .A(n9969), .ZN(n9977) );
  INV_X1 U11027 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10023) );
  AOI22_X1 U11028 ( .A1(n10024), .A2(keyinput51), .B1(keyinput46), .B2(n10023), 
        .ZN(n9971) );
  OAI221_X1 U11029 ( .B1(n10024), .B2(keyinput51), .C1(n10023), .C2(keyinput46), .A(n9971), .ZN(n9976) );
  XOR2_X1 U11030 ( .A(n9972), .B(keyinput9), .Z(n9974) );
  XNOR2_X1 U11031 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput39), .ZN(n9973) );
  NAND2_X1 U11032 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  NOR4_X1 U11033 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n9991)
         );
  INV_X1 U11034 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U11035 ( .A1(n5743), .A2(keyinput36), .B1(keyinput4), .B2(n9998), 
        .ZN(n9979) );
  OAI221_X1 U11036 ( .B1(n5743), .B2(keyinput36), .C1(n9998), .C2(keyinput4), 
        .A(n9979), .ZN(n9989) );
  AOI22_X1 U11037 ( .A1(n9981), .A2(keyinput25), .B1(n10004), .B2(keyinput54), 
        .ZN(n9980) );
  OAI221_X1 U11038 ( .B1(n9981), .B2(keyinput25), .C1(n10004), .C2(keyinput54), 
        .A(n9980), .ZN(n9988) );
  INV_X1 U11039 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11040 ( .A1(n9983), .A2(keyinput56), .B1(keyinput43), .B2(n10005), 
        .ZN(n9982) );
  OAI221_X1 U11041 ( .B1(n9983), .B2(keyinput56), .C1(n10005), .C2(keyinput43), 
        .A(n9982), .ZN(n9987) );
  XOR2_X1 U11042 ( .A(n10003), .B(keyinput38), .Z(n9985) );
  XNOR2_X1 U11043 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput47), .ZN(n9984) );
  NAND2_X1 U11044 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  NOR4_X1 U11045 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n9990)
         );
  NAND4_X1 U11046 ( .A1(n9993), .A2(n9992), .A3(n9991), .A4(n9990), .ZN(n9994)
         );
  NOR2_X1 U11047 ( .A1(n9995), .A2(n9994), .ZN(n10040) );
  NOR4_X1 U11048 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_REG0_REG_3__SCAN_IN), 
        .A3(P2_REG0_REG_29__SCAN_IN), .A4(n7005), .ZN(n10038) );
  NOR4_X1 U11049 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(P1_REG0_REG_27__SCAN_IN), 
        .A3(n9997), .A4(n9996), .ZN(n10037) );
  NAND4_X1 U11050 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .A4(n9998), .ZN(n10000) );
  NAND2_X1 U11051 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P1_REG1_REG_15__SCAN_IN), 
        .ZN(n9999) );
  NOR4_X1 U11052 ( .A1(SI_25_), .A2(P2_D_REG_1__SCAN_IN), .A3(n10000), .A4(
        n9999), .ZN(n10036) );
  NOR4_X1 U11053 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .A3(n10002), .A4(n10001), .ZN(n10034) );
  NOR4_X1 U11054 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10005), .A3(n10004), 
        .A4(n10003), .ZN(n10033) );
  NAND4_X1 U11055 ( .A1(n10006), .A2(n5904), .A3(P1_RD_REG_SCAN_IN), .A4(
        P2_REG3_REG_6__SCAN_IN), .ZN(n10009) );
  NAND4_X1 U11056 ( .A1(n10007), .A2(P2_REG2_REG_4__SCAN_IN), .A3(
        P1_DATAO_REG_6__SCAN_IN), .A4(P1_IR_REG_30__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U11057 ( .A1(n10009), .A2(n10008), .ZN(n10029) );
  NOR2_X1 U11058 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n10022) );
  NOR4_X1 U11059 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(P1_REG2_REG_14__SCAN_IN), 
        .A3(n10011), .A4(n10010), .ZN(n10015) );
  NOR4_X1 U11060 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n10012), .ZN(n10014) );
  NOR4_X1 U11061 ( .A1(SI_2_), .A2(P2_REG1_REG_2__SCAN_IN), .A3(
        P2_REG0_REG_1__SCAN_IN), .A4(n6413), .ZN(n10013) );
  NAND3_X1 U11062 ( .A1(n10015), .A2(n10014), .A3(n10013), .ZN(n10020) );
  NOR4_X1 U11063 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(P1_REG2_REG_15__SCAN_IN), 
        .A3(P1_REG0_REG_1__SCAN_IN), .A4(P2_REG3_REG_25__SCAN_IN), .ZN(n10018)
         );
  NOR4_X1 U11064 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(P1_REG0_REG_6__SCAN_IN), .A4(n10016), .ZN(n10017) );
  NAND2_X1 U11065 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  NOR2_X1 U11066 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND4_X1 U11067 ( .A1(n10022), .A2(P2_IR_REG_26__SCAN_IN), .A3(n10021), .A4(
        n9903), .ZN(n10027) );
  NAND4_X1 U11068 ( .A1(n9972), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10026) );
  NOR2_X1 U11069 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  AND4_X1 U11070 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10032) );
  AND3_X1 U11071 ( .A1(n10034), .A2(n10033), .A3(n10032), .ZN(n10035) );
  NAND4_X1 U11072 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10039) );
  XNOR2_X1 U11073 ( .A(n10040), .B(n10039), .ZN(n10041) );
  XNOR2_X1 U11074 ( .A(n10042), .B(n10041), .ZN(P2_U3405) );
  OAI21_X1 U11075 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(ADD_1068_U50) );
  OAI21_X1 U11076 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(ADD_1068_U51) );
  OAI21_X1 U11077 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(ADD_1068_U47) );
  OAI21_X1 U11078 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(ADD_1068_U49) );
  OAI21_X1 U11079 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(ADD_1068_U48) );
  AOI21_X1 U11080 ( .B1(n10060), .B2(n10059), .A(n10058), .ZN(ADD_1068_U54) );
  AOI21_X1 U11081 ( .B1(n10063), .B2(n10062), .A(n10061), .ZN(ADD_1068_U53) );
  OAI21_X1 U11082 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(ADD_1068_U52) );
  OR2_X1 U7296 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  INV_X1 U4805 ( .A(n7519), .ZN(n7535) );
  AND2_X2 U4838 ( .A1(n5548), .A2(n4299), .ZN(n4982) );
  INV_X2 U4841 ( .A(n5550), .ZN(n5456) );
  CLKBUF_X1 U4884 ( .A(n4992), .Z(n5645) );
  CLKBUF_X1 U5035 ( .A(n4952), .Z(n8615) );
  NAND2_X1 U5043 ( .A1(n5229), .A2(n5228), .ZN(n8448) );
endmodule

