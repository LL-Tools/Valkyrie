

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657;

  CLKBUF_X1 U3403 ( .A(n4403), .Z(n2980) );
  CLKBUF_X2 U3404 ( .A(n3143), .Z(n3865) );
  OR2_X1 U3406 ( .A1(n3189), .A2(n6634), .ZN(n3984) );
  CLKBUF_X2 U3407 ( .A(n3173), .Z(n3867) );
  BUF_X2 U3408 ( .A(n3149), .Z(n3302) );
  AND4_X2 U3409 ( .A1(n4218), .A2(n3202), .A3(n4032), .A4(n2975), .ZN(n2966)
         );
  CLKBUF_X2 U3410 ( .A(n3325), .Z(n3278) );
  CLKBUF_X1 U3411 ( .A(n3150), .Z(n3372) );
  CLKBUF_X2 U3412 ( .A(n3859), .Z(n3846) );
  CLKBUF_X1 U3413 ( .A(n3206), .Z(n3207) );
  AND4_X1 U3414 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n3090)
         );
  AND2_X1 U3415 ( .A1(n3075), .A2(n4408), .ZN(n3149) );
  INV_X1 U3416 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3066) );
  AND2_X4 U3417 ( .A1(n3069), .A2(n4430), .ZN(n3325) );
  AND2_X1 U3419 ( .A1(n4463), .A2(n3443), .ZN(n3055) );
  AOI22_X1 U3420 ( .A1(n6605), .A2(keyinput20), .B1(keyinput46), .B2(n6604), 
        .ZN(n6603) );
  AOI22_X1 U3421 ( .A1(n6572), .A2(keyinput53), .B1(keyinput36), .B2(n6571), 
        .ZN(n6570) );
  OR2_X1 U3422 ( .A1(n3990), .A2(n2965), .ZN(n4249) );
  AND2_X1 U3423 ( .A1(n4083), .A2(n4748), .ZN(n3205) );
  INV_X1 U3424 ( .A(n4180), .ZN(n4172) );
  OAI221_X1 U3425 ( .B1(n6605), .B2(keyinput20), .C1(n6604), .C2(keyinput46), 
        .A(n6603), .ZN(n6613) );
  OAI221_X1 U3426 ( .B1(n6572), .B2(keyinput53), .C1(n6571), .C2(keyinput36), 
        .A(n6570), .ZN(n6585) );
  AND2_X1 U3427 ( .A1(n4083), .A2(n3203), .ZN(n3887) );
  INV_X1 U3428 ( .A(n4527), .ZN(n2967) );
  NAND2_X1 U3429 ( .A1(n2966), .A2(n3203), .ZN(n4070) );
  NAND2_X1 U3430 ( .A1(n3341), .A2(n3340), .ZN(n4463) );
  NAND2_X1 U3431 ( .A1(n4029), .A2(n4028), .ZN(n4865) );
  INV_X1 U3432 ( .A(n5564), .ZN(n5555) );
  INV_X1 U3434 ( .A(n6282), .ZN(n5774) );
  AND2_X2 U3435 ( .A1(n4856), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4851)
         );
  INV_X1 U3436 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6634) );
  INV_X1 U3437 ( .A(n5612), .ZN(n5607) );
  INV_X1 U3438 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3067) );
  INV_X1 U3439 ( .A(n4527), .ZN(n3189) );
  INV_X1 U3440 ( .A(n5616), .ZN(n2955) );
  INV_X1 U3441 ( .A(n2955), .ZN(n2956) );
  INV_X1 U3442 ( .A(n4460), .ZN(n3404) );
  NAND2_X2 U3443 ( .A1(n3938), .A2(n3937), .ZN(n4687) );
  AND4_X2 U3444 ( .A1(n3119), .A2(n3120), .A3(n3118), .A4(n3117), .ZN(n3121)
         );
  NAND2_X2 U34450 ( .A1(n4936), .A2(n3050), .ZN(n4065) );
  AND2_X4 U34460 ( .A1(n4937), .A2(n4938), .ZN(n4936) );
  AND2_X2 U34470 ( .A1(n2960), .A2(n4694), .ZN(n3554) );
  OAI21_X2 U34480 ( .B1(n4780), .B2(n4778), .A(n4776), .ZN(n4812) );
  NAND2_X2 U3449 ( .A1(n2969), .A2(n2963), .ZN(n4780) );
  NAND2_X4 U3450 ( .A1(n3951), .A2(n3950), .ZN(n5414) );
  XNOR2_X1 U34510 ( .A(n4062), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5221)
         );
  BUF_X1 U34520 ( .A(n3884), .Z(n4890) );
  NAND2_X1 U34530 ( .A1(n3471), .A2(n3470), .ZN(n4622) );
  NAND2_X1 U3454 ( .A1(n5414), .A2(n3955), .ZN(n3957) );
  NOR2_X2 U34550 ( .A1(n4561), .A2(n4748), .ZN(n6280) );
  NAND2_X1 U34560 ( .A1(n4073), .A2(n3209), .ZN(n4235) );
  INV_X1 U3457 ( .A(n3201), .ZN(n2957) );
  INV_X2 U3458 ( .A(n4111), .ZN(n4185) );
  INV_X2 U34600 ( .A(n4748), .ZN(n3203) );
  BUF_X2 U34610 ( .A(n3326), .Z(n3743) );
  INV_X2 U34620 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4856) );
  OR2_X1 U34630 ( .A1(n4302), .A2(n5766), .ZN(n4060) );
  MUX2_X1 U34640 ( .A(n5113), .B(n4061), .S(INSTADDRPOINTER_REG_27__SCAN_IN), 
        .Z(n4062) );
  NOR3_X1 U34650 ( .A1(n5134), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4044), .ZN(n4045) );
  NAND2_X1 U3466 ( .A1(n5134), .A2(n3014), .ZN(n4215) );
  OR2_X1 U3467 ( .A1(n5090), .A2(n6282), .ZN(n4067) );
  AND2_X1 U34680 ( .A1(n5133), .A2(n5135), .ZN(n4043) );
  NAND2_X1 U34690 ( .A1(n5151), .A2(n3968), .ZN(n3024) );
  CLKBUF_X1 U34700 ( .A(n5026), .Z(n5027) );
  NAND2_X1 U34710 ( .A1(n5034), .A2(n5035), .ZN(n5026) );
  NAND2_X1 U34720 ( .A1(n4812), .A2(n2985), .ZN(n3005) );
  NAND2_X1 U34730 ( .A1(n4694), .A2(n3057), .ZN(n4733) );
  NOR2_X2 U34740 ( .A1(n4622), .A2(n4698), .ZN(n4694) );
  AOI21_X1 U3475 ( .B1(n2985), .B2(n3008), .A(n2991), .ZN(n3006) );
  AND2_X1 U3476 ( .A1(n3007), .A2(n3963), .ZN(n2985) );
  AND2_X1 U3477 ( .A1(n4453), .A2(n4484), .ZN(n4483) );
  OR2_X1 U3478 ( .A1(n4811), .A2(n3008), .ZN(n3007) );
  AND2_X1 U3479 ( .A1(n3442), .A2(n2962), .ZN(n4453) );
  NAND2_X1 U3480 ( .A1(n3918), .A2(n3917), .ZN(n4443) );
  AOI21_X1 U3481 ( .B1(n3404), .B2(n3592), .A(n4049), .ZN(n4355) );
  NAND2_X1 U3482 ( .A1(n3915), .A2(n3914), .ZN(n3916) );
  NOR2_X1 U3483 ( .A1(n3456), .A2(n3367), .ZN(n3383) );
  NAND2_X1 U3484 ( .A1(n3056), .A2(n3055), .ZN(n3456) );
  NAND2_X1 U3485 ( .A1(n4322), .A2(n4323), .ZN(n4353) );
  NAND2_X1 U3486 ( .A1(n3412), .A2(n3411), .ZN(n4322) );
  MUX2_X1 U3487 ( .A(n3422), .B(n4364), .S(n4363), .Z(n4323) );
  AND2_X1 U3488 ( .A1(n3317), .A2(n3398), .ZN(n3318) );
  CLKBUF_X1 U3489 ( .A(n4462), .Z(n6283) );
  NAND2_X1 U3490 ( .A1(n3418), .A2(n3417), .ZN(n6163) );
  XNOR2_X1 U3491 ( .A(n3408), .B(n3407), .ZN(n4462) );
  NAND2_X1 U3492 ( .A1(n3413), .A2(n3291), .ZN(n3406) );
  AND2_X1 U3493 ( .A1(n3216), .A2(n3292), .ZN(n2973) );
  NAND2_X1 U3494 ( .A1(n3323), .A2(n3322), .ZN(n6170) );
  AOI21_X1 U3495 ( .B1(n3320), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3237), 
        .ZN(n3238) );
  NAND2_X1 U3496 ( .A1(n3255), .A2(n3256), .ZN(n3292) );
  OAI211_X1 U3497 ( .C1(n4070), .C2(n3210), .A(n4282), .B(n4235), .ZN(n3211)
         );
  AND4_X1 U3498 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3231)
         );
  AND3_X1 U3499 ( .A1(n3314), .A2(n3313), .A3(n3312), .ZN(n3397) );
  AND2_X1 U3500 ( .A1(n3197), .A2(n4249), .ZN(n3230) );
  INV_X1 U3501 ( .A(n4013), .ZN(n3379) );
  MUX2_X1 U3502 ( .A(n3310), .B(n3286), .S(n3285), .Z(n3416) );
  OR2_X1 U3503 ( .A1(n4251), .A2(n4228), .ZN(n4282) );
  NAND2_X1 U3504 ( .A1(n2957), .A2(n3142), .ZN(n3599) );
  NOR2_X1 U3505 ( .A1(n3288), .A2(n6634), .ZN(n3286) );
  NAND3_X1 U3506 ( .A1(n3203), .A2(n2967), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4013) );
  NAND2_X1 U3507 ( .A1(n3196), .A2(n4527), .ZN(n3222) );
  OR2_X1 U3508 ( .A1(n3270), .A2(n3269), .ZN(n3952) );
  OR2_X1 U3509 ( .A1(n3308), .A2(n3307), .ZN(n3899) );
  NOR2_X1 U3510 ( .A1(n4562), .A2(n4082), .ZN(n4329) );
  OR2_X1 U3511 ( .A1(n3284), .A2(n3283), .ZN(n3900) );
  INV_X1 U3512 ( .A(n4562), .ZN(n4240) );
  AND4_X2 U3514 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n4527)
         );
  AND4_X2 U3515 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n4748)
         );
  NAND2_X2 U3516 ( .A1(n3140), .A2(n3141), .ZN(n4306) );
  NAND2_X1 U3517 ( .A1(n3064), .A2(n3131), .ZN(n4562) );
  AND4_X1 U3518 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3140)
         );
  AND4_X1 U3519 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3141)
         );
  AND4_X1 U3520 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3081)
         );
  AND4_X1 U3521 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3080)
         );
  AND4_X1 U3522 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n3109)
         );
  AND4_X1 U3523 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3183)
         );
  AND4_X1 U3524 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3185)
         );
  AND4_X1 U3525 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3110)
         );
  AND4_X1 U3526 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3065)
         );
  AND4_X1 U3527 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3111)
         );
  AND4_X1 U3528 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  AND4_X1 U3529 ( .A1(n3095), .A2(n3094), .A3(n3093), .A4(n3092), .ZN(n3112)
         );
  AND4_X1 U3530 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3184)
         );
  BUF_X2 U3531 ( .A(n3245), .Z(n3333) );
  CLKBUF_X1 U3532 ( .A(n3148), .Z(n3859) );
  INV_X2 U3533 ( .A(n5672), .ZN(n5663) );
  BUF_X2 U3534 ( .A(n3295), .Z(n3332) );
  INV_X1 U3535 ( .A(n4035), .ZN(n3321) );
  AND2_X1 U3536 ( .A1(n4327), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3200)
         );
  BUF_X2 U3537 ( .A(n3297), .Z(n3866) );
  NAND2_X2 U3538 ( .A1(n3886), .A2(n6290), .ZN(n6282) );
  BUF_X2 U3539 ( .A(n3276), .Z(n3868) );
  AND2_X1 U3540 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3450), .ZN(n3457)
         );
  BUF_X2 U3541 ( .A(n3277), .Z(n3860) );
  BUF_X2 U3542 ( .A(n3346), .Z(n2958) );
  AND2_X1 U3543 ( .A1(n3066), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3069)
         );
  AND2_X1 U3544 ( .A1(n6468), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4030) );
  AND2_X1 U3545 ( .A1(n3067), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4409)
         );
  AND2_X4 U3546 ( .A1(n4847), .A2(n4430), .ZN(n3151) );
  AND2_X1 U3547 ( .A1(n3067), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2964)
         );
  NOR2_X1 U3548 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3070) );
  AND2_X1 U3549 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4407) );
  INV_X1 U3550 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6466) );
  AND2_X1 U3551 ( .A1(n3631), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3632)
         );
  INV_X1 U3552 ( .A(n3057), .ZN(n2959) );
  NOR2_X1 U3553 ( .A1(n4741), .A2(n2959), .ZN(n2960) );
  INV_X1 U3554 ( .A(n5026), .ZN(n2961) );
  NOR2_X1 U3555 ( .A1(n4472), .A2(n4454), .ZN(n2962) );
  AOI21_X1 U3556 ( .B1(n4891), .B2(n4065), .A(n4890), .ZN(n5110) );
  AND2_X1 U3557 ( .A1(n2970), .A2(n5740), .ZN(n2963) );
  NAND2_X1 U3558 ( .A1(n4527), .A2(n4082), .ZN(n2965) );
  INV_X1 U3559 ( .A(n3990), .ZN(n3196) );
  NAND2_X1 U3560 ( .A1(n3195), .A2(n4306), .ZN(n3990) );
  OR2_X1 U3561 ( .A1(n3194), .A2(n4831), .ZN(n2968) );
  NAND2_X1 U3562 ( .A1(n2968), .A2(n3887), .ZN(n3197) );
  NOR2_X4 U3563 ( .A1(n2979), .A2(n4748), .ZN(n4334) );
  AND2_X1 U3564 ( .A1(n3232), .A2(n3216), .ZN(n3294) );
  AND2_X1 U3565 ( .A1(n3292), .A2(n3259), .ZN(n6052) );
  NAND3_X1 U3566 ( .A1(n3199), .A2(n3198), .A3(n3230), .ZN(n3217) );
  NAND2_X1 U3567 ( .A1(n3004), .A2(n2972), .ZN(n2969) );
  OR2_X1 U3568 ( .A1(n2971), .A2(n4725), .ZN(n2970) );
  INV_X1 U3569 ( .A(n5739), .ZN(n2971) );
  AND2_X1 U3570 ( .A1(n3002), .A2(n5739), .ZN(n2972) );
  NAND2_X1 U3571 ( .A1(n3232), .A2(n2973), .ZN(n3233) );
  NAND2_X1 U3572 ( .A1(n3948), .A2(n3947), .ZN(n2974) );
  INV_X1 U3573 ( .A(n3201), .ZN(n2975) );
  NAND2_X1 U3574 ( .A1(n3442), .A2(n3441), .ZN(n4452) );
  NAND2_X2 U3575 ( .A1(n4818), .A2(n4820), .ZN(n4819) );
  AND2_X2 U3576 ( .A1(n5073), .A2(n5072), .ZN(n4818) );
  NAND2_X1 U3577 ( .A1(n3921), .A2(n3920), .ZN(n2976) );
  NAND2_X1 U3578 ( .A1(n3010), .A2(n3009), .ZN(n2977) );
  NAND2_X1 U3579 ( .A1(n3921), .A2(n3920), .ZN(n4592) );
  NAND2_X1 U3580 ( .A1(n3010), .A2(n3009), .ZN(n5169) );
  CLKBUF_X1 U3581 ( .A(n4421), .Z(n2981) );
  NAND2_X2 U3582 ( .A1(n3959), .A2(n3001), .ZN(n3004) );
  NOR2_X1 U3583 ( .A1(n4043), .A2(n3972), .ZN(n5126) );
  XNOR2_X2 U3584 ( .A(n3294), .B(n3293), .ZN(n4495) );
  NAND2_X2 U3585 ( .A1(n5189), .A2(n3967), .ZN(n5151) );
  INV_X2 U3586 ( .A(n4217), .ZN(n3202) );
  AOI21_X1 U3587 ( .B1(n6163), .B2(n2957), .A(n3391), .ZN(n4364) );
  NAND2_X2 U3588 ( .A1(n3932), .A2(n3931), .ZN(n4552) );
  NAND2_X1 U3589 ( .A1(n3961), .A2(n4725), .ZN(n5741) );
  NAND2_X2 U3590 ( .A1(n3206), .A2(n3204), .ZN(n4328) );
  NAND2_X2 U3591 ( .A1(n3385), .A2(n3158), .ZN(n3201) );
  NAND2_X4 U3592 ( .A1(n3065), .A2(n3121), .ZN(n3158) );
  INV_X1 U3593 ( .A(n3433), .ZN(n3056) );
  OR2_X2 U3594 ( .A1(n5139), .A2(n5138), .ZN(n5182) );
  OAI21_X1 U3595 ( .B1(n3890), .B2(n3990), .A(n3889), .ZN(n3919) );
  OAI21_X1 U3596 ( .B1(n6163), .B2(n3990), .A(n3897), .ZN(n5778) );
  OAI22_X2 U3597 ( .A1(n4421), .A2(STATE2_REG_0__SCAN_IN), .B1(n3891), .B2(
        n3984), .ZN(n3254) );
  NAND2_X2 U3598 ( .A1(n3005), .A2(n3006), .ZN(n5197) );
  AND2_X4 U3599 ( .A1(n4414), .A2(n4408), .ZN(n3143) );
  NAND2_X2 U3600 ( .A1(n3433), .A2(n3403), .ZN(n4460) );
  XNOR2_X2 U3601 ( .A(n3433), .B(n4463), .ZN(n3911) );
  XNOR2_X2 U3602 ( .A(n3916), .B(n4371), .ZN(n4367) );
  OAI22_X2 U3603 ( .A1(n5154), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5165), .B2(n5143), .ZN(n5144) );
  OAI21_X4 U3604 ( .B1(n5197), .B2(n3966), .A(n3965), .ZN(n5189) );
  XNOR2_X1 U3605 ( .A(n3319), .B(n6170), .ZN(n4403) );
  AND2_X1 U3606 ( .A1(n3075), .A2(n4408), .ZN(n2982) );
  AND2_X1 U3607 ( .A1(n3075), .A2(n4408), .ZN(n2983) );
  AND2_X2 U3608 ( .A1(n4959), .A2(n3046), .ZN(n5034) );
  NOR2_X4 U3609 ( .A1(n4819), .A2(n4970), .ZN(n4959) );
  BUF_X1 U3610 ( .A(n3911), .Z(n2984) );
  NAND2_X1 U3611 ( .A1(n3053), .A2(n5006), .ZN(n3052) );
  NOR2_X1 U3612 ( .A1(n4912), .A2(n3054), .ZN(n3053) );
  INV_X1 U3613 ( .A(n4923), .ZN(n3054) );
  OR2_X1 U3614 ( .A1(n6343), .A2(n6634), .ZN(n3880) );
  OAI21_X1 U3615 ( .B1(n4460), .B2(n3990), .A(n3894), .ZN(n3907) );
  OR2_X1 U3616 ( .A1(n4185), .A2(n4186), .ZN(n4178) );
  INV_X1 U3617 ( .A(n4334), .ZN(n4186) );
  NOR2_X1 U3618 ( .A1(n5055), .A2(n5051), .ZN(n5038) );
  INV_X1 U3619 ( .A(n6163), .ZN(n6233) );
  OR2_X1 U3620 ( .A1(n4027), .A2(n4076), .ZN(n4028) );
  NAND2_X1 U3621 ( .A1(n4024), .A2(n4023), .ZN(n4029) );
  NAND2_X1 U3622 ( .A1(n3354), .A2(n3353), .ZN(n3443) );
  XNOR2_X1 U3623 ( .A(n3456), .B(n3455), .ZN(n3922) );
  AND2_X1 U3624 ( .A1(n3716), .A2(n3698), .ZN(n3045) );
  AND2_X1 U3625 ( .A1(n3648), .A2(n4960), .ZN(n3048) );
  NOR2_X1 U3626 ( .A1(n3158), .A2(n3391), .ZN(n3419) );
  INV_X1 U3627 ( .A(n3969), .ZN(n3023) );
  NOR2_X1 U3628 ( .A1(n3036), .A2(n3039), .ZN(n3035) );
  INV_X1 U3629 ( .A(n4723), .ZN(n3039) );
  INV_X1 U3630 ( .A(n3037), .ZN(n3036) );
  INV_X1 U3631 ( .A(n4103), .ZN(n4183) );
  NOR2_X1 U3632 ( .A1(n4373), .A2(n3027), .ZN(n3026) );
  INV_X1 U3633 ( .A(n4358), .ZN(n3027) );
  OR2_X1 U3634 ( .A1(n4082), .A2(n4748), .ZN(n4180) );
  NAND2_X1 U3635 ( .A1(n3063), .A2(n3415), .ZN(n3291) );
  INV_X1 U3636 ( .A(n3397), .ZN(n3405) );
  NAND2_X1 U3637 ( .A1(n3324), .A2(n3984), .ZN(n4020) );
  INV_X1 U3638 ( .A(n4030), .ZN(n4327) );
  OR2_X1 U3639 ( .A1(n6196), .A2(n3235), .ZN(n4543) );
  NOR2_X1 U3640 ( .A1(n4013), .A2(n3990), .ZN(n4025) );
  NAND2_X1 U3641 ( .A1(n4196), .A2(n4227), .ZN(n5597) );
  OR3_X1 U3642 ( .A1(n6484), .A2(n6375), .A3(n4080), .ZN(n5616) );
  NAND2_X1 U3643 ( .A1(n4916), .A2(n3011), .ZN(n4876) );
  AND2_X1 U3644 ( .A1(n4901), .A2(n4275), .ZN(n3011) );
  AND2_X1 U3645 ( .A1(n4916), .A2(n4901), .ZN(n4877) );
  NOR2_X1 U3646 ( .A1(n2987), .A2(n4914), .ZN(n4916) );
  AND2_X1 U3647 ( .A1(n3615), .A2(n3614), .ZN(n4970) );
  INV_X1 U3648 ( .A(n3854), .ZN(n4050) );
  NOR2_X1 U3649 ( .A1(n3052), .A2(n3051), .ZN(n3050) );
  INV_X1 U3650 ( .A(n4066), .ZN(n3051) );
  INV_X1 U3651 ( .A(n3052), .ZN(n3049) );
  NAND2_X1 U3652 ( .A1(n3776), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3793)
         );
  INV_X1 U3653 ( .A(n5028), .ZN(n3698) );
  AND2_X1 U3654 ( .A1(n3058), .A2(n3533), .ZN(n3057) );
  INV_X1 U3655 ( .A(n4735), .ZN(n3533) );
  INV_X1 U3656 ( .A(n3907), .ZN(n3909) );
  AND2_X1 U3657 ( .A1(n4865), .A2(n4839), .ZN(n4609) );
  INV_X1 U3658 ( .A(n3015), .ZN(n3013) );
  AND2_X1 U3659 ( .A1(n5171), .A2(n2993), .ZN(n3009) );
  NAND2_X1 U3660 ( .A1(n5139), .A2(n5138), .ZN(n5181) );
  NAND2_X1 U3661 ( .A1(n5070), .A2(n2994), .ZN(n5055) );
  INV_X1 U3662 ( .A(n4962), .ZN(n3028) );
  NOR2_X1 U3663 ( .A1(n3033), .A2(n3030), .ZN(n3029) );
  INV_X1 U3664 ( .A(n4978), .ZN(n3033) );
  INV_X1 U3665 ( .A(n3031), .ZN(n3030) );
  NOR2_X1 U3666 ( .A1(n4803), .A2(n4804), .ZN(n5070) );
  NAND2_X1 U3667 ( .A1(n4812), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U3668 ( .A1(n4774), .A2(n4775), .ZN(n4803) );
  NOR2_X1 U3669 ( .A1(n3003), .A2(n4726), .ZN(n3002) );
  INV_X1 U3670 ( .A(n3960), .ZN(n3003) );
  NOR2_X1 U3671 ( .A1(n4101), .A2(n4100), .ZN(n4357) );
  NAND2_X1 U3672 ( .A1(n3406), .A2(n3407), .ZN(n3399) );
  OR2_X1 U3673 ( .A1(n4460), .A2(n4461), .ZN(n6225) );
  NAND2_X1 U3674 ( .A1(n6283), .A2(n6233), .ZN(n6128) );
  NOR2_X1 U3675 ( .A1(n6225), .A2(n6283), .ZN(n6204) );
  NAND2_X1 U3676 ( .A1(n6634), .A2(n4502), .ZN(n6024) );
  NAND2_X1 U3677 ( .A1(n4333), .A2(n4332), .ZN(n5076) );
  OR2_X1 U3678 ( .A1(n4399), .A2(n6385), .ZN(n4333) );
  INV_X1 U3679 ( .A(n3158), .ZN(n4831) );
  AND2_X1 U3680 ( .A1(n5081), .A2(n4834), .ZN(n5633) );
  AND2_X1 U3681 ( .A1(n5081), .A2(n5080), .ZN(n5637) );
  AND2_X1 U3682 ( .A1(n5081), .A2(n4612), .ZN(n5102) );
  AOI21_X1 U3683 ( .B1(n5217), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n3019), 
        .ZN(n3018) );
  INV_X1 U3684 ( .A(n4299), .ZN(n3019) );
  XNOR2_X1 U3685 ( .A(n4189), .B(n4188), .ZN(n4297) );
  OR2_X1 U3686 ( .A1(n5126), .A2(n4213), .ZN(n4214) );
  INV_X1 U3687 ( .A(n6290), .ZN(n6278) );
  NAND2_X1 U3688 ( .A1(n3202), .A2(n2967), .ZN(n3190) );
  OR2_X1 U3689 ( .A1(n3378), .A2(n3377), .ZN(n3941) );
  OR2_X1 U3690 ( .A1(n3352), .A2(n3351), .ZN(n3923) );
  OAI21_X1 U3691 ( .B1(n3224), .B2(n4509), .A(n4306), .ZN(n3229) );
  AND2_X1 U3692 ( .A1(n3976), .A2(n3977), .ZN(n4000) );
  OR2_X1 U3693 ( .A1(n3597), .A2(n4826), .ZN(n3598) );
  INV_X1 U3694 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6605) );
  AND2_X1 U3695 ( .A1(n4695), .A2(n4710), .ZN(n3058) );
  INV_X1 U3696 ( .A(n4353), .ZN(n3429) );
  AND2_X1 U3697 ( .A1(n4834), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3434) );
  AND2_X1 U3698 ( .A1(n5124), .A2(n3016), .ZN(n3015) );
  INV_X1 U3699 ( .A(n3972), .ZN(n3016) );
  AND2_X1 U3700 ( .A1(n5414), .A2(n6589), .ZN(n3972) );
  NAND2_X1 U3701 ( .A1(n3042), .A2(n4170), .ZN(n3041) );
  NOR2_X1 U3702 ( .A1(n3043), .A2(n5018), .ZN(n3042) );
  INV_X1 U3703 ( .A(n4952), .ZN(n3043) );
  NOR2_X1 U3704 ( .A1(n4822), .A2(n3032), .ZN(n3031) );
  INV_X1 U3705 ( .A(n5071), .ZN(n3032) );
  INV_X1 U3706 ( .A(n3962), .ZN(n3008) );
  NOR2_X1 U3707 ( .A1(n4714), .A2(n3038), .ZN(n3037) );
  INV_X1 U3708 ( .A(n4680), .ZN(n3038) );
  AND3_X1 U3709 ( .A1(n3026), .A2(n4357), .A3(n2996), .ZN(n4481) );
  INV_X1 U3710 ( .A(n4444), .ZN(n3025) );
  NAND2_X1 U3711 ( .A1(n3922), .A2(n3196), .ZN(n3929) );
  OR2_X1 U3712 ( .A1(n3251), .A2(n3250), .ZN(n3252) );
  INV_X1 U3713 ( .A(n3252), .ZN(n3891) );
  OR2_X1 U3714 ( .A1(n3339), .A2(n3338), .ZN(n3913) );
  INV_X1 U3715 ( .A(n2957), .ZN(n4252) );
  AND2_X2 U3716 ( .A1(n4409), .A2(n4408), .ZN(n3346) );
  INV_X1 U3717 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6558) );
  INV_X1 U3718 ( .A(n3234), .ZN(n3320) );
  OAI21_X1 U3719 ( .B1(n6489), .B2(n4437), .A(n6379), .ZN(n4502) );
  AND2_X1 U3720 ( .A1(n5453), .A2(n4402), .ZN(n4435) );
  AND2_X1 U3721 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  INV_X1 U3722 ( .A(n2978), .ZN(n6488) );
  OR2_X1 U3723 ( .A1(n3583), .A2(n5494), .ZN(n3597) );
  INV_X1 U3724 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U3725 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5616), .ZN(n4743) );
  INV_X1 U3726 ( .A(n4876), .ZN(n4874) );
  XNOR2_X1 U3727 ( .A(n4055), .B(n4194), .ZN(n4755) );
  OR2_X1 U3728 ( .A1(n4054), .A2(n4882), .ZN(n4055) );
  OR2_X1 U3729 ( .A1(n3882), .A2(n5108), .ZN(n4054) );
  OAI21_X1 U3730 ( .B1(n3818), .B2(n5116), .A(n3817), .ZN(n4912) );
  AND2_X1 U3731 ( .A1(n3794), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U3732 ( .A1(n3795), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3833)
         );
  INV_X1 U3733 ( .A(n3778), .ZN(n5006) );
  NOR2_X1 U3734 ( .A1(n3756), .A2(n5157), .ZN(n3776) );
  INV_X1 U3735 ( .A(n4949), .ZN(n3044) );
  INV_X1 U3736 ( .A(n3700), .ZN(n3701) );
  NAND2_X1 U3737 ( .A1(n3702), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3756)
         );
  NOR2_X1 U3738 ( .A1(n3665), .A2(n5383), .ZN(n3666) );
  NAND2_X1 U3739 ( .A1(n3666), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3700)
         );
  NOR2_X1 U3740 ( .A1(n3047), .A2(n5044), .ZN(n3046) );
  INV_X1 U3741 ( .A(n3048), .ZN(n3047) );
  NAND2_X1 U3742 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3632), .ZN(n3665)
         );
  NAND2_X1 U3743 ( .A1(n4959), .A2(n3048), .ZN(n5043) );
  NOR2_X1 U3744 ( .A1(n6605), .A2(n3598), .ZN(n3631) );
  AND2_X1 U3745 ( .A1(n3549), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3550)
         );
  NAND2_X1 U3746 ( .A1(n3550), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3583)
         );
  AND2_X1 U3747 ( .A1(n3534), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3549)
         );
  AND2_X1 U3748 ( .A1(n3548), .A2(n3547), .ZN(n4741) );
  NAND2_X1 U3749 ( .A1(n3512), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3513)
         );
  NOR2_X1 U3750 ( .A1(n6572), .A2(n3513), .ZN(n3534) );
  NOR2_X1 U3751 ( .A1(n6544), .A2(n3482), .ZN(n3512) );
  AND3_X1 U3752 ( .A1(n3487), .A2(n3486), .A3(n3485), .ZN(n4698) );
  AND2_X1 U3753 ( .A1(n3459), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3466)
         );
  AND2_X1 U3754 ( .A1(n3457), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3459)
         );
  AOI21_X1 U3755 ( .B1(n3454), .B2(n3592), .A(n3060), .ZN(n4454) );
  NOR2_X1 U3756 ( .A1(n3435), .A2(n3387), .ZN(n3450) );
  INV_X1 U3757 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U3759 ( .A1(n4184), .A2(n3012), .ZN(n4281) );
  OR2_X1 U3760 ( .A1(n4876), .A2(n4185), .ZN(n3012) );
  AND2_X1 U3761 ( .A1(n3015), .A2(n3973), .ZN(n3014) );
  NOR2_X1 U3762 ( .A1(n5414), .A2(n3021), .ZN(n3020) );
  AOI21_X1 U3763 ( .B1(n5414), .B2(n3970), .A(n3023), .ZN(n3022) );
  NOR2_X1 U3764 ( .A1(n3971), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3021)
         );
  NOR2_X1 U3765 ( .A1(n2986), .A2(n3040), .ZN(n5009) );
  INV_X1 U3766 ( .A(n3042), .ZN(n3040) );
  NOR2_X1 U3767 ( .A1(n2986), .A2(n5018), .ZN(n5019) );
  AND2_X1 U3768 ( .A1(n4148), .A2(n5046), .ZN(n5045) );
  AND2_X1 U3769 ( .A1(n4147), .A2(n4146), .ZN(n5051) );
  OR2_X1 U3770 ( .A1(n5841), .A2(n5320), .ZN(n5288) );
  AND2_X1 U3771 ( .A1(n5414), .A2(n3964), .ZN(n3966) );
  NAND2_X1 U3772 ( .A1(n5070), .A2(n5071), .ZN(n5069) );
  AND2_X1 U3773 ( .A1(n4679), .A2(n2995), .ZN(n4774) );
  INV_X1 U3774 ( .A(n4737), .ZN(n3034) );
  NAND2_X1 U3775 ( .A1(n4679), .A2(n3035), .ZN(n4736) );
  AND2_X1 U3776 ( .A1(n2988), .A2(n3958), .ZN(n3001) );
  NOR2_X1 U3777 ( .A1(n4626), .A2(n4627), .ZN(n4679) );
  NAND2_X1 U3778 ( .A1(n4679), .A2(n4680), .ZN(n4713) );
  INV_X1 U3779 ( .A(n5288), .ZN(n4787) );
  NOR2_X1 U3780 ( .A1(n4787), .A2(n4381), .ZN(n5819) );
  AND2_X1 U3781 ( .A1(n4180), .A2(n4111), .ZN(n4362) );
  AND2_X1 U3782 ( .A1(n4098), .A2(n4097), .ZN(n4361) );
  INV_X1 U3783 ( .A(n3599), .ZN(n3600) );
  AND2_X2 U3784 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4430) );
  NOR3_X1 U3785 ( .A1(n3911), .A2(n3404), .A3(n6283), .ZN(n5879) );
  AND2_X1 U3786 ( .A1(n6056), .A2(n6290), .ZN(n6058) );
  AND2_X1 U3787 ( .A1(n6354), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6196)
         );
  INV_X1 U3788 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6358) );
  INV_X1 U3789 ( .A(n6136), .ZN(n6289) );
  NOR2_X1 U3790 ( .A1(n6468), .A2(n3391), .ZN(n4437) );
  OR2_X1 U3791 ( .A1(n5343), .A2(n4206), .ZN(n4934) );
  INV_X1 U3792 ( .A(n5595), .ZN(n5625) );
  AND2_X1 U3793 ( .A1(n2956), .A2(n4756), .ZN(n5612) );
  AND2_X1 U3794 ( .A1(n4755), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4756) );
  AND2_X1 U3795 ( .A1(n2956), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U3796 ( .A1(n2956), .A2(n5597), .ZN(n4986) );
  INV_X1 U3797 ( .A(n5078), .ZN(n5066) );
  INV_X1 U3798 ( .A(n5068), .ZN(n4807) );
  NAND2_X1 U3799 ( .A1(n6653), .A2(n4610), .ZN(n5081) );
  INV_X1 U3800 ( .A(n5102), .ZN(n4717) );
  AND2_X1 U3801 ( .A1(n4313), .A2(n4312), .ZN(n5670) );
  INV_X1 U3802 ( .A(n5715), .ZN(n5735) );
  OAI21_X1 U3803 ( .B1(n4064), .B2(n4066), .A(n4065), .ZN(n5090) );
  NAND2_X1 U3804 ( .A1(n3699), .A2(n3698), .ZN(n5022) );
  AND2_X1 U3805 ( .A1(n4797), .A2(n4800), .ZN(n5507) );
  INV_X1 U3806 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U3807 ( .A1(n5782), .A2(n4039), .ZN(n5777) );
  INV_X1 U3808 ( .A(n5782), .ZN(n5771) );
  OR2_X1 U3809 ( .A1(n5426), .A2(n4273), .ZN(n5232) );
  AND2_X1 U3810 ( .A1(n3010), .A2(n2993), .ZN(n5170) );
  AND2_X1 U3811 ( .A1(n5140), .A2(n5181), .ZN(n5177) );
  NAND2_X1 U3812 ( .A1(n5070), .A2(n3029), .ZN(n4963) );
  NOR2_X1 U3813 ( .A1(n5309), .A2(n5325), .ZN(n5448) );
  NAND2_X1 U3814 ( .A1(n4810), .A2(n3962), .ZN(n5206) );
  INV_X1 U3815 ( .A(n5791), .ZN(n5325) );
  NAND2_X1 U3816 ( .A1(n3959), .A2(n3958), .ZN(n4719) );
  NAND2_X1 U3817 ( .A1(n4357), .A2(n4358), .ZN(n4372) );
  INV_X1 U3818 ( .A(n4790), .ZN(n5830) );
  OR2_X1 U3819 ( .A1(n6474), .A2(n6391), .ZN(n5845) );
  AND2_X1 U3820 ( .A1(n4284), .A2(n4239), .ZN(n5837) );
  AND2_X1 U3821 ( .A1(n4284), .A2(n6346), .ZN(n5841) );
  INV_X1 U3822 ( .A(n3292), .ZN(n3293) );
  AND2_X1 U3823 ( .A1(n3400), .A2(n3399), .ZN(n3401) );
  INV_X1 U3824 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U3825 ( .A1(n6466), .A2(n6468), .ZN(n6474) );
  INV_X1 U3826 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5454) );
  OAI21_X1 U3827 ( .B1(n5854), .B2(n5878), .A(n5853), .ZN(n5872) );
  OR3_X1 U3828 ( .A1(n3911), .A2(n3404), .A3(n6128), .ZN(n5954) );
  NAND2_X1 U3829 ( .A1(n4639), .A2(n6233), .ZN(n5963) );
  OR2_X1 U3830 ( .A1(n6026), .A2(n6025), .ZN(n6045) );
  INV_X1 U3831 ( .A(n6090), .ZN(n6044) );
  INV_X1 U3832 ( .A(n6162), .ZN(n6154) );
  OR2_X1 U3833 ( .A1(n6174), .A2(n6173), .ZN(n6192) );
  INV_X1 U3834 ( .A(n6168), .ZN(n6191) );
  INV_X1 U3835 ( .A(n6068), .ZN(n6303) );
  INV_X1 U3836 ( .A(n6084), .ZN(n6327) );
  NAND2_X1 U3837 ( .A1(n4865), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6379) );
  INV_X1 U3838 ( .A(n4297), .ZN(n4999) );
  AOI21_X1 U3839 ( .B1(n4297), .B2(n5836), .A(n3017), .ZN(n4301) );
  NAND2_X1 U3840 ( .A1(n4300), .A2(n3018), .ZN(n3017) );
  AND2_X1 U3841 ( .A1(n4294), .A2(n3059), .ZN(n4295) );
  AND2_X1 U3842 ( .A1(n4936), .A2(n3049), .ZN(n4064) );
  INV_X1 U3843 ( .A(n4306), .ZN(n4083) );
  NAND2_X1 U3844 ( .A1(n4922), .A2(n4923), .ZN(n4911) );
  AND2_X2 U3845 ( .A1(n3069), .A2(n4409), .ZN(n3326) );
  INV_X1 U3846 ( .A(n5785), .ZN(n5766) );
  AND2_X2 U3847 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4408) );
  OR2_X1 U3848 ( .A1(n5030), .A2(n5029), .ZN(n2986) );
  INV_X1 U3849 ( .A(n5414), .ZN(n5413) );
  OR3_X1 U3850 ( .A1(n2986), .A2(n3041), .A3(n4927), .ZN(n2987) );
  OR2_X1 U3851 ( .A1(n5414), .A2(n5815), .ZN(n2988) );
  OR2_X1 U3852 ( .A1(n4043), .A2(n3013), .ZN(n4061) );
  AOI21_X1 U3853 ( .B1(n3024), .B2(n3022), .A(n3020), .ZN(n5133) );
  NAND2_X1 U3854 ( .A1(n4959), .A2(n4960), .ZN(n5059) );
  NAND2_X1 U3855 ( .A1(n3699), .A2(n3045), .ZN(n4948) );
  AND2_X1 U3856 ( .A1(n5181), .A2(n5176), .ZN(n2989) );
  NAND2_X1 U3857 ( .A1(n4082), .A2(n4306), .ZN(n4111) );
  AND2_X1 U3858 ( .A1(n4334), .A2(n4185), .ZN(n4103) );
  AND2_X1 U3859 ( .A1(n5070), .A2(n3031), .ZN(n2990) );
  NAND2_X1 U3860 ( .A1(n4694), .A2(n3058), .ZN(n4709) );
  NAND2_X1 U3861 ( .A1(n3004), .A2(n3960), .ZN(n4724) );
  AND2_X1 U3862 ( .A1(n4694), .A2(n4695), .ZN(n4693) );
  AND2_X1 U3863 ( .A1(n5414), .A2(n5321), .ZN(n2991) );
  AND2_X2 U3864 ( .A1(n4408), .A2(n4430), .ZN(n3277) );
  OR2_X1 U3865 ( .A1(n2986), .A2(n3041), .ZN(n2992) );
  OR2_X1 U3866 ( .A1(n5414), .A2(n5141), .ZN(n2993) );
  AND2_X1 U3867 ( .A1(n3029), .A2(n3028), .ZN(n2994) );
  AND2_X1 U3868 ( .A1(n3195), .A2(n3385), .ZN(n4217) );
  AND2_X1 U3869 ( .A1(n3035), .A2(n3034), .ZN(n2995) );
  NOR2_X1 U3870 ( .A1(n4480), .A2(n3025), .ZN(n2996) );
  AND2_X1 U3871 ( .A1(n3044), .A2(n3045), .ZN(n2997) );
  NAND2_X1 U3872 ( .A1(n4284), .A2(n4283), .ZN(n5799) );
  INV_X1 U3873 ( .A(n5799), .ZN(n5836) );
  AND2_X1 U3874 ( .A1(n4679), .A2(n3037), .ZN(n2998) );
  NOR3_X1 U3875 ( .A1(n4234), .A2(n3204), .A3(n2967), .ZN(n2999) );
  AND2_X1 U3876 ( .A1(n3026), .A2(n4357), .ZN(n3000) );
  NAND2_X1 U3877 ( .A1(n3004), .A2(n3002), .ZN(n3961) );
  NAND2_X1 U3878 ( .A1(n5140), .A2(n2989), .ZN(n3010) );
  INV_X1 U3879 ( .A(n2977), .ZN(n5142) );
  AND2_X4 U3880 ( .A1(n4847), .A2(n4414), .ZN(n3150) );
  AND2_X2 U3881 ( .A1(n2964), .A2(n4847), .ZN(n3148) );
  AND2_X4 U3882 ( .A1(n3075), .A2(n4847), .ZN(n3327) );
  NOR2_X4 U3883 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U3884 ( .A1(n4443), .A2(n4442), .ZN(n3921) );
  NAND2_X1 U3885 ( .A1(n3024), .A2(n3969), .ZN(n5139) );
  NAND3_X1 U3886 ( .A1(n3026), .A2(n4357), .A3(n4444), .ZN(n4479) );
  AND2_X2 U3887 ( .A1(n2961), .A2(n2997), .ZN(n4937) );
  AND2_X1 U3888 ( .A1(n4936), .A2(n5006), .ZN(n4922) );
  NAND2_X1 U3889 ( .A1(n3056), .A2(n4463), .ZN(n3445) );
  NAND2_X1 U3890 ( .A1(n3414), .A2(n3287), .ZN(n3418) );
  AOI22_X1 U3891 ( .A1(n3326), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3089) );
  AND2_X1 U3892 ( .A1(n4334), .A2(n4190), .ZN(n5595) );
  AND2_X1 U3893 ( .A1(n4073), .A2(n4072), .ZN(n4867) );
  NAND2_X1 U3894 ( .A1(n4328), .A2(n4527), .ZN(n3194) );
  NAND3_X1 U3895 ( .A1(n3205), .A2(n4329), .A3(n3204), .ZN(n4251) );
  NAND2_X1 U3896 ( .A1(n3456), .A2(n3446), .ZN(n3890) );
  OAI21_X1 U3897 ( .B1(n4890), .B2(n3885), .A(n4053), .ZN(n5084) );
  AOI21_X1 U3898 ( .B1(n4046), .B2(n4298), .A(n4045), .ZN(n4048) );
  OR2_X1 U3899 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3059)
         );
  INV_X1 U3900 ( .A(n3818), .ZN(n3799) );
  NOR2_X1 U3901 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3422) );
  INV_X1 U3902 ( .A(n3422), .ZN(n3818) );
  AND2_X1 U3903 ( .A1(n3453), .A2(n3452), .ZN(n3060) );
  NOR2_X1 U3904 ( .A1(n3066), .A2(n6634), .ZN(n3061) );
  OR2_X1 U3905 ( .A1(n3214), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3062)
         );
  NAND2_X1 U3906 ( .A1(n3287), .A2(n3949), .ZN(n3063) );
  AND4_X1 U3907 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3064)
         );
  INV_X1 U3908 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3908) );
  INV_X1 U3909 ( .A(n3716), .ZN(n5023) );
  NAND2_X1 U3910 ( .A1(n3385), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3582) );
  OAI21_X1 U3911 ( .B1(n3210), .B2(n3142), .A(n4032), .ZN(n3193) );
  INV_X1 U3912 ( .A(n3406), .ZN(n3316) );
  AND2_X1 U3913 ( .A1(n5847), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4016)
         );
  AOI22_X1 U3914 ( .A1(n3149), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3115) );
  OR2_X1 U3915 ( .A1(n5414), .A2(n5321), .ZN(n3963) );
  INV_X1 U3916 ( .A(n3204), .ZN(n3142) );
  AND2_X1 U3917 ( .A1(n6347), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3983)
         );
  OR2_X1 U3918 ( .A1(n4017), .A2(n4016), .ZN(n4019) );
  NAND2_X1 U3919 ( .A1(n3366), .A2(n3365), .ZN(n3455) );
  INV_X1 U3920 ( .A(n3793), .ZN(n3794) );
  INV_X1 U3921 ( .A(n5060), .ZN(n3648) );
  INV_X1 U3922 ( .A(n4798), .ZN(n3566) );
  INV_X1 U3923 ( .A(n4472), .ZN(n3441) );
  INV_X1 U3924 ( .A(n3286), .ZN(n3949) );
  OR2_X1 U3925 ( .A1(n3364), .A2(n3363), .ZN(n3926) );
  AND2_X1 U3926 ( .A1(n5079), .A2(n3159), .ZN(n3161) );
  OR3_X1 U3927 ( .A1(n4017), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n5847), 
        .ZN(n4012) );
  AND2_X1 U3928 ( .A1(n4019), .A2(n4018), .ZN(n4026) );
  INV_X1 U3929 ( .A(n3880), .ZN(n3856) );
  AND2_X1 U3930 ( .A1(n3834), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3835)
         );
  INV_X1 U3931 ( .A(n3419), .ZN(n3854) );
  INV_X1 U3932 ( .A(n4623), .ZN(n3470) );
  OR2_X1 U3933 ( .A1(n5414), .A2(n3964), .ZN(n3965) );
  INV_X1 U3934 ( .A(n4026), .ZN(n4076) );
  NOR2_X1 U3935 ( .A1(n5597), .A2(n4202), .ZN(n4974) );
  NAND2_X1 U3936 ( .A1(n3835), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3882)
         );
  AND2_X1 U3937 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3701), .ZN(n3702)
         );
  INV_X1 U3938 ( .A(n3757), .ZN(n4049) );
  AOI21_X1 U3939 ( .B1(n3939), .B2(n3592), .A(n3469), .ZN(n4623) );
  INV_X1 U3940 ( .A(n3582), .ZN(n3592) );
  INV_X1 U3941 ( .A(n5227), .ZN(n3973) );
  INV_X1 U3942 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6354) );
  AND4_X1 U3943 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3182)
         );
  OR2_X1 U3944 ( .A1(n6474), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4035) );
  INV_X1 U3945 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5383) );
  INV_X1 U3946 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4826) );
  INV_X1 U3947 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6544) );
  INV_X1 U3948 ( .A(n5613), .ZN(n5603) );
  INV_X1 U3949 ( .A(n4743), .ZN(n4751) );
  INV_X1 U3950 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U3951 ( .A1(n4233), .A2(n4232), .ZN(n4284) );
  OR2_X1 U3952 ( .A1(n4865), .A2(n4413), .ZN(n4399) );
  AND2_X1 U3953 ( .A1(n5985), .A2(n4538), .ZN(n4639) );
  INV_X1 U3954 ( .A(n6024), .ZN(n5918) );
  NAND2_X1 U3955 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  NAND2_X1 U3956 ( .A1(n4840), .A2(n4502), .ZN(n4561) );
  INV_X1 U3957 ( .A(n4070), .ZN(n4237) );
  NAND2_X1 U3958 ( .A1(n4317), .A2(n4303), .ZN(n6484) );
  NOR2_X1 U3959 ( .A1(n6437), .A2(n5370), .ZN(n5356) );
  NOR2_X1 U3960 ( .A1(n6432), .A2(n4961), .ZN(n5380) );
  NOR2_X1 U3961 ( .A1(n4755), .A2(n6468), .ZN(n4081) );
  NAND2_X1 U3962 ( .A1(n3466), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3482)
         );
  INV_X1 U3963 ( .A(n5561), .ZN(n5581) );
  INV_X1 U3964 ( .A(n5076), .ZN(n5065) );
  AND2_X1 U3965 ( .A1(n5081), .A2(n4831), .ZN(n4832) );
  INV_X1 U3966 ( .A(n5081), .ZN(n5636) );
  INV_X1 U3967 ( .A(n5737), .ZN(n6649) );
  INV_X1 U3968 ( .A(n5777), .ZN(n5754) );
  AND2_X1 U3969 ( .A1(n4609), .A2(n2999), .ZN(n5785) );
  OR2_X1 U3970 ( .A1(n5264), .A2(n4272), .ZN(n5426) );
  AND2_X1 U3971 ( .A1(n5440), .A2(n5153), .ZN(n5271) );
  NOR2_X1 U3972 ( .A1(n5310), .A2(n4289), .ZN(n5440) );
  AND2_X1 U3973 ( .A1(n4867), .A2(n4306), .ZN(n6346) );
  INV_X1 U3974 ( .A(n5911), .ZN(n5871) );
  OAI21_X1 U3975 ( .B1(n5919), .B2(n5934), .A(n6103), .ZN(n5936) );
  INV_X1 U3976 ( .A(n4500), .ZN(n5943) );
  AND2_X1 U3977 ( .A1(n4639), .A2(n6163), .ZN(n5950) );
  OAI21_X1 U3978 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6466), .A(n5918), 
        .ZN(n6136) );
  INV_X1 U3979 ( .A(n5963), .ZN(n5980) );
  INV_X1 U3980 ( .A(n6048), .ZN(n6039) );
  NOR2_X1 U3981 ( .A1(n4460), .A2(n4463), .ZN(n5985) );
  OAI21_X1 U3982 ( .B1(n6107), .B2(n6133), .A(n6106), .ZN(n6123) );
  OR2_X1 U3983 ( .A1(n6132), .A2(n6283), .ZN(n6049) );
  NAND2_X1 U3984 ( .A1(n3911), .A2(n4460), .ZN(n6132) );
  AND2_X1 U3985 ( .A1(n6204), .A2(n6233), .ZN(n6270) );
  INV_X1 U3986 ( .A(n5875), .ZN(n6336) );
  AND2_X1 U3987 ( .A1(n4030), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4839) );
  INV_X1 U3988 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6468) );
  INV_X1 U3989 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U3990 ( .A1(n4609), .A2(n4237), .ZN(n4317) );
  INV_X1 U3991 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6167) );
  AND2_X1 U3992 ( .A1(n4210), .A2(n4209), .ZN(n4211) );
  NAND2_X1 U3993 ( .A1(n2956), .A2(n4081), .ZN(n5564) );
  NAND2_X1 U3994 ( .A1(n5076), .A2(n3158), .ZN(n5068) );
  INV_X1 U3995 ( .A(n4807), .ZN(n5075) );
  INV_X1 U3996 ( .A(n4784), .ZN(n5518) );
  INV_X1 U3997 ( .A(n5670), .ZN(n5667) );
  INV_X1 U3998 ( .A(n5735), .ZN(n6653) );
  OR3_X1 U3999 ( .A1(n4317), .A2(n2979), .A3(READY_N), .ZN(n5715) );
  NAND2_X1 U4000 ( .A1(n4609), .A2(n4310), .ZN(n5737) );
  OR2_X1 U4001 ( .A1(n5785), .A2(n4036), .ZN(n5782) );
  INV_X1 U4002 ( .A(n5837), .ZN(n5825) );
  INV_X1 U4003 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6347) );
  OR2_X1 U4004 ( .A1(n6225), .A2(n6128), .ZN(n5875) );
  NAND2_X1 U4005 ( .A1(n5879), .A2(n6233), .ZN(n5939) );
  INV_X1 U4006 ( .A(n5944), .ZN(n4537) );
  NAND2_X1 U4007 ( .A1(n5985), .A2(n6226), .ZN(n6011) );
  NAND2_X1 U4008 ( .A1(n5985), .A2(n5984), .ZN(n6048) );
  OR2_X1 U4009 ( .A1(n6049), .A2(n6233), .ZN(n6090) );
  OR2_X1 U4010 ( .A1(n6049), .A2(n6163), .ZN(n6127) );
  OR2_X1 U4011 ( .A1(n6132), .A2(n6128), .ZN(n6168) );
  OR2_X1 U4012 ( .A1(n6132), .A2(n6096), .ZN(n6162) );
  NAND2_X1 U4013 ( .A1(n6204), .A2(n6163), .ZN(n6224) );
  NAND2_X1 U4014 ( .A1(n6284), .A2(n6226), .ZN(n6341) );
  INV_X1 U4015 ( .A(n6380), .ZN(n6489) );
  INV_X1 U4016 ( .A(n6462), .ZN(n6458) );
  INV_X1 U4017 ( .A(n6445), .ZN(n6453) );
  OAI21_X1 U4018 ( .B1(n5112), .B2(n5825), .A(n4295), .ZN(U2989) );
  AOI22_X1 U4019 ( .A1(n3325), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3074) );
  INV_X1 U4020 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3068) );
  AND2_X2 U4021 ( .A1(n3068), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3075)
         );
  NOR2_X4 U4022 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4023 ( .A1(n3327), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3073) );
  AND2_X2 U4024 ( .A1(n3069), .A2(n4414), .ZN(n3276) );
  AND2_X4 U4025 ( .A1(n4851), .A2(n4430), .ZN(n3297) );
  AOI22_X1 U4026 ( .A1(n3276), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3072) );
  AND2_X2 U4027 ( .A1(n4407), .A2(n3070), .ZN(n3271) );
  AOI22_X1 U4028 ( .A1(n3277), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3071) );
  AND2_X4 U4029 ( .A1(n3075), .A2(n4851), .ZN(n3295) );
  AOI22_X1 U4030 ( .A1(n3295), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3079) );
  AND2_X4 U4031 ( .A1(n2964), .A2(n4851), .ZN(n3245) );
  AOI22_X1 U4032 ( .A1(n3245), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3078) );
  AND2_X4 U4033 ( .A1(n4851), .A2(n4414), .ZN(n3173) );
  AOI22_X1 U4034 ( .A1(n3173), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U4035 ( .A1(n3346), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3076) );
  NAND2_X2 U4036 ( .A1(n3081), .A2(n3080), .ZN(n3206) );
  AOI22_X1 U4037 ( .A1(n3276), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3085) );
  AOI22_X1 U4038 ( .A1(n3148), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3084) );
  AOI22_X1 U4039 ( .A1(n3149), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U4040 ( .A1(n3245), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3082) );
  AND4_X2 U4041 ( .A1(n3085), .A2(n3084), .A3(n3083), .A4(n3082), .ZN(n3091)
         );
  AOI22_X1 U4042 ( .A1(n3325), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3088) );
  AOI22_X1 U4043 ( .A1(n3297), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U4044 ( .A1(n3173), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3086) );
  NAND2_X2 U4045 ( .A1(n3090), .A2(n3091), .ZN(n3186) );
  INV_X2 U4046 ( .A(n3186), .ZN(n3204) );
  NAND2_X1 U4047 ( .A1(n3346), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3095)
         );
  NAND2_X1 U4048 ( .A1(n2983), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U4049 ( .A1(n3173), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U4050 ( .A1(n3151), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U4051 ( .A1(n3326), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3099)
         );
  NAND2_X1 U4052 ( .A1(n3295), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U4053 ( .A1(n3245), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U4054 ( .A1(n3148), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4055 ( .A1(n3327), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U4056 ( .A1(n3150), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4057 ( .A1(n3143), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U4058 ( .A1(n3277), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3100)
         );
  NAND2_X1 U4059 ( .A1(n3325), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3108)
         );
  NAND2_X1 U4060 ( .A1(n3276), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4061 ( .A1(n3297), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3106)
         );
  NAND2_X1 U4063 ( .A1(n3271), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3105) );
  INV_X1 U4064 ( .A(n3194), .ZN(n3122) );
  AOI22_X1 U4065 ( .A1(n3295), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4066 ( .A1(n3245), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4067 ( .A1(n3346), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4068 ( .A1(n3325), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4069 ( .A1(n3276), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4070 ( .A1(n3277), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4071 ( .A1(n3327), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U4072 ( .A1(n3122), .A2(n3201), .ZN(n4071) );
  AOI22_X1 U4073 ( .A1(n3149), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3245), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4074 ( .A1(n3148), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4075 ( .A1(n3297), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4076 ( .A1(n3295), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4077 ( .A1(n3325), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4078 ( .A1(n3276), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4079 ( .A1(n3143), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4080 ( .A1(n3346), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4081 ( .A1(n3326), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4082 ( .A1(n3148), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4083 ( .A1(n3245), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4084 ( .A1(n2982), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4085 ( .A1(n3325), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4086 ( .A1(n3277), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4087 ( .A1(n3295), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4088 ( .A1(n3173), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3136) );
  AOI21_X1 U4089 ( .B1(n4071), .B2(n4562), .A(n4306), .ZN(n3164) );
  AOI22_X1 U4090 ( .A1(n3325), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4091 ( .A1(n3276), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4092 ( .A1(n3277), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4093 ( .A1(n3327), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3144) );
  NAND4_X1 U4094 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3157)
         );
  AOI22_X1 U4095 ( .A1(n3295), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4096 ( .A1(n3149), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4097 ( .A1(n3245), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4098 ( .A1(n3346), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3152) );
  NAND4_X1 U4099 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3156)
         );
  OR2_X2 U4100 ( .A1(n3157), .A2(n3156), .ZN(n4082) );
  NAND2_X1 U4101 ( .A1(n3599), .A2(n4082), .ZN(n3163) );
  NAND2_X1 U4102 ( .A1(n3158), .A2(n3204), .ZN(n5079) );
  NAND2_X1 U4103 ( .A1(n3158), .A2(n4562), .ZN(n3159) );
  NAND2_X1 U4104 ( .A1(n2975), .A2(n3189), .ZN(n3160) );
  NAND2_X1 U4105 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  AND2_X2 U4106 ( .A1(n3163), .A2(n3162), .ZN(n4073) );
  NAND2_X1 U4107 ( .A1(n3164), .A2(n4073), .ZN(n3221) );
  NAND2_X1 U4108 ( .A1(n3276), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U4109 ( .A1(n3327), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4110 ( .A1(n3297), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3166)
         );
  NAND2_X1 U4111 ( .A1(n3143), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4112 ( .A1(n3148), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4113 ( .A1(n3295), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4114 ( .A1(n3346), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3170)
         );
  NAND2_X1 U4115 ( .A1(n3151), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U4116 ( .A1(n2982), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U4117 ( .A1(n3245), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4118 ( .A1(n3173), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U4119 ( .A1(n3150), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U4120 ( .A1(n3325), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3181)
         );
  NAND2_X1 U4121 ( .A1(n3326), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3180)
         );
  NAND2_X1 U4122 ( .A1(n3277), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3179)
         );
  NAND2_X1 U4123 ( .A1(n3271), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4124 ( .A1(n3221), .A2(n4748), .ZN(n3199) );
  NAND2_X1 U4125 ( .A1(n4217), .A2(n4527), .ZN(n3188) );
  AND2_X1 U4126 ( .A1(n4328), .A2(n3158), .ZN(n3187) );
  NAND2_X1 U4127 ( .A1(n3188), .A2(n3187), .ZN(n4031) );
  INV_X1 U4128 ( .A(n4031), .ZN(n3191) );
  NAND2_X1 U4129 ( .A1(n3191), .A2(n3190), .ZN(n3224) );
  NAND2_X1 U4130 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6411) );
  OAI21_X1 U4131 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6411), .ZN(n3192) );
  INV_X1 U4132 ( .A(n3192), .ZN(n4191) );
  NOR2_X1 U4133 ( .A1(n4306), .A2(n4191), .ZN(n3210) );
  AND2_X2 U4134 ( .A1(n4240), .A2(n4082), .ZN(n4032) );
  NOR2_X1 U4135 ( .A1(n3224), .A2(n3193), .ZN(n3198) );
  NAND2_X1 U4136 ( .A1(n3217), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3234) );
  XNOR2_X1 U4137 ( .A(n6354), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6227)
         );
  AOI21_X1 U4138 ( .B1(n3321), .B2(n6227), .A(n3200), .ZN(n3213) );
  AND2_X1 U4139 ( .A1(n4328), .A2(n4527), .ZN(n4218) );
  NAND2_X1 U4140 ( .A1(n3158), .A2(n3207), .ZN(n4228) );
  NAND2_X1 U4141 ( .A1(n2979), .A2(n4748), .ZN(n3976) );
  NAND2_X1 U4142 ( .A1(n3205), .A2(n4252), .ZN(n3208) );
  NOR2_X1 U4143 ( .A1(n3208), .A2(n3194), .ZN(n3209) );
  NAND2_X1 U4144 ( .A1(n3211), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3212) );
  OAI211_X2 U4145 ( .C1(n3234), .C2(n4856), .A(n3213), .B(n3212), .ZN(n3232)
         );
  INV_X1 U4146 ( .A(n3212), .ZN(n3215) );
  INV_X1 U4147 ( .A(n3213), .ZN(n3214) );
  NAND2_X1 U4148 ( .A1(n3215), .A2(n3062), .ZN(n3216) );
  NAND2_X1 U4149 ( .A1(n3217), .A2(n3061), .ZN(n3220) );
  MUX2_X1 U4150 ( .A(n4327), .B(n3321), .S(n6347), .Z(n3218) );
  INV_X1 U4151 ( .A(n3218), .ZN(n3219) );
  NAND2_X1 U4152 ( .A1(n3220), .A2(n3219), .ZN(n3255) );
  AND2_X1 U4153 ( .A1(n3221), .A2(n4748), .ZN(n3223) );
  NAND2_X1 U4154 ( .A1(n3223), .A2(n3222), .ZN(n4248) );
  INV_X1 U4155 ( .A(n4082), .ZN(n4509) );
  OR2_X1 U4156 ( .A1(n6474), .A2(n6634), .ZN(n6386) );
  INV_X1 U4157 ( .A(n6386), .ZN(n3228) );
  INV_X1 U4158 ( .A(n4329), .ZN(n4250) );
  OAI21_X1 U4159 ( .B1(n4250), .B2(n4252), .A(n4748), .ZN(n3226) );
  NAND2_X1 U4160 ( .A1(n4032), .A2(n3202), .ZN(n3225) );
  NAND2_X1 U4161 ( .A1(n4240), .A2(n4306), .ZN(n4394) );
  NAND3_X1 U4162 ( .A1(n3226), .A2(n3225), .A3(n4394), .ZN(n3227) );
  NAND2_X1 U4163 ( .A1(n3231), .A2(n4248), .ZN(n3256) );
  NAND2_X1 U4164 ( .A1(n3233), .A2(n3232), .ZN(n3239) );
  NOR2_X1 U4165 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6354), .ZN(n6097)
         );
  NAND2_X1 U4166 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6097), .ZN(n6129) );
  OAI21_X1 U4167 ( .B1(n6558), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6129), 
        .ZN(n3235) );
  NAND2_X1 U4168 ( .A1(n3321), .A2(n4543), .ZN(n3236) );
  OAI21_X1 U4169 ( .B1(n4030), .B2(n6558), .A(n3236), .ZN(n3237) );
  NAND2_X1 U4170 ( .A1(n3239), .A2(n3238), .ZN(n3240) );
  OR2_X2 U4171 ( .A1(n3239), .A2(n3238), .ZN(n3319) );
  NAND2_X1 U4172 ( .A1(n3240), .A2(n3319), .ZN(n4421) );
  AOI22_X1 U4173 ( .A1(n3278), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4174 ( .A1(n3868), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4175 ( .A1(n3277), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3242) );
  BUF_X1 U4176 ( .A(n3327), .Z(n3296) );
  AOI22_X1 U4177 ( .A1(n3296), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3241) );
  NAND4_X1 U4178 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(n3251)
         );
  AOI22_X1 U4179 ( .A1(n3332), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4180 ( .A1(n3302), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3248) );
  INV_X1 U4181 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6633) );
  AOI22_X1 U4182 ( .A1(n3333), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4183 ( .A1(n2958), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4184 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  NAND2_X1 U4185 ( .A1(n4748), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3324) );
  INV_X1 U4186 ( .A(n3324), .ZN(n3311) );
  AOI22_X1 U4187 ( .A1(n3311), .A2(n3252), .B1(n3379), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3253) );
  XNOR2_X2 U4188 ( .A(n3254), .B(n3253), .ZN(n3396) );
  INV_X1 U4189 ( .A(n3255), .ZN(n3258) );
  INV_X1 U4190 ( .A(n3256), .ZN(n3257) );
  NAND2_X1 U4191 ( .A1(n3258), .A2(n3257), .ZN(n3259) );
  NAND2_X1 U4192 ( .A1(n6052), .A2(n6634), .ZN(n3413) );
  AOI22_X1 U4193 ( .A1(n3278), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4194 ( .A1(n3276), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3263) );
  BUF_X1 U4195 ( .A(n3271), .Z(n3260) );
  AOI22_X1 U4196 ( .A1(n3277), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4197 ( .A1(n3296), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3261) );
  NAND4_X1 U4198 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3270)
         );
  AOI22_X1 U4199 ( .A1(n3332), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4200 ( .A1(n2983), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4201 ( .A1(n3333), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4202 ( .A1(n2958), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U4203 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3269)
         );
  NOR2_X1 U4204 ( .A1(n3984), .A2(n3952), .ZN(n3310) );
  NAND2_X1 U4205 ( .A1(n4527), .A2(n3952), .ZN(n3288) );
  AOI22_X1 U4206 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3332), .B1(n3297), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4207 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3302), .B1(n2958), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4208 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3333), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4209 ( .A1(n3326), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3272) );
  NAND4_X1 U4210 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3284)
         );
  AOI22_X1 U4211 ( .A1(n3868), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4212 ( .A1(n3859), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4213 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3867), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4214 ( .A1(n3278), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3279) );
  NAND4_X1 U4215 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3283)
         );
  INV_X1 U4216 ( .A(n3900), .ZN(n3285) );
  INV_X1 U4217 ( .A(n3416), .ZN(n3287) );
  INV_X1 U4218 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3290) );
  AOI21_X1 U4219 ( .B1(n4748), .B2(n3900), .A(n6634), .ZN(n3289) );
  OAI211_X1 U4220 ( .C1(n4013), .C2(n3290), .A(n3289), .B(n3288), .ZN(n3415)
         );
  INV_X1 U4221 ( .A(n3984), .ZN(n4604) );
  AOI22_X1 U4222 ( .A1(n3278), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3868), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4223 ( .A1(n3296), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4224 ( .A1(n3333), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4225 ( .A1(n3866), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4226 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3308)
         );
  AOI22_X1 U4227 ( .A1(n3743), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4228 ( .A1(n3302), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4229 ( .A1(n3867), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4230 ( .A1(n2958), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3303) );
  NAND4_X1 U4231 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3307)
         );
  NAND2_X1 U4232 ( .A1(n4604), .A2(n3899), .ZN(n3309) );
  OAI21_X2 U4233 ( .B1(n4495), .B2(STATE2_REG_0__SCAN_IN), .A(n3309), .ZN(
        n3407) );
  INV_X1 U4234 ( .A(n3310), .ZN(n3314) );
  NAND2_X1 U4235 ( .A1(n3379), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4236 ( .A1(n3311), .A2(n3899), .ZN(n3312) );
  NAND2_X1 U4237 ( .A1(n3399), .A2(n3397), .ZN(n3317) );
  INV_X1 U4238 ( .A(n3407), .ZN(n3315) );
  NAND2_X1 U4239 ( .A1(n3316), .A2(n3315), .ZN(n3398) );
  NAND2_X2 U4240 ( .A1(n3396), .A2(n3318), .ZN(n3433) );
  NAND2_X1 U4241 ( .A1(n3320), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3323) );
  NOR3_X1 U4242 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6558), .A3(n6354), 
        .ZN(n5993) );
  NAND2_X1 U4243 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5993), .ZN(n5986) );
  NAND3_X1 U4244 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6281) );
  NOR2_X1 U4245 ( .A1(n6347), .A2(n6281), .ZN(n6332) );
  AOI21_X1 U4246 ( .B1(n5986), .B2(n6358), .A(n6332), .ZN(n6019) );
  AOI22_X1 U4247 ( .A1(n6019), .A2(n3321), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4327), .ZN(n3322) );
  NAND2_X1 U4248 ( .A1(n4403), .A2(n6634), .ZN(n3341) );
  AOI22_X1 U4249 ( .A1(n3278), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4250 ( .A1(n3868), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4251 ( .A1(n3860), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4252 ( .A1(n3296), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3328) );
  NAND4_X1 U4253 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3339)
         );
  AOI22_X1 U4254 ( .A1(n3332), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4255 ( .A1(n3302), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4256 ( .A1(n3333), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4257 ( .A1(n2958), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3334) );
  NAND4_X1 U4258 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3338)
         );
  AOI22_X1 U4259 ( .A1(n4020), .A2(n3913), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3379), .ZN(n3340) );
  AOI22_X1 U4260 ( .A1(n3278), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3345) );
  INV_X1 U4261 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6632) );
  AOI22_X1 U4262 ( .A1(n3868), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4263 ( .A1(n3860), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4264 ( .A1(n3296), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3143), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4265 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3352)
         );
  AOI22_X1 U4266 ( .A1(n3332), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4267 ( .A1(n3302), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4268 ( .A1(n3333), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4269 ( .A1(n2958), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3347) );
  NAND4_X1 U4270 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3351)
         );
  NAND2_X1 U4271 ( .A1(n4020), .A2(n3923), .ZN(n3354) );
  NAND2_X1 U4272 ( .A1(n3379), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4273 ( .A1(n3278), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4274 ( .A1(n3846), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4275 ( .A1(n3302), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4276 ( .A1(n3743), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3355) );
  NAND4_X1 U4277 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3364)
         );
  AOI22_X1 U4278 ( .A1(n3333), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4279 ( .A1(n3332), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4280 ( .A1(n3296), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4281 ( .A1(n3868), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4282 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3363)
         );
  NAND2_X1 U4283 ( .A1(n4020), .A2(n3926), .ZN(n3366) );
  NAND2_X1 U4284 ( .A1(n3379), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3365) );
  INV_X1 U4285 ( .A(n3455), .ZN(n3367) );
  AOI22_X1 U4286 ( .A1(n3278), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4287 ( .A1(n3868), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4288 ( .A1(n3860), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4289 ( .A1(n3296), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4290 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3378)
         );
  AOI22_X1 U4291 ( .A1(n3332), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3376) );
  INV_X1 U4292 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U4293 ( .A1(n3302), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4294 ( .A1(n3333), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4295 ( .A1(n2958), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4296 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3377)
         );
  NAND2_X1 U4297 ( .A1(n4020), .A2(n3941), .ZN(n3381) );
  NAND2_X1 U4298 ( .A1(n3379), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4299 ( .A1(n3381), .A2(n3380), .ZN(n3382) );
  OR2_X1 U4300 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  NAND2_X1 U4301 ( .A1(n3383), .A2(n3382), .ZN(n3951) );
  NAND2_X1 U4302 ( .A1(n3384), .A2(n3951), .ZN(n3935) );
  INV_X1 U4303 ( .A(n3935), .ZN(n3386) );
  NAND2_X1 U4304 ( .A1(n3386), .A2(n3592), .ZN(n3395) );
  INV_X1 U4305 ( .A(n3466), .ZN(n3390) );
  INV_X1 U4306 ( .A(n3459), .ZN(n3388) );
  INV_X1 U4307 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U4308 ( .A1(n3388), .A2(n5563), .ZN(n3389) );
  NAND2_X1 U4309 ( .A1(n3390), .A2(n3389), .ZN(n5570) );
  INV_X1 U4310 ( .A(n5570), .ZN(n3393) );
  INV_X2 U4311 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4312 ( .A1(n4050), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3391), .ZN(n3392) );
  MUX2_X1 U4313 ( .A(n3393), .B(n3392), .S(n3818), .Z(n3394) );
  NAND2_X1 U4314 ( .A1(n3395), .A2(n3394), .ZN(n4488) );
  INV_X1 U4315 ( .A(n3396), .ZN(n3402) );
  NAND2_X1 U4316 ( .A1(n3398), .A2(n3405), .ZN(n3400) );
  NAND2_X1 U4317 ( .A1(n3402), .A2(n3401), .ZN(n3403) );
  NAND2_X1 U4318 ( .A1(n3391), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3757) );
  XNOR2_X1 U4319 ( .A(n3406), .B(n3405), .ZN(n3408) );
  NAND2_X1 U4320 ( .A1(n4462), .A2(n3592), .ZN(n3412) );
  AOI22_X1 U4321 ( .A1(n3419), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n3391), .ZN(n3410) );
  INV_X1 U4322 ( .A(n4228), .ZN(n4834) );
  NAND2_X1 U4323 ( .A1(n3434), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3409) );
  AND2_X1 U4324 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  NAND2_X1 U4325 ( .A1(n3413), .A2(n3415), .ZN(n3414) );
  INV_X1 U4326 ( .A(n6052), .ZN(n6345) );
  AOI22_X1 U4327 ( .A1(n3419), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n3391), .ZN(n3421) );
  NAND2_X1 U4328 ( .A1(n3434), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3420) );
  OAI211_X1 U4329 ( .C1(n6345), .C2(n3582), .A(n3421), .B(n3420), .ZN(n4363)
         );
  NAND2_X1 U4330 ( .A1(n3434), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3427) );
  INV_X1 U4331 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3424) );
  OAI21_X1 U4332 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3435), .ZN(n5770) );
  NAND2_X1 U4333 ( .A1(n3422), .A2(n5770), .ZN(n3423) );
  OAI21_X1 U4334 ( .B1(n3757), .B2(n3424), .A(n3423), .ZN(n3425) );
  AOI21_X1 U4335 ( .B1(n4050), .B2(EAX_REG_2__SCAN_IN), .A(n3425), .ZN(n3426)
         );
  AND2_X1 U4336 ( .A1(n3427), .A2(n3426), .ZN(n4354) );
  INV_X1 U4337 ( .A(n4354), .ZN(n3428) );
  NAND2_X1 U4338 ( .A1(n3429), .A2(n3428), .ZN(n3430) );
  NAND2_X1 U4339 ( .A1(n4355), .A2(n3430), .ZN(n3432) );
  NAND2_X1 U4340 ( .A1(n4353), .A2(n4354), .ZN(n3431) );
  NAND2_X1 U4341 ( .A1(n3432), .A2(n3431), .ZN(n4352) );
  INV_X1 U4342 ( .A(n4352), .ZN(n3442) );
  INV_X1 U4343 ( .A(n3434), .ZN(n3449) );
  INV_X1 U4344 ( .A(n3435), .ZN(n3437) );
  INV_X1 U4345 ( .A(n3450), .ZN(n3436) );
  OAI21_X1 U4346 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3437), .A(n3436), 
        .ZN(n4760) );
  AOI22_X1 U4347 ( .A1(n3422), .A2(n4760), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4348 ( .A1(n4050), .A2(EAX_REG_3__SCAN_IN), .ZN(n3438) );
  OAI211_X1 U4349 ( .C1(n3449), .C2(n3068), .A(n3439), .B(n3438), .ZN(n3440)
         );
  AOI21_X1 U4350 ( .B1(n2984), .B2(n3592), .A(n3440), .ZN(n4472) );
  INV_X1 U4351 ( .A(n3443), .ZN(n3444) );
  NAND2_X1 U4352 ( .A1(n3445), .A2(n3444), .ZN(n3446) );
  INV_X1 U4353 ( .A(n3890), .ZN(n3454) );
  OAI21_X1 U4354 ( .B1(n6167), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3391), 
        .ZN(n3448) );
  NAND2_X1 U4355 ( .A1(n4050), .A2(EAX_REG_4__SCAN_IN), .ZN(n3447) );
  OAI211_X1 U4356 ( .C1(n3449), .C2(n5454), .A(n3448), .B(n3447), .ZN(n3453)
         );
  NOR2_X1 U4357 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3450), .ZN(n3451)
         );
  NOR2_X1 U4358 ( .A1(n3457), .A2(n3451), .ZN(n5587) );
  NAND2_X1 U4359 ( .A1(n5587), .A2(n3422), .ZN(n3452) );
  NAND2_X1 U4360 ( .A1(n3922), .A2(n3592), .ZN(n3462) );
  NOR2_X1 U4361 ( .A1(n3457), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3458)
         );
  NOR2_X1 U4362 ( .A1(n3459), .A2(n3458), .ZN(n5755) );
  INV_X1 U4363 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5760) );
  OAI22_X1 U4364 ( .A1(n5755), .A2(n3818), .B1(n3757), .B2(n5760), .ZN(n3460)
         );
  AOI21_X1 U4365 ( .B1(n4050), .B2(EAX_REG_5__SCAN_IN), .A(n3460), .ZN(n3461)
         );
  NAND2_X1 U4366 ( .A1(n3462), .A2(n3461), .ZN(n4484) );
  NAND2_X1 U4367 ( .A1(n4488), .A2(n4483), .ZN(n4487) );
  INV_X1 U4368 ( .A(n4487), .ZN(n3471) );
  INV_X1 U4369 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U4370 ( .A1(n4020), .A2(n3952), .ZN(n3463) );
  OAI21_X1 U4371 ( .B1(n3464), .B2(n4013), .A(n3463), .ZN(n3465) );
  XNOR2_X1 U4372 ( .A(n3951), .B(n3465), .ZN(n3939) );
  INV_X1 U4373 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3468) );
  OAI21_X1 U4374 ( .B1(n3466), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3482), 
        .ZN(n5747) );
  AOI22_X1 U4375 ( .A1(n5747), .A2(n3799), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3467) );
  OAI21_X1 U4376 ( .B1(n3854), .B2(n3468), .A(n3467), .ZN(n3469) );
  AOI22_X1 U4377 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3296), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4378 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3867), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4379 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n2958), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4380 ( .A1(n3743), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4381 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3481)
         );
  AOI22_X1 U4382 ( .A1(n3868), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4383 ( .A1(n3302), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4384 ( .A1(n3278), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4385 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3846), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4386 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3480)
         );
  OAI21_X1 U4387 ( .B1(n3481), .B2(n3480), .A(n3592), .ZN(n3487) );
  INV_X1 U4388 ( .A(n3482), .ZN(n3484) );
  INV_X1 U4389 ( .A(n3512), .ZN(n3483) );
  OAI21_X1 U4390 ( .B1(PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n3484), .A(n3483), 
        .ZN(n5544) );
  AOI22_X1 U4391 ( .A1(n3799), .A2(n5544), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3486) );
  NAND2_X1 U4392 ( .A1(n4050), .A2(EAX_REG_8__SCAN_IN), .ZN(n3485) );
  INV_X1 U4393 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5534) );
  XNOR2_X1 U4394 ( .A(n5534), .B(n3512), .ZN(n5532) );
  AOI22_X1 U4395 ( .A1(n3278), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4396 ( .A1(n3333), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4397 ( .A1(n3743), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4398 ( .A1(n3846), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4399 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3497)
         );
  AOI22_X1 U4400 ( .A1(n3868), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4401 ( .A1(n3302), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4402 ( .A1(n3867), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4403 ( .A1(n3866), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4404 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3496)
         );
  OR2_X1 U4405 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  AOI22_X1 U4406 ( .A1(n3592), .A2(n3498), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U4407 ( .A1(n4050), .A2(EAX_REG_9__SCAN_IN), .ZN(n3499) );
  OAI211_X1 U4408 ( .C1(n5532), .C2(n3818), .A(n3500), .B(n3499), .ZN(n4695)
         );
  AOI22_X1 U4409 ( .A1(n3302), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4410 ( .A1(n3332), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4411 ( .A1(n3278), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4412 ( .A1(n3743), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4413 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3511)
         );
  AOI22_X1 U4414 ( .A1(n3868), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4415 ( .A1(n3867), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4416 ( .A1(n2958), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4417 ( .A1(n3296), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3506) );
  NAND4_X1 U4418 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3510)
         );
  NOR2_X1 U4419 ( .A1(n3511), .A2(n3510), .ZN(n3517) );
  AOI21_X1 U4420 ( .B1(n6572), .B2(n3513), .A(n3534), .ZN(n4992) );
  OAI22_X1 U4421 ( .A1(n4992), .A2(n3818), .B1(n3757), .B2(n6572), .ZN(n3514)
         );
  INV_X1 U4422 ( .A(n3514), .ZN(n3516) );
  NAND2_X1 U4423 ( .A1(n4050), .A2(EAX_REG_10__SCAN_IN), .ZN(n3515) );
  OAI211_X1 U4424 ( .C1(n3582), .C2(n3517), .A(n3516), .B(n3515), .ZN(n4710)
         );
  INV_X1 U4425 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5527) );
  XNOR2_X1 U4426 ( .A(n5527), .B(n3534), .ZN(n5743) );
  INV_X1 U4427 ( .A(n5743), .ZN(n3532) );
  AOI22_X1 U4428 ( .A1(n3332), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4429 ( .A1(n3868), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4430 ( .A1(n3296), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4431 ( .A1(n3743), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3518) );
  NAND4_X1 U4432 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3518), .ZN(n3527)
         );
  AOI22_X1 U4433 ( .A1(n3278), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4434 ( .A1(n3302), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4435 ( .A1(n3372), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4436 ( .A1(n2958), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4437 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3526)
         );
  OAI21_X1 U4438 ( .B1(n3527), .B2(n3526), .A(n3592), .ZN(n3530) );
  NAND2_X1 U4439 ( .A1(n4050), .A2(EAX_REG_11__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4440 ( .A1(n4049), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3528)
         );
  NAND3_X1 U4441 ( .A1(n3530), .A2(n3529), .A3(n3528), .ZN(n3531) );
  AOI21_X1 U4442 ( .B1(n3532), .B2(n3799), .A(n3531), .ZN(n4735) );
  INV_X1 U4443 ( .A(n3549), .ZN(n3535) );
  XNOR2_X1 U4444 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3535), .ZN(n5520)
         );
  INV_X1 U4445 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4782) );
  OAI22_X1 U4446 ( .A1(n5520), .A2(n3818), .B1(n3757), .B2(n4782), .ZN(n3536)
         );
  AOI21_X1 U4447 ( .B1(n4050), .B2(EAX_REG_12__SCAN_IN), .A(n3536), .ZN(n3548)
         );
  AOI22_X1 U4448 ( .A1(n3278), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4449 ( .A1(n3846), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4450 ( .A1(n3868), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4451 ( .A1(n3296), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3537) );
  NAND4_X1 U4452 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(n3546)
         );
  AOI22_X1 U4453 ( .A1(n3302), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4454 ( .A1(n3332), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4455 ( .A1(n3333), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4456 ( .A1(n3743), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4457 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3545)
         );
  OAI21_X1 U4458 ( .B1(n3546), .B2(n3545), .A(n3592), .ZN(n3547) );
  NAND2_X1 U4459 ( .A1(n4050), .A2(EAX_REG_13__SCAN_IN), .ZN(n3552) );
  OAI21_X1 U4460 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3550), .A(n3583), 
        .ZN(n5513) );
  AOI22_X1 U4461 ( .A1(n3799), .A2(n5513), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4462 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  NAND2_X1 U4463 ( .A1(n3554), .A2(n3553), .ZN(n3568) );
  OAI21_X1 U4464 ( .B1(n3554), .B2(n3553), .A(n3568), .ZN(n4799) );
  INV_X1 U4465 ( .A(n4799), .ZN(n3567) );
  AOI22_X1 U4466 ( .A1(n3278), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4467 ( .A1(n3332), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4468 ( .A1(n2958), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4469 ( .A1(n3860), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4470 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3564)
         );
  AOI22_X1 U4471 ( .A1(n3302), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4472 ( .A1(n3296), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4473 ( .A1(n3868), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4474 ( .A1(n3867), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4475 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3563)
         );
  OR2_X1 U4476 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  NAND2_X1 U4477 ( .A1(n3592), .A2(n3565), .ZN(n4798) );
  NAND2_X1 U4478 ( .A1(n3567), .A2(n3566), .ZN(n4797) );
  NAND2_X1 U4479 ( .A1(n4797), .A2(n3568), .ZN(n5073) );
  AOI22_X1 U4480 ( .A1(n3332), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4481 ( .A1(n3333), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4482 ( .A1(n3866), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4483 ( .A1(n2958), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3569) );
  NAND4_X1 U4484 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(n3578)
         );
  AOI22_X1 U4485 ( .A1(n3278), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3868), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4486 ( .A1(n3743), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4487 ( .A1(n3327), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4488 ( .A1(n3846), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4489 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  NOR2_X1 U4490 ( .A1(n3578), .A2(n3577), .ZN(n3581) );
  XNOR2_X1 U4491 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3583), .ZN(n5496)
         );
  INV_X1 U4492 ( .A(n5496), .ZN(n5208) );
  AOI22_X1 U4493 ( .A1(n4049), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3799), 
        .B2(n5208), .ZN(n3580) );
  NAND2_X1 U4494 ( .A1(n4050), .A2(EAX_REG_14__SCAN_IN), .ZN(n3579) );
  OAI211_X1 U4495 ( .C1(n3582), .C2(n3581), .A(n3580), .B(n3579), .ZN(n5072)
         );
  XNOR2_X1 U4496 ( .A(n3597), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5199)
         );
  AOI22_X1 U4497 ( .A1(n3419), .A2(EAX_REG_15__SCAN_IN), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4498 ( .A1(n3278), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4499 ( .A1(n3866), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4500 ( .A1(n3327), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4501 ( .A1(n3860), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3584) );
  NAND4_X1 U4502 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3594)
         );
  AOI22_X1 U4503 ( .A1(n3302), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4504 ( .A1(n2958), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4505 ( .A1(n3868), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4506 ( .A1(n3332), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4507 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3593)
         );
  OAI21_X1 U4508 ( .B1(n3594), .B2(n3593), .A(n3592), .ZN(n3595) );
  OAI211_X1 U4509 ( .C1(n5199), .C2(n3818), .A(n3596), .B(n3595), .ZN(n4820)
         );
  AOI21_X1 U4510 ( .B1(n6605), .B2(n3598), .A(n3631), .ZN(n4977) );
  OR2_X1 U4511 ( .A1(n4977), .A2(n3818), .ZN(n3615) );
  NAND2_X1 U4512 ( .A1(n3600), .A2(n2967), .ZN(n6343) );
  AOI22_X1 U4513 ( .A1(n3743), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4514 ( .A1(n3296), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4515 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3333), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4516 ( .A1(n3868), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3601) );
  NAND4_X1 U4517 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3610)
         );
  AOI22_X1 U4518 ( .A1(n3278), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4519 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n2958), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4520 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3150), .B1(n3505), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4521 ( .A1(n3866), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3605) );
  NAND4_X1 U4522 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3609)
         );
  NOR2_X1 U4523 ( .A1(n3610), .A2(n3609), .ZN(n3612) );
  AOI22_X1 U4524 ( .A1(n4050), .A2(EAX_REG_16__SCAN_IN), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3611) );
  OAI21_X1 U4525 ( .B1(n3880), .B2(n3612), .A(n3611), .ZN(n3613) );
  INV_X1 U4526 ( .A(n3613), .ZN(n3614) );
  INV_X1 U4527 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3616) );
  XNOR2_X1 U4528 ( .A(n3631), .B(n3616), .ZN(n5418) );
  AOI22_X1 U4529 ( .A1(n4050), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3391), .ZN(n3630) );
  AOI22_X1 U4530 ( .A1(n3868), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4531 ( .A1(n3866), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4532 ( .A1(n3327), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4533 ( .A1(n3333), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4534 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3628)
         );
  AOI22_X1 U4535 ( .A1(n3332), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4536 ( .A1(n3743), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4537 ( .A1(n3278), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3624) );
  AOI21_X1 U4538 ( .B1(n3260), .B2(INSTQUEUE_REG_9__1__SCAN_IN), .A(n3799), 
        .ZN(n3622) );
  NAND2_X1 U4539 ( .A1(n3372), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3621) );
  AND2_X1 U4540 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  NAND4_X1 U4541 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  NAND2_X1 U4542 ( .A1(n3880), .A2(n3818), .ZN(n3691) );
  OAI21_X1 U4543 ( .B1(n3628), .B2(n3627), .A(n3691), .ZN(n3629) );
  AOI22_X1 U4544 ( .A1(n5418), .A2(n3799), .B1(n3630), .B2(n3629), .ZN(n4960)
         );
  OR2_X1 U4545 ( .A1(n3632), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3633)
         );
  NAND2_X1 U4546 ( .A1(n3633), .A2(n3665), .ZN(n5483) );
  AOI22_X1 U4547 ( .A1(n3278), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4548 ( .A1(n3332), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4549 ( .A1(n3333), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4550 ( .A1(n3302), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4551 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4552 ( .A1(n3743), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4553 ( .A1(n2958), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4554 ( .A1(n3372), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4555 ( .A1(n3868), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4556 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  NOR2_X1 U4557 ( .A1(n3643), .A2(n3642), .ZN(n3646) );
  OAI21_X1 U4558 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6167), .A(n3391), 
        .ZN(n3645) );
  NAND2_X1 U4559 ( .A1(n3419), .A2(EAX_REG_18__SCAN_IN), .ZN(n3644) );
  OAI211_X1 U4560 ( .C1(n3880), .C2(n3646), .A(n3645), .B(n3644), .ZN(n3647)
         );
  OAI21_X1 U4561 ( .B1(n5483), .B2(n3818), .A(n3647), .ZN(n5060) );
  AOI22_X1 U4562 ( .A1(n3743), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3868), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4563 ( .A1(n3332), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4564 ( .A1(n3333), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4565 ( .A1(n3325), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4566 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3660)
         );
  AOI22_X1 U4567 ( .A1(n3327), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4568 ( .A1(n3846), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4569 ( .A1(n3302), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3656) );
  AOI21_X1 U4570 ( .B1(n3260), .B2(INSTQUEUE_REG_9__3__SCAN_IN), .A(n3799), 
        .ZN(n3654) );
  NAND2_X1 U4571 ( .A1(n3150), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3653) );
  AND2_X1 U4572 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  NAND4_X1 U4573 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3659)
         );
  OAI21_X1 U4574 ( .B1(n3660), .B2(n3659), .A(n3691), .ZN(n3662) );
  AOI22_X1 U4575 ( .A1(n4050), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3391), .ZN(n3661) );
  NAND2_X1 U4576 ( .A1(n3662), .A2(n3661), .ZN(n3664) );
  XNOR2_X1 U4577 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3665), .ZN(n5381)
         );
  NAND2_X1 U4578 ( .A1(n5381), .A2(n3799), .ZN(n3663) );
  NAND2_X1 U4579 ( .A1(n3664), .A2(n3663), .ZN(n5044) );
  OR2_X1 U4580 ( .A1(n3666), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3667)
         );
  NAND2_X1 U4581 ( .A1(n3667), .A2(n3700), .ZN(n5371) );
  AOI22_X1 U4582 ( .A1(n3743), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3868), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4583 ( .A1(n2958), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4584 ( .A1(n3325), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4585 ( .A1(n3332), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4586 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3677)
         );
  AOI22_X1 U4587 ( .A1(n3302), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4588 ( .A1(n3333), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4589 ( .A1(n3866), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4590 ( .A1(n3296), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3672) );
  NAND4_X1 U4591 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3676)
         );
  NOR2_X1 U4592 ( .A1(n3677), .A2(n3676), .ZN(n3679) );
  AOI22_X1 U4593 ( .A1(n4050), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3391), .ZN(n3678) );
  OAI21_X1 U4594 ( .B1(n3880), .B2(n3679), .A(n3678), .ZN(n3680) );
  MUX2_X1 U4595 ( .A(n5371), .B(n3680), .S(n3818), .Z(n5035) );
  INV_X1 U4596 ( .A(n5026), .ZN(n3699) );
  AOI22_X1 U4597 ( .A1(n3743), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4598 ( .A1(n3868), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4599 ( .A1(n3333), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4600 ( .A1(n3866), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4601 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3693)
         );
  AOI22_X1 U4602 ( .A1(n3325), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4603 ( .A1(n2958), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4604 ( .A1(n3867), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3688) );
  AOI21_X1 U4605 ( .B1(n3260), .B2(INSTQUEUE_REG_9__5__SCAN_IN), .A(n3799), 
        .ZN(n3686) );
  NAND2_X1 U4606 ( .A1(n3150), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3685) );
  AND2_X1 U4607 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  NAND4_X1 U4608 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3692)
         );
  OAI21_X1 U4609 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3695) );
  AOI22_X1 U4610 ( .A1(n3419), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n3391), .ZN(n3694) );
  NAND2_X1 U4611 ( .A1(n3695), .A2(n3694), .ZN(n3697) );
  XNOR2_X1 U4612 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3700), .ZN(n5362)
         );
  NAND2_X1 U4613 ( .A1(n5362), .A2(n3799), .ZN(n3696) );
  NAND2_X1 U4614 ( .A1(n3697), .A2(n3696), .ZN(n5028) );
  OAI21_X1 U4615 ( .B1(n3702), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3756), 
        .ZN(n5350) );
  AOI22_X1 U4616 ( .A1(n3327), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4617 ( .A1(n3302), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4618 ( .A1(n3743), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4619 ( .A1(n2958), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4620 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3712)
         );
  AOI22_X1 U4621 ( .A1(n3325), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3868), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4622 ( .A1(n3867), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4623 ( .A1(n3846), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4624 ( .A1(n3860), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4625 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3711)
         );
  NOR2_X1 U4626 ( .A1(n3712), .A2(n3711), .ZN(n3714) );
  AOI22_X1 U4627 ( .A1(n4050), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n3391), .ZN(n3713) );
  OAI21_X1 U4628 ( .B1(n3880), .B2(n3714), .A(n3713), .ZN(n3715) );
  MUX2_X1 U4629 ( .A(n5350), .B(n3715), .S(n3818), .Z(n3716) );
  XNOR2_X1 U4630 ( .A(n3756), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5161)
         );
  AOI22_X1 U4631 ( .A1(n3278), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4632 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3868), .B1(n3866), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4633 ( .A1(n3860), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4634 ( .A1(n3296), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4635 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3726)
         );
  AOI22_X1 U4636 ( .A1(n3332), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4637 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3302), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4638 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3333), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4639 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n2958), .B1(n3505), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4640 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3725)
         );
  NOR2_X1 U4641 ( .A1(n3726), .A2(n3725), .ZN(n3742) );
  AOI22_X1 U4642 ( .A1(n3302), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4643 ( .A1(n3846), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4644 ( .A1(n3743), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4645 ( .A1(n3296), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3727) );
  NAND4_X1 U4646 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(n3736)
         );
  AOI22_X1 U4647 ( .A1(n3278), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4648 ( .A1(n3332), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4649 ( .A1(n3333), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4650 ( .A1(n3868), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3731) );
  NAND4_X1 U4651 ( .A1(n3734), .A2(n3733), .A3(n3732), .A4(n3731), .ZN(n3735)
         );
  NOR2_X1 U4652 ( .A1(n3736), .A2(n3735), .ZN(n3741) );
  XOR2_X1 U4653 ( .A(n3742), .B(n3741), .Z(n3739) );
  INV_X1 U4654 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3737) );
  INV_X1 U4655 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U4656 ( .A1(n3854), .A2(n3737), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5157), .ZN(n3738) );
  AOI21_X1 U4657 ( .B1(n3856), .B2(n3739), .A(n3738), .ZN(n3740) );
  MUX2_X1 U4658 ( .A(n5161), .B(n3740), .S(n3818), .Z(n4949) );
  NOR2_X1 U4659 ( .A1(n3742), .A2(n3741), .ZN(n3762) );
  AOI22_X1 U4660 ( .A1(n3278), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4661 ( .A1(n3868), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4662 ( .A1(n3860), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4663 ( .A1(n3296), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4664 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4665 ( .A1(n3332), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4666 ( .A1(n3302), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4667 ( .A1(n3333), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4668 ( .A1(n2958), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4669 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OR2_X1 U4670 ( .A1(n3753), .A2(n3752), .ZN(n3761) );
  INV_X1 U4671 ( .A(n3761), .ZN(n3754) );
  XNOR2_X1 U4672 ( .A(n3762), .B(n3754), .ZN(n3755) );
  NAND2_X1 U4673 ( .A1(n3755), .A2(n3856), .ZN(n3760) );
  INV_X1 U4674 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5145) );
  XNOR2_X1 U4675 ( .A(n3776), .B(n5145), .ZN(n5149) );
  OAI22_X1 U4676 ( .A1(n5149), .A2(n3818), .B1(n5145), .B2(n3757), .ZN(n3758)
         );
  AOI21_X1 U4677 ( .B1(n4050), .B2(EAX_REG_24__SCAN_IN), .A(n3758), .ZN(n3759)
         );
  NAND2_X1 U4678 ( .A1(n3760), .A2(n3759), .ZN(n4938) );
  NAND2_X1 U4679 ( .A1(n3762), .A2(n3761), .ZN(n3779) );
  AOI22_X1 U4680 ( .A1(n3278), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4681 ( .A1(n3302), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4682 ( .A1(n3866), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4683 ( .A1(n2958), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4684 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3772)
         );
  AOI22_X1 U4685 ( .A1(n3868), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4686 ( .A1(n3867), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4687 ( .A1(n3846), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4688 ( .A1(n3296), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4689 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  NOR2_X1 U4690 ( .A1(n3772), .A2(n3771), .ZN(n3780) );
  XOR2_X1 U4691 ( .A(n3779), .B(n3780), .Z(n3775) );
  INV_X1 U4692 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3773) );
  INV_X1 U4693 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5131) );
  OAI22_X1 U4694 ( .A1(n3854), .A2(n3773), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5131), .ZN(n3774) );
  AOI21_X1 U4695 ( .B1(n3775), .B2(n3856), .A(n3774), .ZN(n3777) );
  XNOR2_X1 U4696 ( .A(n3793), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5341)
         );
  MUX2_X1 U4697 ( .A(n3777), .B(n5341), .S(n3799), .Z(n3778) );
  NOR2_X1 U4698 ( .A1(n3780), .A2(n3779), .ZN(n3802) );
  AOI22_X1 U4699 ( .A1(n3278), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4700 ( .A1(n3868), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4701 ( .A1(n3860), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4702 ( .A1(n3327), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4703 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AOI22_X1 U4704 ( .A1(n3332), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4705 ( .A1(n3302), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4706 ( .A1(n3333), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4707 ( .A1(n2958), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4708 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  OR2_X1 U4709 ( .A1(n3790), .A2(n3789), .ZN(n3801) );
  XNOR2_X1 U4710 ( .A(n3802), .B(n3801), .ZN(n3792) );
  AOI22_X1 U4711 ( .A1(n3419), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n3391), .ZN(n3791) );
  OAI21_X1 U4712 ( .B1(n3792), .B2(n3880), .A(n3791), .ZN(n3800) );
  INV_X1 U4713 ( .A(n3795), .ZN(n3797) );
  INV_X1 U4714 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4715 ( .A1(n3797), .A2(n3796), .ZN(n3798) );
  NAND2_X1 U4716 ( .A1(n3833), .A2(n3798), .ZN(n5121) );
  MUX2_X1 U4717 ( .A(n3800), .B(n5121), .S(n3799), .Z(n4923) );
  XOR2_X1 U4718 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n3833), .Z(n5116) );
  INV_X1 U4719 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4720 ( .A1(n3802), .A2(n3801), .ZN(n3819) );
  AOI22_X1 U4721 ( .A1(n3325), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4722 ( .A1(n3333), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4723 ( .A1(n3866), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4724 ( .A1(n3860), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4725 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4726 ( .A1(n3868), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4727 ( .A1(n3846), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4728 ( .A1(n3302), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4729 ( .A1(n3332), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4730 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  NOR2_X1 U4731 ( .A1(n3812), .A2(n3811), .ZN(n3820) );
  XOR2_X1 U4732 ( .A(n3819), .B(n3820), .Z(n3813) );
  NAND2_X1 U4733 ( .A1(n3813), .A2(n3856), .ZN(n3815) );
  OAI21_X1 U4734 ( .B1(n6167), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n3391), 
        .ZN(n3814) );
  OAI211_X1 U4735 ( .C1(n3854), .C2(n3816), .A(n3815), .B(n3814), .ZN(n3817)
         );
  NOR2_X1 U4736 ( .A1(n3820), .A2(n3819), .ZN(n3841) );
  AOI22_X1 U4737 ( .A1(n3325), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4738 ( .A1(n3868), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4739 ( .A1(n3860), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4740 ( .A1(n3327), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4741 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3830)
         );
  AOI22_X1 U4742 ( .A1(n3332), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3859), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4743 ( .A1(n3302), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4744 ( .A1(n3333), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4745 ( .A1(n2958), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4746 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  OR2_X1 U4747 ( .A1(n3830), .A2(n3829), .ZN(n3840) );
  XNOR2_X1 U4748 ( .A(n3841), .B(n3840), .ZN(n3832) );
  AOI22_X1 U4749 ( .A1(n4050), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n3391), .ZN(n3831) );
  OAI21_X1 U4750 ( .B1(n3832), .B2(n3880), .A(n3831), .ZN(n3839) );
  INV_X1 U4751 ( .A(n3833), .ZN(n3834) );
  INV_X1 U4752 ( .A(n3835), .ZN(n3837) );
  INV_X1 U4753 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4754 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  NAND2_X1 U4755 ( .A1(n3882), .A2(n3838), .ZN(n4903) );
  MUX2_X1 U4756 ( .A(n3839), .B(n4903), .S(n3799), .Z(n4066) );
  NAND2_X1 U4757 ( .A1(n3841), .A2(n3840), .ZN(n3875) );
  AOI22_X1 U4758 ( .A1(n3332), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4759 ( .A1(n3333), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4760 ( .A1(n3866), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4761 ( .A1(n3743), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4762 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3852)
         );
  AOI22_X1 U4763 ( .A1(n3868), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4764 ( .A1(n3302), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4765 ( .A1(n3325), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4766 ( .A1(n3846), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4767 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  NOR2_X1 U4768 ( .A1(n3852), .A2(n3851), .ZN(n3876) );
  XOR2_X1 U4769 ( .A(n3875), .B(n3876), .Z(n3857) );
  INV_X1 U4770 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3853) );
  INV_X1 U4771 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5108) );
  OAI22_X1 U4772 ( .A1(n3854), .A2(n3853), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5108), .ZN(n3855) );
  AOI21_X1 U4773 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3858) );
  XNOR2_X1 U4774 ( .A(n3882), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5105)
         );
  MUX2_X1 U4775 ( .A(n3858), .B(n5105), .S(n3799), .Z(n4891) );
  NOR2_X2 U4776 ( .A1(n4065), .A2(n4891), .ZN(n3884) );
  AOI22_X1 U4777 ( .A1(n3743), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4778 ( .A1(n3302), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4779 ( .A1(n3859), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2958), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4780 ( .A1(n3325), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4781 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3874)
         );
  AOI22_X1 U4782 ( .A1(n3866), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4783 ( .A1(n3867), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4784 ( .A1(n3332), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4785 ( .A1(n3868), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4786 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  NOR2_X1 U4787 ( .A1(n3874), .A2(n3873), .ZN(n3878) );
  NOR2_X1 U4788 ( .A1(n3876), .A2(n3875), .ZN(n3877) );
  XOR2_X1 U4789 ( .A(n3878), .B(n3877), .Z(n3881) );
  AOI22_X1 U4790 ( .A1(n3419), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n3391), .ZN(n3879) );
  OAI21_X1 U4791 ( .B1(n3881), .B2(n3880), .A(n3879), .ZN(n3883) );
  INV_X1 U4792 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4882) );
  XNOR2_X1 U4793 ( .A(n4054), .B(n4882), .ZN(n4881) );
  MUX2_X1 U4794 ( .A(n3883), .B(n4881), .S(n3799), .Z(n3885) );
  NAND2_X1 U4795 ( .A1(n3884), .A2(n3885), .ZN(n4053) );
  NAND3_X1 U4796 ( .A1(n6634), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6392) );
  INV_X1 U4797 ( .A(n6392), .ZN(n3886) );
  NOR2_X2 U4798 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6290) );
  NAND2_X1 U4799 ( .A1(n3899), .A2(n3900), .ZN(n3898) );
  NAND2_X1 U4800 ( .A1(n3898), .A2(n3891), .ZN(n3912) );
  NAND2_X1 U4801 ( .A1(n3912), .A2(n3913), .ZN(n3925) );
  XNOR2_X1 U4802 ( .A(n3925), .B(n3923), .ZN(n3888) );
  NAND2_X1 U4803 ( .A1(n3888), .A2(n2978), .ZN(n3889) );
  INV_X1 U4804 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U4805 ( .A(n3919), .B(n6539), .ZN(n4442) );
  OAI21_X1 U4806 ( .B1(n3891), .B2(n3898), .A(n3912), .ZN(n3893) );
  NAND2_X1 U4807 ( .A1(n4748), .A2(n4082), .ZN(n3895) );
  INV_X1 U4808 ( .A(n3895), .ZN(n3892) );
  AOI21_X1 U4809 ( .B1(n3893), .B2(n2978), .A(n3892), .ZN(n3894) );
  NAND2_X1 U4810 ( .A1(n3907), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5761)
         );
  OAI21_X1 U4811 ( .B1(n6488), .B2(n3900), .A(n3895), .ZN(n3896) );
  INV_X1 U4812 ( .A(n3896), .ZN(n3897) );
  NAND2_X1 U4813 ( .A1(n5778), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3905)
         );
  XNOR2_X1 U4814 ( .A(n3905), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4377)
         );
  NAND2_X1 U4815 ( .A1(n4462), .A2(n3196), .ZN(n3904) );
  OAI21_X1 U4816 ( .B1(n3900), .B2(n3899), .A(n3898), .ZN(n3901) );
  OAI211_X1 U4817 ( .C1(n3901), .C2(n6488), .A(n4032), .B(n3142), .ZN(n3902)
         );
  INV_X1 U4818 ( .A(n3902), .ZN(n3903) );
  NAND2_X1 U4819 ( .A1(n3904), .A2(n3903), .ZN(n4376) );
  NAND2_X1 U4820 ( .A1(n4377), .A2(n4376), .ZN(n4378) );
  INV_X1 U4821 ( .A(n3905), .ZN(n5779) );
  NAND2_X1 U4822 ( .A1(n5779), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3906)
         );
  AND2_X1 U4823 ( .A1(n4378), .A2(n3906), .ZN(n5763) );
  NAND2_X1 U4824 ( .A1(n5761), .A2(n5763), .ZN(n3910) );
  NAND2_X1 U4825 ( .A1(n3909), .A2(n3908), .ZN(n5762) );
  AND2_X1 U4826 ( .A1(n3910), .A2(n5762), .ZN(n4368) );
  NAND2_X1 U4827 ( .A1(n3911), .A2(n3196), .ZN(n3915) );
  OAI211_X1 U4828 ( .C1(n3913), .C2(n3912), .A(n3925), .B(n2978), .ZN(n3914)
         );
  INV_X1 U4829 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U4830 ( .A1(n4368), .A2(n4367), .ZN(n3918) );
  NAND2_X1 U4831 ( .A1(n3916), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3917)
         );
  NAND2_X1 U4832 ( .A1(n3919), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3920)
         );
  INV_X1 U4833 ( .A(n3923), .ZN(n3924) );
  NOR2_X1 U4834 ( .A1(n3925), .A2(n3924), .ZN(n3927) );
  NAND2_X1 U4835 ( .A1(n3927), .A2(n3926), .ZN(n3940) );
  OAI211_X1 U4836 ( .C1(n3927), .C2(n3926), .A(n3940), .B(n2978), .ZN(n3928)
         );
  NAND2_X1 U4837 ( .A1(n3929), .A2(n3928), .ZN(n3930) );
  INV_X1 U4838 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4599) );
  XNOR2_X1 U4839 ( .A(n3930), .B(n4599), .ZN(n4593) );
  NAND2_X1 U4840 ( .A1(n4592), .A2(n4593), .ZN(n3932) );
  NAND2_X1 U4841 ( .A1(n3930), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3931)
         );
  XNOR2_X1 U4842 ( .A(n3940), .B(n3941), .ZN(n3933) );
  NAND2_X1 U4843 ( .A1(n3933), .A2(n2978), .ZN(n3934) );
  OAI21_X1 U4844 ( .B1(n3935), .B2(n3990), .A(n3934), .ZN(n3936) );
  INV_X1 U4845 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6511) );
  XNOR2_X1 U4846 ( .A(n3936), .B(n6511), .ZN(n4553) );
  NAND2_X1 U4847 ( .A1(n4552), .A2(n4553), .ZN(n3938) );
  NAND2_X1 U4848 ( .A1(n3936), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3937)
         );
  NAND2_X1 U4849 ( .A1(n3939), .A2(n3196), .ZN(n3945) );
  INV_X1 U4850 ( .A(n3940), .ZN(n3942) );
  NAND2_X1 U4851 ( .A1(n3942), .A2(n3941), .ZN(n3954) );
  XNOR2_X1 U4852 ( .A(n3954), .B(n3952), .ZN(n3943) );
  NAND2_X1 U4853 ( .A1(n3943), .A2(n2978), .ZN(n3944) );
  NAND2_X1 U4854 ( .A1(n3945), .A2(n3944), .ZN(n3946) );
  INV_X1 U4855 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4114) );
  XNOR2_X1 U4856 ( .A(n3946), .B(n4114), .ZN(n4688) );
  NAND2_X1 U4857 ( .A1(n4687), .A2(n4688), .ZN(n3948) );
  NAND2_X1 U4858 ( .A1(n3946), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3947)
         );
  NAND2_X1 U4859 ( .A1(n3948), .A2(n3947), .ZN(n4676) );
  NOR2_X1 U4860 ( .A1(n3949), .A2(n3990), .ZN(n3950) );
  NAND2_X1 U4861 ( .A1(n2978), .A2(n3952), .ZN(n3953) );
  OR2_X1 U4862 ( .A1(n3954), .A2(n3953), .ZN(n3955) );
  INV_X1 U4863 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3956) );
  XNOR2_X1 U4864 ( .A(n3957), .B(n3956), .ZN(n4675) );
  NAND2_X1 U4865 ( .A1(n4676), .A2(n4675), .ZN(n3959) );
  NAND2_X1 U4866 ( .A1(n3957), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3958)
         );
  INV_X1 U4867 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U4868 ( .A1(n5414), .A2(n5815), .ZN(n3960) );
  INV_X1 U4869 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5807) );
  AND2_X1 U4870 ( .A1(n5414), .A2(n5807), .ZN(n4726) );
  OR2_X1 U4871 ( .A1(n5414), .A2(n5807), .ZN(n4725) );
  INV_X1 U4872 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U4873 ( .A1(n5414), .A2(n5790), .ZN(n5739) );
  OR2_X1 U4874 ( .A1(n5414), .A2(n5790), .ZN(n5740) );
  INV_X1 U4875 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4128) );
  NOR2_X1 U4876 ( .A1(n5414), .A2(n4128), .ZN(n4778) );
  NAND2_X1 U4877 ( .A1(n5414), .A2(n4128), .ZN(n4776) );
  XNOR2_X1 U4878 ( .A(n5414), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4811)
         );
  INV_X1 U4879 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U4880 ( .A1(n5414), .A2(n5318), .ZN(n3962) );
  INV_X1 U4881 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5321) );
  INV_X1 U4882 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3964) );
  INV_X1 U4883 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U4884 ( .A1(n5414), .A2(n5412), .ZN(n3967) );
  INV_X1 U4885 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U4886 ( .A1(n5412), .A2(n5439), .ZN(n5406) );
  OAI21_X1 U4887 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5406), .A(n5413), 
        .ZN(n3968) );
  NAND2_X1 U4888 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U4889 ( .A1(n5414), .A2(n5301), .ZN(n3969) );
  INV_X1 U4890 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5138) );
  NOR2_X1 U4891 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5273) );
  INV_X1 U4892 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5255) );
  INV_X1 U4893 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5141) );
  INV_X1 U4894 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5265) );
  NAND4_X1 U4895 ( .A1(n5273), .A2(n5255), .A3(n5141), .A4(n5265), .ZN(n3971)
         );
  NAND2_X1 U4896 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U4897 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4270) );
  NOR2_X1 U4898 ( .A1(n5152), .A2(n4270), .ZN(n4290) );
  AND2_X1 U4899 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U4900 ( .A1(n4290), .A2(n5286), .ZN(n3970) );
  XNOR2_X1 U4901 ( .A(n5414), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5135)
         );
  INV_X1 U4902 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6589) );
  INV_X1 U4903 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5243) );
  NOR2_X1 U4904 ( .A1(n5413), .A2(n5243), .ZN(n5124) );
  NAND2_X1 U4905 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5227) );
  INV_X1 U4906 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6498) );
  AND2_X1 U4907 ( .A1(n5413), .A2(n5243), .ZN(n5123) );
  NOR2_X1 U4908 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5226) );
  NAND3_X1 U4909 ( .A1(n5123), .A2(n5226), .A3(n6498), .ZN(n4044) );
  OAI22_X1 U4910 ( .A1(n4215), .A2(n6498), .B1(n5126), .B2(n4044), .ZN(n3975)
         );
  XNOR2_X1 U4911 ( .A(n3975), .B(n3974), .ZN(n5211) );
  NAND2_X1 U4912 ( .A1(n2979), .A2(n3142), .ZN(n3977) );
  XNOR2_X1 U4913 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U4914 ( .A1(n3983), .A2(n3980), .ZN(n3979) );
  NAND2_X1 U4915 ( .A1(n6354), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U4916 ( .A1(n3979), .A2(n3978), .ZN(n4003) );
  XNOR2_X1 U4917 ( .A(n3067), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4001)
         );
  XNOR2_X1 U4918 ( .A(n4003), .B(n4001), .ZN(n4075) );
  NAND2_X1 U4919 ( .A1(n4020), .A2(n4075), .ZN(n3999) );
  AOI21_X1 U4920 ( .B1(n4020), .B2(n4306), .A(n3204), .ZN(n3995) );
  INV_X1 U4921 ( .A(n3980), .ZN(n3981) );
  XNOR2_X1 U4922 ( .A(n3981), .B(n3983), .ZN(n4074) );
  NAND2_X1 U4923 ( .A1(n4074), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3994) );
  AND2_X1 U4924 ( .A1(n3066), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3982)
         );
  NOR2_X1 U4925 ( .A1(n3983), .A2(n3982), .ZN(n3987) );
  OAI21_X1 U4926 ( .B1(n3204), .B2(n3984), .A(n3987), .ZN(n3985) );
  NAND2_X1 U4927 ( .A1(n3985), .A2(n3203), .ZN(n3986) );
  AOI22_X1 U4928 ( .A1(n3995), .A2(n3994), .B1(n4000), .B2(n3986), .ZN(n3988)
         );
  NAND3_X1 U4929 ( .A1(n3988), .A2(n3987), .A3(n4020), .ZN(n3993) );
  INV_X1 U4930 ( .A(n3988), .ZN(n3989) );
  NAND2_X1 U4931 ( .A1(n3989), .A2(n4074), .ZN(n3991) );
  NAND2_X1 U4932 ( .A1(n3991), .A2(n4025), .ZN(n3992) );
  OAI211_X1 U4933 ( .C1(n3995), .C2(n3994), .A(n3993), .B(n3992), .ZN(n3997)
         );
  OAI211_X1 U4934 ( .C1(n4075), .C2(n4013), .A(n3999), .B(n4000), .ZN(n3996)
         );
  NAND2_X1 U4935 ( .A1(n3997), .A2(n3996), .ZN(n3998) );
  OAI21_X1 U4936 ( .B1(n4000), .B2(n3999), .A(n3998), .ZN(n4015) );
  INV_X1 U4937 ( .A(n4001), .ZN(n4002) );
  NAND2_X1 U4938 ( .A1(n4003), .A2(n4002), .ZN(n4005) );
  NAND2_X1 U4939 ( .A1(n6558), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4004) );
  NAND2_X1 U4940 ( .A1(n4005), .A2(n4004), .ZN(n4010) );
  XNOR2_X1 U4941 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U4942 ( .A1(n4010), .A2(n4008), .ZN(n4007) );
  NAND2_X1 U4943 ( .A1(n6358), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4944 ( .A1(n4007), .A2(n4006), .ZN(n4017) );
  INV_X1 U4945 ( .A(n4008), .ZN(n4009) );
  XNOR2_X1 U4946 ( .A(n4010), .B(n4009), .ZN(n4011) );
  NAND2_X1 U4947 ( .A1(n4012), .A2(n4011), .ZN(n4078) );
  NAND2_X1 U4948 ( .A1(n4013), .A2(n4078), .ZN(n4014) );
  NAND2_X1 U4949 ( .A1(n4015), .A2(n4014), .ZN(n4024) );
  NAND2_X1 U4950 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5454), .ZN(n4018) );
  AOI22_X1 U4951 ( .A1(n4020), .A2(n4026), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6634), .ZN(n4022) );
  NAND2_X1 U4952 ( .A1(n4025), .A2(n4078), .ZN(n4021) );
  INV_X1 U4953 ( .A(n4025), .ZN(n4027) );
  NAND2_X1 U4954 ( .A1(n6343), .A2(n4748), .ZN(n4034) );
  INV_X1 U4955 ( .A(n4032), .ZN(n4242) );
  NOR2_X1 U4956 ( .A1(n4031), .A2(n4242), .ZN(n4033) );
  NAND2_X1 U4957 ( .A1(n4034), .A2(n4033), .ZN(n4234) );
  NAND2_X1 U4958 ( .A1(n5211), .A2(n5785), .ZN(n4042) );
  NAND2_X1 U4959 ( .A1(n6278), .A2(n4035), .ZN(n6485) );
  AND2_X1 U4960 ( .A1(n6485), .A2(n6634), .ZN(n4036) );
  NAND2_X1 U4961 ( .A1(n6634), .A2(n3391), .ZN(n6391) );
  INV_X1 U4962 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U4963 ( .A1(n5845), .A2(n6454), .ZN(n5215) );
  NAND2_X1 U4964 ( .A1(n6634), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U4965 ( .A1(n6167), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4037) );
  AND2_X1 U4966 ( .A1(n4038), .A2(n4037), .ZN(n5783) );
  INV_X1 U4967 ( .A(n5783), .ZN(n4039) );
  NOR2_X1 U4968 ( .A1(n5777), .A2(n4881), .ZN(n4040) );
  AOI211_X1 U4969 ( .C1(PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n5771), .A(n5215), 
        .B(n4040), .ZN(n4041) );
  OAI211_X1 U4970 ( .C1(n5084), .C2(n6282), .A(n4042), .B(n4041), .ZN(U2956)
         );
  INV_X1 U4971 ( .A(n4215), .ZN(n4046) );
  AND2_X1 U4972 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4298) );
  INV_X1 U4973 ( .A(n4043), .ZN(n5134) );
  INV_X1 U4974 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4047) );
  XNOR2_X1 U4975 ( .A(n4048), .B(n4047), .ZN(n4302) );
  AOI22_X1 U4976 ( .A1(n4050), .A2(EAX_REG_31__SCAN_IN), .B1(n4049), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4051) );
  INV_X1 U4977 ( .A(n4051), .ZN(n4052) );
  XNOR2_X2 U4978 ( .A(n4053), .B(n4052), .ZN(n4833) );
  NAND2_X1 U4979 ( .A1(n4833), .A2(n5774), .ZN(n4059) );
  INV_X1 U4980 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4194) );
  INV_X2 U4981 ( .A(n5845), .ZN(n5817) );
  NAND2_X1 U4982 ( .A1(n5817), .A2(REIP_REG_31__SCAN_IN), .ZN(n4299) );
  NAND2_X1 U4983 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4056)
         );
  OAI211_X1 U4984 ( .C1(n5777), .C2(n4755), .A(n4299), .B(n4056), .ZN(n4057)
         );
  INV_X1 U4985 ( .A(n4057), .ZN(n4058) );
  NAND3_X1 U4986 ( .A1(n4060), .A2(n4059), .A3(n4058), .ZN(U2955) );
  NAND2_X1 U4987 ( .A1(n4043), .A2(n5123), .ZN(n5113) );
  NAND2_X1 U4988 ( .A1(n5221), .A2(n5785), .ZN(n4069) );
  INV_X1 U4989 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6449) );
  NOR2_X1 U4990 ( .A1(n5845), .A2(n6449), .ZN(n5225) );
  NOR2_X1 U4991 ( .A1(n5777), .A2(n4903), .ZN(n4063) );
  AOI211_X1 U4992 ( .C1(n5771), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5225), 
        .B(n4063), .ZN(n4068) );
  NAND3_X1 U4993 ( .A1(n4069), .A2(n4068), .A3(n4067), .ZN(U2958) );
  NOR2_X1 U4994 ( .A1(n4071), .A2(n3203), .ZN(n4072) );
  NAND2_X1 U4995 ( .A1(n4075), .A2(n4074), .ZN(n4077) );
  OAI21_X1 U4996 ( .B1(n4078), .B2(n4077), .A(n4076), .ZN(n4861) );
  INV_X1 U4997 ( .A(n4861), .ZN(n4866) );
  NAND3_X1 U4998 ( .A1(n4867), .A2(n4839), .A3(n4866), .ZN(n4303) );
  NAND2_X1 U4999 ( .A1(n6468), .A2(n3391), .ZN(n6380) );
  NOR3_X1 U5000 ( .A1(n6634), .A2(n6466), .A3(n6380), .ZN(n6375) );
  NOR3_X1 U5001 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6391), .A3(n6468), .ZN(
        n6387) );
  INV_X1 U5002 ( .A(n6387), .ZN(n4079) );
  NAND2_X1 U5003 ( .A1(n5845), .A2(n4079), .ZN(n4080) );
  NAND2_X1 U5004 ( .A1(n4833), .A2(n5555), .ZN(n4212) );
  INV_X1 U5005 ( .A(n4362), .ZN(n4187) );
  NAND2_X1 U5006 ( .A1(n4187), .A2(EBX_REG_30__SCAN_IN), .ZN(n4085) );
  NAND2_X1 U5007 ( .A1(n4186), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4084) );
  AND2_X1 U5008 ( .A1(n4085), .A2(n4084), .ZN(n4875) );
  INV_X1 U5009 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4086) );
  NAND2_X1 U5010 ( .A1(n4334), .A2(n4086), .ZN(n4087) );
  OAI211_X1 U5011 ( .C1(n4185), .C2(n3964), .A(n4087), .B(n4180), .ZN(n4088)
         );
  OAI21_X1 U5012 ( .B1(n4178), .B2(EBX_REG_15__SCAN_IN), .A(n4088), .ZN(n4822)
         );
  INV_X1 U5013 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4715) );
  INV_X1 U5014 ( .A(n4178), .ZN(n4166) );
  AOI22_X1 U5015 ( .A1(n4166), .A2(n4715), .B1(n4362), .B2(n5815), .ZN(n4089)
         );
  OAI21_X1 U5016 ( .B1(n4111), .B2(n4715), .A(n4089), .ZN(n4714) );
  NAND2_X1 U5017 ( .A1(n4185), .A2(EBX_REG_5__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5018 ( .A1(n4362), .A2(n4599), .ZN(n4090) );
  OAI211_X1 U5019 ( .C1(EBX_REG_5__SCAN_IN), .C2(n4178), .A(n4091), .B(n4090), 
        .ZN(n4480) );
  NAND2_X1 U5020 ( .A1(n4185), .A2(EBX_REG_3__SCAN_IN), .ZN(n4093) );
  NAND2_X1 U5021 ( .A1(n4362), .A2(n4371), .ZN(n4092) );
  OAI211_X1 U5022 ( .C1(EBX_REG_3__SCAN_IN), .C2(n4178), .A(n4093), .B(n4092), 
        .ZN(n4373) );
  INV_X1 U5023 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4335) );
  NAND2_X1 U5024 ( .A1(n4103), .A2(n4335), .ZN(n4096) );
  NAND2_X1 U5025 ( .A1(n4334), .A2(n4335), .ZN(n4094) );
  OAI211_X1 U5026 ( .C1(n4172), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4094), 
        .B(n4111), .ZN(n4095) );
  NAND2_X1 U5027 ( .A1(n4096), .A2(n4095), .ZN(n4099) );
  INV_X1 U5028 ( .A(n4099), .ZN(n4101) );
  NAND2_X1 U5029 ( .A1(n4180), .A2(EBX_REG_0__SCAN_IN), .ZN(n4098) );
  INV_X1 U5030 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5031 ( .A1(n4111), .A2(n4365), .ZN(n4097) );
  XNOR2_X1 U5032 ( .A(n4099), .B(n4361), .ZN(n5626) );
  NOR2_X1 U5033 ( .A1(n5626), .A2(n4186), .ZN(n4100) );
  OR2_X1 U5034 ( .A1(n4334), .A2(n3908), .ZN(n4106) );
  NAND2_X1 U5035 ( .A1(n4172), .A2(n4186), .ZN(n4159) );
  NAND2_X1 U5036 ( .A1(n4172), .A2(EBX_REG_2__SCAN_IN), .ZN(n4102) );
  AND2_X1 U5037 ( .A1(n4159), .A2(n4102), .ZN(n4105) );
  INV_X1 U5038 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U5039 ( .A1(n4103), .A2(n4359), .ZN(n4104) );
  NAND3_X1 U5040 ( .A1(n4106), .A2(n4105), .A3(n4104), .ZN(n4358) );
  INV_X1 U5041 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U5042 ( .A1(n4103), .A2(n5585), .ZN(n4109) );
  NAND2_X1 U5043 ( .A1(n4334), .A2(n5585), .ZN(n4107) );
  OAI211_X1 U5044 ( .C1(n4172), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4107), 
        .B(n4111), .ZN(n4108) );
  NAND2_X1 U5045 ( .A1(n4109), .A2(n4108), .ZN(n4444) );
  INV_X1 U5046 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4110) );
  NAND2_X1 U5047 ( .A1(n4334), .A2(n4110), .ZN(n4112) );
  OAI211_X1 U5048 ( .C1(n4172), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4112), 
        .B(n4111), .ZN(n4113) );
  OAI21_X1 U5049 ( .B1(n4183), .B2(EBX_REG_6__SCAN_IN), .A(n4113), .ZN(n4490)
         );
  NAND2_X1 U5050 ( .A1(n4481), .A2(n4490), .ZN(n4626) );
  NAND2_X1 U5051 ( .A1(n4185), .A2(EBX_REG_7__SCAN_IN), .ZN(n4116) );
  NAND2_X1 U5052 ( .A1(n4362), .A2(n4114), .ZN(n4115) );
  OAI211_X1 U5053 ( .C1(EBX_REG_7__SCAN_IN), .C2(n4178), .A(n4116), .B(n4115), 
        .ZN(n4627) );
  INV_X1 U5054 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5055 ( .A1(n4103), .A2(n4699), .ZN(n4119) );
  NAND2_X1 U5056 ( .A1(n4334), .A2(n4699), .ZN(n4117) );
  OAI211_X1 U5057 ( .C1(n4172), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4117), 
        .B(n4111), .ZN(n4118) );
  NAND2_X1 U5058 ( .A1(n4119), .A2(n4118), .ZN(n4680) );
  OR2_X1 U5059 ( .A1(n4334), .A2(n5807), .ZN(n4124) );
  NAND2_X1 U5060 ( .A1(n4172), .A2(EBX_REG_10__SCAN_IN), .ZN(n4120) );
  AND2_X1 U5061 ( .A1(n4159), .A2(n4120), .ZN(n4123) );
  INV_X1 U5062 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4121) );
  NAND2_X1 U5063 ( .A1(n4103), .A2(n4121), .ZN(n4122) );
  NAND3_X1 U5064 ( .A1(n4124), .A2(n4123), .A3(n4122), .ZN(n4723) );
  INV_X1 U5065 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4125) );
  NAND2_X1 U5066 ( .A1(n4334), .A2(n4125), .ZN(n4126) );
  OAI211_X1 U5067 ( .C1(n4185), .C2(n5790), .A(n4126), .B(n4180), .ZN(n4127)
         );
  OAI21_X1 U5068 ( .B1(n4178), .B2(EBX_REG_11__SCAN_IN), .A(n4127), .ZN(n4737)
         );
  OR2_X1 U5069 ( .A1(n4334), .A2(n4128), .ZN(n4132) );
  NAND2_X1 U5070 ( .A1(n4172), .A2(EBX_REG_12__SCAN_IN), .ZN(n4129) );
  AND2_X1 U5071 ( .A1(n4159), .A2(n4129), .ZN(n4131) );
  INV_X1 U5072 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U5073 ( .A1(n4103), .A2(n5514), .ZN(n4130) );
  NAND3_X1 U5074 ( .A1(n4132), .A2(n4131), .A3(n4130), .ZN(n4775) );
  INV_X1 U5075 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U5076 ( .A1(n4334), .A2(n4805), .ZN(n4133) );
  OAI211_X1 U5077 ( .C1(n4185), .C2(n5318), .A(n4133), .B(n4180), .ZN(n4134)
         );
  OAI21_X1 U5078 ( .B1(n4178), .B2(EBX_REG_13__SCAN_IN), .A(n4134), .ZN(n4804)
         );
  OR2_X1 U5079 ( .A1(n4334), .A2(n5321), .ZN(n4138) );
  NAND2_X1 U5080 ( .A1(n4172), .A2(EBX_REG_14__SCAN_IN), .ZN(n4135) );
  AND2_X1 U5081 ( .A1(n4159), .A2(n4135), .ZN(n4137) );
  INV_X1 U5082 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5083 ( .A1(n4103), .A2(n5077), .ZN(n4136) );
  NAND3_X1 U5084 ( .A1(n4138), .A2(n4137), .A3(n4136), .ZN(n5071) );
  INV_X1 U5085 ( .A(n4159), .ZN(n4139) );
  AOI21_X1 U5086 ( .B1(n4172), .B2(EBX_REG_16__SCAN_IN), .A(n4139), .ZN(n4141)
         );
  NAND2_X1 U5087 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4186), .ZN(n4140) );
  OAI211_X1 U5088 ( .C1(EBX_REG_16__SCAN_IN), .C2(n4183), .A(n4141), .B(n4140), 
        .ZN(n4978) );
  NAND2_X1 U5089 ( .A1(n4111), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4142) );
  OAI211_X1 U5090 ( .C1(n4186), .C2(EBX_REG_17__SCAN_IN), .A(n4180), .B(n4142), 
        .ZN(n4143) );
  OAI21_X1 U5091 ( .B1(n4178), .B2(EBX_REG_17__SCAN_IN), .A(n4143), .ZN(n4962)
         );
  INV_X1 U5092 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U5093 ( .A1(n4103), .A2(n4144), .ZN(n4147) );
  NAND2_X1 U5094 ( .A1(n4180), .A2(n5138), .ZN(n4145) );
  OAI211_X1 U5095 ( .C1(n4186), .C2(EBX_REG_19__SCAN_IN), .A(n4111), .B(n4145), 
        .ZN(n4146) );
  INV_X1 U5096 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4153) );
  INV_X1 U5097 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U5098 ( .A1(n4362), .A2(n5436), .ZN(n4148) );
  OR2_X1 U5099 ( .A1(n4186), .A2(EBX_REG_18__SCAN_IN), .ZN(n5046) );
  OR2_X1 U5100 ( .A1(n4186), .A2(EBX_REG_20__SCAN_IN), .ZN(n4149) );
  OAI21_X1 U5101 ( .B1(n4187), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n4149), 
        .ZN(n5039) );
  NAND2_X1 U5102 ( .A1(n5045), .A2(n5039), .ZN(n4152) );
  INV_X1 U5103 ( .A(n5045), .ZN(n4150) );
  NAND2_X1 U5104 ( .A1(n4150), .A2(n4111), .ZN(n4151) );
  OAI211_X1 U5105 ( .C1(n4111), .C2(n4153), .A(n4152), .B(n4151), .ZN(n4154)
         );
  INV_X1 U5106 ( .A(n4154), .ZN(n4155) );
  NAND2_X1 U5107 ( .A1(n5038), .A2(n4155), .ZN(n5030) );
  NAND2_X1 U5108 ( .A1(n4111), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4156) );
  OAI211_X1 U5109 ( .C1(n4186), .C2(EBX_REG_21__SCAN_IN), .A(n4180), .B(n4156), 
        .ZN(n4157) );
  OAI21_X1 U5110 ( .B1(n4178), .B2(EBX_REG_21__SCAN_IN), .A(n4157), .ZN(n5029)
         );
  NAND2_X1 U5111 ( .A1(n4172), .A2(EBX_REG_22__SCAN_IN), .ZN(n4158) );
  AND2_X1 U5112 ( .A1(n4159), .A2(n4158), .ZN(n4161) );
  NAND2_X1 U5113 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n4186), .ZN(n4160) );
  OAI211_X1 U5114 ( .C1(n4183), .C2(EBX_REG_22__SCAN_IN), .A(n4161), .B(n4160), 
        .ZN(n4162) );
  INV_X1 U5115 ( .A(n4162), .ZN(n5018) );
  INV_X1 U5116 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U5117 ( .A1(n4166), .A2(n4951), .ZN(n4165) );
  NAND2_X1 U5118 ( .A1(n4111), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4163) );
  OAI211_X1 U5119 ( .C1(n4186), .C2(EBX_REG_23__SCAN_IN), .A(n4180), .B(n4163), 
        .ZN(n4164) );
  AND2_X1 U5120 ( .A1(n4165), .A2(n4164), .ZN(n4952) );
  AOI22_X1 U5121 ( .A1(n4362), .A2(n6589), .B1(EBX_REG_25__SCAN_IN), .B2(n4185), .ZN(n4168) );
  INV_X1 U5122 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5123 ( .A1(n4166), .A2(n5014), .ZN(n4167) );
  AND2_X1 U5124 ( .A1(n4168), .A2(n4167), .ZN(n5010) );
  AOI22_X1 U5125 ( .A1(n4172), .A2(EBX_REG_24__SCAN_IN), .B1(n4186), .B2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4169) );
  OAI21_X1 U5126 ( .B1(n4183), .B2(EBX_REG_24__SCAN_IN), .A(n4169), .ZN(n5008)
         );
  AND2_X1 U5127 ( .A1(n5010), .A2(n5008), .ZN(n4170) );
  INV_X1 U5128 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U5129 ( .A1(n4103), .A2(n4171), .ZN(n4174) );
  AOI22_X1 U5130 ( .A1(n4172), .A2(EBX_REG_26__SCAN_IN), .B1(n4186), .B2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4173) );
  AND2_X1 U5131 ( .A1(n4174), .A2(n4173), .ZN(n4927) );
  INV_X1 U5132 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5238) );
  INV_X1 U5133 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4175) );
  NOR2_X1 U5134 ( .A1(n4111), .A2(n4175), .ZN(n4176) );
  AOI21_X1 U5135 ( .B1(n4362), .B2(n5238), .A(n4176), .ZN(n4177) );
  OAI21_X1 U5136 ( .B1(n4178), .B2(EBX_REG_27__SCAN_IN), .A(n4177), .ZN(n4914)
         );
  INV_X1 U5137 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4179) );
  NAND2_X1 U5138 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  OAI211_X1 U5139 ( .C1(n4186), .C2(EBX_REG_28__SCAN_IN), .A(n4111), .B(n4181), 
        .ZN(n4182) );
  OAI21_X1 U5140 ( .B1(n4183), .B2(EBX_REG_28__SCAN_IN), .A(n4182), .ZN(n4901)
         );
  INV_X1 U5141 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U5142 ( .A1(n4362), .A2(n6498), .B1(n4334), .B2(n4893), .ZN(n4275)
         );
  NOR2_X1 U5143 ( .A1(n4183), .A2(EBX_REG_29__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U5144 ( .A1(n4877), .A2(n4276), .ZN(n4184) );
  NOR2_X1 U5145 ( .A1(n4874), .A2(n4185), .ZN(n4880) );
  AOI21_X1 U5146 ( .B1(n4875), .B2(n4281), .A(n4880), .ZN(n4189) );
  OAI22_X1 U5147 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4187), .B1(n4186), .B2(EBX_REG_31__SCAN_IN), .ZN(n4188) );
  NOR2_X1 U5148 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4746) );
  NAND2_X1 U5149 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4751), .ZN(n4193) );
  NOR2_X1 U5150 ( .A1(n4746), .A2(n4193), .ZN(n4190) );
  NAND2_X1 U5151 ( .A1(n4191), .A2(n6405), .ZN(n6398) );
  INV_X1 U5152 ( .A(n4746), .ZN(n4192) );
  OR2_X1 U5153 ( .A1(n6398), .A2(n4192), .ZN(n6369) );
  NAND2_X1 U5154 ( .A1(n2978), .A2(n6369), .ZN(n4750) );
  OAI22_X1 U5155 ( .A1(n5603), .A2(n4194), .B1(n4193), .B2(n4750), .ZN(n4201)
         );
  INV_X1 U5156 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6437) );
  INV_X1 U5157 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U5158 ( .A1(n4746), .A2(n4751), .ZN(n4195) );
  NOR2_X1 U5159 ( .A1(n4748), .A2(n4195), .ZN(n4196) );
  NAND2_X1 U5160 ( .A1(n2979), .A2(n6398), .ZN(n4227) );
  INV_X1 U5161 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6517) );
  NAND3_X1 U5162 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4990) );
  NAND3_X1 U5163 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U5164 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5524) );
  NOR3_X1 U5165 ( .A1(n4990), .A2(n4985), .A3(n5524), .ZN(n4197) );
  NAND4_X1 U5166 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        REIP_REG_4__SCAN_IN), .A4(n4197), .ZN(n5508) );
  NOR2_X1 U5167 ( .A1(n6517), .A2(n5508), .ZN(n5491) );
  NAND3_X1 U5168 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        n5491), .ZN(n4202) );
  NAND3_X1 U5169 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n4974), .ZN(n4961) );
  NAND3_X1 U5170 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        n5380), .ZN(n5370) );
  NAND4_X1 U5171 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5356), .ZN(n4940) );
  NAND3_X1 U5172 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4913) );
  INV_X1 U5173 ( .A(n4913), .ZN(n4198) );
  NAND2_X1 U5174 ( .A1(REIP_REG_27__SCAN_IN), .A2(n4198), .ZN(n4199) );
  NOR2_X1 U5175 ( .A1(n4940), .A2(n4199), .ZN(n4900) );
  NAND2_X1 U5176 ( .A1(n4900), .A2(REIP_REG_28__SCAN_IN), .ZN(n4208) );
  INV_X1 U5177 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6452) );
  NOR4_X1 U5178 ( .A1(n4208), .A2(REIP_REG_31__SCAN_IN), .A3(n6454), .A4(n6452), .ZN(n4200) );
  AOI211_X1 U5179 ( .C1(n4297), .C2(n5595), .A(n4201), .B(n4200), .ZN(n4210)
         );
  INV_X1 U5180 ( .A(n5597), .ZN(n5492) );
  NAND2_X1 U5181 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4207) );
  INV_X1 U5182 ( .A(n4986), .ZN(n4989) );
  INV_X1 U5183 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6435) );
  INV_X1 U5184 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6434) );
  NOR2_X1 U5185 ( .A1(n6435), .A2(n6434), .ZN(n4203) );
  NAND2_X1 U5186 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4973) );
  OAI21_X1 U5187 ( .B1(n4202), .B2(n2955), .A(n4986), .ZN(n5500) );
  INV_X1 U5188 ( .A(n5500), .ZN(n4972) );
  AOI221_X1 U5189 ( .B1(n6432), .B2(n4986), .C1(n4973), .C2(n4986), .A(n4972), 
        .ZN(n5480) );
  OAI221_X1 U5190 ( .B1(n4989), .B2(REIP_REG_20__SCAN_IN), .C1(n4989), .C2(
        n4203), .A(n5480), .ZN(n5361) );
  INV_X1 U5191 ( .A(n5361), .ZN(n5369) );
  INV_X1 U5192 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6442) );
  INV_X1 U5193 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6440) );
  INV_X1 U5194 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6438) );
  OR3_X1 U5195 ( .A1(n6442), .A2(n6440), .A3(n6438), .ZN(n4204) );
  NAND2_X1 U5196 ( .A1(n4986), .A2(n4204), .ZN(n4205) );
  NAND2_X1 U5197 ( .A1(n5369), .A2(n4205), .ZN(n5343) );
  AND2_X1 U5198 ( .A1(n4986), .A2(n4913), .ZN(n4206) );
  AOI21_X1 U5199 ( .B1(n5492), .B2(n4207), .A(n4934), .ZN(n4892) );
  OR2_X1 U5200 ( .A1(n4208), .A2(REIP_REG_29__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U5201 ( .A1(n4892), .A2(n4896), .ZN(n4888) );
  NOR3_X1 U5202 ( .A1(n4208), .A2(REIP_REG_30__SCAN_IN), .A3(n6452), .ZN(n4887) );
  OAI21_X1 U5203 ( .B1(n4888), .B2(n4887), .A(REIP_REG_31__SCAN_IN), .ZN(n4209) );
  NAND2_X1 U5204 ( .A1(n4212), .A2(n4211), .ZN(U2796) );
  NAND2_X1 U5205 ( .A1(n5123), .A2(n5226), .ZN(n4213) );
  NAND2_X1 U5206 ( .A1(n4215), .A2(n4214), .ZN(n4216) );
  XNOR2_X1 U5207 ( .A(n4216), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5112)
         );
  NOR2_X1 U5208 ( .A1(n6343), .A2(n4394), .ZN(n4255) );
  INV_X1 U5209 ( .A(n4255), .ZN(n4225) );
  OR2_X1 U5210 ( .A1(n4217), .A2(n4831), .ZN(n4611) );
  INV_X1 U5211 ( .A(n4611), .ZN(n4612) );
  NAND2_X1 U5212 ( .A1(n4612), .A2(n4218), .ZN(n4220) );
  OAI21_X1 U5213 ( .B1(n4217), .B2(n4748), .A(n6488), .ZN(n4219) );
  NAND2_X1 U5214 ( .A1(n4220), .A2(n4219), .ZN(n4246) );
  INV_X1 U5215 ( .A(n4246), .ZN(n4222) );
  INV_X1 U5216 ( .A(n4867), .ZN(n4221) );
  OAI21_X1 U5217 ( .B1(n4222), .B2(n4234), .A(n4221), .ZN(n4393) );
  NAND2_X1 U5218 ( .A1(n4306), .A2(n6398), .ZN(n4223) );
  NOR2_X1 U5219 ( .A1(READY_N), .A2(n4861), .ZN(n4391) );
  NAND3_X1 U5220 ( .A1(n4223), .A2(n4391), .A3(n4562), .ZN(n4224) );
  OAI211_X1 U5221 ( .C1(n4865), .C2(n4225), .A(n4393), .B(n4224), .ZN(n4226)
         );
  NAND2_X1 U5222 ( .A1(n4226), .A2(n4839), .ZN(n4233) );
  INV_X1 U5223 ( .A(n2966), .ZN(n4404) );
  INV_X1 U5224 ( .A(READY_N), .ZN(n6486) );
  AND2_X1 U5225 ( .A1(n4227), .A2(n6486), .ZN(n4388) );
  NAND2_X1 U5226 ( .A1(n2966), .A2(n4388), .ZN(n4230) );
  AND2_X1 U5227 ( .A1(n3203), .A2(n4228), .ZN(n4229) );
  AOI21_X1 U5228 ( .B1(n4230), .B2(n4229), .A(n4562), .ZN(n4231) );
  NAND2_X1 U5229 ( .A1(n4609), .A2(n4231), .ZN(n4232) );
  NOR2_X1 U5230 ( .A1(n4234), .A2(n3976), .ZN(n4608) );
  NOR2_X1 U5231 ( .A1(n4608), .A2(n2999), .ZN(n4859) );
  OAI21_X1 U5232 ( .B1(n4527), .B2(n4282), .A(n4235), .ZN(n4236) );
  AOI21_X1 U5233 ( .B1(n4237), .B2(n4306), .A(n4236), .ZN(n4238) );
  NAND2_X1 U5234 ( .A1(n4859), .A2(n4238), .ZN(n4239) );
  AOI21_X1 U5235 ( .B1(n4834), .B2(n4748), .A(n4240), .ZN(n4241) );
  AOI21_X1 U5236 ( .B1(n4031), .B2(n4185), .A(n4241), .ZN(n4245) );
  NAND2_X1 U5237 ( .A1(n4362), .A2(n4394), .ZN(n4243) );
  NAND2_X1 U5238 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  AND3_X1 U5239 ( .A1(n4246), .A2(n4245), .A3(n4244), .ZN(n4247) );
  NAND2_X1 U5240 ( .A1(n4248), .A2(n4247), .ZN(n4406) );
  OR3_X1 U5241 ( .A1(n6343), .A2(n3203), .A3(n4250), .ZN(n4424) );
  OR2_X1 U5242 ( .A1(n4251), .A2(n4252), .ZN(n4253) );
  OAI211_X1 U5243 ( .C1(n4249), .C2(n3203), .A(n4424), .B(n4253), .ZN(n4254)
         );
  NOR2_X1 U5244 ( .A1(n4406), .A2(n4254), .ZN(n4256) );
  NAND2_X1 U5245 ( .A1(n4256), .A2(n4255), .ZN(n4413) );
  INV_X1 U5246 ( .A(n4413), .ZN(n4860) );
  NAND2_X1 U5247 ( .A1(n4284), .A2(n4860), .ZN(n4790) );
  INV_X1 U5248 ( .A(n4284), .ZN(n4257) );
  NOR2_X1 U5249 ( .A1(n4257), .A2(n4256), .ZN(n5320) );
  NOR2_X1 U5250 ( .A1(n5830), .A2(n5320), .ZN(n5839) );
  OAI22_X1 U5251 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5839), .B1(n5817), 
        .B2(n4284), .ZN(n5840) );
  NOR2_X1 U5252 ( .A1(n5830), .A2(n5840), .ZN(n5291) );
  NOR2_X1 U5253 ( .A1(n5790), .A2(n4128), .ZN(n4813) );
  NAND2_X1 U5254 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4813), .ZN(n5324) );
  OR2_X1 U5255 ( .A1(n5321), .A2(n5324), .ZN(n5309) );
  NAND2_X1 U5256 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5310) );
  NOR2_X1 U5257 ( .A1(n5309), .A2(n5310), .ZN(n4261) );
  NAND2_X1 U5258 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U5259 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5804) );
  NOR2_X1 U5260 ( .A1(n5803), .A2(n5804), .ZN(n4260) );
  NAND2_X1 U5261 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4446) );
  NAND2_X1 U5262 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4369) );
  NOR2_X1 U5263 ( .A1(n4446), .A2(n4369), .ZN(n4594) );
  AND3_X1 U5264 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4594), .ZN(n4677) );
  AND2_X1 U5265 ( .A1(n4260), .A2(n4677), .ZN(n4786) );
  NAND2_X1 U5266 ( .A1(n4261), .A2(n4786), .ZN(n5287) );
  INV_X1 U5267 ( .A(n5287), .ZN(n4258) );
  NAND2_X1 U5268 ( .A1(n5291), .A2(n4258), .ZN(n4263) );
  AOI21_X1 U5269 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4370) );
  NOR2_X1 U5270 ( .A1(n4370), .A2(n4446), .ZN(n4554) );
  NAND2_X1 U5271 ( .A1(n5830), .A2(n4554), .ZN(n4598) );
  NAND2_X1 U5272 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4259) );
  NOR2_X1 U5273 ( .A1(n4598), .A2(n4259), .ZN(n4678) );
  NAND2_X1 U5274 ( .A1(n4678), .A2(n4260), .ZN(n4288) );
  INV_X1 U5275 ( .A(n4288), .ZN(n5319) );
  AND2_X1 U5276 ( .A1(n5319), .A2(n4261), .ZN(n5290) );
  INV_X1 U5277 ( .A(n5290), .ZN(n4262) );
  NAND2_X1 U5278 ( .A1(n4263), .A2(n4262), .ZN(n4265) );
  INV_X1 U5279 ( .A(n5301), .ZN(n4264) );
  AND2_X1 U5280 ( .A1(n4264), .A2(n5286), .ZN(n5153) );
  NAND2_X1 U5281 ( .A1(n4265), .A2(n5153), .ZN(n4267) );
  NAND2_X1 U5282 ( .A1(n5291), .A2(n4787), .ZN(n4266) );
  NAND2_X1 U5283 ( .A1(n4267), .A2(n4266), .ZN(n5269) );
  INV_X1 U5284 ( .A(n5841), .ZN(n4268) );
  NAND2_X1 U5285 ( .A1(n5839), .A2(n4268), .ZN(n5797) );
  NAND2_X1 U5286 ( .A1(n5797), .A2(n5152), .ZN(n4269) );
  NAND2_X1 U5287 ( .A1(n5269), .A2(n4269), .ZN(n5264) );
  NOR2_X1 U5288 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5841), .ZN(n4381)
         );
  OAI21_X1 U5289 ( .B1(n5819), .B2(n5830), .A(n4270), .ZN(n4271) );
  INV_X1 U5290 ( .A(n4271), .ZN(n4272) );
  AND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4291) );
  INV_X1 U5292 ( .A(n4291), .ZN(n5247) );
  AND2_X1 U5293 ( .A1(n5797), .A2(n5247), .ZN(n4273) );
  AND2_X1 U5294 ( .A1(n5797), .A2(n5227), .ZN(n4274) );
  NOR2_X1 U5295 ( .A1(n5232), .A2(n4274), .ZN(n4296) );
  NAND2_X1 U5296 ( .A1(n4275), .A2(n4111), .ZN(n4278) );
  INV_X1 U5297 ( .A(n4276), .ZN(n4277) );
  NAND2_X1 U5298 ( .A1(n4278), .A2(n4277), .ZN(n4279) );
  NOR2_X1 U5299 ( .A1(n4877), .A2(n4279), .ZN(n4280) );
  NOR2_X1 U5300 ( .A1(n4281), .A2(n4280), .ZN(n5001) );
  NAND2_X1 U5301 ( .A1(n2966), .A2(n2978), .ZN(n6370) );
  OAI21_X1 U5302 ( .B1(n4282), .B2(n2967), .A(n6370), .ZN(n4283) );
  NAND2_X1 U5303 ( .A1(n5817), .A2(REIP_REG_29__SCAN_IN), .ZN(n5106) );
  INV_X1 U5304 ( .A(n5106), .ZN(n4285) );
  AOI21_X1 U5305 ( .B1(n5001), .B2(n5836), .A(n4285), .ZN(n4286) );
  OAI21_X1 U5306 ( .B1(n4296), .B2(n6498), .A(n4286), .ZN(n4287) );
  INV_X1 U5307 ( .A(n4287), .ZN(n4294) );
  NAND2_X1 U5308 ( .A1(n4786), .A2(n5819), .ZN(n4789) );
  NAND2_X1 U5309 ( .A1(n4288), .A2(n4789), .ZN(n5791) );
  INV_X1 U5310 ( .A(n5448), .ZN(n4289) );
  NAND2_X1 U5311 ( .A1(n5271), .A2(n4290), .ZN(n5432) );
  NAND2_X1 U5312 ( .A1(n3973), .A2(n4291), .ZN(n4292) );
  NOR2_X1 U5313 ( .A1(n5432), .A2(n4292), .ZN(n5213) );
  INV_X1 U5314 ( .A(n5213), .ZN(n4293) );
  INV_X1 U5315 ( .A(n5797), .ZN(n5292) );
  OAI21_X1 U5316 ( .B1(n4298), .B2(n5292), .A(n4296), .ZN(n5217) );
  NAND3_X1 U5317 ( .A1(n5213), .A2(n4298), .A3(n4047), .ZN(n4300) );
  OAI21_X1 U5318 ( .B1(n4302), .B2(n5825), .A(n4301), .ZN(U2987) );
  INV_X1 U5319 ( .A(n4303), .ZN(n4305) );
  INV_X1 U5320 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6577) );
  NOR2_X1 U5321 ( .A1(n6278), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4824) );
  INV_X1 U5322 ( .A(n4824), .ZN(n4304) );
  OAI211_X1 U5323 ( .C1(n4305), .C2(n6577), .A(n4317), .B(n4304), .ZN(U2788)
         );
  INV_X1 U5324 ( .A(n6484), .ZN(n4309) );
  AND2_X1 U5325 ( .A1(n4748), .A2(n4306), .ZN(n4745) );
  INV_X1 U5326 ( .A(n4745), .ZN(n4307) );
  NAND2_X1 U5327 ( .A1(n6488), .A2(n4307), .ZN(n4871) );
  OAI21_X1 U5328 ( .B1(n4824), .B2(READREQUEST_REG_SCAN_IN), .A(n4309), .ZN(
        n4308) );
  OAI21_X1 U5329 ( .B1(n4309), .B2(n4871), .A(n4308), .ZN(U3474) );
  INV_X1 U5330 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4315) );
  INV_X1 U5331 ( .A(n6370), .ZN(n4310) );
  NAND2_X1 U5332 ( .A1(n4609), .A2(n6346), .ZN(n4311) );
  NAND2_X1 U5333 ( .A1(n5737), .A2(n4311), .ZN(n4313) );
  INV_X1 U5334 ( .A(n6398), .ZN(n4312) );
  NAND2_X1 U5335 ( .A1(n5670), .A2(n3203), .ZN(n5640) );
  NAND2_X1 U5336 ( .A1(n6634), .A2(n4437), .ZN(n5672) );
  NOR2_X4 U5337 ( .A1(n5670), .A2(n5663), .ZN(n5669) );
  AOI22_X1 U5338 ( .A1(DATAO_REG_18__SCAN_IN), .A2(n5669), .B1(n5663), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4314) );
  OAI21_X1 U5339 ( .B1(n4315), .B2(n5640), .A(n4314), .ZN(U2905) );
  NOR2_X1 U5340 ( .A1(n2978), .A2(n6486), .ZN(n4316) );
  NOR2_X1 U5341 ( .A1(n4317), .A2(n4316), .ZN(n5673) );
  INV_X1 U5342 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U5343 ( .A1(n6649), .A2(EAX_REG_14__SCAN_IN), .ZN(n4319) );
  INV_X1 U5344 ( .A(DATAI_14_), .ZN(n4318) );
  OR2_X1 U5345 ( .A1(n6653), .A2(n4318), .ZN(n5697) );
  OAI211_X1 U5346 ( .C1(n5673), .C2(n6574), .A(n4319), .B(n5697), .ZN(U2953)
         );
  INV_X1 U5347 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6538) );
  INV_X1 U5348 ( .A(DATAI_8_), .ZN(n4320) );
  OR2_X1 U5349 ( .A1(n6653), .A2(n4320), .ZN(n5717) );
  NAND2_X1 U5350 ( .A1(n6649), .A2(EAX_REG_24__SCAN_IN), .ZN(n4321) );
  OAI211_X1 U5351 ( .C1(n5673), .C2(n6538), .A(n5717), .B(n4321), .ZN(U2932)
         );
  INV_X1 U5352 ( .A(n4322), .ZN(n4325) );
  INV_X1 U5353 ( .A(n4323), .ZN(n4324) );
  NAND2_X1 U5354 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  AND2_X1 U5355 ( .A1(n4326), .A2(n4353), .ZN(n5773) );
  INV_X1 U5356 ( .A(n4839), .ZN(n6385) );
  NOR2_X1 U5357 ( .A1(n3158), .A2(n4327), .ZN(n4603) );
  AND2_X1 U5358 ( .A1(n4603), .A2(n4604), .ZN(n4331) );
  INV_X1 U5359 ( .A(n4328), .ZN(n4330) );
  NAND4_X1 U5360 ( .A1(n4331), .A2(n4334), .A3(n4330), .A4(n4329), .ZN(n4332)
         );
  NAND2_X1 U5361 ( .A1(n5076), .A2(n4831), .ZN(n5078) );
  XNOR2_X1 U5362 ( .A(n5626), .B(n4334), .ZN(n4380) );
  OAI22_X1 U5363 ( .A1(n5078), .A2(n4380), .B1(n4335), .B2(n5076), .ZN(n4336)
         );
  AOI21_X1 U5364 ( .B1(n5773), .B2(n4807), .A(n4336), .ZN(n4337) );
  INV_X1 U5365 ( .A(n4337), .ZN(U2858) );
  INV_X1 U5366 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5699) );
  AOI22_X1 U5367 ( .A1(n5663), .A2(UWORD_REG_14__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4338) );
  OAI21_X1 U5368 ( .B1(n5699), .B2(n5640), .A(n4338), .ZN(U2893) );
  INV_X1 U5369 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U5370 ( .A1(n5663), .A2(UWORD_REG_0__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4339) );
  OAI21_X1 U5371 ( .B1(n4340), .B2(n5640), .A(n4339), .ZN(U2907) );
  INV_X1 U5372 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5373 ( .A1(n5663), .A2(UWORD_REG_1__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4341) );
  OAI21_X1 U5374 ( .B1(n4342), .B2(n5640), .A(n4341), .ZN(U2906) );
  INV_X1 U5375 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6526) );
  AOI22_X1 U5376 ( .A1(n5663), .A2(UWORD_REG_3__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4343) );
  OAI21_X1 U5377 ( .B1(n6526), .B2(n5640), .A(n4343), .ZN(U2904) );
  INV_X1 U5378 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5692) );
  AOI22_X1 U5379 ( .A1(n5663), .A2(UWORD_REG_12__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4344) );
  OAI21_X1 U5380 ( .B1(n5692), .B2(n5640), .A(n4344), .ZN(U2895) );
  INV_X1 U5381 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U5382 ( .A1(n5663), .A2(UWORD_REG_5__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4345) );
  OAI21_X1 U5383 ( .B1(n4346), .B2(n5640), .A(n4345), .ZN(U2902) );
  INV_X1 U5384 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5687) );
  AOI22_X1 U5385 ( .A1(n5663), .A2(UWORD_REG_10__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4347) );
  OAI21_X1 U5386 ( .B1(n5687), .B2(n5640), .A(n4347), .ZN(U2897) );
  AOI22_X1 U5387 ( .A1(n5663), .A2(UWORD_REG_7__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5388 ( .B1(n3737), .B2(n5640), .A(n4348), .ZN(U2900) );
  AOI22_X1 U5389 ( .A1(n5663), .A2(UWORD_REG_9__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5390 ( .B1(n3773), .B2(n5640), .A(n4349), .ZN(U2898) );
  AOI22_X1 U5391 ( .A1(n5663), .A2(UWORD_REG_11__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4350) );
  OAI21_X1 U5392 ( .B1(n3816), .B2(n5640), .A(n4350), .ZN(U2896) );
  AOI22_X1 U5393 ( .A1(n5663), .A2(UWORD_REG_13__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4351) );
  OAI21_X1 U5394 ( .B1(n3853), .B2(n5640), .A(n4351), .ZN(U2894) );
  NAND3_X1 U5395 ( .A1(n4355), .A2(n4354), .A3(n4353), .ZN(n4356) );
  NAND2_X1 U5396 ( .A1(n4352), .A2(n4356), .ZN(n5765) );
  XOR2_X1 U5397 ( .A(n4358), .B(n4357), .Z(n5818) );
  INV_X1 U5398 ( .A(n5818), .ZN(n4360) );
  OAI222_X1 U5399 ( .A1(n5765), .A2(n5075), .B1(n5078), .B2(n4360), .C1(n5076), 
        .C2(n4359), .ZN(U2857) );
  INV_X1 U5400 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5780) );
  AOI21_X1 U5401 ( .B1(n4362), .B2(n5780), .A(n4361), .ZN(n5835) );
  INV_X1 U5402 ( .A(n5835), .ZN(n4366) );
  XNOR2_X1 U5403 ( .A(n4364), .B(n4363), .ZN(n5788) );
  OAI222_X1 U5404 ( .A1(n4366), .A2(n5078), .B1(n5076), .B2(n4365), .C1(n5075), 
        .C2(n5788), .ZN(U2859) );
  XNOR2_X1 U5405 ( .A(n4368), .B(n4367), .ZN(n4478) );
  AOI22_X1 U5406 ( .A1(n4790), .A2(n5840), .B1(n5288), .B2(n4369), .ZN(n5822)
         );
  NAND2_X1 U5407 ( .A1(n5830), .A2(n4370), .ZN(n5832) );
  NAND2_X1 U5408 ( .A1(n5822), .A2(n5832), .ZN(n4450) );
  INV_X1 U5409 ( .A(n4369), .ZN(n5829) );
  AOI21_X1 U5410 ( .B1(n5829), .B2(n5819), .A(n5830), .ZN(n4557) );
  NOR2_X1 U5411 ( .A1(n4370), .A2(n4557), .ZN(n4447) );
  AOI22_X1 U5412 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4450), .B1(n4447), 
        .B2(n4371), .ZN(n4375) );
  AOI21_X1 U5413 ( .B1(n4373), .B2(n4372), .A(n3000), .ZN(n4759) );
  INV_X1 U5414 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4763) );
  NOR2_X1 U5415 ( .A1(n5845), .A2(n4763), .ZN(n4474) );
  AOI21_X1 U5416 ( .B1(n5836), .B2(n4759), .A(n4474), .ZN(n4374) );
  OAI211_X1 U5417 ( .C1(n4478), .C2(n5825), .A(n4375), .B(n4374), .ZN(U3015)
         );
  OR2_X1 U5418 ( .A1(n4377), .A2(n4376), .ZN(n4379) );
  AND2_X1 U5419 ( .A1(n4379), .A2(n4378), .ZN(n5772) );
  INV_X1 U5420 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5615) );
  OAI22_X1 U5421 ( .A1(n5799), .A2(n4380), .B1(n5845), .B2(n5615), .ZN(n4384)
         );
  NOR2_X1 U5422 ( .A1(n5292), .A2(n4381), .ZN(n4382) );
  MUX2_X1 U5423 ( .A(n4382), .B(n5840), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4383) );
  AOI211_X1 U5424 ( .C1(n5837), .C2(n5772), .A(n4384), .B(n4383), .ZN(n4385)
         );
  INV_X1 U5425 ( .A(n4385), .ZN(U3017) );
  INV_X1 U5426 ( .A(n6170), .ZN(n5988) );
  NOR2_X1 U5427 ( .A1(n3319), .A2(n5988), .ZN(n4386) );
  XNOR2_X1 U5428 ( .A(n4386), .B(n5454), .ZN(n5583) );
  NOR2_X1 U5429 ( .A1(n4235), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U5430 ( .A1(n5583), .A2(n4387), .ZN(n5453) );
  INV_X1 U5431 ( .A(n4388), .ZN(n4389) );
  AOI21_X1 U5432 ( .B1(n4070), .B2(n6398), .A(n4389), .ZN(n4390) );
  OAI211_X1 U5433 ( .C1(n2966), .C2(n6346), .A(n4865), .B(n4390), .ZN(n4398)
         );
  INV_X1 U5434 ( .A(n4235), .ZN(n4392) );
  NAND2_X1 U5435 ( .A1(n4392), .A2(n4391), .ZN(n4606) );
  OAI211_X1 U5436 ( .C1(n4394), .C2(n3203), .A(n4393), .B(n4606), .ZN(n4395)
         );
  INV_X1 U5437 ( .A(n4395), .ZN(n4397) );
  NAND2_X1 U5438 ( .A1(n4865), .A2(n4608), .ZN(n4396) );
  NAND4_X1 U5439 ( .A1(n4399), .A2(n4398), .A3(n4397), .A4(n4396), .ZN(n4838)
         );
  MUX2_X1 U5440 ( .A(n4838), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4400) );
  INV_X1 U5441 ( .A(n4400), .ZN(n4401) );
  NAND2_X1 U5442 ( .A1(n4401), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4402) );
  INV_X1 U5443 ( .A(n4838), .ZN(n6351) );
  NAND4_X1 U5444 ( .A1(n4404), .A2(n4249), .A3(n4235), .A4(n4251), .ZN(n4405)
         );
  NOR2_X1 U5445 ( .A1(n4406), .A2(n4405), .ZN(n6344) );
  INV_X1 U5446 ( .A(n6344), .ZN(n4419) );
  INV_X1 U5447 ( .A(n6346), .ZN(n4411) );
  XNOR2_X1 U5448 ( .A(n4407), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4410)
         );
  INV_X1 U5449 ( .A(n4408), .ZN(n4841) );
  AOI211_X1 U5450 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n4841), .A(n2964), .B(n3302), .ZN(n5337) );
  OAI22_X1 U5451 ( .A1(n4411), .A2(n4410), .B1(n5337), .B2(n4424), .ZN(n4418)
         );
  INV_X1 U5452 ( .A(n4608), .ZN(n4412) );
  NAND2_X1 U5453 ( .A1(n4413), .A2(n4412), .ZN(n4427) );
  INV_X1 U5454 ( .A(n4427), .ZN(n4416) );
  MUX2_X1 U5455 ( .A(n4414), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4408), 
        .Z(n4415) );
  NOR3_X1 U5456 ( .A1(n4416), .A2(n4430), .A3(n4415), .ZN(n4417) );
  AOI211_X1 U5457 ( .C1(n2980), .C2(n4419), .A(n4418), .B(n4417), .ZN(n5338)
         );
  NAND2_X1 U5458 ( .A1(n6351), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4420) );
  OAI21_X1 U5459 ( .B1(n6351), .B2(n5338), .A(n4420), .ZN(n6360) );
  XNOR2_X1 U5460 ( .A(n4408), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4426)
         );
  XNOR2_X1 U5461 ( .A(n4856), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4422)
         );
  NAND2_X1 U5462 ( .A1(n6346), .A2(n4422), .ZN(n4423) );
  OAI21_X1 U5463 ( .B1(n4426), .B2(n4424), .A(n4423), .ZN(n4425) );
  AOI21_X1 U5464 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n4428) );
  OAI21_X1 U5465 ( .B1(n2981), .B2(n6344), .A(n4428), .ZN(n4844) );
  NOR2_X1 U5466 ( .A1(n4838), .A2(n3067), .ZN(n4429) );
  AOI21_X1 U5467 ( .B1(n4844), .B2(n4838), .A(n4429), .ZN(n6357) );
  NOR2_X1 U5468 ( .A1(n6357), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4434) );
  INV_X1 U5469 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5464) );
  NAND2_X1 U5470 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5464), .ZN(n4432) );
  INV_X1 U5471 ( .A(n4430), .ZN(n4431) );
  OAI21_X1 U5472 ( .B1(n4432), .B2(n4431), .A(n4435), .ZN(n4433) );
  AOI21_X1 U5473 ( .B1(n6360), .B2(n4434), .A(n4433), .ZN(n6366) );
  AOI21_X1 U5474 ( .B1(n4435), .B2(n4847), .A(n6366), .ZN(n4439) );
  NOR2_X1 U5475 ( .A1(n4439), .A2(FLUSH_REG_SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5476 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4437), .ZN(n6463) );
  OAI21_X1 U5477 ( .B1(n4436), .B2(n6463), .A(n6024), .ZN(n5846) );
  INV_X1 U5478 ( .A(n4437), .ZN(n4438) );
  NOR2_X1 U5479 ( .A1(n4439), .A2(n4438), .ZN(n6376) );
  NAND2_X1 U5480 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6466), .ZN(n4464) );
  INV_X1 U5481 ( .A(n4464), .ZN(n5334) );
  OAI22_X1 U5482 ( .A1(n6163), .A2(n6278), .B1(n6345), .B2(n5334), .ZN(n4440)
         );
  OAI21_X1 U5483 ( .B1(n6376), .B2(n4440), .A(n5846), .ZN(n4441) );
  OAI21_X1 U5484 ( .B1(n5846), .B2(n6347), .A(n4441), .ZN(U3465) );
  XNOR2_X1 U5485 ( .A(n4442), .B(n4443), .ZN(n4459) );
  OR2_X1 U5486 ( .A1(n4444), .A2(n3000), .ZN(n4445) );
  NAND2_X1 U5487 ( .A1(n4445), .A2(n4479), .ZN(n5578) );
  OAI211_X1 U5488 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4447), .B(n4446), .ZN(n4448) );
  INV_X1 U5489 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6418) );
  OR2_X1 U5490 ( .A1(n5845), .A2(n6418), .ZN(n4455) );
  OAI211_X1 U5491 ( .C1(n5799), .C2(n5578), .A(n4448), .B(n4455), .ZN(n4449)
         );
  AOI21_X1 U5492 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4450), .A(n4449), 
        .ZN(n4451) );
  OAI21_X1 U5493 ( .B1(n5825), .B2(n4459), .A(n4451), .ZN(U3014) );
  AOI21_X1 U5494 ( .B1(n4454), .B2(n4452), .A(n4453), .ZN(n4468) );
  INV_X1 U5495 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U5496 ( .A1(n5754), .A2(n5587), .ZN(n4456) );
  OAI211_X1 U5497 ( .C1(n5782), .C2(n5579), .A(n4456), .B(n4455), .ZN(n4457)
         );
  AOI21_X1 U5498 ( .B1(n4468), .B2(n5774), .A(n4457), .ZN(n4458) );
  OAI21_X1 U5499 ( .B1(n5766), .B2(n4459), .A(n4458), .ZN(U2982) );
  INV_X1 U5500 ( .A(n5846), .ZN(n4467) );
  INV_X1 U5501 ( .A(n4463), .ZN(n4461) );
  NOR2_X1 U5502 ( .A1(n6225), .A2(n6167), .ZN(n6232) );
  INV_X1 U5503 ( .A(n6283), .ZN(n4538) );
  NAND2_X1 U5504 ( .A1(n6232), .A2(n4538), .ZN(n6200) );
  NAND2_X1 U5505 ( .A1(n6283), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6131) );
  INV_X1 U5506 ( .A(n6131), .ZN(n4492) );
  NAND2_X1 U5507 ( .A1(n5985), .A2(n4492), .ZN(n5987) );
  NAND3_X1 U5508 ( .A1(n6200), .A2(n6132), .A3(n5987), .ZN(n4494) );
  AND2_X1 U5509 ( .A1(n6290), .A2(n6167), .ZN(n6286) );
  AOI222_X1 U5510 ( .A1(n4494), .A2(n6290), .B1(n2980), .B2(n4464), .C1(n3911), 
        .C2(n6286), .ZN(n4466) );
  NAND2_X1 U5511 ( .A1(n4467), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4465) );
  OAI21_X1 U5512 ( .B1(n4467), .B2(n4466), .A(n4465), .ZN(U3462) );
  INV_X1 U5513 ( .A(n4468), .ZN(n5589) );
  INV_X1 U5514 ( .A(n5578), .ZN(n4469) );
  AOI22_X1 U5515 ( .A1(n5066), .A2(n4469), .B1(n5065), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4470) );
  OAI21_X1 U5516 ( .B1(n5589), .B2(n5075), .A(n4470), .ZN(U2855) );
  INV_X1 U5517 ( .A(n4452), .ZN(n4471) );
  AOI21_X1 U5518 ( .B1(n4472), .B2(n4352), .A(n4471), .ZN(n4772) );
  INV_X1 U5519 ( .A(n4772), .ZN(n4615) );
  AOI22_X1 U5520 ( .A1(n5066), .A2(n4759), .B1(n5065), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4473) );
  OAI21_X1 U5521 ( .B1(n4615), .B2(n5068), .A(n4473), .ZN(U2856) );
  AOI21_X1 U5522 ( .B1(n5771), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4474), 
        .ZN(n4475) );
  OAI21_X1 U5523 ( .B1(n4760), .B2(n5777), .A(n4475), .ZN(n4476) );
  AOI21_X1 U5524 ( .B1(n4772), .B2(n5774), .A(n4476), .ZN(n4477) );
  OAI21_X1 U5525 ( .B1(n4478), .B2(n5766), .A(n4477), .ZN(U2983) );
  NAND2_X1 U5526 ( .A1(n4480), .A2(n4479), .ZN(n4482) );
  INV_X1 U5527 ( .A(n4481), .ZN(n4489) );
  NAND2_X1 U5528 ( .A1(n4482), .A2(n4489), .ZN(n5571) );
  INV_X1 U5529 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5530 ( .A1(n4453), .A2(n4484), .ZN(n4485) );
  OR2_X1 U5531 ( .A1(n4483), .A2(n4485), .ZN(n5573) );
  OAI222_X1 U5532 ( .A1(n5571), .A2(n5078), .B1(n4486), .B2(n5076), .C1(n5075), 
        .C2(n5573), .ZN(U2854) );
  OAI21_X1 U5533 ( .B1(n4483), .B2(n4488), .A(n4487), .ZN(n5565) );
  XNOR2_X1 U5534 ( .A(n4490), .B(n4489), .ZN(n5560) );
  AOI22_X1 U5535 ( .A1(n5066), .A2(n5560), .B1(n5065), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4491) );
  OAI21_X1 U5536 ( .B1(n5565), .B2(n5068), .A(n4491), .ZN(U2853) );
  NAND2_X1 U5537 ( .A1(n4492), .A2(n4460), .ZN(n4493) );
  OAI21_X1 U5538 ( .B1(n4494), .B2(n4493), .A(n6290), .ZN(n4499) );
  INV_X1 U5539 ( .A(n4495), .ZN(n5955) );
  NAND2_X1 U5540 ( .A1(n2981), .A2(n5955), .ZN(n6099) );
  NOR2_X1 U5541 ( .A1(n2980), .A2(n6099), .ZN(n5913) );
  NOR2_X1 U5542 ( .A1(n6129), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5942)
         );
  AOI21_X1 U5543 ( .B1(n5913), .B2(n6052), .A(n5942), .ZN(n4496) );
  NAND2_X1 U5544 ( .A1(n6097), .A2(n6358), .ZN(n5912) );
  OAI22_X1 U5545 ( .A1(n4499), .A2(n4496), .B1(n5912), .B2(n3391), .ZN(n5944)
         );
  INV_X1 U5546 ( .A(DATAI_7_), .ZN(n5714) );
  NOR2_X2 U5547 ( .A1(n5714), .A2(n6024), .ZN(n6335) );
  INV_X1 U5548 ( .A(n6335), .ZN(n4506) );
  INV_X1 U5549 ( .A(n4496), .ZN(n4498) );
  AOI21_X1 U5550 ( .B1(n5912), .B2(n6278), .A(n6136), .ZN(n4497) );
  OAI21_X1 U5551 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n5945) );
  INV_X1 U5552 ( .A(DATAI_23_), .ZN(n6592) );
  OR2_X1 U5553 ( .A1(n6282), .A2(n6592), .ZN(n6275) );
  NAND2_X1 U5554 ( .A1(n6283), .A2(n6163), .ZN(n6096) );
  OR3_X1 U5555 ( .A1(n3911), .A2(n3404), .A3(n6096), .ZN(n4500) );
  INV_X1 U5556 ( .A(DATAI_31_), .ZN(n4501) );
  OR2_X1 U5557 ( .A1(n6282), .A2(n4501), .ZN(n6342) );
  INV_X1 U5558 ( .A(n6342), .ZN(n6271) );
  NOR2_X1 U5559 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6466), .ZN(n4840) );
  NOR2_X2 U5560 ( .A1(n4561), .A2(n4831), .ZN(n6333) );
  AOI22_X1 U5561 ( .A1(n5943), .A2(n6271), .B1(n6333), .B2(n5942), .ZN(n4503)
         );
  OAI21_X1 U5562 ( .B1(n6275), .B2(n5954), .A(n4503), .ZN(n4504) );
  AOI21_X1 U5563 ( .B1(n5945), .B2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4504), 
        .ZN(n4505) );
  OAI21_X1 U5564 ( .B1(n4537), .B2(n4506), .A(n4505), .ZN(U3051) );
  INV_X1 U5565 ( .A(DATAI_3_), .ZN(n5707) );
  NOR2_X2 U5566 ( .A1(n5707), .A2(n6024), .ZN(n6308) );
  INV_X1 U5567 ( .A(n6308), .ZN(n4513) );
  INV_X1 U5568 ( .A(DATAI_19_), .ZN(n4507) );
  OR2_X1 U5569 ( .A1(n6282), .A2(n4507), .ZN(n6255) );
  INV_X1 U5570 ( .A(DATAI_27_), .ZN(n4508) );
  OR2_X1 U5571 ( .A1(n6282), .A2(n4508), .ZN(n6313) );
  INV_X1 U5572 ( .A(n6313), .ZN(n6252) );
  NOR2_X2 U5573 ( .A1(n4561), .A2(n4509), .ZN(n6309) );
  AOI22_X1 U5574 ( .A1(n5943), .A2(n6252), .B1(n6309), .B2(n5942), .ZN(n4510)
         );
  OAI21_X1 U5575 ( .B1(n6255), .B2(n5954), .A(n4510), .ZN(n4511) );
  AOI21_X1 U5576 ( .B1(n5945), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4511), 
        .ZN(n4512) );
  OAI21_X1 U5577 ( .B1(n4537), .B2(n4513), .A(n4512), .ZN(U3047) );
  INV_X1 U5578 ( .A(DATAI_0_), .ZN(n5701) );
  NOR2_X2 U5579 ( .A1(n5701), .A2(n6024), .ZN(n6279) );
  INV_X1 U5580 ( .A(n6279), .ZN(n4519) );
  INV_X1 U5581 ( .A(DATAI_16_), .ZN(n4514) );
  OR2_X1 U5582 ( .A1(n6282), .A2(n4514), .ZN(n6243) );
  INV_X1 U5583 ( .A(DATAI_24_), .ZN(n4515) );
  OR2_X1 U5584 ( .A1(n6282), .A2(n4515), .ZN(n6295) );
  INV_X1 U5585 ( .A(n6295), .ZN(n6240) );
  AOI22_X1 U5586 ( .A1(n5943), .A2(n6240), .B1(n6280), .B2(n5942), .ZN(n4516)
         );
  OAI21_X1 U5587 ( .B1(n6243), .B2(n5954), .A(n4516), .ZN(n4517) );
  AOI21_X1 U5588 ( .B1(n5945), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4517), 
        .ZN(n4518) );
  OAI21_X1 U5589 ( .B1(n4537), .B2(n4519), .A(n4518), .ZN(U3044) );
  INV_X1 U5590 ( .A(DATAI_5_), .ZN(n5710) );
  NOR2_X2 U5591 ( .A1(n5710), .A2(n6024), .ZN(n6320) );
  INV_X1 U5592 ( .A(n6320), .ZN(n4524) );
  INV_X1 U5593 ( .A(DATAI_21_), .ZN(n6496) );
  OR2_X1 U5594 ( .A1(n6282), .A2(n6496), .ZN(n6263) );
  INV_X1 U5595 ( .A(DATAI_29_), .ZN(n4520) );
  OR2_X1 U5596 ( .A1(n6282), .A2(n4520), .ZN(n6325) );
  INV_X1 U5597 ( .A(n6325), .ZN(n6260) );
  NOR2_X2 U5598 ( .A1(n4561), .A2(n3204), .ZN(n6321) );
  AOI22_X1 U5599 ( .A1(n5943), .A2(n6260), .B1(n6321), .B2(n5942), .ZN(n4521)
         );
  OAI21_X1 U5600 ( .B1(n6263), .B2(n5954), .A(n4521), .ZN(n4522) );
  AOI21_X1 U5601 ( .B1(n5945), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4522), 
        .ZN(n4523) );
  OAI21_X1 U5602 ( .B1(n4537), .B2(n4524), .A(n4523), .ZN(U3049) );
  INV_X1 U5603 ( .A(DATAI_4_), .ZN(n6621) );
  NOR2_X2 U5604 ( .A1(n6621), .A2(n6024), .ZN(n6314) );
  INV_X1 U5605 ( .A(n6314), .ZN(n4531) );
  INV_X1 U5606 ( .A(DATAI_20_), .ZN(n4525) );
  OR2_X1 U5607 ( .A1(n6282), .A2(n4525), .ZN(n6259) );
  INV_X1 U5608 ( .A(DATAI_28_), .ZN(n4526) );
  OR2_X1 U5609 ( .A1(n6282), .A2(n4526), .ZN(n6319) );
  INV_X1 U5610 ( .A(n6319), .ZN(n6256) );
  NOR2_X2 U5611 ( .A1(n4561), .A2(n4527), .ZN(n6315) );
  AOI22_X1 U5612 ( .A1(n5943), .A2(n6256), .B1(n6315), .B2(n5942), .ZN(n4528)
         );
  OAI21_X1 U5613 ( .B1(n6259), .B2(n5954), .A(n4528), .ZN(n4529) );
  AOI21_X1 U5614 ( .B1(n5945), .B2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n4529), 
        .ZN(n4530) );
  OAI21_X1 U5615 ( .B1(n4537), .B2(n4531), .A(n4530), .ZN(U3048) );
  INV_X1 U5616 ( .A(DATAI_1_), .ZN(n5703) );
  NOR2_X2 U5617 ( .A1(n5703), .A2(n6024), .ZN(n6296) );
  INV_X1 U5618 ( .A(n6296), .ZN(n4536) );
  INV_X1 U5619 ( .A(DATAI_17_), .ZN(n4532) );
  OR2_X1 U5620 ( .A1(n6282), .A2(n4532), .ZN(n6247) );
  INV_X1 U5621 ( .A(DATAI_25_), .ZN(n5389) );
  OR2_X1 U5622 ( .A1(n6282), .A2(n5389), .ZN(n6301) );
  INV_X1 U5623 ( .A(n6301), .ZN(n6244) );
  NOR2_X2 U5624 ( .A1(n4561), .A2(n2979), .ZN(n6297) );
  AOI22_X1 U5625 ( .A1(n5943), .A2(n6244), .B1(n6297), .B2(n5942), .ZN(n4533)
         );
  OAI21_X1 U5626 ( .B1(n6247), .B2(n5954), .A(n4533), .ZN(n4534) );
  AOI21_X1 U5627 ( .B1(n5945), .B2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4534), 
        .ZN(n4535) );
  OAI21_X1 U5628 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(U3045) );
  INV_X1 U5629 ( .A(n5954), .ZN(n4539) );
  NOR3_X1 U5630 ( .A1(n5950), .A2(n4539), .A3(n6278), .ZN(n4540) );
  NOR2_X1 U5631 ( .A1(n2981), .A2(n5955), .ZN(n6195) );
  NAND2_X1 U5632 ( .A1(n6195), .A2(n5988), .ZN(n4631) );
  OAI21_X1 U5633 ( .B1(n4540), .B2(n6286), .A(n4631), .ZN(n4542) );
  NAND2_X1 U5634 ( .A1(n6196), .A2(n6358), .ZN(n4636) );
  NOR2_X1 U5635 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4636), .ZN(n5949)
         );
  INV_X1 U5636 ( .A(n5949), .ZN(n4572) );
  NOR2_X1 U5637 ( .A1(n4543), .A2(n3391), .ZN(n6105) );
  OR2_X1 U5638 ( .A1(n6019), .A2(n6227), .ZN(n5848) );
  INV_X1 U5639 ( .A(n5848), .ZN(n4544) );
  OAI21_X1 U5640 ( .B1(n4544), .B2(n3391), .A(n5918), .ZN(n5851) );
  AOI211_X1 U5641 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4572), .A(n6105), .B(
        n5851), .ZN(n4541) );
  NAND2_X1 U5642 ( .A1(n4542), .A2(n4541), .ZN(n5951) );
  INV_X1 U5643 ( .A(n5951), .ZN(n4551) );
  INV_X1 U5644 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5645 ( .A1(n6195), .A2(n6290), .ZN(n6166) );
  OR2_X1 U5646 ( .A1(n6166), .A2(n2980), .ZN(n4546) );
  NAND2_X1 U5647 ( .A1(n4543), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6164) );
  INV_X1 U5648 ( .A(n6164), .ZN(n6228) );
  NAND2_X1 U5649 ( .A1(n4544), .A2(n6228), .ZN(n4545) );
  NAND2_X1 U5650 ( .A1(n4546), .A2(n4545), .ZN(n5948) );
  INV_X1 U5651 ( .A(n6275), .ZN(n6337) );
  AOI22_X1 U5652 ( .A1(n5950), .A2(n6337), .B1(n6333), .B2(n5949), .ZN(n4547)
         );
  OAI21_X1 U5653 ( .B1(n5954), .B2(n6342), .A(n4547), .ZN(n4548) );
  AOI21_X1 U5654 ( .B1(n6335), .B2(n5948), .A(n4548), .ZN(n4549) );
  OAI21_X1 U5655 ( .B1(n4551), .B2(n4550), .A(n4549), .ZN(U3059) );
  XNOR2_X1 U5656 ( .A(n4553), .B(n4552), .ZN(n4621) );
  NAND2_X1 U5657 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4554), .ZN(n4556)
         );
  INV_X1 U5658 ( .A(n4556), .ZN(n4555) );
  OAI21_X1 U5659 ( .B1(n5292), .B2(n4555), .A(n5822), .ZN(n4596) );
  NOR2_X1 U5660 ( .A1(n4557), .A2(n4556), .ZN(n4682) );
  AOI22_X1 U5661 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4596), .B1(n4682), 
        .B2(n6511), .ZN(n4559) );
  INV_X1 U5662 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U5663 ( .A1(n5845), .A2(n6419), .ZN(n4616) );
  AOI21_X1 U5664 ( .B1(n5836), .B2(n5560), .A(n4616), .ZN(n4558) );
  OAI211_X1 U5665 ( .C1(n4621), .C2(n5825), .A(n4559), .B(n4558), .ZN(U3012)
         );
  INV_X1 U5666 ( .A(DATAI_26_), .ZN(n4560) );
  OR2_X1 U5667 ( .A1(n6282), .A2(n4560), .ZN(n6307) );
  NAND2_X1 U5668 ( .A1(n5951), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4566) );
  INV_X1 U5669 ( .A(DATAI_18_), .ZN(n6565) );
  OR2_X1 U5670 ( .A1(n6282), .A2(n6565), .ZN(n6251) );
  INV_X1 U5671 ( .A(n6251), .ZN(n6304) );
  INV_X1 U5672 ( .A(n4561), .ZN(n4569) );
  NAND2_X1 U5673 ( .A1(n4569), .A2(n4562), .ZN(n6068) );
  INV_X1 U5674 ( .A(n5948), .ZN(n4571) );
  INV_X1 U5675 ( .A(DATAI_2_), .ZN(n5705) );
  NOR2_X2 U5676 ( .A1(n5705), .A2(n6024), .ZN(n6302) );
  INV_X1 U5677 ( .A(n6302), .ZN(n4563) );
  OAI22_X1 U5678 ( .A1(n6068), .A2(n4572), .B1(n4571), .B2(n4563), .ZN(n4564)
         );
  AOI21_X1 U5679 ( .B1(n5950), .B2(n6304), .A(n4564), .ZN(n4565) );
  OAI211_X1 U5680 ( .C1(n5954), .C2(n6307), .A(n4566), .B(n4565), .ZN(U3054)
         );
  INV_X1 U5681 ( .A(DATAI_30_), .ZN(n4567) );
  OR2_X1 U5682 ( .A1(n6282), .A2(n4567), .ZN(n6331) );
  NAND2_X1 U5683 ( .A1(n5951), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4575) );
  INV_X1 U5684 ( .A(DATAI_22_), .ZN(n4568) );
  OR2_X1 U5685 ( .A1(n6282), .A2(n4568), .ZN(n6267) );
  INV_X1 U5686 ( .A(n6267), .ZN(n6328) );
  NAND2_X1 U5687 ( .A1(n4569), .A2(n3207), .ZN(n6084) );
  INV_X1 U5688 ( .A(DATAI_6_), .ZN(n5712) );
  NOR2_X2 U5689 ( .A1(n5712), .A2(n6024), .ZN(n6326) );
  INV_X1 U5690 ( .A(n6326), .ZN(n4570) );
  OAI22_X1 U5691 ( .A1(n6084), .A2(n4572), .B1(n4571), .B2(n4570), .ZN(n4573)
         );
  AOI21_X1 U5692 ( .B1(n5950), .B2(n6328), .A(n4573), .ZN(n4574) );
  OAI211_X1 U5693 ( .C1(n5954), .C2(n6331), .A(n4575), .B(n4574), .ZN(U3058)
         );
  INV_X1 U5694 ( .A(n6263), .ZN(n6322) );
  NAND2_X1 U5695 ( .A1(n5950), .A2(n6322), .ZN(n4577) );
  AOI22_X1 U5696 ( .A1(n6321), .A2(n5949), .B1(n6320), .B2(n5948), .ZN(n4576)
         );
  OAI211_X1 U5697 ( .C1(n6325), .C2(n5954), .A(n4577), .B(n4576), .ZN(n4578)
         );
  AOI21_X1 U5698 ( .B1(n5951), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n4578), 
        .ZN(n4579) );
  INV_X1 U5699 ( .A(n4579), .ZN(U3057) );
  INV_X1 U5700 ( .A(n6243), .ZN(n6292) );
  NAND2_X1 U5701 ( .A1(n5950), .A2(n6292), .ZN(n4581) );
  AOI22_X1 U5702 ( .A1(n6280), .A2(n5949), .B1(n6279), .B2(n5948), .ZN(n4580)
         );
  OAI211_X1 U5703 ( .C1(n6295), .C2(n5954), .A(n4581), .B(n4580), .ZN(n4582)
         );
  AOI21_X1 U5704 ( .B1(n5951), .B2(INSTQUEUE_REG_4__0__SCAN_IN), .A(n4582), 
        .ZN(n4583) );
  INV_X1 U5705 ( .A(n4583), .ZN(U3052) );
  INV_X1 U5706 ( .A(n6247), .ZN(n6298) );
  NAND2_X1 U5707 ( .A1(n5950), .A2(n6298), .ZN(n4585) );
  AOI22_X1 U5708 ( .A1(n6297), .A2(n5949), .B1(n6296), .B2(n5948), .ZN(n4584)
         );
  OAI211_X1 U5709 ( .C1(n6301), .C2(n5954), .A(n4585), .B(n4584), .ZN(n4586)
         );
  AOI21_X1 U5710 ( .B1(n5951), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n4586), 
        .ZN(n4587) );
  INV_X1 U5711 ( .A(n4587), .ZN(U3053) );
  INV_X1 U5712 ( .A(n6255), .ZN(n6310) );
  NAND2_X1 U5713 ( .A1(n5950), .A2(n6310), .ZN(n4589) );
  AOI22_X1 U5714 ( .A1(n6309), .A2(n5949), .B1(n6308), .B2(n5948), .ZN(n4588)
         );
  OAI211_X1 U5715 ( .C1(n6313), .C2(n5954), .A(n4589), .B(n4588), .ZN(n4590)
         );
  AOI21_X1 U5716 ( .B1(n5951), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n4590), 
        .ZN(n4591) );
  INV_X1 U5717 ( .A(n4591), .ZN(U3055) );
  XOR2_X1 U5718 ( .A(n4593), .B(n2976), .Z(n5757) );
  NAND3_X1 U5719 ( .A1(n4594), .A2(n5819), .A3(n4599), .ZN(n4595) );
  NAND2_X1 U5720 ( .A1(n5817), .A2(REIP_REG_5__SCAN_IN), .ZN(n5758) );
  OAI211_X1 U5721 ( .C1(n5799), .C2(n5571), .A(n4595), .B(n5758), .ZN(n4601)
         );
  INV_X1 U5722 ( .A(n4596), .ZN(n4597) );
  AOI21_X1 U5723 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n4600) );
  AOI211_X1 U5724 ( .C1(n5757), .C2(n5837), .A(n4601), .B(n4600), .ZN(n4602)
         );
  INV_X1 U5725 ( .A(n4602), .ZN(U3013) );
  NAND3_X1 U5726 ( .A1(n4604), .A2(n4603), .A3(n3207), .ZN(n4605) );
  OAI22_X1 U5727 ( .A1(n4606), .A2(n6385), .B1(n4251), .B2(n4605), .ZN(n4607)
         );
  AOI21_X1 U5728 ( .B1(n4609), .B2(n4608), .A(n4607), .ZN(n4610) );
  NAND2_X2 U5729 ( .A1(n5081), .A2(n4611), .ZN(n5395) );
  INV_X1 U5730 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4613) );
  OAI222_X1 U5731 ( .A1(n5395), .A2(n5788), .B1(n4717), .B2(n5701), .C1(n5081), 
        .C2(n4613), .ZN(U2891) );
  INV_X1 U5732 ( .A(n5773), .ZN(n4614) );
  INV_X1 U5733 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5668) );
  OAI222_X1 U5734 ( .A1(n4614), .A2(n5395), .B1(n4717), .B2(n5703), .C1(n5081), 
        .C2(n5668), .ZN(U2890) );
  INV_X1 U5735 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5662) );
  OAI222_X1 U5736 ( .A1(n4615), .A2(n5395), .B1(n4717), .B2(n5707), .C1(n5081), 
        .C2(n5662), .ZN(U2888) );
  INV_X1 U5737 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6499) );
  OAI222_X1 U5738 ( .A1(n5565), .A2(n5395), .B1(n4717), .B2(n5712), .C1(n5081), 
        .C2(n6499), .ZN(U2885) );
  INV_X1 U5739 ( .A(n5565), .ZN(n4619) );
  AOI21_X1 U5740 ( .B1(n5771), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4616), 
        .ZN(n4617) );
  OAI21_X1 U5741 ( .B1(n5570), .B2(n5777), .A(n4617), .ZN(n4618) );
  AOI21_X1 U5742 ( .B1(n4619), .B2(n5774), .A(n4618), .ZN(n4620) );
  OAI21_X1 U5743 ( .B1(n5766), .B2(n4621), .A(n4620), .ZN(U2980) );
  NAND2_X1 U5744 ( .A1(n4487), .A2(n4623), .ZN(n4624) );
  AND2_X1 U5745 ( .A1(n4622), .A2(n4624), .ZN(n5749) );
  INV_X1 U5746 ( .A(n5749), .ZN(n4629) );
  AOI22_X1 U5747 ( .A1(n5102), .A2(DATAI_7_), .B1(n5636), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5748 ( .B1(n4629), .B2(n5395), .A(n4625), .ZN(U2884) );
  XNOR2_X1 U5749 ( .A(n4627), .B(n4626), .ZN(n5553) );
  INV_X1 U5750 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4628) );
  OAI222_X1 U5751 ( .A1(n4629), .A2(n5075), .B1(n5078), .B2(n5553), .C1(n5076), 
        .C2(n4628), .ZN(U2852) );
  INV_X1 U5752 ( .A(n4639), .ZN(n4630) );
  OAI21_X1 U5753 ( .B1(n4630), .B2(n6167), .A(n6290), .ZN(n4638) );
  OR2_X1 U5754 ( .A1(n4631), .A2(n6345), .ZN(n4633) );
  NOR2_X1 U5755 ( .A1(n6347), .A2(n4636), .ZN(n4668) );
  INV_X1 U5756 ( .A(n4668), .ZN(n4632) );
  NAND2_X1 U5757 ( .A1(n4633), .A2(n4632), .ZN(n4635) );
  NOR2_X1 U5758 ( .A1(n4638), .A2(n4635), .ZN(n4634) );
  AOI211_X2 U5759 ( .C1(n6278), .C2(n4636), .A(n6136), .B(n4634), .ZN(n4674)
         );
  INV_X1 U5760 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4643) );
  INV_X1 U5761 ( .A(n4635), .ZN(n4637) );
  OAI22_X1 U5762 ( .A1(n4638), .A2(n4637), .B1(n3391), .B2(n4636), .ZN(n4671)
         );
  INV_X1 U5763 ( .A(n6307), .ZN(n6248) );
  AOI22_X1 U5764 ( .A1(n5950), .A2(n6248), .B1(n6303), .B2(n4668), .ZN(n4640)
         );
  OAI21_X1 U5765 ( .B1(n6251), .B2(n5963), .A(n4640), .ZN(n4641) );
  AOI21_X1 U5766 ( .B1(n4671), .B2(n6302), .A(n4641), .ZN(n4642) );
  OAI21_X1 U5767 ( .B1(n4674), .B2(n4643), .A(n4642), .ZN(U3062) );
  INV_X1 U5768 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5769 ( .A1(n5950), .A2(n6256), .B1(n6315), .B2(n4668), .ZN(n4644)
         );
  OAI21_X1 U5770 ( .B1(n6259), .B2(n5963), .A(n4644), .ZN(n4645) );
  AOI21_X1 U5771 ( .B1(n4671), .B2(n6314), .A(n4645), .ZN(n4646) );
  OAI21_X1 U5772 ( .B1(n4674), .B2(n4647), .A(n4646), .ZN(U3064) );
  INV_X1 U5773 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4651) );
  AOI22_X1 U5774 ( .A1(n5950), .A2(n6240), .B1(n6280), .B2(n4668), .ZN(n4648)
         );
  OAI21_X1 U5775 ( .B1(n6243), .B2(n5963), .A(n4648), .ZN(n4649) );
  AOI21_X1 U5776 ( .B1(n4671), .B2(n6279), .A(n4649), .ZN(n4650) );
  OAI21_X1 U5777 ( .B1(n4674), .B2(n4651), .A(n4650), .ZN(U3060) );
  INV_X1 U5778 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5779 ( .A1(n5950), .A2(n6260), .B1(n6321), .B2(n4668), .ZN(n4652)
         );
  OAI21_X1 U5780 ( .B1(n6263), .B2(n5963), .A(n4652), .ZN(n4653) );
  AOI21_X1 U5781 ( .B1(n4671), .B2(n6320), .A(n4653), .ZN(n4654) );
  OAI21_X1 U5782 ( .B1(n4674), .B2(n4655), .A(n4654), .ZN(U3065) );
  INV_X1 U5783 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5784 ( .A1(n5950), .A2(n6244), .B1(n6297), .B2(n4668), .ZN(n4656)
         );
  OAI21_X1 U5785 ( .B1(n6247), .B2(n5963), .A(n4656), .ZN(n4657) );
  AOI21_X1 U5786 ( .B1(n4671), .B2(n6296), .A(n4657), .ZN(n4658) );
  OAI21_X1 U5787 ( .B1(n4674), .B2(n4659), .A(n4658), .ZN(U3061) );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5789 ( .A1(n5950), .A2(n6271), .B1(n6333), .B2(n4668), .ZN(n4660)
         );
  OAI21_X1 U5790 ( .B1(n6275), .B2(n5963), .A(n4660), .ZN(n4661) );
  AOI21_X1 U5791 ( .B1(n4671), .B2(n6335), .A(n4661), .ZN(n4662) );
  OAI21_X1 U5792 ( .B1(n4674), .B2(n4663), .A(n4662), .ZN(U3067) );
  INV_X1 U5793 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4667) );
  INV_X1 U5794 ( .A(n6331), .ZN(n6264) );
  AOI22_X1 U5795 ( .A1(n5950), .A2(n6264), .B1(n6327), .B2(n4668), .ZN(n4664)
         );
  OAI21_X1 U5796 ( .B1(n6267), .B2(n5963), .A(n4664), .ZN(n4665) );
  AOI21_X1 U5797 ( .B1(n4671), .B2(n6326), .A(n4665), .ZN(n4666) );
  OAI21_X1 U5798 ( .B1(n4674), .B2(n4667), .A(n4666), .ZN(U3066) );
  INV_X1 U5799 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5800 ( .A1(n5950), .A2(n6252), .B1(n6309), .B2(n4668), .ZN(n4669)
         );
  OAI21_X1 U5801 ( .B1(n6255), .B2(n5963), .A(n4669), .ZN(n4670) );
  AOI21_X1 U5802 ( .B1(n4671), .B2(n6308), .A(n4670), .ZN(n4672) );
  OAI21_X1 U5803 ( .B1(n4674), .B2(n4673), .A(n4672), .ZN(U3063) );
  XNOR2_X1 U5804 ( .A(n4675), .B(n2974), .ZN(n4708) );
  OAI22_X1 U5805 ( .A1(n5291), .A2(n4678), .B1(n4787), .B2(n4677), .ZN(n5796)
         );
  OR2_X1 U5806 ( .A1(n4680), .A2(n4679), .ZN(n4681) );
  NAND2_X1 U5807 ( .A1(n4681), .A2(n4713), .ZN(n5542) );
  NAND2_X1 U5808 ( .A1(n5817), .A2(REIP_REG_8__SCAN_IN), .ZN(n4705) );
  OAI21_X1 U5809 ( .B1(n5799), .B2(n5542), .A(n4705), .ZN(n4685) );
  NAND2_X1 U5810 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4682), .ZN(n5802)
         );
  OAI21_X1 U5811 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5803), .ZN(n4683) );
  NOR2_X1 U5812 ( .A1(n5802), .A2(n4683), .ZN(n4684) );
  AOI211_X1 U5813 ( .C1(n5796), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4685), 
        .B(n4684), .ZN(n4686) );
  OAI21_X1 U5814 ( .B1(n4708), .B2(n5825), .A(n4686), .ZN(U3010) );
  XOR2_X1 U5815 ( .A(n4687), .B(n4688), .Z(n5750) );
  INV_X1 U5816 ( .A(n5750), .ZN(n4692) );
  NAND2_X1 U5817 ( .A1(n5817), .A2(REIP_REG_7__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U5818 ( .B1(n5799), .B2(n5553), .A(n5751), .ZN(n4690) );
  NOR2_X1 U5819 ( .A1(n5802), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4689)
         );
  AOI211_X1 U5820 ( .C1(n5796), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4690), 
        .B(n4689), .ZN(n4691) );
  OAI21_X1 U5821 ( .B1(n4692), .B2(n5825), .A(n4691), .ZN(U3011) );
  NOR2_X1 U5822 ( .A1(n4694), .A2(n4695), .ZN(n4696) );
  OR2_X1 U5823 ( .A1(n4693), .A2(n4696), .ZN(n5536) );
  AOI22_X1 U5824 ( .A1(n5102), .A2(DATAI_9_), .B1(n5636), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4697) );
  OAI21_X1 U5825 ( .B1(n5536), .B2(n5395), .A(n4697), .ZN(U2882) );
  XOR2_X1 U5826 ( .A(n4622), .B(n4698), .Z(n5546) );
  OAI22_X1 U5827 ( .A1(n5078), .A2(n5542), .B1(n4699), .B2(n5076), .ZN(n4700)
         );
  AOI21_X1 U5828 ( .B1(n5546), .B2(n4807), .A(n4700), .ZN(n4701) );
  INV_X1 U5829 ( .A(n4701), .ZN(U2851) );
  INV_X1 U5830 ( .A(n5546), .ZN(n4703) );
  AOI22_X1 U5831 ( .A1(n5102), .A2(DATAI_8_), .B1(n5636), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4702) );
  OAI21_X1 U5832 ( .B1(n4703), .B2(n5395), .A(n4702), .ZN(U2883) );
  NAND2_X1 U5833 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4704)
         );
  OAI211_X1 U5834 ( .C1(n5777), .C2(n5544), .A(n4705), .B(n4704), .ZN(n4706)
         );
  AOI21_X1 U5835 ( .B1(n5546), .B2(n5774), .A(n4706), .ZN(n4707) );
  OAI21_X1 U5836 ( .B1(n4708), .B2(n5766), .A(n4707), .ZN(U2978) );
  OR2_X1 U5837 ( .A1(n4693), .A2(n4710), .ZN(n4711) );
  NAND2_X1 U5838 ( .A1(n4709), .A2(n4711), .ZN(n4983) );
  AOI22_X1 U5839 ( .A1(n5102), .A2(DATAI_10_), .B1(n5636), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4712) );
  OAI21_X1 U5840 ( .B1(n4983), .B2(n5395), .A(n4712), .ZN(U2881) );
  AOI21_X1 U5841 ( .B1(n4714), .B2(n4713), .A(n2998), .ZN(n5810) );
  INV_X1 U5842 ( .A(n5810), .ZN(n4716) );
  OAI222_X1 U5843 ( .A1(n4716), .A2(n5078), .B1(n4715), .B2(n5076), .C1(n5075), 
        .C2(n5536), .ZN(U2850) );
  INV_X1 U5844 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5660) );
  OAI222_X1 U5845 ( .A1(n5589), .A2(n5395), .B1(n4717), .B2(n6621), .C1(n5660), 
        .C2(n5081), .ZN(U2887) );
  INV_X1 U5846 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5658) );
  OAI222_X1 U5847 ( .A1(n5573), .A2(n5395), .B1(n4717), .B2(n5710), .C1(n5081), 
        .C2(n5658), .ZN(U2886) );
  INV_X1 U5848 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5665) );
  OAI222_X1 U5849 ( .A1(n5765), .A2(n5395), .B1(n4717), .B2(n5705), .C1(n5081), 
        .C2(n5665), .ZN(U2889) );
  XNOR2_X1 U5850 ( .A(n5414), .B(n5815), .ZN(n4718) );
  XNOR2_X1 U5851 ( .A(n4719), .B(n4718), .ZN(n5812) );
  NAND2_X1 U5852 ( .A1(n5812), .A2(n5785), .ZN(n4722) );
  NAND2_X1 U5853 ( .A1(n5817), .A2(REIP_REG_9__SCAN_IN), .ZN(n5808) );
  OAI21_X1 U5854 ( .B1(n5782), .B2(n5534), .A(n5808), .ZN(n4720) );
  AOI21_X1 U5855 ( .B1(n5754), .B2(n5532), .A(n4720), .ZN(n4721) );
  OAI211_X1 U5856 ( .C1(n6282), .C2(n5536), .A(n4722), .B(n4721), .ZN(U2977)
         );
  OAI21_X1 U5857 ( .B1(n4723), .B2(n2998), .A(n4736), .ZN(n5798) );
  OAI222_X1 U5858 ( .A1(n5798), .A2(n5078), .B1(n5076), .B2(n4121), .C1(n5075), 
        .C2(n4983), .ZN(U2849) );
  INV_X1 U5859 ( .A(n4725), .ZN(n4727) );
  NOR2_X1 U5860 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  XNOR2_X1 U5861 ( .A(n4724), .B(n4728), .ZN(n5801) );
  NAND2_X1 U5862 ( .A1(n5801), .A2(n5785), .ZN(n4732) );
  INV_X1 U5863 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4729) );
  OAI22_X1 U5864 ( .A1(n5782), .A2(n6572), .B1(n5845), .B2(n4729), .ZN(n4730)
         );
  AOI21_X1 U5865 ( .B1(n5754), .B2(n4992), .A(n4730), .ZN(n4731) );
  OAI211_X1 U5866 ( .C1(n6282), .C2(n4983), .A(n4732), .B(n4731), .ZN(U2976)
         );
  INV_X1 U5867 ( .A(n4733), .ZN(n4734) );
  AOI21_X1 U5868 ( .B1(n4735), .B2(n4709), .A(n4734), .ZN(n5744) );
  INV_X1 U5869 ( .A(n5744), .ZN(n4740) );
  AOI21_X1 U5870 ( .B1(n4737), .B2(n4736), .A(n4774), .ZN(n5789) );
  AOI22_X1 U5871 ( .A1(n5066), .A2(n5789), .B1(n5065), .B2(EBX_REG_11__SCAN_IN), .ZN(n4738) );
  OAI21_X1 U5872 ( .B1(n4740), .B2(n5068), .A(n4738), .ZN(U2848) );
  AOI22_X1 U5873 ( .A1(n5102), .A2(DATAI_11_), .B1(n5636), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4739) );
  OAI21_X1 U5874 ( .B1(n4740), .B2(n5395), .A(n4739), .ZN(U2880) );
  XOR2_X1 U5875 ( .A(n4741), .B(n4733), .Z(n4784) );
  AOI22_X1 U5876 ( .A1(n5102), .A2(DATAI_12_), .B1(n5636), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U5877 ( .B1(n5518), .B2(n5395), .A(n4742), .ZN(U2879) );
  OR2_X1 U5878 ( .A1(n3976), .A2(n4743), .ZN(n4744) );
  NAND2_X1 U5879 ( .A1(n5564), .A2(n4744), .ZN(n5622) );
  INV_X1 U5880 ( .A(n5622), .ZN(n5596) );
  AND2_X1 U5881 ( .A1(n4745), .A2(n4751), .ZN(n5598) );
  INV_X1 U5882 ( .A(n5598), .ZN(n5614) );
  OR2_X1 U5883 ( .A1(n4746), .A2(EBX_REG_31__SCAN_IN), .ZN(n4747) );
  OR2_X1 U5884 ( .A1(n4748), .A2(n4747), .ZN(n4749) );
  NAND2_X1 U5885 ( .A1(n4750), .A2(n4749), .ZN(n4752) );
  AND2_X2 U5886 ( .A1(n4752), .A2(n4751), .ZN(n5610) );
  AOI22_X1 U5887 ( .A1(n5835), .A2(n5595), .B1(n5610), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4753) );
  OAI21_X1 U5888 ( .B1(n6345), .B2(n5614), .A(n4753), .ZN(n4754) );
  AOI21_X1 U5889 ( .B1(n4986), .B2(REIP_REG_0__SCAN_IN), .A(n4754), .ZN(n4758)
         );
  OAI21_X1 U5890 ( .B1(n5613), .B2(n5612), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4757) );
  OAI211_X1 U5891 ( .C1(n5788), .C2(n5596), .A(n4758), .B(n4757), .ZN(U2827)
         );
  AOI22_X1 U5892 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n5598), 
        .B2(n2980), .ZN(n4770) );
  AOI22_X1 U5893 ( .A1(n4759), .A2(n5595), .B1(n5610), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4769) );
  INV_X1 U5894 ( .A(n4760), .ZN(n4761) );
  NAND2_X1 U5895 ( .A1(n5612), .A2(n4761), .ZN(n4768) );
  OR2_X1 U5896 ( .A1(n5597), .A2(REIP_REG_1__SCAN_IN), .ZN(n5608) );
  AND2_X1 U5897 ( .A1(n5608), .A2(REIP_REG_2__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U5898 ( .A1(n2956), .A2(n4762), .ZN(n5600) );
  NAND2_X1 U5899 ( .A1(n5600), .A2(n4763), .ZN(n4766) );
  INV_X1 U5900 ( .A(n4990), .ZN(n4764) );
  OR2_X1 U5901 ( .A1(n5597), .A2(n4764), .ZN(n4765) );
  NAND2_X1 U5902 ( .A1(n2956), .A2(n4765), .ZN(n5582) );
  NAND2_X1 U5903 ( .A1(n4766), .A2(n5582), .ZN(n4767) );
  NAND4_X1 U5904 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4771)
         );
  AOI21_X1 U5905 ( .B1(n4772), .B2(n5622), .A(n4771), .ZN(n4773) );
  INV_X1 U5906 ( .A(n4773), .ZN(U2824) );
  OAI21_X1 U5907 ( .B1(n4775), .B2(n4774), .A(n4803), .ZN(n5523) );
  OAI222_X1 U5908 ( .A1(n5523), .A2(n5078), .B1(n5076), .B2(n5514), .C1(n5075), 
        .C2(n5518), .ZN(U2847) );
  INV_X1 U5909 ( .A(n4776), .ZN(n4777) );
  NOR2_X1 U5910 ( .A1(n4778), .A2(n4777), .ZN(n4779) );
  XNOR2_X1 U5911 ( .A(n4780), .B(n4779), .ZN(n4796) );
  NAND2_X1 U5912 ( .A1(n5754), .A2(n5520), .ZN(n4781) );
  NAND2_X1 U5913 ( .A1(n5817), .A2(REIP_REG_12__SCAN_IN), .ZN(n4791) );
  OAI211_X1 U5914 ( .C1(n5782), .C2(n4782), .A(n4781), .B(n4791), .ZN(n4783)
         );
  AOI21_X1 U5915 ( .B1(n4784), .B2(n5774), .A(n4783), .ZN(n4785) );
  OAI21_X1 U5916 ( .B1(n4796), .B2(n5766), .A(n4785), .ZN(U2974) );
  OAI22_X1 U5917 ( .A1(n5291), .A2(n5319), .B1(n4787), .B2(n4786), .ZN(n5792)
         );
  INV_X1 U5918 ( .A(n5792), .ZN(n4788) );
  OAI221_X1 U5919 ( .B1(n4813), .B2(n4790), .C1(n4813), .C2(n4789), .A(n4788), 
        .ZN(n4794) );
  OAI21_X1 U5920 ( .B1(n5325), .B2(n5790), .A(n4128), .ZN(n4793) );
  OAI21_X1 U5921 ( .B1(n5799), .B2(n5523), .A(n4791), .ZN(n4792) );
  AOI21_X1 U5922 ( .B1(n4794), .B2(n4793), .A(n4792), .ZN(n4795) );
  OAI21_X1 U5923 ( .B1(n4796), .B2(n5825), .A(n4795), .ZN(U3006) );
  NAND2_X1 U5924 ( .A1(n4799), .A2(n4798), .ZN(n4800) );
  INV_X1 U5925 ( .A(n5507), .ZN(n4802) );
  AOI22_X1 U5926 ( .A1(n5102), .A2(DATAI_13_), .B1(n5636), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4801) );
  OAI21_X1 U5927 ( .B1(n4802), .B2(n5395), .A(n4801), .ZN(U2878) );
  XNOR2_X1 U5928 ( .A(n4804), .B(n4803), .ZN(n5505) );
  OAI22_X1 U5929 ( .A1(n5078), .A2(n5505), .B1(n4805), .B2(n5076), .ZN(n4806)
         );
  AOI21_X1 U5930 ( .B1(n5507), .B2(n4807), .A(n4806), .ZN(n4808) );
  INV_X1 U5931 ( .A(n4808), .ZN(U2846) );
  NOR2_X1 U5932 ( .A1(n5839), .A2(n4813), .ZN(n4809) );
  AOI211_X1 U5933 ( .C1(n5841), .C2(n5324), .A(n4809), .B(n5792), .ZN(n5323)
         );
  OAI21_X1 U5934 ( .B1(n4812), .B2(n4811), .A(n4810), .ZN(n5422) );
  NAND2_X1 U5935 ( .A1(n5422), .A2(n5837), .ZN(n4817) );
  AND2_X1 U5936 ( .A1(n5318), .A2(n4813), .ZN(n4815) );
  NAND2_X1 U5937 ( .A1(n5817), .A2(REIP_REG_13__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U5938 ( .B1(n5799), .B2(n5505), .A(n5423), .ZN(n4814) );
  AOI21_X1 U5939 ( .B1(n5791), .B2(n4815), .A(n4814), .ZN(n4816) );
  OAI211_X1 U5940 ( .C1(n5323), .C2(n5318), .A(n4817), .B(n4816), .ZN(U3005)
         );
  OAI21_X1 U5941 ( .B1(n4818), .B2(n4820), .A(n4819), .ZN(n5204) );
  AOI22_X1 U5942 ( .A1(n5102), .A2(DATAI_15_), .B1(n5636), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4821) );
  OAI21_X1 U5943 ( .B1(n5204), .B2(n5395), .A(n4821), .ZN(U2876) );
  AOI21_X1 U5944 ( .B1(n4822), .B2(n5069), .A(n2990), .ZN(n5447) );
  INV_X1 U5945 ( .A(n5447), .ZN(n4823) );
  INV_X1 U5946 ( .A(n5610), .ZN(n5584) );
  OAI22_X1 U5947 ( .A1(n4823), .A2(n5625), .B1(n5584), .B2(n4086), .ZN(n4828)
         );
  INV_X1 U5948 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6430) );
  AOI22_X1 U5949 ( .A1(REIP_REG_15__SCAN_IN), .A2(n4972), .B1(n4974), .B2(
        n6430), .ZN(n4825) );
  NAND2_X1 U5950 ( .A1(n4824), .A2(n2956), .ZN(n5561) );
  OAI211_X1 U5951 ( .C1(n5603), .C2(n4826), .A(n4825), .B(n5561), .ZN(n4827)
         );
  AOI211_X1 U5952 ( .C1(n5612), .C2(n5199), .A(n4828), .B(n4827), .ZN(n4829)
         );
  OAI21_X1 U5953 ( .B1(n5204), .B2(n5564), .A(n4829), .ZN(U2812) );
  AOI22_X1 U5954 ( .A1(n5066), .A2(n5447), .B1(n5065), .B2(EBX_REG_15__SCAN_IN), .ZN(n4830) );
  OAI21_X1 U5955 ( .B1(n5204), .B2(n5068), .A(n4830), .ZN(U2844) );
  NAND2_X1 U5956 ( .A1(n4833), .A2(n4832), .ZN(n4836) );
  AOI22_X1 U5957 ( .A1(n5633), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5636), .ZN(n4835) );
  NAND2_X1 U5958 ( .A1(n4836), .A2(n4835), .ZN(U2860) );
  INV_X1 U5959 ( .A(n6379), .ZN(n4850) );
  INV_X1 U5960 ( .A(n6463), .ZN(n4837) );
  AOI22_X1 U5961 ( .A1(n4839), .A2(n4838), .B1(FLUSH_REG_SCAN_IN), .B2(n4837), 
        .ZN(n5456) );
  INV_X1 U5962 ( .A(n4840), .ZN(n6464) );
  NAND2_X1 U5963 ( .A1(n5456), .A2(n6464), .ZN(n6472) );
  INV_X1 U5964 ( .A(n6472), .ZN(n4858) );
  AOI21_X1 U5965 ( .B1(n4850), .B2(n4841), .A(n4858), .ZN(n4846) );
  INV_X1 U5966 ( .A(n6474), .ZN(n4854) );
  INV_X1 U5967 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5821) );
  AOI22_X1 U5968 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4047), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5821), .ZN(n4853) );
  NOR3_X1 U5969 ( .A1(n6468), .A2(n5780), .A3(n4853), .ZN(n4843) );
  NOR3_X1 U5970 ( .A1(n6379), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4841), 
        .ZN(n4842) );
  AOI211_X1 U5971 ( .C1(n4844), .C2(n4854), .A(n4843), .B(n4842), .ZN(n4845)
         );
  OAI22_X1 U5972 ( .A1(n4846), .A2(n3067), .B1(n4845), .B2(n4858), .ZN(U3459)
         );
  NOR3_X1 U5973 ( .A1(n6343), .A2(n4408), .A3(n4847), .ZN(n4848) );
  AOI21_X1 U5974 ( .B1(n6346), .B2(n4856), .A(n4848), .ZN(n4849) );
  OAI21_X1 U5975 ( .B1(n4495), .B2(n6344), .A(n4849), .ZN(n6349) );
  NOR2_X1 U5976 ( .A1(n6468), .A2(n5780), .ZN(n4852) );
  AOI222_X1 U5977 ( .A1(n6349), .A2(n4854), .B1(n4853), .B2(n4852), .C1(n4851), 
        .C2(n4850), .ZN(n4857) );
  OAI21_X1 U5978 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6379), .A(n6472), 
        .ZN(n6470) );
  INV_X1 U5979 ( .A(n6470), .ZN(n4855) );
  OAI22_X1 U5980 ( .A1(n4858), .A2(n4857), .B1(n4856), .B2(n4855), .ZN(U3460)
         );
  AND2_X1 U5981 ( .A1(n4070), .A2(n4859), .ZN(n4864) );
  NAND2_X1 U5982 ( .A1(n4860), .A2(n4865), .ZN(n4863) );
  NAND2_X1 U5983 ( .A1(n4867), .A2(n4861), .ZN(n4862) );
  OAI211_X1 U5984 ( .C1(n4864), .C2(n4865), .A(n4863), .B(n4862), .ZN(n6364)
         );
  OR2_X1 U5985 ( .A1(n4865), .A2(n3205), .ZN(n4870) );
  NAND2_X1 U5986 ( .A1(n4867), .A2(n4866), .ZN(n4868) );
  NAND2_X1 U5987 ( .A1(n4868), .A2(n4070), .ZN(n4869) );
  NAND2_X1 U5988 ( .A1(n4870), .A2(n4869), .ZN(n5458) );
  AOI21_X1 U5989 ( .B1(n4871), .B2(n6398), .A(READY_N), .ZN(n6487) );
  NOR2_X1 U5990 ( .A1(n5458), .A2(n6487), .ZN(n6361) );
  OR2_X1 U5991 ( .A1(n6361), .A2(n6385), .ZN(n5463) );
  MUX2_X1 U5992 ( .A(n6364), .B(MORE_REG_SCAN_IN), .S(n5463), .Z(U3471) );
  INV_X1 U5993 ( .A(n4877), .ZN(n4873) );
  INV_X1 U5994 ( .A(n4875), .ZN(n4872) );
  OAI21_X1 U5995 ( .B1(n4874), .B2(n4873), .A(n4872), .ZN(n4879) );
  OAI211_X1 U5996 ( .C1(n4877), .C2(n4111), .A(n4876), .B(n4875), .ZN(n4878)
         );
  OAI21_X1 U5997 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n5212) );
  INV_X1 U5998 ( .A(n4881), .ZN(n4884) );
  INV_X1 U5999 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5000) );
  OAI22_X1 U6000 ( .A1(n5603), .A2(n4882), .B1(n5000), .B2(n5584), .ZN(n4883)
         );
  AOI21_X1 U6001 ( .B1(n4884), .B2(n5612), .A(n4883), .ZN(n4885) );
  OAI21_X1 U6002 ( .B1(n5212), .B2(n5625), .A(n4885), .ZN(n4886) );
  AOI211_X1 U6003 ( .C1(n4888), .C2(REIP_REG_30__SCAN_IN), .A(n4887), .B(n4886), .ZN(n4889) );
  OAI21_X1 U6004 ( .B1(n5084), .B2(n5564), .A(n4889), .ZN(U2797) );
  INV_X1 U6005 ( .A(n5110), .ZN(n5087) );
  INV_X1 U6006 ( .A(n4892), .ZN(n4909) );
  INV_X1 U6007 ( .A(n5001), .ZN(n4897) );
  OAI22_X1 U6008 ( .A1(n5603), .A2(n5108), .B1(n5584), .B2(n4893), .ZN(n4894)
         );
  AOI21_X1 U6009 ( .B1(n5105), .B2(n5612), .A(n4894), .ZN(n4895) );
  OAI211_X1 U6010 ( .C1(n4897), .C2(n5625), .A(n4896), .B(n4895), .ZN(n4898)
         );
  AOI21_X1 U6011 ( .B1(n4909), .B2(REIP_REG_29__SCAN_IN), .A(n4898), .ZN(n4899) );
  OAI21_X1 U6012 ( .B1(n5087), .B2(n5564), .A(n4899), .ZN(U2798) );
  INV_X1 U6013 ( .A(n4900), .ZN(n4907) );
  AOI22_X1 U6014 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .B1(n5610), 
        .B2(EBX_REG_28__SCAN_IN), .ZN(n4906) );
  INV_X1 U6015 ( .A(n4901), .ZN(n4902) );
  XNOR2_X1 U6016 ( .A(n4916), .B(n4902), .ZN(n5222) );
  INV_X1 U6017 ( .A(n4903), .ZN(n4904) );
  AOI22_X1 U6018 ( .A1(n5222), .A2(n5595), .B1(n4904), .B2(n5612), .ZN(n4905)
         );
  OAI211_X1 U6019 ( .C1(n4907), .C2(REIP_REG_28__SCAN_IN), .A(n4906), .B(n4905), .ZN(n4908) );
  AOI21_X1 U6020 ( .B1(n4909), .B2(REIP_REG_28__SCAN_IN), .A(n4908), .ZN(n4910) );
  OAI21_X1 U6021 ( .B1(n5090), .B2(n5564), .A(n4910), .ZN(U2799) );
  AOI21_X1 U6022 ( .B1(n4912), .B2(n4911), .A(n4064), .ZN(n5118) );
  INV_X1 U6023 ( .A(n5118), .ZN(n5093) );
  NOR3_X1 U6024 ( .A1(n4940), .A2(REIP_REG_27__SCAN_IN), .A3(n4913), .ZN(n4920) );
  AND2_X1 U6025 ( .A1(n2987), .A2(n4914), .ZN(n4915) );
  NOR2_X1 U6026 ( .A1(n4916), .A2(n4915), .ZN(n5234) );
  AOI22_X1 U6027 ( .A1(n5234), .A2(n5595), .B1(n5610), .B2(EBX_REG_27__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6028 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4917)
         );
  OAI211_X1 U6029 ( .C1(n5607), .C2(n5116), .A(n4918), .B(n4917), .ZN(n4919)
         );
  AOI211_X1 U6030 ( .C1(n4934), .C2(REIP_REG_27__SCAN_IN), .A(n4920), .B(n4919), .ZN(n4921) );
  OAI21_X1 U6031 ( .B1(n5093), .B2(n5564), .A(n4921), .ZN(U2800) );
  OAI21_X1 U6032 ( .B1(n4922), .B2(n4923), .A(n4911), .ZN(n5129) );
  INV_X1 U6033 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4924) );
  NOR2_X1 U6034 ( .A1(n4924), .A2(n4940), .ZN(n5340) );
  NAND2_X1 U6035 ( .A1(n5340), .A2(REIP_REG_25__SCAN_IN), .ZN(n4925) );
  INV_X1 U6036 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6037 ( .A1(n4925), .A2(n5120), .ZN(n4933) );
  NAND2_X1 U6038 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4931)
         );
  INV_X1 U6039 ( .A(n5121), .ZN(n4926) );
  NAND2_X1 U6040 ( .A1(n5612), .A2(n4926), .ZN(n4930) );
  NAND2_X1 U6041 ( .A1(n2992), .A2(n4927), .ZN(n4928) );
  AND2_X1 U6042 ( .A1(n2987), .A2(n4928), .ZN(n5246) );
  AOI22_X1 U6043 ( .A1(n5246), .A2(n5595), .B1(n5610), .B2(EBX_REG_26__SCAN_IN), .ZN(n4929) );
  NAND3_X1 U6044 ( .A1(n4931), .A2(n4930), .A3(n4929), .ZN(n4932) );
  AOI21_X1 U6045 ( .B1(n4934), .B2(n4933), .A(n4932), .ZN(n4935) );
  OAI21_X1 U6046 ( .B1(n5129), .B2(n5564), .A(n4935), .ZN(U2801) );
  NOR2_X1 U6047 ( .A1(n4937), .A2(n4938), .ZN(n4939) );
  OR2_X1 U6048 ( .A1(n4936), .A2(n4939), .ZN(n5146) );
  NOR2_X1 U6049 ( .A1(REIP_REG_24__SCAN_IN), .A2(n4940), .ZN(n5344) );
  INV_X1 U6050 ( .A(n5344), .ZN(n4945) );
  INV_X1 U6051 ( .A(n5008), .ZN(n4941) );
  XNOR2_X1 U6052 ( .A(n5009), .B(n4941), .ZN(n5258) );
  AOI22_X1 U6053 ( .A1(n5258), .A2(n5595), .B1(EBX_REG_24__SCAN_IN), .B2(n5610), .ZN(n4942) );
  OAI21_X1 U6054 ( .B1(n5603), .B2(n5145), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6055 ( .B1(n5149), .B2(n5612), .A(n4943), .ZN(n4944) );
  NAND2_X1 U6056 ( .A1(n4945), .A2(n4944), .ZN(n4946) );
  AOI21_X1 U6057 ( .B1(n5343), .B2(REIP_REG_24__SCAN_IN), .A(n4946), .ZN(n4947) );
  OAI21_X1 U6058 ( .B1(n5146), .B2(n5564), .A(n4947), .ZN(U2803) );
  AND2_X1 U6059 ( .A1(n4948), .A2(n4949), .ZN(n4950) );
  OR2_X1 U6060 ( .A1(n4950), .A2(n4937), .ZN(n5158) );
  OAI22_X1 U6061 ( .A1(n4951), .A2(n5584), .B1(n5157), .B2(n5603), .ZN(n4955)
         );
  NOR2_X1 U6062 ( .A1(n5019), .A2(n4952), .ZN(n4953) );
  OR2_X1 U6063 ( .A1(n5009), .A2(n4953), .ZN(n5262) );
  NOR2_X1 U6064 ( .A1(n5262), .A2(n5625), .ZN(n4954) );
  AOI211_X1 U6065 ( .C1(n5612), .C2(n5161), .A(n4955), .B(n4954), .ZN(n4958)
         );
  NAND2_X1 U6066 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5356), .ZN(n5349) );
  OAI21_X1 U6067 ( .B1(n6440), .B2(n5349), .A(n6442), .ZN(n4956) );
  NAND2_X1 U6068 ( .A1(n5343), .A2(n4956), .ZN(n4957) );
  OAI211_X1 U6069 ( .C1(n5158), .C2(n5564), .A(n4958), .B(n4957), .ZN(U2804)
         );
  XOR2_X1 U6070 ( .A(n4960), .B(n4959), .Z(n5630) );
  INV_X1 U6071 ( .A(n5630), .ZN(n5064) );
  AOI21_X1 U6072 ( .B1(n6432), .B2(n4961), .A(n5480), .ZN(n4968) );
  OAI21_X1 U6073 ( .B1(n5603), .B2(n3616), .A(n5561), .ZN(n4967) );
  INV_X1 U6074 ( .A(n5418), .ZN(n4965) );
  INV_X1 U6075 ( .A(n5055), .ZN(n5050) );
  AOI21_X1 U6076 ( .B1(n4963), .B2(n4962), .A(n5050), .ZN(n5441) );
  AOI22_X1 U6077 ( .A1(n5441), .A2(n5595), .B1(n5610), .B2(EBX_REG_17__SCAN_IN), .ZN(n4964) );
  OAI21_X1 U6078 ( .B1(n5607), .B2(n4965), .A(n4964), .ZN(n4966) );
  NOR3_X1 U6079 ( .A1(n4968), .A2(n4967), .A3(n4966), .ZN(n4969) );
  OAI21_X1 U6080 ( .B1(n5064), .B2(n5564), .A(n4969), .ZN(U2810) );
  AND2_X1 U6081 ( .A1(n4819), .A2(n4970), .ZN(n4971) );
  OR2_X1 U6082 ( .A1(n4971), .A2(n4959), .ZN(n5191) );
  AOI22_X1 U6083 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5610), .B1(n4972), .B2(
        REIP_REG_16__SCAN_IN), .ZN(n4976) );
  OAI211_X1 U6084 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n4974), .B(n4973), .ZN(n4975) );
  NAND2_X1 U6085 ( .A1(n4976), .A2(n4975), .ZN(n4981) );
  INV_X1 U6086 ( .A(n4977), .ZN(n5194) );
  XOR2_X1 U6087 ( .A(n2990), .B(n4978), .Z(n5314) );
  AOI22_X1 U6088 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5595), 
        .B2(n5314), .ZN(n4979) );
  OAI21_X1 U6089 ( .B1(n5607), .B2(n5194), .A(n4979), .ZN(n4980) );
  NOR3_X1 U6090 ( .A1(n4981), .A2(n5581), .A3(n4980), .ZN(n4982) );
  OAI21_X1 U6091 ( .B1(n5191), .B2(n5564), .A(n4982), .ZN(U2811) );
  NOR2_X1 U6092 ( .A1(n4983), .A2(n5564), .ZN(n4984) );
  AOI211_X1 U6093 ( .C1(n5613), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5581), 
        .B(n4984), .ZN(n4997) );
  INV_X1 U6094 ( .A(n4985), .ZN(n4988) );
  NAND2_X1 U6095 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .ZN(
        n4987) );
  AOI21_X1 U6096 ( .B1(n4987), .B2(n4986), .A(n5582), .ZN(n5577) );
  OAI21_X1 U6097 ( .B1(n4989), .B2(n4988), .A(n5577), .ZN(n5541) );
  INV_X1 U6098 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6424) );
  NOR2_X1 U6099 ( .A1(n5597), .A2(n4990), .ZN(n5592) );
  NAND3_X1 U6100 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n5592), .ZN(n5559) );
  NOR2_X1 U6101 ( .A1(n6419), .A2(n5559), .ZN(n5551) );
  NAND3_X1 U6102 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n5551), .ZN(n5540) );
  AOI21_X1 U6103 ( .B1(n4729), .B2(n6424), .A(n5540), .ZN(n4991) );
  AOI22_X1 U6104 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5541), .B1(n4991), .B2(
        n5524), .ZN(n4996) );
  AOI22_X1 U6105 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5610), .B1(n4992), .B2(n5612), .ZN(n4993) );
  OAI21_X1 U6106 ( .B1(n5625), .B2(n5798), .A(n4993), .ZN(n4994) );
  INV_X1 U6107 ( .A(n4994), .ZN(n4995) );
  NAND3_X1 U6108 ( .A1(n4997), .A2(n4996), .A3(n4995), .ZN(U2817) );
  INV_X1 U6109 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4998) );
  OAI22_X1 U6110 ( .A1(n4999), .A2(n5078), .B1(n4998), .B2(n5076), .ZN(U2828)
         );
  OAI222_X1 U6111 ( .A1(n5068), .A2(n5084), .B1(n5076), .B2(n5000), .C1(n5212), 
        .C2(n5078), .ZN(U2829) );
  AOI22_X1 U6112 ( .A1(n5001), .A2(n5066), .B1(n5065), .B2(EBX_REG_29__SCAN_IN), .ZN(n5002) );
  OAI21_X1 U6113 ( .B1(n5087), .B2(n5068), .A(n5002), .ZN(U2830) );
  AOI22_X1 U6114 ( .A1(n5222), .A2(n5066), .B1(EBX_REG_28__SCAN_IN), .B2(n5065), .ZN(n5003) );
  OAI21_X1 U6115 ( .B1(n5090), .B2(n5068), .A(n5003), .ZN(U2831) );
  AOI22_X1 U6116 ( .A1(n5234), .A2(n5066), .B1(n5065), .B2(EBX_REG_27__SCAN_IN), .ZN(n5004) );
  OAI21_X1 U6117 ( .B1(n5093), .B2(n5068), .A(n5004), .ZN(U2832) );
  AOI22_X1 U6118 ( .A1(n5246), .A2(n5066), .B1(n5065), .B2(EBX_REG_26__SCAN_IN), .ZN(n5005) );
  OAI21_X1 U6119 ( .B1(n5129), .B2(n5068), .A(n5005), .ZN(U2833) );
  NOR2_X1 U6120 ( .A1(n4936), .A2(n5006), .ZN(n5007) );
  OR2_X1 U6121 ( .A1(n4922), .A2(n5007), .ZN(n5391) );
  NAND2_X1 U6122 ( .A1(n5009), .A2(n5008), .ZN(n5012) );
  INV_X1 U6123 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6124 ( .A1(n5012), .A2(n5011), .ZN(n5013) );
  NAND2_X1 U6125 ( .A1(n5013), .A2(n2992), .ZN(n5427) );
  OAI222_X1 U6126 ( .A1(n5068), .A2(n5391), .B1(n5076), .B2(n5014), .C1(n5427), 
        .C2(n5078), .ZN(U2834) );
  AOI22_X1 U6127 ( .A1(n5066), .A2(n5258), .B1(EBX_REG_24__SCAN_IN), .B2(n5065), .ZN(n5015) );
  OAI21_X1 U6128 ( .B1(n5146), .B2(n5068), .A(n5015), .ZN(U2835) );
  INV_X1 U6129 ( .A(n5262), .ZN(n5016) );
  AOI22_X1 U6130 ( .A1(n5066), .A2(n5016), .B1(n5065), .B2(EBX_REG_23__SCAN_IN), .ZN(n5017) );
  OAI21_X1 U6131 ( .B1(n5158), .B2(n5075), .A(n5017), .ZN(U2836) );
  AND2_X1 U6132 ( .A1(n2986), .A2(n5018), .ZN(n5020) );
  OR2_X1 U6133 ( .A1(n5020), .A2(n5019), .ZN(n5360) );
  INV_X1 U6134 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5025) );
  INV_X1 U6135 ( .A(n4948), .ZN(n5021) );
  AOI21_X1 U6136 ( .B1(n5023), .B2(n5022), .A(n5021), .ZN(n5396) );
  INV_X1 U6137 ( .A(n5396), .ZN(n5024) );
  OAI222_X1 U6138 ( .A1(n5078), .A2(n5360), .B1(n5076), .B2(n5025), .C1(n5024), 
        .C2(n5075), .ZN(U2837) );
  XNOR2_X1 U6139 ( .A(n5027), .B(n5028), .ZN(n5399) );
  NAND2_X1 U6140 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  NAND2_X1 U6141 ( .A1(n2986), .A2(n5031), .ZN(n5363) );
  INV_X1 U6142 ( .A(n5363), .ZN(n5032) );
  AOI22_X1 U6143 ( .A1(n5066), .A2(n5032), .B1(n5065), .B2(EBX_REG_21__SCAN_IN), .ZN(n5033) );
  OAI21_X1 U6144 ( .B1(n5399), .B2(n5075), .A(n5033), .ZN(U2838) );
  OR2_X1 U6145 ( .A1(n5034), .A2(n5035), .ZN(n5036) );
  AND2_X1 U6146 ( .A1(n5027), .A2(n5036), .ZN(n5403) );
  INV_X1 U6147 ( .A(n5403), .ZN(n5042) );
  NAND2_X1 U6148 ( .A1(n5038), .A2(n5045), .ZN(n5037) );
  OAI21_X1 U6149 ( .B1(n5038), .B2(n4111), .A(n5037), .ZN(n5041) );
  INV_X1 U6150 ( .A(n5039), .ZN(n5040) );
  XNOR2_X1 U6151 ( .A(n5041), .B(n5040), .ZN(n5375) );
  OAI222_X1 U6152 ( .A1(n5068), .A2(n5042), .B1(n5078), .B2(n5375), .C1(n5076), 
        .C2(n4153), .ZN(U2839) );
  AOI21_X1 U6153 ( .B1(n5044), .B2(n5043), .A(n5034), .ZN(n5187) );
  INV_X1 U6154 ( .A(n5187), .ZN(n5385) );
  NAND2_X1 U6155 ( .A1(n5045), .A2(n4111), .ZN(n5049) );
  INV_X1 U6156 ( .A(n5046), .ZN(n5047) );
  NAND2_X1 U6157 ( .A1(n5047), .A2(n4185), .ZN(n5048) );
  NAND2_X1 U6158 ( .A1(n5049), .A2(n5048), .ZN(n5054) );
  NAND2_X1 U6159 ( .A1(n5050), .A2(n5054), .ZN(n5058) );
  XNOR2_X1 U6160 ( .A(n5058), .B(n5051), .ZN(n5384) );
  INV_X1 U6161 ( .A(n5384), .ZN(n5052) );
  AOI22_X1 U6162 ( .A1(n5066), .A2(n5052), .B1(n5065), .B2(EBX_REG_19__SCAN_IN), .ZN(n5053) );
  OAI21_X1 U6163 ( .B1(n5385), .B2(n5068), .A(n5053), .ZN(U2840) );
  INV_X1 U6164 ( .A(n5054), .ZN(n5056) );
  NAND2_X1 U6165 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  NAND2_X1 U6166 ( .A1(n5058), .A2(n5057), .ZN(n5490) );
  INV_X1 U6167 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U6168 ( .A1(n5059), .A2(n5060), .ZN(n5061) );
  AND2_X1 U6169 ( .A1(n5043), .A2(n5061), .ZN(n5627) );
  INV_X1 U6170 ( .A(n5627), .ZN(n5062) );
  OAI222_X1 U6171 ( .A1(n5490), .A2(n5078), .B1(n5076), .B2(n6602), .C1(n5062), 
        .C2(n5075), .ZN(U2841) );
  AOI22_X1 U6172 ( .A1(n5066), .A2(n5441), .B1(n5065), .B2(EBX_REG_17__SCAN_IN), .ZN(n5063) );
  OAI21_X1 U6173 ( .B1(n5064), .B2(n5068), .A(n5063), .ZN(U2842) );
  AOI22_X1 U6174 ( .A1(n5066), .A2(n5314), .B1(n5065), .B2(EBX_REG_16__SCAN_IN), .ZN(n5067) );
  OAI21_X1 U6175 ( .B1(n5191), .B2(n5068), .A(n5067), .ZN(U2843) );
  OAI21_X1 U6176 ( .B1(n5071), .B2(n5070), .A(n5069), .ZN(n5493) );
  NOR2_X1 U6177 ( .A1(n5073), .A2(n5072), .ZN(n5074) );
  NOR2_X1 U6178 ( .A1(n4818), .A2(n5074), .ZN(n5497) );
  INV_X1 U6179 ( .A(n5497), .ZN(n5104) );
  OAI222_X1 U6180 ( .A1(n5493), .A2(n5078), .B1(n5077), .B2(n5076), .C1(n5075), 
        .C2(n5104), .ZN(U2845) );
  AOI22_X1 U6181 ( .A1(n5633), .A2(DATAI_30_), .B1(n5636), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5083) );
  INV_X1 U6182 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6183 ( .A1(n5637), .A2(DATAI_14_), .ZN(n5082) );
  OAI211_X1 U6184 ( .C1(n5084), .C2(n5395), .A(n5083), .B(n5082), .ZN(U2861)
         );
  AOI22_X1 U6185 ( .A1(n5633), .A2(DATAI_29_), .B1(n5636), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6186 ( .A1(n5637), .A2(DATAI_13_), .ZN(n5085) );
  OAI211_X1 U6187 ( .C1(n5087), .C2(n5395), .A(n5086), .B(n5085), .ZN(U2862)
         );
  AOI22_X1 U6188 ( .A1(n5633), .A2(DATAI_28_), .B1(n5636), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6189 ( .A1(n5637), .A2(DATAI_12_), .ZN(n5088) );
  OAI211_X1 U6190 ( .C1(n5090), .C2(n5395), .A(n5089), .B(n5088), .ZN(U2863)
         );
  AOI22_X1 U6191 ( .A1(n5633), .A2(DATAI_27_), .B1(n5636), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6192 ( .A1(n5637), .A2(DATAI_11_), .ZN(n5091) );
  OAI211_X1 U6193 ( .C1(n5093), .C2(n5395), .A(n5092), .B(n5091), .ZN(U2864)
         );
  AOI22_X1 U6194 ( .A1(n5633), .A2(DATAI_26_), .B1(n5636), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6195 ( .A1(n5637), .A2(DATAI_10_), .ZN(n5094) );
  OAI211_X1 U6196 ( .C1(n5129), .C2(n5395), .A(n5095), .B(n5094), .ZN(U2865)
         );
  AOI22_X1 U6197 ( .A1(n5633), .A2(DATAI_24_), .B1(n5636), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6198 ( .A1(n5637), .A2(DATAI_8_), .ZN(n5096) );
  OAI211_X1 U6199 ( .C1(n5146), .C2(n5395), .A(n5097), .B(n5096), .ZN(U2867)
         );
  AOI22_X1 U6200 ( .A1(n5633), .A2(DATAI_23_), .B1(n5636), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6201 ( .A1(n5637), .A2(DATAI_7_), .ZN(n5098) );
  OAI211_X1 U6202 ( .C1(n5158), .C2(n5395), .A(n5099), .B(n5098), .ZN(U2868)
         );
  AOI22_X1 U6203 ( .A1(n5633), .A2(DATAI_19_), .B1(n5636), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6204 ( .A1(n5637), .A2(DATAI_3_), .ZN(n5100) );
  OAI211_X1 U6205 ( .C1(n5385), .C2(n5395), .A(n5101), .B(n5100), .ZN(U2872)
         );
  AOI22_X1 U6206 ( .A1(n5102), .A2(DATAI_14_), .B1(n5636), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5103) );
  OAI21_X1 U6207 ( .B1(n5104), .B2(n5395), .A(n5103), .ZN(U2877) );
  NAND2_X1 U6208 ( .A1(n5754), .A2(n5105), .ZN(n5107) );
  OAI211_X1 U6209 ( .C1(n5782), .C2(n5108), .A(n5107), .B(n5106), .ZN(n5109)
         );
  AOI21_X1 U6210 ( .B1(n5110), .B2(n5774), .A(n5109), .ZN(n5111) );
  OAI21_X1 U6211 ( .B1(n5112), .B2(n5766), .A(n5111), .ZN(U2957) );
  NAND2_X1 U6212 ( .A1(n4061), .A2(n5113), .ZN(n5114) );
  XNOR2_X1 U6213 ( .A(n5114), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5241)
         );
  INV_X1 U6214 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6448) );
  NOR2_X1 U6215 ( .A1(n5845), .A2(n6448), .ZN(n5233) );
  AOI21_X1 U6216 ( .B1(n5771), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5233), 
        .ZN(n5115) );
  OAI21_X1 U6217 ( .B1(n5116), .B2(n5777), .A(n5115), .ZN(n5117) );
  AOI21_X1 U6218 ( .B1(n5118), .B2(n5774), .A(n5117), .ZN(n5119) );
  OAI21_X1 U6219 ( .B1(n5241), .B2(n5766), .A(n5119), .ZN(U2959) );
  NOR2_X1 U6220 ( .A1(n5845), .A2(n5120), .ZN(n5245) );
  NOR2_X1 U6221 ( .A1(n5777), .A2(n5121), .ZN(n5122) );
  AOI211_X1 U6222 ( .C1(n5771), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5245), 
        .B(n5122), .ZN(n5128) );
  NOR2_X1 U6223 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  XNOR2_X1 U6224 ( .A(n5126), .B(n5125), .ZN(n5242) );
  NAND2_X1 U6225 ( .A1(n5242), .A2(n5785), .ZN(n5127) );
  OAI211_X1 U6226 ( .C1(n5129), .C2(n6282), .A(n5128), .B(n5127), .ZN(U2960)
         );
  INV_X1 U6227 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5130) );
  OAI22_X1 U6228 ( .A1(n5782), .A2(n5131), .B1(n5845), .B2(n5130), .ZN(n5132)
         );
  AOI21_X1 U6229 ( .B1(n5754), .B2(n5341), .A(n5132), .ZN(n5137) );
  OAI21_X1 U6230 ( .B1(n5135), .B2(n5133), .A(n5134), .ZN(n5429) );
  NAND2_X1 U6231 ( .A1(n5429), .A2(n5785), .ZN(n5136) );
  OAI211_X1 U6232 ( .C1(n5391), .C2(n6282), .A(n5137), .B(n5136), .ZN(U2961)
         );
  NAND2_X1 U6233 ( .A1(n5182), .A2(n5414), .ZN(n5140) );
  XNOR2_X1 U6234 ( .A(n5414), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5176)
         );
  XNOR2_X1 U6235 ( .A(n5414), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5171)
         );
  NOR2_X1 U6236 ( .A1(n5414), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5163)
         );
  NAND2_X1 U6237 ( .A1(n5142), .A2(n5163), .ZN(n5154) );
  OAI21_X1 U6238 ( .B1(n5413), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5169), 
        .ZN(n5165) );
  NAND3_X1 U6239 ( .A1(n5414), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5143) );
  XNOR2_X1 U6240 ( .A(n5144), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5260)
         );
  NAND2_X1 U6241 ( .A1(n5817), .A2(REIP_REG_24__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U6242 ( .B1(n5782), .B2(n5145), .A(n5252), .ZN(n5148) );
  NOR2_X1 U6243 ( .A1(n5146), .A2(n6282), .ZN(n5147) );
  AOI211_X1 U6244 ( .C1(n5754), .C2(n5149), .A(n5148), .B(n5147), .ZN(n5150)
         );
  OAI21_X1 U6245 ( .B1(n5260), .B2(n5766), .A(n5150), .ZN(U2962) );
  INV_X1 U6246 ( .A(n5152), .ZN(n5272) );
  NAND3_X1 U6247 ( .A1(n5414), .A2(n5272), .A3(n5153), .ZN(n5155) );
  OAI21_X1 U6248 ( .B1(n5151), .B2(n5155), .A(n5154), .ZN(n5156) );
  XNOR2_X1 U6249 ( .A(n5156), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5268)
         );
  NAND2_X1 U6250 ( .A1(n5817), .A2(REIP_REG_23__SCAN_IN), .ZN(n5261) );
  OAI21_X1 U6251 ( .B1(n5782), .B2(n5157), .A(n5261), .ZN(n5160) );
  NOR2_X1 U6252 ( .A1(n5158), .A2(n6282), .ZN(n5159) );
  AOI211_X1 U6253 ( .C1(n5754), .C2(n5161), .A(n5160), .B(n5159), .ZN(n5162)
         );
  OAI21_X1 U6254 ( .B1(n5268), .B2(n5766), .A(n5162), .ZN(U2963) );
  AOI21_X1 U6255 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5414), .A(n5163), 
        .ZN(n5164) );
  XNOR2_X1 U6256 ( .A(n5165), .B(n5164), .ZN(n5277) );
  NAND2_X1 U6257 ( .A1(n5817), .A2(REIP_REG_22__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6258 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5166)
         );
  OAI211_X1 U6259 ( .C1(n5777), .C2(n5350), .A(n5270), .B(n5166), .ZN(n5167)
         );
  AOI21_X1 U6260 ( .B1(n5396), .B2(n5774), .A(n5167), .ZN(n5168) );
  OAI21_X1 U6261 ( .B1(n5277), .B2(n5766), .A(n5168), .ZN(U2964) );
  OAI21_X1 U6262 ( .B1(n5171), .B2(n5170), .A(n2977), .ZN(n5278) );
  NAND2_X1 U6263 ( .A1(n5278), .A2(n5785), .ZN(n5175) );
  INV_X1 U6264 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5172) );
  OAI22_X1 U6265 ( .A1(n5782), .A2(n5172), .B1(n5845), .B2(n6438), .ZN(n5173)
         );
  AOI21_X1 U6266 ( .B1(n5754), .B2(n5362), .A(n5173), .ZN(n5174) );
  OAI211_X1 U6267 ( .C1(n6282), .C2(n5399), .A(n5175), .B(n5174), .ZN(U2965)
         );
  XNOR2_X1 U6268 ( .A(n5177), .B(n5176), .ZN(n5299) );
  NAND2_X1 U6269 ( .A1(n5817), .A2(REIP_REG_20__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6270 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5178)
         );
  OAI211_X1 U6271 ( .C1(n5371), .C2(n5777), .A(n5294), .B(n5178), .ZN(n5179)
         );
  AOI21_X1 U6272 ( .B1(n5403), .B2(n5774), .A(n5179), .ZN(n5180) );
  OAI21_X1 U6273 ( .B1(n5299), .B2(n5766), .A(n5180), .ZN(U2966) );
  NAND2_X1 U6274 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  XNOR2_X1 U6275 ( .A(n5183), .B(n5414), .ZN(n5308) );
  INV_X1 U6276 ( .A(n5381), .ZN(n5185) );
  NAND2_X1 U6277 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5184)
         );
  NAND2_X1 U6278 ( .A1(n5817), .A2(REIP_REG_19__SCAN_IN), .ZN(n5304) );
  OAI211_X1 U6279 ( .C1(n5777), .C2(n5185), .A(n5184), .B(n5304), .ZN(n5186)
         );
  AOI21_X1 U6280 ( .B1(n5187), .B2(n5774), .A(n5186), .ZN(n5188) );
  OAI21_X1 U6281 ( .B1(n5766), .B2(n5308), .A(n5188), .ZN(U2967) );
  XNOR2_X1 U6282 ( .A(n5414), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5190)
         );
  XNOR2_X1 U6283 ( .A(n5189), .B(n5190), .ZN(n5317) );
  INV_X1 U6284 ( .A(n5191), .ZN(n5635) );
  INV_X1 U6285 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5192) );
  NOR2_X1 U6286 ( .A1(n5845), .A2(n5192), .ZN(n5313) );
  AOI21_X1 U6287 ( .B1(n5771), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5313), 
        .ZN(n5193) );
  OAI21_X1 U6288 ( .B1(n5194), .B2(n5777), .A(n5193), .ZN(n5195) );
  AOI21_X1 U6289 ( .B1(n5635), .B2(n5774), .A(n5195), .ZN(n5196) );
  OAI21_X1 U6290 ( .B1(n5317), .B2(n5766), .A(n5196), .ZN(U2970) );
  XNOR2_X1 U6291 ( .A(n5414), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5198)
         );
  XNOR2_X1 U6292 ( .A(n5197), .B(n5198), .ZN(n5449) );
  NAND2_X1 U6293 ( .A1(n5449), .A2(n5785), .ZN(n5203) );
  NOR2_X1 U6294 ( .A1(n5845), .A2(n6430), .ZN(n5446) );
  INV_X1 U6295 ( .A(n5199), .ZN(n5200) );
  NOR2_X1 U6296 ( .A1(n5777), .A2(n5200), .ZN(n5201) );
  AOI211_X1 U6297 ( .C1(n5771), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5446), 
        .B(n5201), .ZN(n5202) );
  OAI211_X1 U6298 ( .C1(n6282), .C2(n5204), .A(n5203), .B(n5202), .ZN(U2971)
         );
  XNOR2_X1 U6299 ( .A(n5414), .B(n5321), .ZN(n5205) );
  XNOR2_X1 U6300 ( .A(n5206), .B(n5205), .ZN(n5331) );
  NAND2_X1 U6301 ( .A1(n5817), .A2(REIP_REG_14__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6302 ( .A1(n5771), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5207)
         );
  OAI211_X1 U6303 ( .C1(n5777), .C2(n5208), .A(n5326), .B(n5207), .ZN(n5209)
         );
  AOI21_X1 U6304 ( .B1(n5497), .B2(n5774), .A(n5209), .ZN(n5210) );
  OAI21_X1 U6305 ( .B1(n5766), .B2(n5331), .A(n5210), .ZN(U2972) );
  INV_X1 U6306 ( .A(n5211), .ZN(n5220) );
  INV_X1 U6307 ( .A(n5212), .ZN(n5216) );
  NOR3_X1 U6308 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6498), 
        .ZN(n5214) );
  AOI211_X1 U6309 ( .C1(n5836), .C2(n5216), .A(n5215), .B(n5214), .ZN(n5219)
         );
  NAND2_X1 U6310 ( .A1(n5217), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5218) );
  OAI211_X1 U6311 ( .C1(n5220), .C2(n5825), .A(n5219), .B(n5218), .ZN(U2988)
         );
  INV_X1 U6312 ( .A(n5221), .ZN(n5231) );
  INV_X1 U6313 ( .A(n5222), .ZN(n5223) );
  NOR2_X1 U6314 ( .A1(n5223), .A2(n5799), .ZN(n5224) );
  AOI211_X1 U6315 ( .C1(n5232), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5225), .B(n5224), .ZN(n5230) );
  NOR2_X1 U6316 ( .A1(n5432), .A2(n5247), .ZN(n5239) );
  INV_X1 U6317 ( .A(n5226), .ZN(n5228) );
  NAND3_X1 U6318 ( .A1(n5239), .A2(n5228), .A3(n5227), .ZN(n5229) );
  OAI211_X1 U6319 ( .C1(n5231), .C2(n5825), .A(n5230), .B(n5229), .ZN(U2990)
         );
  INV_X1 U6320 ( .A(n5232), .ZN(n5236) );
  AOI21_X1 U6321 ( .B1(n5234), .B2(n5836), .A(n5233), .ZN(n5235) );
  OAI21_X1 U6322 ( .B1(n5236), .B2(n5238), .A(n5235), .ZN(n5237) );
  AOI21_X1 U6323 ( .B1(n5239), .B2(n5238), .A(n5237), .ZN(n5240) );
  OAI21_X1 U6324 ( .B1(n5241), .B2(n5825), .A(n5240), .ZN(U2991) );
  INV_X1 U6325 ( .A(n5242), .ZN(n5251) );
  INV_X1 U6326 ( .A(n5426), .ZN(n5253) );
  NOR2_X1 U6327 ( .A1(n5253), .A2(n5243), .ZN(n5244) );
  AOI211_X1 U6328 ( .C1(n5836), .C2(n5246), .A(n5245), .B(n5244), .ZN(n5250)
         );
  INV_X1 U6329 ( .A(n5432), .ZN(n5248) );
  OAI211_X1 U6330 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5248), .B(n5247), .ZN(n5249) );
  OAI211_X1 U6331 ( .C1(n5251), .C2(n5825), .A(n5250), .B(n5249), .ZN(U2992)
         );
  INV_X1 U6332 ( .A(n5252), .ZN(n5257) );
  NAND3_X1 U6333 ( .A1(n5271), .A2(n5272), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5254) );
  AOI21_X1 U6334 ( .B1(n5255), .B2(n5254), .A(n5253), .ZN(n5256) );
  AOI211_X1 U6335 ( .C1(n5836), .C2(n5258), .A(n5257), .B(n5256), .ZN(n5259)
         );
  OAI21_X1 U6336 ( .B1(n5260), .B2(n5825), .A(n5259), .ZN(U2994) );
  OAI21_X1 U6337 ( .B1(n5799), .B2(n5262), .A(n5261), .ZN(n5263) );
  AOI21_X1 U6338 ( .B1(n5264), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5263), 
        .ZN(n5267) );
  NAND3_X1 U6339 ( .A1(n5271), .A2(n5272), .A3(n5265), .ZN(n5266) );
  OAI211_X1 U6340 ( .C1(n5268), .C2(n5825), .A(n5267), .B(n5266), .ZN(U2995)
         );
  INV_X1 U6341 ( .A(n5269), .ZN(n5281) );
  OAI21_X1 U6342 ( .B1(n5799), .B2(n5360), .A(n5270), .ZN(n5275) );
  INV_X1 U6343 ( .A(n5271), .ZN(n5284) );
  NOR3_X1 U6344 ( .A1(n5284), .A2(n5273), .A3(n5272), .ZN(n5274) );
  AOI211_X1 U6345 ( .C1(n5281), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5275), .B(n5274), .ZN(n5276) );
  OAI21_X1 U6346 ( .B1(n5277), .B2(n5825), .A(n5276), .ZN(U2996) );
  NAND2_X1 U6347 ( .A1(n5278), .A2(n5837), .ZN(n5283) );
  NAND2_X1 U6348 ( .A1(n5817), .A2(REIP_REG_21__SCAN_IN), .ZN(n5279) );
  OAI21_X1 U6349 ( .B1(n5799), .B2(n5363), .A(n5279), .ZN(n5280) );
  AOI21_X1 U6350 ( .B1(n5281), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5280), 
        .ZN(n5282) );
  OAI211_X1 U6351 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5284), .A(n5283), .B(n5282), .ZN(U2997) );
  NOR2_X1 U6352 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5285) );
  INV_X1 U6353 ( .A(n5440), .ZN(n5300) );
  NOR3_X1 U6354 ( .A1(n5285), .A2(n5301), .A3(n5300), .ZN(n5297) );
  INV_X1 U6355 ( .A(n5286), .ZN(n5296) );
  NAND2_X1 U6356 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  OAI221_X1 U6357 ( .B1(n5291), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n5291), .C2(n5290), .A(n5289), .ZN(n5442) );
  AOI21_X1 U6358 ( .B1(n5819), .B2(n5439), .A(n5442), .ZN(n5433) );
  OAI21_X1 U6359 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5292), .A(n5433), 
        .ZN(n5302) );
  NAND2_X1 U6360 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n5302), .ZN(n5293) );
  OAI211_X1 U6361 ( .C1(n5799), .C2(n5375), .A(n5294), .B(n5293), .ZN(n5295)
         );
  AOI21_X1 U6362 ( .B1(n5297), .B2(n5296), .A(n5295), .ZN(n5298) );
  OAI21_X1 U6363 ( .B1(n5299), .B2(n5825), .A(n5298), .ZN(U2998) );
  NOR2_X1 U6364 ( .A1(n5301), .A2(n5300), .ZN(n5306) );
  NAND2_X1 U6365 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5302), .ZN(n5303) );
  OAI211_X1 U6366 ( .C1(n5799), .C2(n5384), .A(n5304), .B(n5303), .ZN(n5305)
         );
  AOI21_X1 U6367 ( .B1(n5306), .B2(n5138), .A(n5305), .ZN(n5307) );
  OAI21_X1 U6368 ( .B1(n5308), .B2(n5825), .A(n5307), .ZN(U2999) );
  AOI21_X1 U6369 ( .B1(n5309), .B2(n5797), .A(n5792), .ZN(n5452) );
  NAND2_X1 U6370 ( .A1(n5448), .A2(n5310), .ZN(n5311) );
  OAI21_X1 U6371 ( .B1(n5452), .B2(n5412), .A(n5311), .ZN(n5312) );
  OAI21_X1 U6372 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5312), .ZN(n5316) );
  AOI21_X1 U6373 ( .B1(n5836), .B2(n5314), .A(n5313), .ZN(n5315) );
  OAI211_X1 U6374 ( .C1(n5317), .C2(n5825), .A(n5316), .B(n5315), .ZN(U3002)
         );
  OAI21_X1 U6375 ( .B1(n5320), .B2(n5319), .A(n5318), .ZN(n5322) );
  AOI21_X1 U6376 ( .B1(n5323), .B2(n5322), .A(n5321), .ZN(n5329) );
  NOR3_X1 U6377 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5325), .A3(n5324), 
        .ZN(n5328) );
  OAI21_X1 U6378 ( .B1(n5799), .B2(n5493), .A(n5326), .ZN(n5327) );
  NOR3_X1 U6379 ( .A1(n5329), .A2(n5328), .A3(n5327), .ZN(n5330) );
  OAI21_X1 U6380 ( .B1(n5331), .B2(n5825), .A(n5330), .ZN(U3004) );
  OAI211_X1 U6381 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6283), .A(n6131), .B(
        n6290), .ZN(n5332) );
  OAI21_X1 U6382 ( .B1(n5334), .B2(n4495), .A(n5332), .ZN(n5333) );
  MUX2_X1 U6383 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5333), .S(n5846), 
        .Z(U3464) );
  XNOR2_X1 U6384 ( .A(n4460), .B(n6131), .ZN(n5335) );
  OAI22_X1 U6385 ( .A1(n5335), .A2(n6278), .B1(n2981), .B2(n5334), .ZN(n5336)
         );
  MUX2_X1 U6386 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5336), .S(n5846), 
        .Z(U3463) );
  OAI22_X1 U6387 ( .A1(n5338), .A2(n6474), .B1(n5337), .B2(n6379), .ZN(n5339)
         );
  MUX2_X1 U6388 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5339), .S(n6472), 
        .Z(U3456) );
  AND2_X1 U6389 ( .A1(n5669), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6390 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5610), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5613), .ZN(n5348) );
  AOI22_X1 U6391 ( .A1(n5341), .A2(n5612), .B1(n5340), .B2(n5130), .ZN(n5347)
         );
  OAI22_X1 U6392 ( .A1(n5391), .A2(n5564), .B1(n5625), .B2(n5427), .ZN(n5342)
         );
  INV_X1 U6393 ( .A(n5342), .ZN(n5346) );
  OAI21_X1 U6394 ( .B1(n5344), .B2(n5343), .A(REIP_REG_25__SCAN_IN), .ZN(n5345) );
  NAND4_X1 U6395 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(U2802)
         );
  NOR2_X1 U6396 ( .A1(n5349), .A2(REIP_REG_22__SCAN_IN), .ZN(n5355) );
  INV_X1 U6397 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5353) );
  INV_X1 U6398 ( .A(n5350), .ZN(n5351) );
  AOI22_X1 U6399 ( .A1(n5612), .A2(n5351), .B1(n5610), .B2(EBX_REG_22__SCAN_IN), .ZN(n5352) );
  OAI21_X1 U6400 ( .B1(n5603), .B2(n5353), .A(n5352), .ZN(n5354) );
  AOI211_X1 U6401 ( .C1(n5396), .C2(n5555), .A(n5355), .B(n5354), .ZN(n5359)
         );
  NAND2_X1 U6402 ( .A1(n6438), .A2(n5356), .ZN(n5365) );
  INV_X1 U6403 ( .A(n5365), .ZN(n5357) );
  OAI21_X1 U6404 ( .B1(n5357), .B2(n5361), .A(REIP_REG_22__SCAN_IN), .ZN(n5358) );
  OAI211_X1 U6405 ( .C1(n5625), .C2(n5360), .A(n5359), .B(n5358), .ZN(U2805)
         );
  AOI22_X1 U6406 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5610), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5613), .ZN(n5368) );
  AOI22_X1 U6407 ( .A1(n5362), .A2(n5612), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5361), .ZN(n5367) );
  OAI22_X1 U6408 ( .A1(n5399), .A2(n5564), .B1(n5625), .B2(n5363), .ZN(n5364)
         );
  INV_X1 U6409 ( .A(n5364), .ZN(n5366) );
  NAND4_X1 U6410 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(U2806)
         );
  AOI21_X1 U6411 ( .B1(n6437), .B2(n5370), .A(n5369), .ZN(n5374) );
  INV_X1 U6412 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5372) );
  OAI22_X1 U6413 ( .A1(n5372), .A2(n5603), .B1(n5371), .B2(n5607), .ZN(n5373)
         );
  AOI211_X1 U6414 ( .C1(n5610), .C2(EBX_REG_20__SCAN_IN), .A(n5374), .B(n5373), 
        .ZN(n5378) );
  NOR2_X1 U6415 ( .A1(n5375), .A2(n5625), .ZN(n5376) );
  AOI21_X1 U6416 ( .B1(n5403), .B2(n5555), .A(n5376), .ZN(n5377) );
  NAND2_X1 U6417 ( .A1(n5378), .A2(n5377), .ZN(U2807) );
  NAND2_X1 U6418 ( .A1(n5380), .A2(n6434), .ZN(n5481) );
  NOR2_X1 U6419 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6434), .ZN(n5379) );
  AOI22_X1 U6420 ( .A1(n5381), .A2(n5612), .B1(n5380), .B2(n5379), .ZN(n5382)
         );
  OAI211_X1 U6421 ( .C1(n5603), .C2(n5383), .A(n5382), .B(n5561), .ZN(n5387)
         );
  OAI22_X1 U6422 ( .A1(n5385), .A2(n5564), .B1(n5384), .B2(n5625), .ZN(n5386)
         );
  AOI211_X1 U6423 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5610), .A(n5387), .B(n5386), 
        .ZN(n5388) );
  OAI221_X1 U6424 ( .B1(n6435), .B2(n5480), .C1(n6435), .C2(n5481), .A(n5388), 
        .ZN(U2808) );
  INV_X1 U6425 ( .A(n5633), .ZN(n5390) );
  OAI22_X1 U6426 ( .A1(n5391), .A2(n5395), .B1(n5390), .B2(n5389), .ZN(n5392)
         );
  INV_X1 U6427 ( .A(n5392), .ZN(n5394) );
  AOI22_X1 U6428 ( .A1(n5637), .A2(DATAI_9_), .B1(n5636), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6429 ( .A1(n5394), .A2(n5393), .ZN(U2866) );
  INV_X1 U6430 ( .A(n5395), .ZN(n5634) );
  AOI22_X1 U6431 ( .A1(n5396), .A2(n5634), .B1(n5633), .B2(DATAI_22_), .ZN(
        n5398) );
  AOI22_X1 U6432 ( .A1(n5637), .A2(DATAI_6_), .B1(n5636), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6433 ( .A1(n5398), .A2(n5397), .ZN(U2869) );
  INV_X1 U6434 ( .A(n5399), .ZN(n5400) );
  AOI22_X1 U6435 ( .A1(n5400), .A2(n5634), .B1(n5633), .B2(DATAI_21_), .ZN(
        n5402) );
  AOI22_X1 U6436 ( .A1(n5637), .A2(DATAI_5_), .B1(n5636), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6437 ( .A1(n5402), .A2(n5401), .ZN(U2870) );
  AOI22_X1 U6438 ( .A1(n5403), .A2(n5634), .B1(n5633), .B2(DATAI_20_), .ZN(
        n5405) );
  AOI22_X1 U6439 ( .A1(n5637), .A2(DATAI_4_), .B1(n5636), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6440 ( .A1(n5405), .A2(n5404), .ZN(U2871) );
  AOI22_X1 U6441 ( .A1(n5817), .A2(REIP_REG_18__SCAN_IN), .B1(n5771), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5411) );
  NOR2_X1 U6442 ( .A1(n5189), .A2(n5406), .ZN(n5408) );
  NOR2_X1 U6443 ( .A1(n5151), .A2(n5439), .ZN(n5407) );
  MUX2_X1 U6444 ( .A(n5408), .B(n5407), .S(n5414), .Z(n5409) );
  XOR2_X1 U6445 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5409), .Z(n5435) );
  AOI22_X1 U6446 ( .A1(n5435), .A2(n5785), .B1(n5774), .B2(n5627), .ZN(n5410)
         );
  OAI211_X1 U6447 ( .C1(n5777), .C2(n5483), .A(n5411), .B(n5410), .ZN(U2968)
         );
  NAND2_X1 U6448 ( .A1(n5413), .A2(n5412), .ZN(n5416) );
  NAND3_X1 U6449 ( .A1(n5189), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5414), .ZN(n5415) );
  OAI21_X1 U6450 ( .B1(n5189), .B2(n5416), .A(n5415), .ZN(n5417) );
  XNOR2_X1 U6451 ( .A(n5417), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5445)
         );
  AOI22_X1 U6452 ( .A1(n5817), .A2(REIP_REG_17__SCAN_IN), .B1(n5771), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5420) );
  AOI22_X1 U6453 ( .A1(n5630), .A2(n5774), .B1(n5418), .B2(n5754), .ZN(n5419)
         );
  OAI211_X1 U6454 ( .C1(n5445), .C2(n5766), .A(n5420), .B(n5419), .ZN(U2969)
         );
  INV_X1 U6455 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5425) );
  INV_X1 U6456 ( .A(n5513), .ZN(n5421) );
  AOI222_X1 U6457 ( .A1(n5422), .A2(n5785), .B1(n5421), .B2(n5754), .C1(n5774), 
        .C2(n5507), .ZN(n5424) );
  OAI211_X1 U6458 ( .C1(n5425), .C2(n5782), .A(n5424), .B(n5423), .ZN(U2973)
         );
  AOI22_X1 U6459 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5426), .B1(n5817), .B2(REIP_REG_25__SCAN_IN), .ZN(n5431) );
  INV_X1 U6460 ( .A(n5427), .ZN(n5428) );
  AOI22_X1 U6461 ( .A1(n5429), .A2(n5837), .B1(n5836), .B2(n5428), .ZN(n5430)
         );
  OAI211_X1 U6462 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5432), .A(n5431), .B(n5430), .ZN(U2993) );
  OAI22_X1 U6463 ( .A1(n5799), .A2(n5490), .B1(n5436), .B2(n5433), .ZN(n5434)
         );
  AOI21_X1 U6464 ( .B1(n5837), .B2(n5435), .A(n5434), .ZN(n5438) );
  NAND3_X1 U6465 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5440), .A3(n5436), .ZN(n5437) );
  OAI211_X1 U6466 ( .C1(n6434), .C2(n5845), .A(n5438), .B(n5437), .ZN(U3000)
         );
  AOI22_X1 U6467 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5817), .B1(n5440), .B2(
        n5439), .ZN(n5444) );
  AOI22_X1 U6468 ( .A1(n5442), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n5836), .B2(n5441), .ZN(n5443) );
  OAI211_X1 U6469 ( .C1(n5445), .C2(n5825), .A(n5444), .B(n5443), .ZN(U3001)
         );
  AOI21_X1 U6470 ( .B1(n5836), .B2(n5447), .A(n5446), .ZN(n5451) );
  AOI22_X1 U6471 ( .A1(n5449), .A2(n5837), .B1(n3964), .B2(n5448), .ZN(n5450)
         );
  OAI211_X1 U6472 ( .C1(n5452), .C2(n3964), .A(n5451), .B(n5450), .ZN(U3003)
         );
  OR2_X1 U6473 ( .A1(n5453), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5455) );
  OAI22_X1 U6474 ( .A1(n5456), .A2(n5455), .B1(n5454), .B2(n6472), .ZN(U3455)
         );
  INV_X1 U6475 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6403) );
  AOI21_X1 U6476 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6403), .A(n6405), .ZN(n5461) );
  INV_X1 U6477 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5457) );
  INV_X1 U6478 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6563) );
  NOR2_X2 U6479 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6563), .ZN(n6494) );
  AOI21_X1 U6480 ( .B1(n5461), .B2(n5457), .A(n6494), .ZN(U2789) );
  OAI21_X1 U6481 ( .B1(n5458), .B2(n6385), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5459) );
  OAI21_X1 U6482 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6386), .A(n5459), .ZN(
        U2790) );
  INV_X2 U6483 ( .A(n6494), .ZN(n6483) );
  NOR2_X1 U6484 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5462) );
  OAI21_X1 U6485 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5462), .A(n6483), .ZN(n5460)
         );
  OAI21_X1 U6486 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6483), .A(n5460), .ZN(
        U2791) );
  NOR2_X1 U6487 ( .A1(n6494), .A2(n5461), .ZN(n6462) );
  OAI21_X1 U6488 ( .B1(BS16_N), .B2(n5462), .A(n6462), .ZN(n6460) );
  OAI21_X1 U6489 ( .B1(n6462), .B2(n6167), .A(n6460), .ZN(U2792) );
  INV_X1 U6490 ( .A(n5463), .ZN(n5465) );
  OAI21_X1 U6491 ( .B1(n5465), .B2(n5464), .A(n5766), .ZN(U2793) );
  NOR4_X1 U6492 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5469) );
  NOR4_X1 U6493 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5468) );
  NOR4_X1 U6494 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5467) );
  NOR4_X1 U6495 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5466) );
  NAND4_X1 U6496 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n5475)
         );
  NOR4_X1 U6497 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5473) );
  AOI211_X1 U6498 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_25__SCAN_IN), .B(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5472) );
  NOR4_X1 U6499 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n5471) );
  NOR4_X1 U6500 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5470) );
  NAND4_X1 U6501 ( .A1(n5473), .A2(n5472), .A3(n5471), .A4(n5470), .ZN(n5474)
         );
  NOR2_X1 U6502 ( .A1(n5475), .A2(n5474), .ZN(n6479) );
  INV_X1 U6503 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5477) );
  NOR3_X1 U6504 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5478) );
  OAI21_X1 U6505 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5478), .A(n6479), .ZN(n5476)
         );
  OAI21_X1 U6506 ( .B1(n6479), .B2(n5477), .A(n5476), .ZN(U2794) );
  INV_X1 U6507 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6461) );
  AOI21_X1 U6508 ( .B1(n5615), .B2(n6461), .A(n5478), .ZN(n5479) );
  INV_X1 U6509 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6607) );
  INV_X1 U6510 ( .A(n6479), .ZN(n6481) );
  AOI22_X1 U6511 ( .A1(n6479), .A2(n5479), .B1(n6607), .B2(n6481), .ZN(U2795)
         );
  OR2_X1 U6512 ( .A1(n5480), .A2(n6434), .ZN(n5487) );
  AOI22_X1 U6513 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5610), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5613), .ZN(n5482) );
  NAND3_X1 U6514 ( .A1(n5482), .A2(n5481), .A3(n5561), .ZN(n5485) );
  NOR2_X1 U6515 ( .A1(n5607), .A2(n5483), .ZN(n5484) );
  NOR2_X1 U6516 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  NAND2_X1 U6517 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  AOI21_X1 U6518 ( .B1(n5627), .B2(n5555), .A(n5488), .ZN(n5489) );
  OAI21_X1 U6519 ( .B1(n5625), .B2(n5490), .A(n5489), .ZN(U2809) );
  AND2_X1 U6520 ( .A1(n5492), .A2(n5491), .ZN(n5502) );
  AOI21_X1 U6521 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5502), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5501) );
  OAI22_X1 U6522 ( .A1(n5494), .A2(n5603), .B1(n5625), .B2(n5493), .ZN(n5495)
         );
  AOI211_X1 U6523 ( .C1(n5610), .C2(EBX_REG_14__SCAN_IN), .A(n5581), .B(n5495), 
        .ZN(n5499) );
  AOI22_X1 U6524 ( .A1(n5497), .A2(n5555), .B1(n5612), .B2(n5496), .ZN(n5498)
         );
  OAI211_X1 U6525 ( .C1(n5501), .C2(n5500), .A(n5499), .B(n5498), .ZN(U2813)
         );
  INV_X1 U6526 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U6527 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5610), .B1(n5502), .B2(n6561), .ZN(n5504) );
  AOI21_X1 U6528 ( .B1(n5613), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5581), 
        .ZN(n5503) );
  OAI211_X1 U6529 ( .C1(n5505), .C2(n5625), .A(n5504), .B(n5503), .ZN(n5506)
         );
  AOI21_X1 U6530 ( .B1(n5507), .B2(n5555), .A(n5506), .ZN(n5512) );
  INV_X1 U6531 ( .A(n5508), .ZN(n5509) );
  OAI21_X1 U6532 ( .B1(n5509), .B2(n5597), .A(n2956), .ZN(n5525) );
  NAND2_X1 U6533 ( .A1(n5509), .A2(n6517), .ZN(n5510) );
  NOR2_X1 U6534 ( .A1(n5597), .A2(n5510), .ZN(n5516) );
  OAI21_X1 U6535 ( .B1(n5525), .B2(n5516), .A(REIP_REG_13__SCAN_IN), .ZN(n5511) );
  OAI211_X1 U6536 ( .C1(n5607), .C2(n5513), .A(n5512), .B(n5511), .ZN(U2814)
         );
  AOI21_X1 U6537 ( .B1(n5613), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5581), 
        .ZN(n5522) );
  NOR2_X1 U6538 ( .A1(n5584), .A2(n5514), .ZN(n5515) );
  AOI211_X1 U6539 ( .C1(n5525), .C2(REIP_REG_12__SCAN_IN), .A(n5516), .B(n5515), .ZN(n5517) );
  OAI21_X1 U6540 ( .B1(n5518), .B2(n5564), .A(n5517), .ZN(n5519) );
  AOI21_X1 U6541 ( .B1(n5520), .B2(n5612), .A(n5519), .ZN(n5521) );
  OAI211_X1 U6542 ( .C1(n5625), .C2(n5523), .A(n5522), .B(n5521), .ZN(U2815)
         );
  AOI22_X1 U6543 ( .A1(n5744), .A2(n5555), .B1(n5612), .B2(n5743), .ZN(n5531)
         );
  NOR3_X1 U6544 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5524), .A3(n5540), .ZN(n5529) );
  AOI22_X1 U6545 ( .A1(n5595), .A2(n5789), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5525), .ZN(n5526) );
  OAI211_X1 U6546 ( .C1(n5603), .C2(n5527), .A(n5526), .B(n5561), .ZN(n5528)
         );
  AOI211_X1 U6547 ( .C1(n5610), .C2(EBX_REG_11__SCAN_IN), .A(n5529), .B(n5528), 
        .ZN(n5530) );
  NAND2_X1 U6548 ( .A1(n5531), .A2(n5530), .ZN(U2816) );
  AOI22_X1 U6549 ( .A1(n5532), .A2(n5612), .B1(n5595), .B2(n5810), .ZN(n5533)
         );
  OAI211_X1 U6550 ( .C1(n5603), .C2(n5534), .A(n5533), .B(n5561), .ZN(n5535)
         );
  AOI21_X1 U6551 ( .B1(EBX_REG_9__SCAN_IN), .B2(n5610), .A(n5535), .ZN(n5539)
         );
  INV_X1 U6552 ( .A(n5536), .ZN(n5537) );
  AOI22_X1 U6553 ( .A1(n5537), .A2(n5555), .B1(REIP_REG_9__SCAN_IN), .B2(n5541), .ZN(n5538) );
  OAI211_X1 U6554 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5540), .A(n5539), .B(n5538), 
        .ZN(U2818) );
  INV_X1 U6555 ( .A(n5541), .ZN(n5550) );
  AOI21_X1 U6556 ( .B1(REIP_REG_7__SCAN_IN), .B2(n5551), .A(
        REIP_REG_8__SCAN_IN), .ZN(n5549) );
  OAI22_X1 U6557 ( .A1(n6544), .A2(n5603), .B1(n5625), .B2(n5542), .ZN(n5543)
         );
  AOI211_X1 U6558 ( .C1(n5610), .C2(EBX_REG_8__SCAN_IN), .A(n5581), .B(n5543), 
        .ZN(n5548) );
  INV_X1 U6559 ( .A(n5544), .ZN(n5545) );
  AOI22_X1 U6560 ( .A1(n5546), .A2(n5555), .B1(n5545), .B2(n5612), .ZN(n5547)
         );
  OAI211_X1 U6561 ( .C1(n5550), .C2(n5549), .A(n5548), .B(n5547), .ZN(U2819)
         );
  INV_X1 U6562 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6421) );
  AOI22_X1 U6563 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5610), .B1(n5551), .B2(n6421), 
        .ZN(n5552) );
  OAI21_X1 U6564 ( .B1(n5625), .B2(n5553), .A(n5552), .ZN(n5554) );
  AOI211_X1 U6565 ( .C1(n5613), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5581), 
        .B(n5554), .ZN(n5558) );
  OAI21_X1 U6566 ( .B1(REIP_REG_6__SCAN_IN), .B2(n5559), .A(n5577), .ZN(n5556)
         );
  AOI22_X1 U6567 ( .A1(n5556), .A2(REIP_REG_7__SCAN_IN), .B1(n5749), .B2(n5555), .ZN(n5557) );
  OAI211_X1 U6568 ( .C1(n5747), .C2(n5607), .A(n5558), .B(n5557), .ZN(U2820)
         );
  NOR2_X1 U6569 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5559), .ZN(n5568) );
  AOI22_X1 U6570 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5610), .B1(n5595), .B2(n5560), 
        .ZN(n5562) );
  OAI211_X1 U6571 ( .C1(n5603), .C2(n5563), .A(n5562), .B(n5561), .ZN(n5567)
         );
  OAI22_X1 U6572 ( .A1(n5565), .A2(n5564), .B1(n6419), .B2(n5577), .ZN(n5566)
         );
  NOR3_X1 U6573 ( .A1(n5568), .A2(n5567), .A3(n5566), .ZN(n5569) );
  OAI21_X1 U6574 ( .B1(n5570), .B2(n5607), .A(n5569), .ZN(U2821) );
  AOI21_X1 U6575 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5592), .A(
        REIP_REG_5__SCAN_IN), .ZN(n5576) );
  OAI22_X1 U6576 ( .A1(n5760), .A2(n5603), .B1(n5625), .B2(n5571), .ZN(n5572)
         );
  AOI211_X1 U6577 ( .C1(n5610), .C2(EBX_REG_5__SCAN_IN), .A(n5581), .B(n5572), 
        .ZN(n5575) );
  INV_X1 U6578 ( .A(n5573), .ZN(n5756) );
  AOI22_X1 U6579 ( .A1(n5756), .A2(n5622), .B1(n5755), .B2(n5612), .ZN(n5574)
         );
  OAI211_X1 U6580 ( .C1(n5577), .C2(n5576), .A(n5575), .B(n5574), .ZN(U2822)
         );
  OAI22_X1 U6581 ( .A1(n5579), .A2(n5603), .B1(n5625), .B2(n5578), .ZN(n5580)
         );
  AOI211_X1 U6582 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5582), .A(n5581), .B(n5580), 
        .ZN(n5594) );
  INV_X1 U6583 ( .A(n5583), .ZN(n5586) );
  OAI22_X1 U6584 ( .A1(n5586), .A2(n5614), .B1(n5585), .B2(n5584), .ZN(n5591)
         );
  INV_X1 U6585 ( .A(n5587), .ZN(n5588) );
  OAI22_X1 U6586 ( .A1(n5589), .A2(n5596), .B1(n5588), .B2(n5607), .ZN(n5590)
         );
  AOI211_X1 U6587 ( .C1(n5592), .C2(n6418), .A(n5591), .B(n5590), .ZN(n5593)
         );
  NAND2_X1 U6588 ( .A1(n5594), .A2(n5593), .ZN(U2823) );
  AOI22_X1 U6589 ( .A1(EBX_REG_2__SCAN_IN), .A2(n5610), .B1(n5595), .B2(n5818), 
        .ZN(n5606) );
  OR2_X1 U6590 ( .A1(n5765), .A2(n5596), .ZN(n5602) );
  INV_X1 U6591 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6415) );
  OAI21_X1 U6592 ( .B1(n5597), .B2(n5615), .A(n6415), .ZN(n5599) );
  INV_X1 U6593 ( .A(n2981), .ZN(n5956) );
  AOI22_X1 U6594 ( .A1(n5600), .A2(n5599), .B1(n5956), .B2(n5598), .ZN(n5601)
         );
  OAI211_X1 U6595 ( .C1(n3424), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5604)
         );
  INV_X1 U6596 ( .A(n5604), .ZN(n5605) );
  OAI211_X1 U6597 ( .C1(n5770), .C2(n5607), .A(n5606), .B(n5605), .ZN(U2825)
         );
  INV_X1 U6598 ( .A(n5608), .ZN(n5609) );
  AOI21_X1 U6599 ( .B1(n5610), .B2(EBX_REG_1__SCAN_IN), .A(n5609), .ZN(n5624)
         );
  INV_X1 U6600 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6601 ( .A1(n5612), .A2(n5611), .ZN(n5620) );
  NAND2_X1 U6602 ( .A1(n5613), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5619)
         );
  OAI22_X1 U6603 ( .A1(n2956), .A2(n5615), .B1(n4495), .B2(n5614), .ZN(n5617)
         );
  INV_X1 U6604 ( .A(n5617), .ZN(n5618) );
  NAND3_X1 U6605 ( .A1(n5620), .A2(n5619), .A3(n5618), .ZN(n5621) );
  AOI21_X1 U6606 ( .B1(n5773), .B2(n5622), .A(n5621), .ZN(n5623) );
  OAI211_X1 U6607 ( .C1(n5626), .C2(n5625), .A(n5624), .B(n5623), .ZN(U2826)
         );
  AOI22_X1 U6608 ( .A1(n5627), .A2(n5634), .B1(n5633), .B2(DATAI_18_), .ZN(
        n5629) );
  AOI22_X1 U6609 ( .A1(n5637), .A2(DATAI_2_), .B1(n5636), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U6610 ( .A1(n5629), .A2(n5628), .ZN(U2873) );
  AOI22_X1 U6611 ( .A1(n5630), .A2(n5634), .B1(n5633), .B2(DATAI_17_), .ZN(
        n5632) );
  AOI22_X1 U6612 ( .A1(n5637), .A2(DATAI_1_), .B1(n5636), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6613 ( .A1(n5632), .A2(n5631), .ZN(U2874) );
  AOI22_X1 U6614 ( .A1(n5635), .A2(n5634), .B1(n5633), .B2(DATAI_16_), .ZN(
        n5639) );
  AOI22_X1 U6615 ( .A1(n5637), .A2(DATAI_0_), .B1(n5636), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6616 ( .A1(n5639), .A2(n5638), .ZN(U2875) );
  INV_X1 U6617 ( .A(n5640), .ZN(n5643) );
  AOI22_X1 U6618 ( .A1(n5669), .A2(DATAO_REG_24__SCAN_IN), .B1(n5643), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5641) );
  OAI21_X1 U6619 ( .B1(n6538), .B2(n5672), .A(n5641), .ZN(U2899) );
  INV_X1 U6620 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6545) );
  AOI22_X1 U6621 ( .A1(n5669), .A2(DATAO_REG_22__SCAN_IN), .B1(n5643), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5642) );
  OAI21_X1 U6622 ( .B1(n6545), .B2(n5672), .A(n5642), .ZN(U2901) );
  INV_X1 U6623 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6610) );
  AOI22_X1 U6624 ( .A1(n5669), .A2(DATAO_REG_20__SCAN_IN), .B1(n5643), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5644) );
  OAI21_X1 U6625 ( .B1(n6610), .B2(n5672), .A(n5644), .ZN(U2903) );
  INV_X1 U6626 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5738) );
  AOI22_X1 U6627 ( .A1(n5663), .A2(LWORD_REG_15__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5645) );
  OAI21_X1 U6628 ( .B1(n5738), .B2(n5667), .A(n5645), .ZN(U2908) );
  AOI22_X1 U6629 ( .A1(EAX_REG_14__SCAN_IN), .A2(n5670), .B1(n5669), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U6630 ( .B1(n6574), .B2(n5672), .A(n5646), .ZN(U2909) );
  INV_X1 U6631 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5734) );
  AOI22_X1 U6632 ( .A1(n5663), .A2(LWORD_REG_13__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5647) );
  OAI21_X1 U6633 ( .B1(n5734), .B2(n5667), .A(n5647), .ZN(U2910) );
  INV_X1 U6634 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5730) );
  AOI22_X1 U6635 ( .A1(n5663), .A2(LWORD_REG_12__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5648) );
  OAI21_X1 U6636 ( .B1(n5730), .B2(n5667), .A(n5648), .ZN(U2911) );
  INV_X1 U6637 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5650) );
  AOI22_X1 U6638 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n5663), .B1(n5669), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5649) );
  OAI21_X1 U6639 ( .B1(n5650), .B2(n5667), .A(n5649), .ZN(U2912) );
  INV_X1 U6640 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5726) );
  AOI22_X1 U6641 ( .A1(n5663), .A2(LWORD_REG_10__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U6642 ( .B1(n5726), .B2(n5667), .A(n5651), .ZN(U2913) );
  INV_X1 U6643 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5722) );
  AOI22_X1 U6644 ( .A1(n5663), .A2(LWORD_REG_9__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5652) );
  OAI21_X1 U6645 ( .B1(n5722), .B2(n5667), .A(n5652), .ZN(U2914) );
  INV_X1 U6646 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6513) );
  INV_X1 U6647 ( .A(n5669), .ZN(n5654) );
  AOI22_X1 U6648 ( .A1(EAX_REG_8__SCAN_IN), .A2(n5670), .B1(n5663), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5653) );
  OAI21_X1 U6649 ( .B1(n6513), .B2(n5654), .A(n5653), .ZN(U2915) );
  AOI22_X1 U6650 ( .A1(n5663), .A2(LWORD_REG_7__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5655) );
  OAI21_X1 U6651 ( .B1(n3468), .B2(n5667), .A(n5655), .ZN(U2916) );
  AOI22_X1 U6652 ( .A1(n5663), .A2(LWORD_REG_6__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5656) );
  OAI21_X1 U6653 ( .B1(n6499), .B2(n5667), .A(n5656), .ZN(U2917) );
  AOI22_X1 U6654 ( .A1(n5663), .A2(LWORD_REG_5__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5657) );
  OAI21_X1 U6655 ( .B1(n5658), .B2(n5667), .A(n5657), .ZN(U2918) );
  AOI22_X1 U6656 ( .A1(n5663), .A2(LWORD_REG_4__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U6657 ( .B1(n5660), .B2(n5667), .A(n5659), .ZN(U2919) );
  AOI22_X1 U6658 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n5663), .B1(n5669), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5661) );
  OAI21_X1 U6659 ( .B1(n5662), .B2(n5667), .A(n5661), .ZN(U2920) );
  AOI22_X1 U6660 ( .A1(n5663), .A2(LWORD_REG_2__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5664) );
  OAI21_X1 U6661 ( .B1(n5665), .B2(n5667), .A(n5664), .ZN(U2921) );
  AOI22_X1 U6662 ( .A1(n5663), .A2(LWORD_REG_1__SCAN_IN), .B1(n5669), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5666) );
  OAI21_X1 U6663 ( .B1(n5668), .B2(n5667), .A(n5666), .ZN(U2922) );
  INV_X1 U6664 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6518) );
  AOI22_X1 U6665 ( .A1(EAX_REG_0__SCAN_IN), .A2(n5670), .B1(n5669), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5671) );
  OAI21_X1 U6666 ( .B1(n6518), .B2(n5672), .A(n5671), .ZN(U2923) );
  INV_X2 U6667 ( .A(n5673), .ZN(n6650) );
  AOI22_X1 U6668 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5674) );
  OAI21_X1 U6669 ( .B1(n6653), .B2(n5701), .A(n5674), .ZN(U2924) );
  AOI22_X1 U6670 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5675) );
  OAI21_X1 U6671 ( .B1(n5715), .B2(n5703), .A(n5675), .ZN(U2925) );
  AOI22_X1 U6672 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5676) );
  OAI21_X1 U6673 ( .B1(n6653), .B2(n5705), .A(n5676), .ZN(U2926) );
  AOI22_X1 U6674 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U6675 ( .B1(n5715), .B2(n5707), .A(n5677), .ZN(U2927) );
  AOI22_X1 U6676 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5678) );
  OAI21_X1 U6677 ( .B1(n6653), .B2(n6621), .A(n5678), .ZN(U2928) );
  AOI22_X1 U6678 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5679) );
  OAI21_X1 U6679 ( .B1(n6653), .B2(n5710), .A(n5679), .ZN(U2929) );
  AOI22_X1 U6680 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5680) );
  OAI21_X1 U6681 ( .B1(n5715), .B2(n5712), .A(n5680), .ZN(U2930) );
  AOI22_X1 U6682 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5681) );
  OAI21_X1 U6683 ( .B1(n6653), .B2(n5714), .A(n5681), .ZN(U2931) );
  INV_X1 U6684 ( .A(DATAI_9_), .ZN(n5682) );
  NOR2_X1 U6685 ( .A1(n6653), .A2(n5682), .ZN(n5720) );
  AOI21_X1 U6686 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6650), .A(n5720), .ZN(n5683) );
  OAI21_X1 U6687 ( .B1(n3773), .B2(n5737), .A(n5683), .ZN(U2933) );
  INV_X1 U6688 ( .A(DATAI_10_), .ZN(n5684) );
  OR2_X1 U6689 ( .A1(n6653), .A2(n5684), .ZN(n5724) );
  NAND2_X1 U6690 ( .A1(n6650), .A2(UWORD_REG_10__SCAN_IN), .ZN(n5685) );
  AND2_X1 U6691 ( .A1(n5724), .A2(n5685), .ZN(n5686) );
  OAI21_X1 U6692 ( .B1(n5687), .B2(n5737), .A(n5686), .ZN(U2934) );
  INV_X1 U6693 ( .A(DATAI_11_), .ZN(n6652) );
  AOI22_X1 U6694 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5688) );
  OAI21_X1 U6695 ( .B1(n6653), .B2(n6652), .A(n5688), .ZN(U2935) );
  INV_X1 U6696 ( .A(DATAI_12_), .ZN(n5689) );
  OR2_X1 U6697 ( .A1(n6653), .A2(n5689), .ZN(n5728) );
  NAND2_X1 U6698 ( .A1(n6650), .A2(UWORD_REG_12__SCAN_IN), .ZN(n5690) );
  AND2_X1 U6699 ( .A1(n5728), .A2(n5690), .ZN(n5691) );
  OAI21_X1 U6700 ( .B1(n5692), .B2(n5737), .A(n5691), .ZN(U2936) );
  INV_X1 U6701 ( .A(DATAI_13_), .ZN(n5693) );
  OR2_X1 U6702 ( .A1(n6653), .A2(n5693), .ZN(n5732) );
  NAND2_X1 U6703 ( .A1(n6650), .A2(UWORD_REG_13__SCAN_IN), .ZN(n5694) );
  AND2_X1 U6704 ( .A1(n5732), .A2(n5694), .ZN(n5695) );
  OAI21_X1 U6705 ( .B1(n3853), .B2(n5737), .A(n5695), .ZN(U2937) );
  NAND2_X1 U6706 ( .A1(n6650), .A2(UWORD_REG_14__SCAN_IN), .ZN(n5696) );
  AND2_X1 U6707 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  OAI21_X1 U6708 ( .B1(n5699), .B2(n5737), .A(n5698), .ZN(U2938) );
  AOI22_X1 U6709 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n5700) );
  OAI21_X1 U6710 ( .B1(n6653), .B2(n5701), .A(n5700), .ZN(U2939) );
  AOI22_X1 U6711 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U6712 ( .B1(n6653), .B2(n5703), .A(n5702), .ZN(U2940) );
  AOI22_X1 U6713 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n5704) );
  OAI21_X1 U6714 ( .B1(n6653), .B2(n5705), .A(n5704), .ZN(U2941) );
  AOI22_X1 U6715 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n5706) );
  OAI21_X1 U6716 ( .B1(n5715), .B2(n5707), .A(n5706), .ZN(U2942) );
  AOI22_X1 U6717 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n5708) );
  OAI21_X1 U6718 ( .B1(n5715), .B2(n6621), .A(n5708), .ZN(U2943) );
  AOI22_X1 U6719 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n5709) );
  OAI21_X1 U6720 ( .B1(n6653), .B2(n5710), .A(n5709), .ZN(U2944) );
  AOI22_X1 U6721 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n5711) );
  OAI21_X1 U6722 ( .B1(n5715), .B2(n5712), .A(n5711), .ZN(U2945) );
  AOI22_X1 U6723 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5713) );
  OAI21_X1 U6724 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(U2946) );
  INV_X1 U6725 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6726 ( .A1(n6650), .A2(LWORD_REG_8__SCAN_IN), .ZN(n5716) );
  AND2_X1 U6727 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  OAI21_X1 U6728 ( .B1(n5719), .B2(n5737), .A(n5718), .ZN(U2947) );
  AOI21_X1 U6729 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6650), .A(n5720), .ZN(n5721) );
  OAI21_X1 U6730 ( .B1(n5722), .B2(n5737), .A(n5721), .ZN(U2948) );
  NAND2_X1 U6731 ( .A1(n6650), .A2(LWORD_REG_10__SCAN_IN), .ZN(n5723) );
  AND2_X1 U6732 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  OAI21_X1 U6733 ( .B1(n5726), .B2(n5737), .A(n5725), .ZN(U2949) );
  NAND2_X1 U6734 ( .A1(n6650), .A2(LWORD_REG_12__SCAN_IN), .ZN(n5727) );
  AND2_X1 U6735 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  OAI21_X1 U6736 ( .B1(n5730), .B2(n5737), .A(n5729), .ZN(U2951) );
  NAND2_X1 U6737 ( .A1(n6650), .A2(LWORD_REG_13__SCAN_IN), .ZN(n5731) );
  AND2_X1 U6738 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  OAI21_X1 U6739 ( .B1(n5734), .B2(n5737), .A(n5733), .ZN(U2952) );
  AOI22_X1 U6740 ( .A1(n5735), .A2(DATAI_15_), .B1(LWORD_REG_15__SCAN_IN), 
        .B2(n6650), .ZN(n5736) );
  OAI21_X1 U6741 ( .B1(n5738), .B2(n5737), .A(n5736), .ZN(U2954) );
  NAND2_X1 U6742 ( .A1(n5740), .A2(n5739), .ZN(n5742) );
  XOR2_X1 U6743 ( .A(n5742), .B(n5741), .Z(n5795) );
  AOI22_X1 U6744 ( .A1(n5817), .A2(REIP_REG_11__SCAN_IN), .B1(n5771), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5746) );
  AOI22_X1 U6745 ( .A1(n5744), .A2(n5774), .B1(n5754), .B2(n5743), .ZN(n5745)
         );
  OAI211_X1 U6746 ( .C1(n5795), .C2(n5766), .A(n5746), .B(n5745), .ZN(U2975)
         );
  INV_X1 U6747 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5753) );
  INV_X1 U6748 ( .A(n5747), .ZN(n5748) );
  AOI222_X1 U6749 ( .A1(n5750), .A2(n5785), .B1(n5774), .B2(n5749), .C1(n5748), 
        .C2(n5754), .ZN(n5752) );
  OAI211_X1 U6750 ( .C1(n5753), .C2(n5782), .A(n5752), .B(n5751), .ZN(U2979)
         );
  AOI222_X1 U6751 ( .A1(n5757), .A2(n5785), .B1(n5756), .B2(n5774), .C1(n5755), 
        .C2(n5754), .ZN(n5759) );
  OAI211_X1 U6752 ( .C1(n5760), .C2(n5782), .A(n5759), .B(n5758), .ZN(U2981)
         );
  AOI22_X1 U6753 ( .A1(n5817), .A2(REIP_REG_2__SCAN_IN), .B1(n5771), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6754 ( .A1(n5762), .A2(n5761), .ZN(n5764) );
  XNOR2_X1 U6755 ( .A(n5764), .B(n5763), .ZN(n5826) );
  OAI22_X1 U6756 ( .A1(n5826), .A2(n5766), .B1(n5765), .B2(n6282), .ZN(n5767)
         );
  INV_X1 U6757 ( .A(n5767), .ZN(n5768) );
  OAI211_X1 U6758 ( .C1(n5777), .C2(n5770), .A(n5769), .B(n5768), .ZN(U2984)
         );
  AOI22_X1 U6759 ( .A1(n5817), .A2(REIP_REG_1__SCAN_IN), .B1(n5771), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5776) );
  AOI22_X1 U6760 ( .A1(n5774), .A2(n5773), .B1(n5772), .B2(n5785), .ZN(n5775)
         );
  OAI211_X1 U6761 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5777), .A(n5776), 
        .B(n5775), .ZN(U2985) );
  INV_X1 U6762 ( .A(n5778), .ZN(n5781) );
  AOI21_X1 U6763 ( .B1(n5781), .B2(n5780), .A(n5779), .ZN(n5838) );
  NAND2_X1 U6764 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  AOI22_X1 U6765 ( .A1(n5785), .A2(n5838), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5784), .ZN(n5787) );
  NAND2_X1 U6766 ( .A1(n5817), .A2(REIP_REG_0__SCAN_IN), .ZN(n5786) );
  OAI211_X1 U6767 ( .C1(n5788), .C2(n6282), .A(n5787), .B(n5786), .ZN(U2986)
         );
  AOI22_X1 U6768 ( .A1(n5836), .A2(n5789), .B1(n5817), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5794) );
  AOI22_X1 U6769 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5792), .B1(n5791), .B2(n5790), .ZN(n5793) );
  OAI211_X1 U6770 ( .C1(n5795), .C2(n5825), .A(n5794), .B(n5793), .ZN(U3007)
         );
  AOI21_X1 U6771 ( .B1(n5803), .B2(n5797), .A(n5796), .ZN(n5816) );
  OAI22_X1 U6772 ( .A1(n5799), .A2(n5798), .B1(n4729), .B2(n5845), .ZN(n5800)
         );
  AOI21_X1 U6773 ( .B1(n5801), .B2(n5837), .A(n5800), .ZN(n5806) );
  NOR2_X1 U6774 ( .A1(n5803), .A2(n5802), .ZN(n5811) );
  OAI211_X1 U6775 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5811), .B(n5804), .ZN(n5805) );
  OAI211_X1 U6776 ( .C1(n5816), .C2(n5807), .A(n5806), .B(n5805), .ZN(U3008)
         );
  INV_X1 U6777 ( .A(n5808), .ZN(n5809) );
  AOI21_X1 U6778 ( .B1(n5836), .B2(n5810), .A(n5809), .ZN(n5814) );
  AOI22_X1 U6779 ( .A1(n5812), .A2(n5837), .B1(n5811), .B2(n5815), .ZN(n5813)
         );
  OAI211_X1 U6780 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5813), .ZN(U3009)
         );
  AOI22_X1 U6781 ( .A1(n5818), .A2(n5836), .B1(n5817), .B2(REIP_REG_2__SCAN_IN), .ZN(n5834) );
  INV_X1 U6782 ( .A(n5819), .ZN(n5820) );
  NOR2_X1 U6783 ( .A1(n5821), .A2(n5820), .ZN(n5824) );
  INV_X1 U6784 ( .A(n5822), .ZN(n5823) );
  MUX2_X1 U6785 ( .A(n5824), .B(n5823), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n5828) );
  NOR2_X1 U6786 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  NOR2_X1 U6787 ( .A1(n5828), .A2(n5827), .ZN(n5833) );
  NAND3_X1 U6788 ( .A1(n5830), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5829), 
        .ZN(n5831) );
  NAND4_X1 U6789 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(U3016)
         );
  INV_X1 U6790 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6527) );
  AOI22_X1 U6791 ( .A1(n5838), .A2(n5837), .B1(n5836), .B2(n5835), .ZN(n5844)
         );
  INV_X1 U6792 ( .A(n5839), .ZN(n5842) );
  OAI22_X1 U6793 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5842), .B1(n5841), 
        .B2(n5840), .ZN(n5843) );
  OAI211_X1 U6794 ( .C1(n6527), .C2(n5845), .A(n5844), .B(n5843), .ZN(U3018)
         );
  NOR2_X1 U6795 ( .A1(n5847), .A2(n5846), .ZN(U3019) );
  NAND3_X1 U6796 ( .A1(n6358), .A2(n6558), .A3(n6354), .ZN(n5882) );
  NOR2_X1 U6797 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5882), .ZN(n5869)
         );
  NAND2_X1 U6798 ( .A1(n2981), .A2(n4495), .ZN(n6053) );
  NOR2_X1 U6799 ( .A1(n2980), .A2(n6053), .ZN(n5878) );
  INV_X1 U6800 ( .A(n5878), .ZN(n5849) );
  INV_X1 U6801 ( .A(n6105), .ZN(n6172) );
  OAI22_X1 U6802 ( .A1(n5849), .A2(n6278), .B1(n6172), .B2(n5848), .ZN(n5870)
         );
  AOI22_X1 U6803 ( .A1(n6280), .A2(n5869), .B1(n6279), .B2(n5870), .ZN(n5856)
         );
  NAND2_X1 U6804 ( .A1(n5879), .A2(n6163), .ZN(n5911) );
  NOR3_X1 U6805 ( .A1(n5871), .A2(n6336), .A3(n6278), .ZN(n5850) );
  NOR2_X1 U6806 ( .A1(n5850), .A2(n6286), .ZN(n5854) );
  INV_X1 U6807 ( .A(n5869), .ZN(n5852) );
  AOI211_X1 U6808 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5852), .A(n6228), .B(
        n5851), .ZN(n5853) );
  AOI22_X1 U6809 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5872), .B1(n6292), 
        .B2(n5871), .ZN(n5855) );
  OAI211_X1 U6810 ( .C1(n6295), .C2(n5875), .A(n5856), .B(n5855), .ZN(U3020)
         );
  AOI22_X1 U6811 ( .A1(n6297), .A2(n5869), .B1(n6296), .B2(n5870), .ZN(n5858)
         );
  AOI22_X1 U6812 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5872), .B1(n6298), 
        .B2(n5871), .ZN(n5857) );
  OAI211_X1 U6813 ( .C1(n6301), .C2(n5875), .A(n5858), .B(n5857), .ZN(U3021)
         );
  AOI22_X1 U6814 ( .A1(n6303), .A2(n5869), .B1(n6302), .B2(n5870), .ZN(n5860)
         );
  AOI22_X1 U6815 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5872), .B1(n6304), 
        .B2(n5871), .ZN(n5859) );
  OAI211_X1 U6816 ( .C1(n6307), .C2(n5875), .A(n5860), .B(n5859), .ZN(U3022)
         );
  AOI22_X1 U6817 ( .A1(n6309), .A2(n5869), .B1(n6308), .B2(n5870), .ZN(n5862)
         );
  AOI22_X1 U6818 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5872), .B1(n6310), 
        .B2(n5871), .ZN(n5861) );
  OAI211_X1 U6819 ( .C1(n6313), .C2(n5875), .A(n5862), .B(n5861), .ZN(U3023)
         );
  AOI22_X1 U6820 ( .A1(n6315), .A2(n5869), .B1(n6314), .B2(n5870), .ZN(n5864)
         );
  INV_X1 U6821 ( .A(n6259), .ZN(n6316) );
  AOI22_X1 U6822 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5872), .B1(n6316), 
        .B2(n5871), .ZN(n5863) );
  OAI211_X1 U6823 ( .C1(n6319), .C2(n5875), .A(n5864), .B(n5863), .ZN(U3024)
         );
  AOI22_X1 U6824 ( .A1(n6321), .A2(n5869), .B1(n6320), .B2(n5870), .ZN(n5866)
         );
  AOI22_X1 U6825 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5872), .B1(n6322), 
        .B2(n5871), .ZN(n5865) );
  OAI211_X1 U6826 ( .C1(n6325), .C2(n5875), .A(n5866), .B(n5865), .ZN(U3025)
         );
  AOI22_X1 U6827 ( .A1(n6327), .A2(n5869), .B1(n6326), .B2(n5870), .ZN(n5868)
         );
  AOI22_X1 U6828 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5872), .B1(n6328), 
        .B2(n5871), .ZN(n5867) );
  OAI211_X1 U6829 ( .C1(n6331), .C2(n5875), .A(n5868), .B(n5867), .ZN(U3026)
         );
  AOI22_X1 U6830 ( .A1(n6335), .A2(n5870), .B1(n6333), .B2(n5869), .ZN(n5874)
         );
  AOI22_X1 U6831 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5872), .B1(n6337), 
        .B2(n5871), .ZN(n5873) );
  OAI211_X1 U6832 ( .C1(n6342), .C2(n5875), .A(n5874), .B(n5873), .ZN(U3027)
         );
  INV_X1 U6833 ( .A(n6280), .ZN(n6050) );
  NOR2_X1 U6834 ( .A1(n6347), .A2(n5882), .ZN(n5877) );
  INV_X1 U6835 ( .A(n5877), .ZN(n5905) );
  OAI22_X1 U6836 ( .A1(n5911), .A2(n6295), .B1(n6050), .B2(n5905), .ZN(n5876)
         );
  INV_X1 U6837 ( .A(n5876), .ZN(n5886) );
  AOI21_X1 U6838 ( .B1(n5878), .B2(n6052), .A(n5877), .ZN(n5883) );
  AOI21_X1 U6839 ( .B1(n5879), .B2(STATEBS16_REG_SCAN_IN), .A(n6278), .ZN(
        n5881) );
  AOI22_X1 U6840 ( .A1(n5883), .A2(n5881), .B1(n6278), .B2(n5882), .ZN(n5880)
         );
  NAND2_X1 U6841 ( .A1(n6289), .A2(n5880), .ZN(n5908) );
  INV_X1 U6842 ( .A(n5881), .ZN(n5884) );
  OAI22_X1 U6843 ( .A1(n5884), .A2(n5883), .B1(n3391), .B2(n5882), .ZN(n5907)
         );
  AOI22_X1 U6844 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5908), .B1(n6279), 
        .B2(n5907), .ZN(n5885) );
  OAI211_X1 U6845 ( .C1(n5939), .C2(n6243), .A(n5886), .B(n5885), .ZN(U3028)
         );
  INV_X1 U6846 ( .A(n6297), .ZN(n6064) );
  OAI22_X1 U6847 ( .A1(n5939), .A2(n6247), .B1(n6064), .B2(n5905), .ZN(n5887)
         );
  INV_X1 U6848 ( .A(n5887), .ZN(n5889) );
  AOI22_X1 U6849 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5908), .B1(n6296), 
        .B2(n5907), .ZN(n5888) );
  OAI211_X1 U6850 ( .C1(n6301), .C2(n5911), .A(n5889), .B(n5888), .ZN(U3029)
         );
  OAI22_X1 U6851 ( .A1(n5911), .A2(n6307), .B1(n6068), .B2(n5905), .ZN(n5890)
         );
  INV_X1 U6852 ( .A(n5890), .ZN(n5892) );
  AOI22_X1 U6853 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5908), .B1(n6302), 
        .B2(n5907), .ZN(n5891) );
  OAI211_X1 U6854 ( .C1(n5939), .C2(n6251), .A(n5892), .B(n5891), .ZN(U3030)
         );
  INV_X1 U6855 ( .A(n6309), .ZN(n6072) );
  OAI22_X1 U6856 ( .A1(n5939), .A2(n6255), .B1(n6072), .B2(n5905), .ZN(n5893)
         );
  INV_X1 U6857 ( .A(n5893), .ZN(n5895) );
  AOI22_X1 U6858 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5908), .B1(n6308), 
        .B2(n5907), .ZN(n5894) );
  OAI211_X1 U6859 ( .C1(n6313), .C2(n5911), .A(n5895), .B(n5894), .ZN(U3031)
         );
  INV_X1 U6860 ( .A(n6315), .ZN(n6076) );
  OAI22_X1 U6861 ( .A1(n5939), .A2(n6259), .B1(n6076), .B2(n5905), .ZN(n5896)
         );
  INV_X1 U6862 ( .A(n5896), .ZN(n5898) );
  AOI22_X1 U6863 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5908), .B1(n6314), 
        .B2(n5907), .ZN(n5897) );
  OAI211_X1 U6864 ( .C1(n6319), .C2(n5911), .A(n5898), .B(n5897), .ZN(U3032)
         );
  INV_X1 U6865 ( .A(n6321), .ZN(n6080) );
  OAI22_X1 U6866 ( .A1(n5939), .A2(n6263), .B1(n6080), .B2(n5905), .ZN(n5899)
         );
  INV_X1 U6867 ( .A(n5899), .ZN(n5901) );
  AOI22_X1 U6868 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5908), .B1(n6320), 
        .B2(n5907), .ZN(n5900) );
  OAI211_X1 U6869 ( .C1(n6325), .C2(n5911), .A(n5901), .B(n5900), .ZN(U3033)
         );
  OAI22_X1 U6870 ( .A1(n5911), .A2(n6331), .B1(n6084), .B2(n5905), .ZN(n5902)
         );
  INV_X1 U6871 ( .A(n5902), .ZN(n5904) );
  AOI22_X1 U6872 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5908), .B1(n6326), 
        .B2(n5907), .ZN(n5903) );
  OAI211_X1 U6873 ( .C1(n5939), .C2(n6267), .A(n5904), .B(n5903), .ZN(U3034)
         );
  INV_X1 U6874 ( .A(n6333), .ZN(n6089) );
  OAI22_X1 U6875 ( .A1(n5939), .A2(n6275), .B1(n6089), .B2(n5905), .ZN(n5906)
         );
  INV_X1 U6876 ( .A(n5906), .ZN(n5910) );
  AOI22_X1 U6877 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5908), .B1(n6335), 
        .B2(n5907), .ZN(n5909) );
  OAI211_X1 U6878 ( .C1(n6342), .C2(n5911), .A(n5910), .B(n5909), .ZN(U3035)
         );
  NOR2_X1 U6879 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5912), .ZN(n5934)
         );
  INV_X1 U6880 ( .A(n5913), .ZN(n5916) );
  NAND3_X1 U6881 ( .A1(n6105), .A2(n6227), .A3(n6358), .ZN(n5914) );
  OAI21_X1 U6882 ( .B1(n5916), .B2(n6278), .A(n5914), .ZN(n5935) );
  AOI22_X1 U6883 ( .A1(n6280), .A2(n5934), .B1(n6279), .B2(n5935), .ZN(n5921)
         );
  INV_X1 U6884 ( .A(n5939), .ZN(n5915) );
  INV_X1 U6885 ( .A(n6286), .ZN(n6022) );
  OAI21_X1 U6886 ( .B1(n5915), .B2(n5943), .A(n6022), .ZN(n5917) );
  AOI21_X1 U6887 ( .B1(n5917), .B2(n5916), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5919) );
  OAI21_X1 U6888 ( .B1(n6227), .B2(n3391), .A(n5918), .ZN(n5958) );
  NOR2_X1 U6889 ( .A1(n6228), .A2(n5958), .ZN(n6103) );
  AOI22_X1 U6890 ( .A1(n5936), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5943), 
        .B2(n6292), .ZN(n5920) );
  OAI211_X1 U6891 ( .C1(n6295), .C2(n5939), .A(n5921), .B(n5920), .ZN(U3036)
         );
  AOI22_X1 U6892 ( .A1(n6297), .A2(n5934), .B1(n6296), .B2(n5935), .ZN(n5923)
         );
  AOI22_X1 U6893 ( .A1(n5936), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5943), 
        .B2(n6298), .ZN(n5922) );
  OAI211_X1 U6894 ( .C1(n5939), .C2(n6301), .A(n5923), .B(n5922), .ZN(U3037)
         );
  AOI22_X1 U6895 ( .A1(n6303), .A2(n5934), .B1(n6302), .B2(n5935), .ZN(n5925)
         );
  AOI22_X1 U6896 ( .A1(n5936), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5943), 
        .B2(n6304), .ZN(n5924) );
  OAI211_X1 U6897 ( .C1(n5939), .C2(n6307), .A(n5925), .B(n5924), .ZN(U3038)
         );
  AOI22_X1 U6898 ( .A1(n6309), .A2(n5934), .B1(n6308), .B2(n5935), .ZN(n5927)
         );
  AOI22_X1 U6899 ( .A1(n5936), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5943), 
        .B2(n6310), .ZN(n5926) );
  OAI211_X1 U6900 ( .C1(n5939), .C2(n6313), .A(n5927), .B(n5926), .ZN(U3039)
         );
  AOI22_X1 U6901 ( .A1(n6315), .A2(n5934), .B1(n6314), .B2(n5935), .ZN(n5929)
         );
  AOI22_X1 U6902 ( .A1(n5936), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5943), 
        .B2(n6316), .ZN(n5928) );
  OAI211_X1 U6903 ( .C1(n5939), .C2(n6319), .A(n5929), .B(n5928), .ZN(U3040)
         );
  AOI22_X1 U6904 ( .A1(n6321), .A2(n5934), .B1(n6320), .B2(n5935), .ZN(n5931)
         );
  AOI22_X1 U6905 ( .A1(n5936), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5943), 
        .B2(n6322), .ZN(n5930) );
  OAI211_X1 U6906 ( .C1(n5939), .C2(n6325), .A(n5931), .B(n5930), .ZN(U3041)
         );
  AOI22_X1 U6907 ( .A1(n6327), .A2(n5934), .B1(n6326), .B2(n5935), .ZN(n5933)
         );
  AOI22_X1 U6908 ( .A1(n5936), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5943), 
        .B2(n6328), .ZN(n5932) );
  OAI211_X1 U6909 ( .C1(n5939), .C2(n6331), .A(n5933), .B(n5932), .ZN(U3042)
         );
  AOI22_X1 U6910 ( .A1(n6335), .A2(n5935), .B1(n6333), .B2(n5934), .ZN(n5938)
         );
  AOI22_X1 U6911 ( .A1(n5936), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5943), 
        .B2(n6337), .ZN(n5937) );
  OAI211_X1 U6912 ( .C1(n5939), .C2(n6342), .A(n5938), .B(n5937), .ZN(U3043)
         );
  AOI22_X1 U6913 ( .A1(n5943), .A2(n6248), .B1(n6303), .B2(n5942), .ZN(n5941)
         );
  AOI22_X1 U6914 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5945), .B1(n6302), 
        .B2(n5944), .ZN(n5940) );
  OAI211_X1 U6915 ( .C1(n6251), .C2(n5954), .A(n5941), .B(n5940), .ZN(U3046)
         );
  AOI22_X1 U6916 ( .A1(n5943), .A2(n6264), .B1(n6327), .B2(n5942), .ZN(n5947)
         );
  AOI22_X1 U6917 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5945), .B1(n6326), 
        .B2(n5944), .ZN(n5946) );
  OAI211_X1 U6918 ( .C1(n6267), .C2(n5954), .A(n5947), .B(n5946), .ZN(U3050)
         );
  AOI22_X1 U6919 ( .A1(n6315), .A2(n5949), .B1(n6314), .B2(n5948), .ZN(n5953)
         );
  AOI22_X1 U6920 ( .A1(n5951), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6316), 
        .B2(n5950), .ZN(n5952) );
  OAI211_X1 U6921 ( .C1(n6319), .C2(n5954), .A(n5953), .B(n5952), .ZN(U3056)
         );
  INV_X1 U6922 ( .A(n6096), .ZN(n6226) );
  INV_X1 U6923 ( .A(n5993), .ZN(n5994) );
  NOR2_X1 U6924 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5994), .ZN(n5978)
         );
  NAND2_X1 U6925 ( .A1(n5956), .A2(n5955), .ZN(n6235) );
  INV_X1 U6926 ( .A(n6235), .ZN(n6277) );
  NAND2_X1 U6927 ( .A1(n6277), .A2(n6290), .ZN(n6231) );
  NAND3_X1 U6928 ( .A1(n6228), .A2(n6227), .A3(n6358), .ZN(n5957) );
  OAI21_X1 U6929 ( .B1(n6231), .B2(n2980), .A(n5957), .ZN(n5979) );
  AOI22_X1 U6930 ( .A1(n6280), .A2(n5978), .B1(n6279), .B2(n5979), .ZN(n5965)
         );
  AOI21_X1 U6931 ( .B1(n5963), .B2(n6011), .A(n6167), .ZN(n5962) );
  NAND2_X1 U6932 ( .A1(n6290), .A2(n6235), .ZN(n5961) );
  NOR2_X1 U6933 ( .A1(n6105), .A2(n5958), .ZN(n6238) );
  INV_X1 U6934 ( .A(n5978), .ZN(n5959) );
  AOI21_X1 U6935 ( .B1(n5959), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5960) );
  OAI211_X1 U6936 ( .C1(n5962), .C2(n5961), .A(n6238), .B(n5960), .ZN(n5981)
         );
  AOI22_X1 U6937 ( .A1(n5981), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6240), 
        .B2(n5980), .ZN(n5964) );
  OAI211_X1 U6938 ( .C1(n6243), .C2(n6011), .A(n5965), .B(n5964), .ZN(U3068)
         );
  AOI22_X1 U6939 ( .A1(n6297), .A2(n5978), .B1(n6296), .B2(n5979), .ZN(n5967)
         );
  AOI22_X1 U6940 ( .A1(n5981), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6244), 
        .B2(n5980), .ZN(n5966) );
  OAI211_X1 U6941 ( .C1(n6247), .C2(n6011), .A(n5967), .B(n5966), .ZN(U3069)
         );
  AOI22_X1 U6942 ( .A1(n6303), .A2(n5978), .B1(n6302), .B2(n5979), .ZN(n5969)
         );
  AOI22_X1 U6943 ( .A1(n5981), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6248), 
        .B2(n5980), .ZN(n5968) );
  OAI211_X1 U6944 ( .C1(n6251), .C2(n6011), .A(n5969), .B(n5968), .ZN(U3070)
         );
  AOI22_X1 U6945 ( .A1(n6309), .A2(n5978), .B1(n6308), .B2(n5979), .ZN(n5971)
         );
  AOI22_X1 U6946 ( .A1(n5981), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6252), 
        .B2(n5980), .ZN(n5970) );
  OAI211_X1 U6947 ( .C1(n6255), .C2(n6011), .A(n5971), .B(n5970), .ZN(U3071)
         );
  AOI22_X1 U6948 ( .A1(n6315), .A2(n5978), .B1(n6314), .B2(n5979), .ZN(n5973)
         );
  AOI22_X1 U6949 ( .A1(n5981), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6256), 
        .B2(n5980), .ZN(n5972) );
  OAI211_X1 U6950 ( .C1(n6259), .C2(n6011), .A(n5973), .B(n5972), .ZN(U3072)
         );
  AOI22_X1 U6951 ( .A1(n6321), .A2(n5978), .B1(n6320), .B2(n5979), .ZN(n5975)
         );
  AOI22_X1 U6952 ( .A1(n5981), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6260), 
        .B2(n5980), .ZN(n5974) );
  OAI211_X1 U6953 ( .C1(n6263), .C2(n6011), .A(n5975), .B(n5974), .ZN(U3073)
         );
  AOI22_X1 U6954 ( .A1(n6327), .A2(n5978), .B1(n6326), .B2(n5979), .ZN(n5977)
         );
  AOI22_X1 U6955 ( .A1(n5981), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6264), 
        .B2(n5980), .ZN(n5976) );
  OAI211_X1 U6956 ( .C1(n6267), .C2(n6011), .A(n5977), .B(n5976), .ZN(U3074)
         );
  AOI22_X1 U6957 ( .A1(n6335), .A2(n5979), .B1(n6333), .B2(n5978), .ZN(n5983)
         );
  AOI22_X1 U6958 ( .A1(n5981), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6271), 
        .B2(n5980), .ZN(n5982) );
  OAI211_X1 U6959 ( .C1(n6275), .C2(n6011), .A(n5983), .B(n5982), .ZN(U3075)
         );
  INV_X1 U6960 ( .A(n6128), .ZN(n5984) );
  INV_X1 U6961 ( .A(n5986), .ZN(n6012) );
  AOI22_X1 U6962 ( .A1(n6039), .A2(n6292), .B1(n6280), .B2(n6012), .ZN(n5998)
         );
  NAND2_X1 U6963 ( .A1(n5987), .A2(n6290), .ZN(n5996) );
  INV_X1 U6964 ( .A(n5996), .ZN(n5991) );
  NAND2_X1 U6965 ( .A1(n6052), .A2(n5988), .ZN(n5989) );
  OR2_X1 U6966 ( .A1(n6235), .A2(n5989), .ZN(n5990) );
  AND2_X1 U6967 ( .A1(n5990), .A2(n5986), .ZN(n5995) );
  NAND2_X1 U6968 ( .A1(n5991), .A2(n5995), .ZN(n5992) );
  OAI211_X1 U6969 ( .C1(n5993), .C2(n6290), .A(n6289), .B(n5992), .ZN(n6015)
         );
  OAI22_X1 U6970 ( .A1(n5996), .A2(n5995), .B1(n5994), .B2(n3391), .ZN(n6014)
         );
  AOI22_X1 U6971 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6015), .B1(n6279), 
        .B2(n6014), .ZN(n5997) );
  OAI211_X1 U6972 ( .C1(n6295), .C2(n6011), .A(n5998), .B(n5997), .ZN(U3076)
         );
  INV_X1 U6973 ( .A(n6011), .ZN(n6013) );
  AOI22_X1 U6974 ( .A1(n6013), .A2(n6244), .B1(n6297), .B2(n6012), .ZN(n6000)
         );
  AOI22_X1 U6975 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6015), .B1(n6296), 
        .B2(n6014), .ZN(n5999) );
  OAI211_X1 U6976 ( .C1(n6247), .C2(n6048), .A(n6000), .B(n5999), .ZN(U3077)
         );
  AOI22_X1 U6977 ( .A1(n6013), .A2(n6248), .B1(n6303), .B2(n6012), .ZN(n6002)
         );
  AOI22_X1 U6978 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6015), .B1(n6302), 
        .B2(n6014), .ZN(n6001) );
  OAI211_X1 U6979 ( .C1(n6251), .C2(n6048), .A(n6002), .B(n6001), .ZN(U3078)
         );
  AOI22_X1 U6980 ( .A1(n6013), .A2(n6252), .B1(n6309), .B2(n6012), .ZN(n6004)
         );
  AOI22_X1 U6981 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6015), .B1(n6308), 
        .B2(n6014), .ZN(n6003) );
  OAI211_X1 U6982 ( .C1(n6255), .C2(n6048), .A(n6004), .B(n6003), .ZN(U3079)
         );
  AOI22_X1 U6983 ( .A1(n6013), .A2(n6256), .B1(n6315), .B2(n6012), .ZN(n6006)
         );
  AOI22_X1 U6984 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6015), .B1(n6314), 
        .B2(n6014), .ZN(n6005) );
  OAI211_X1 U6985 ( .C1(n6259), .C2(n6048), .A(n6006), .B(n6005), .ZN(U3080)
         );
  AOI22_X1 U6986 ( .A1(n6039), .A2(n6322), .B1(n6321), .B2(n6012), .ZN(n6008)
         );
  AOI22_X1 U6987 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6015), .B1(n6320), 
        .B2(n6014), .ZN(n6007) );
  OAI211_X1 U6988 ( .C1(n6325), .C2(n6011), .A(n6008), .B(n6007), .ZN(U3081)
         );
  AOI22_X1 U6989 ( .A1(n6039), .A2(n6328), .B1(n6327), .B2(n6012), .ZN(n6010)
         );
  AOI22_X1 U6990 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6015), .B1(n6326), 
        .B2(n6014), .ZN(n6009) );
  OAI211_X1 U6991 ( .C1(n6331), .C2(n6011), .A(n6010), .B(n6009), .ZN(U3082)
         );
  AOI22_X1 U6992 ( .A1(n6013), .A2(n6271), .B1(n6333), .B2(n6012), .ZN(n6017)
         );
  AOI22_X1 U6993 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6015), .B1(n6335), 
        .B2(n6014), .ZN(n6016) );
  OAI211_X1 U6994 ( .C1(n6275), .C2(n6048), .A(n6017), .B(n6016), .ZN(U3083)
         );
  NAND3_X1 U6995 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6558), .A3(n6354), .ZN(n6059) );
  NOR2_X1 U6996 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6059), .ZN(n6042)
         );
  INV_X1 U6997 ( .A(n2980), .ZN(n6230) );
  NOR2_X1 U6998 ( .A1(n6230), .A2(n6053), .ZN(n6021) );
  INV_X1 U6999 ( .A(n6021), .ZN(n6020) );
  INV_X1 U7000 ( .A(n6227), .ZN(n6018) );
  NAND2_X1 U7001 ( .A1(n6019), .A2(n6018), .ZN(n6165) );
  OAI22_X1 U7002 ( .A1(n6020), .A2(n6278), .B1(n6172), .B2(n6165), .ZN(n6043)
         );
  AOI22_X1 U7003 ( .A1(n6280), .A2(n6042), .B1(n6279), .B2(n6043), .ZN(n6028)
         );
  NAND3_X1 U7004 ( .A1(n6090), .A2(n6290), .A3(n6048), .ZN(n6023) );
  AOI21_X1 U7005 ( .B1(n6023), .B2(n6022), .A(n6021), .ZN(n6026) );
  AOI21_X1 U7006 ( .B1(n6165), .B2(STATE2_REG_2__SCAN_IN), .A(n6024), .ZN(
        n6171) );
  OAI211_X1 U7007 ( .C1(n6466), .C2(n6042), .A(n6164), .B(n6171), .ZN(n6025)
         );
  AOI22_X1 U7008 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n6045), .B1(n6240), 
        .B2(n6039), .ZN(n6027) );
  OAI211_X1 U7009 ( .C1(n6243), .C2(n6090), .A(n6028), .B(n6027), .ZN(U3084)
         );
  AOI22_X1 U7010 ( .A1(n6297), .A2(n6042), .B1(n6296), .B2(n6043), .ZN(n6030)
         );
  AOI22_X1 U7011 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n6045), .B1(n6298), 
        .B2(n6044), .ZN(n6029) );
  OAI211_X1 U7012 ( .C1(n6301), .C2(n6048), .A(n6030), .B(n6029), .ZN(U3085)
         );
  AOI22_X1 U7013 ( .A1(n6303), .A2(n6042), .B1(n6302), .B2(n6043), .ZN(n6032)
         );
  AOI22_X1 U7014 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n6045), .B1(n6248), 
        .B2(n6039), .ZN(n6031) );
  OAI211_X1 U7015 ( .C1(n6251), .C2(n6090), .A(n6032), .B(n6031), .ZN(U3086)
         );
  AOI22_X1 U7016 ( .A1(n6309), .A2(n6042), .B1(n6308), .B2(n6043), .ZN(n6034)
         );
  AOI22_X1 U7017 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n6045), .B1(n6310), 
        .B2(n6044), .ZN(n6033) );
  OAI211_X1 U7018 ( .C1(n6313), .C2(n6048), .A(n6034), .B(n6033), .ZN(U3087)
         );
  AOI22_X1 U7019 ( .A1(n6315), .A2(n6042), .B1(n6314), .B2(n6043), .ZN(n6036)
         );
  AOI22_X1 U7020 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6045), .B1(n6316), 
        .B2(n6044), .ZN(n6035) );
  OAI211_X1 U7021 ( .C1(n6319), .C2(n6048), .A(n6036), .B(n6035), .ZN(U3088)
         );
  AOI22_X1 U7022 ( .A1(n6321), .A2(n6042), .B1(n6320), .B2(n6043), .ZN(n6038)
         );
  AOI22_X1 U7023 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n6045), .B1(n6322), 
        .B2(n6044), .ZN(n6037) );
  OAI211_X1 U7024 ( .C1(n6325), .C2(n6048), .A(n6038), .B(n6037), .ZN(U3089)
         );
  AOI22_X1 U7025 ( .A1(n6327), .A2(n6042), .B1(n6326), .B2(n6043), .ZN(n6041)
         );
  AOI22_X1 U7026 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n6045), .B1(n6264), 
        .B2(n6039), .ZN(n6040) );
  OAI211_X1 U7027 ( .C1(n6267), .C2(n6090), .A(n6041), .B(n6040), .ZN(U3090)
         );
  AOI22_X1 U7028 ( .A1(n6335), .A2(n6043), .B1(n6333), .B2(n6042), .ZN(n6047)
         );
  AOI22_X1 U7029 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n6045), .B1(n6337), 
        .B2(n6044), .ZN(n6046) );
  OAI211_X1 U7030 ( .C1(n6342), .C2(n6048), .A(n6047), .B(n6046), .ZN(U3091)
         );
  NOR2_X1 U7031 ( .A1(n6347), .A2(n6059), .ZN(n6054) );
  INV_X1 U7032 ( .A(n6054), .ZN(n6088) );
  OAI22_X1 U7033 ( .A1(n6090), .A2(n6295), .B1(n6050), .B2(n6088), .ZN(n6051)
         );
  INV_X1 U7034 ( .A(n6051), .ZN(n6063) );
  AND2_X1 U7035 ( .A1(n6052), .A2(n2980), .ZN(n6276) );
  INV_X1 U7036 ( .A(n6053), .ZN(n6055) );
  AOI21_X1 U7037 ( .B1(n6276), .B2(n6055), .A(n6054), .ZN(n6061) );
  OR3_X1 U7038 ( .A1(n6132), .A2(n6283), .A3(n6167), .ZN(n6056) );
  AOI22_X1 U7039 ( .A1(n6061), .A2(n6058), .B1(n6278), .B2(n6059), .ZN(n6057)
         );
  NAND2_X1 U7040 ( .A1(n6289), .A2(n6057), .ZN(n6093) );
  INV_X1 U7041 ( .A(n6058), .ZN(n6060) );
  OAI22_X1 U7042 ( .A1(n6061), .A2(n6060), .B1(n3391), .B2(n6059), .ZN(n6092)
         );
  AOI22_X1 U7043 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6093), .B1(n6279), 
        .B2(n6092), .ZN(n6062) );
  OAI211_X1 U7044 ( .C1(n6243), .C2(n6127), .A(n6063), .B(n6062), .ZN(U3092)
         );
  OAI22_X1 U7045 ( .A1(n6090), .A2(n6301), .B1(n6064), .B2(n6088), .ZN(n6065)
         );
  INV_X1 U7046 ( .A(n6065), .ZN(n6067) );
  AOI22_X1 U7047 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6093), .B1(n6296), 
        .B2(n6092), .ZN(n6066) );
  OAI211_X1 U7048 ( .C1(n6247), .C2(n6127), .A(n6067), .B(n6066), .ZN(U3093)
         );
  OAI22_X1 U7049 ( .A1(n6127), .A2(n6251), .B1(n6068), .B2(n6088), .ZN(n6069)
         );
  INV_X1 U7050 ( .A(n6069), .ZN(n6071) );
  AOI22_X1 U7051 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6093), .B1(n6302), 
        .B2(n6092), .ZN(n6070) );
  OAI211_X1 U7052 ( .C1(n6307), .C2(n6090), .A(n6071), .B(n6070), .ZN(U3094)
         );
  OAI22_X1 U7053 ( .A1(n6090), .A2(n6313), .B1(n6072), .B2(n6088), .ZN(n6073)
         );
  INV_X1 U7054 ( .A(n6073), .ZN(n6075) );
  AOI22_X1 U7055 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6093), .B1(n6308), 
        .B2(n6092), .ZN(n6074) );
  OAI211_X1 U7056 ( .C1(n6255), .C2(n6127), .A(n6075), .B(n6074), .ZN(U3095)
         );
  OAI22_X1 U7057 ( .A1(n6127), .A2(n6259), .B1(n6076), .B2(n6088), .ZN(n6077)
         );
  INV_X1 U7058 ( .A(n6077), .ZN(n6079) );
  AOI22_X1 U7059 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6093), .B1(n6314), 
        .B2(n6092), .ZN(n6078) );
  OAI211_X1 U7060 ( .C1(n6319), .C2(n6090), .A(n6079), .B(n6078), .ZN(U3096)
         );
  OAI22_X1 U7061 ( .A1(n6090), .A2(n6325), .B1(n6080), .B2(n6088), .ZN(n6081)
         );
  INV_X1 U7062 ( .A(n6081), .ZN(n6083) );
  AOI22_X1 U7063 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6093), .B1(n6320), 
        .B2(n6092), .ZN(n6082) );
  OAI211_X1 U7064 ( .C1(n6263), .C2(n6127), .A(n6083), .B(n6082), .ZN(U3097)
         );
  OAI22_X1 U7065 ( .A1(n6090), .A2(n6331), .B1(n6084), .B2(n6088), .ZN(n6085)
         );
  INV_X1 U7066 ( .A(n6085), .ZN(n6087) );
  AOI22_X1 U7067 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6093), .B1(n6326), 
        .B2(n6092), .ZN(n6086) );
  OAI211_X1 U7068 ( .C1(n6267), .C2(n6127), .A(n6087), .B(n6086), .ZN(U3098)
         );
  OAI22_X1 U7069 ( .A1(n6090), .A2(n6342), .B1(n6089), .B2(n6088), .ZN(n6091)
         );
  INV_X1 U7070 ( .A(n6091), .ZN(n6095) );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6093), .B1(n6335), 
        .B2(n6092), .ZN(n6094) );
  OAI211_X1 U7072 ( .C1(n6275), .C2(n6127), .A(n6095), .B(n6094), .ZN(U3099)
         );
  NAND2_X1 U7073 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6097), .ZN(n6139) );
  NOR2_X1 U7074 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6139), .ZN(n6122)
         );
  AOI22_X1 U7075 ( .A1(n6154), .A2(n6292), .B1(n6280), .B2(n6122), .ZN(n6109)
         );
  AOI21_X1 U7076 ( .B1(n6127), .B2(n6162), .A(n6167), .ZN(n6098) );
  NOR2_X1 U7077 ( .A1(n6098), .A2(n6278), .ZN(n6104) );
  INV_X1 U7078 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7079 ( .A1(n6100), .A2(n2980), .ZN(n6133) );
  INV_X1 U7080 ( .A(n6122), .ZN(n6101) );
  AOI22_X1 U7081 ( .A1(n6104), .A2(n6133), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6101), .ZN(n6102) );
  OAI211_X1 U7082 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n3391), .A(n6103), .B(n6102), .ZN(n6124) );
  INV_X1 U7083 ( .A(n6104), .ZN(n6107) );
  NAND3_X1 U7084 ( .A1(n6105), .A2(n6227), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6106) );
  AOI22_X1 U7085 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6124), .B1(n6279), 
        .B2(n6123), .ZN(n6108) );
  OAI211_X1 U7086 ( .C1(n6295), .C2(n6127), .A(n6109), .B(n6108), .ZN(U3100)
         );
  AOI22_X1 U7087 ( .A1(n6154), .A2(n6298), .B1(n6297), .B2(n6122), .ZN(n6111)
         );
  AOI22_X1 U7088 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6124), .B1(n6296), 
        .B2(n6123), .ZN(n6110) );
  OAI211_X1 U7089 ( .C1(n6301), .C2(n6127), .A(n6111), .B(n6110), .ZN(U3101)
         );
  AOI22_X1 U7090 ( .A1(n6154), .A2(n6304), .B1(n6303), .B2(n6122), .ZN(n6113)
         );
  AOI22_X1 U7091 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6124), .B1(n6302), 
        .B2(n6123), .ZN(n6112) );
  OAI211_X1 U7092 ( .C1(n6307), .C2(n6127), .A(n6113), .B(n6112), .ZN(U3102)
         );
  AOI22_X1 U7093 ( .A1(n6154), .A2(n6310), .B1(n6309), .B2(n6122), .ZN(n6115)
         );
  AOI22_X1 U7094 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6124), .B1(n6308), 
        .B2(n6123), .ZN(n6114) );
  OAI211_X1 U7095 ( .C1(n6313), .C2(n6127), .A(n6115), .B(n6114), .ZN(U3103)
         );
  AOI22_X1 U7096 ( .A1(n6154), .A2(n6316), .B1(n6315), .B2(n6122), .ZN(n6117)
         );
  AOI22_X1 U7097 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6124), .B1(n6314), 
        .B2(n6123), .ZN(n6116) );
  OAI211_X1 U7098 ( .C1(n6319), .C2(n6127), .A(n6117), .B(n6116), .ZN(U3104)
         );
  AOI22_X1 U7099 ( .A1(n6154), .A2(n6322), .B1(n6321), .B2(n6122), .ZN(n6119)
         );
  AOI22_X1 U7100 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6124), .B1(n6320), 
        .B2(n6123), .ZN(n6118) );
  OAI211_X1 U7101 ( .C1(n6325), .C2(n6127), .A(n6119), .B(n6118), .ZN(U3105)
         );
  AOI22_X1 U7102 ( .A1(n6154), .A2(n6328), .B1(n6327), .B2(n6122), .ZN(n6121)
         );
  AOI22_X1 U7103 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6124), .B1(n6326), 
        .B2(n6123), .ZN(n6120) );
  OAI211_X1 U7104 ( .C1(n6331), .C2(n6127), .A(n6121), .B(n6120), .ZN(U3106)
         );
  AOI22_X1 U7105 ( .A1(n6154), .A2(n6337), .B1(n6333), .B2(n6122), .ZN(n6126)
         );
  AOI22_X1 U7106 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6124), .B1(n6335), 
        .B2(n6123), .ZN(n6125) );
  OAI211_X1 U7107 ( .C1(n6342), .C2(n6127), .A(n6126), .B(n6125), .ZN(U3107)
         );
  INV_X1 U7108 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7109 ( .A1(n6130), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6134) );
  INV_X1 U7110 ( .A(n6134), .ZN(n6157) );
  AOI22_X1 U7111 ( .A1(n6191), .A2(n6292), .B1(n6280), .B2(n6157), .ZN(n6143)
         );
  OAI21_X1 U7112 ( .B1(n6132), .B2(n6131), .A(n6290), .ZN(n6141) );
  OR2_X1 U7113 ( .A1(n6133), .A2(n6345), .ZN(n6135) );
  NAND2_X1 U7114 ( .A1(n6135), .A2(n6134), .ZN(n6138) );
  AOI21_X1 U7115 ( .B1(n6139), .B2(n6278), .A(n6136), .ZN(n6137) );
  OAI21_X1 U7116 ( .B1(n6141), .B2(n6138), .A(n6137), .ZN(n6159) );
  INV_X1 U7117 ( .A(n6138), .ZN(n6140) );
  OAI22_X1 U7118 ( .A1(n6141), .A2(n6140), .B1(n6139), .B2(n3391), .ZN(n6158)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6159), .B1(n6279), 
        .B2(n6158), .ZN(n6142) );
  OAI211_X1 U7120 ( .C1(n6295), .C2(n6162), .A(n6143), .B(n6142), .ZN(U3108)
         );
  AOI22_X1 U7121 ( .A1(n6191), .A2(n6298), .B1(n6297), .B2(n6157), .ZN(n6145)
         );
  AOI22_X1 U7122 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6159), .B1(n6296), 
        .B2(n6158), .ZN(n6144) );
  OAI211_X1 U7123 ( .C1(n6301), .C2(n6162), .A(n6145), .B(n6144), .ZN(U3109)
         );
  AOI22_X1 U7124 ( .A1(n6154), .A2(n6248), .B1(n6303), .B2(n6157), .ZN(n6147)
         );
  AOI22_X1 U7125 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6159), .B1(n6302), 
        .B2(n6158), .ZN(n6146) );
  OAI211_X1 U7126 ( .C1(n6251), .C2(n6168), .A(n6147), .B(n6146), .ZN(U3110)
         );
  AOI22_X1 U7127 ( .A1(n6191), .A2(n6310), .B1(n6309), .B2(n6157), .ZN(n6149)
         );
  AOI22_X1 U7128 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6159), .B1(n6308), 
        .B2(n6158), .ZN(n6148) );
  OAI211_X1 U7129 ( .C1(n6313), .C2(n6162), .A(n6149), .B(n6148), .ZN(U3111)
         );
  AOI22_X1 U7130 ( .A1(n6191), .A2(n6316), .B1(n6315), .B2(n6157), .ZN(n6151)
         );
  AOI22_X1 U7131 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6159), .B1(n6314), 
        .B2(n6158), .ZN(n6150) );
  OAI211_X1 U7132 ( .C1(n6319), .C2(n6162), .A(n6151), .B(n6150), .ZN(U3112)
         );
  AOI22_X1 U7133 ( .A1(n6191), .A2(n6322), .B1(n6321), .B2(n6157), .ZN(n6153)
         );
  AOI22_X1 U7134 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6159), .B1(n6320), 
        .B2(n6158), .ZN(n6152) );
  OAI211_X1 U7135 ( .C1(n6325), .C2(n6162), .A(n6153), .B(n6152), .ZN(U3113)
         );
  AOI22_X1 U7136 ( .A1(n6154), .A2(n6264), .B1(n6327), .B2(n6157), .ZN(n6156)
         );
  AOI22_X1 U7137 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6159), .B1(n6326), 
        .B2(n6158), .ZN(n6155) );
  OAI211_X1 U7138 ( .C1(n6267), .C2(n6168), .A(n6156), .B(n6155), .ZN(U3114)
         );
  AOI22_X1 U7139 ( .A1(n6191), .A2(n6337), .B1(n6333), .B2(n6157), .ZN(n6161)
         );
  AOI22_X1 U7140 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6159), .B1(n6335), 
        .B2(n6158), .ZN(n6160) );
  OAI211_X1 U7141 ( .C1(n6342), .C2(n6162), .A(n6161), .B(n6160), .ZN(U3115)
         );
  NAND2_X1 U7142 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6196), .ZN(n6199) );
  NOR2_X1 U7143 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6199), .ZN(n6189)
         );
  OAI22_X1 U7144 ( .A1(n6166), .A2(n6230), .B1(n6165), .B2(n6164), .ZN(n6190)
         );
  AOI22_X1 U7145 ( .A1(n6280), .A2(n6189), .B1(n6279), .B2(n6190), .ZN(n6176)
         );
  AOI21_X1 U7146 ( .B1(n6224), .B2(n6168), .A(n6167), .ZN(n6169) );
  AOI211_X1 U7147 ( .C1(n6195), .C2(n6170), .A(n6278), .B(n6169), .ZN(n6174)
         );
  OAI211_X1 U7148 ( .C1(n6466), .C2(n6189), .A(n6172), .B(n6171), .ZN(n6173)
         );
  AOI22_X1 U7149 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6192), .B1(n6240), 
        .B2(n6191), .ZN(n6175) );
  OAI211_X1 U7150 ( .C1(n6243), .C2(n6224), .A(n6176), .B(n6175), .ZN(U3116)
         );
  AOI22_X1 U7151 ( .A1(n6297), .A2(n6189), .B1(n6296), .B2(n6190), .ZN(n6178)
         );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6192), .B1(n6244), 
        .B2(n6191), .ZN(n6177) );
  OAI211_X1 U7153 ( .C1(n6247), .C2(n6224), .A(n6178), .B(n6177), .ZN(U3117)
         );
  AOI22_X1 U7154 ( .A1(n6303), .A2(n6189), .B1(n6302), .B2(n6190), .ZN(n6180)
         );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6192), .B1(n6248), 
        .B2(n6191), .ZN(n6179) );
  OAI211_X1 U7156 ( .C1(n6251), .C2(n6224), .A(n6180), .B(n6179), .ZN(U3118)
         );
  AOI22_X1 U7157 ( .A1(n6309), .A2(n6189), .B1(n6308), .B2(n6190), .ZN(n6182)
         );
  AOI22_X1 U7158 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6192), .B1(n6252), 
        .B2(n6191), .ZN(n6181) );
  OAI211_X1 U7159 ( .C1(n6255), .C2(n6224), .A(n6182), .B(n6181), .ZN(U3119)
         );
  AOI22_X1 U7160 ( .A1(n6315), .A2(n6189), .B1(n6314), .B2(n6190), .ZN(n6184)
         );
  AOI22_X1 U7161 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6192), .B1(n6256), 
        .B2(n6191), .ZN(n6183) );
  OAI211_X1 U7162 ( .C1(n6259), .C2(n6224), .A(n6184), .B(n6183), .ZN(U3120)
         );
  AOI22_X1 U7163 ( .A1(n6321), .A2(n6189), .B1(n6320), .B2(n6190), .ZN(n6186)
         );
  AOI22_X1 U7164 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6192), .B1(n6260), 
        .B2(n6191), .ZN(n6185) );
  OAI211_X1 U7165 ( .C1(n6263), .C2(n6224), .A(n6186), .B(n6185), .ZN(U3121)
         );
  AOI22_X1 U7166 ( .A1(n6327), .A2(n6189), .B1(n6326), .B2(n6190), .ZN(n6188)
         );
  AOI22_X1 U7167 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6192), .B1(n6264), 
        .B2(n6191), .ZN(n6187) );
  OAI211_X1 U7168 ( .C1(n6267), .C2(n6224), .A(n6188), .B(n6187), .ZN(U3122)
         );
  AOI22_X1 U7169 ( .A1(n6335), .A2(n6190), .B1(n6333), .B2(n6189), .ZN(n6194)
         );
  AOI22_X1 U7170 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6192), .B1(n6271), 
        .B2(n6191), .ZN(n6193) );
  OAI211_X1 U7171 ( .C1(n6275), .C2(n6224), .A(n6194), .B(n6193), .ZN(U3123)
         );
  NOR2_X1 U7172 ( .A1(n6347), .A2(n6199), .ZN(n6219) );
  AOI21_X1 U7173 ( .B1(n6276), .B2(n6195), .A(n6219), .ZN(n6201) );
  NAND2_X1 U7174 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6198) );
  INV_X1 U7175 ( .A(n6196), .ZN(n6197) );
  OAI22_X1 U7176 ( .A1(n6201), .A2(n6278), .B1(n6198), .B2(n6197), .ZN(n6220)
         );
  AOI22_X1 U7177 ( .A1(n6280), .A2(n6219), .B1(n6279), .B2(n6220), .ZN(n6206)
         );
  INV_X1 U7178 ( .A(n6199), .ZN(n6203) );
  NAND2_X1 U7179 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  OAI221_X1 U7180 ( .B1(n6290), .B2(n6203), .C1(n6278), .C2(n6202), .A(n6289), 
        .ZN(n6221) );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6221), .B1(n6292), 
        .B2(n6270), .ZN(n6205) );
  OAI211_X1 U7182 ( .C1(n6295), .C2(n6224), .A(n6206), .B(n6205), .ZN(U3124)
         );
  AOI22_X1 U7183 ( .A1(n6297), .A2(n6219), .B1(n6296), .B2(n6220), .ZN(n6208)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6221), .B1(n6298), 
        .B2(n6270), .ZN(n6207) );
  OAI211_X1 U7185 ( .C1(n6301), .C2(n6224), .A(n6208), .B(n6207), .ZN(U3125)
         );
  AOI22_X1 U7186 ( .A1(n6303), .A2(n6219), .B1(n6302), .B2(n6220), .ZN(n6210)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6221), .B1(n6304), 
        .B2(n6270), .ZN(n6209) );
  OAI211_X1 U7188 ( .C1(n6307), .C2(n6224), .A(n6210), .B(n6209), .ZN(U3126)
         );
  AOI22_X1 U7189 ( .A1(n6309), .A2(n6219), .B1(n6308), .B2(n6220), .ZN(n6212)
         );
  AOI22_X1 U7190 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6221), .B1(n6310), 
        .B2(n6270), .ZN(n6211) );
  OAI211_X1 U7191 ( .C1(n6313), .C2(n6224), .A(n6212), .B(n6211), .ZN(U3127)
         );
  AOI22_X1 U7192 ( .A1(n6315), .A2(n6219), .B1(n6314), .B2(n6220), .ZN(n6214)
         );
  AOI22_X1 U7193 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6221), .B1(n6316), 
        .B2(n6270), .ZN(n6213) );
  OAI211_X1 U7194 ( .C1(n6319), .C2(n6224), .A(n6214), .B(n6213), .ZN(U3128)
         );
  AOI22_X1 U7195 ( .A1(n6321), .A2(n6219), .B1(n6320), .B2(n6220), .ZN(n6216)
         );
  AOI22_X1 U7196 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6221), .B1(n6322), 
        .B2(n6270), .ZN(n6215) );
  OAI211_X1 U7197 ( .C1(n6325), .C2(n6224), .A(n6216), .B(n6215), .ZN(U3129)
         );
  AOI22_X1 U7198 ( .A1(n6327), .A2(n6219), .B1(n6326), .B2(n6220), .ZN(n6218)
         );
  AOI22_X1 U7199 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6221), .B1(n6328), 
        .B2(n6270), .ZN(n6217) );
  OAI211_X1 U7200 ( .C1(n6331), .C2(n6224), .A(n6218), .B(n6217), .ZN(U3130)
         );
  AOI22_X1 U7201 ( .A1(n6335), .A2(n6220), .B1(n6333), .B2(n6219), .ZN(n6223)
         );
  AOI22_X1 U7202 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6221), .B1(n6337), 
        .B2(n6270), .ZN(n6222) );
  OAI211_X1 U7203 ( .C1(n6342), .C2(n6224), .A(n6223), .B(n6222), .ZN(U3131)
         );
  INV_X1 U7204 ( .A(n6225), .ZN(n6284) );
  NOR2_X1 U7205 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6281), .ZN(n6268)
         );
  NAND3_X1 U7206 ( .A1(n6228), .A2(n6227), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7207 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(n6269) );
  AOI22_X1 U7208 ( .A1(n6280), .A2(n6268), .B1(n6279), .B2(n6269), .ZN(n6242)
         );
  OAI21_X1 U7209 ( .B1(n6233), .B2(n6283), .A(n6232), .ZN(n6234) );
  NAND3_X1 U7210 ( .A1(n6235), .A2(n6290), .A3(n6234), .ZN(n6239) );
  INV_X1 U7211 ( .A(n6268), .ZN(n6236) );
  AOI21_X1 U7212 ( .B1(n6236), .B2(STATE2_REG_3__SCAN_IN), .A(n6358), .ZN(
        n6237) );
  NAND3_X1 U7213 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6272) );
  AOI22_X1 U7214 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6272), .B1(n6240), 
        .B2(n6270), .ZN(n6241) );
  OAI211_X1 U7215 ( .C1(n6243), .C2(n6341), .A(n6242), .B(n6241), .ZN(U3132)
         );
  AOI22_X1 U7216 ( .A1(n6297), .A2(n6268), .B1(n6296), .B2(n6269), .ZN(n6246)
         );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6272), .B1(n6244), 
        .B2(n6270), .ZN(n6245) );
  OAI211_X1 U7218 ( .C1(n6247), .C2(n6341), .A(n6246), .B(n6245), .ZN(U3133)
         );
  AOI22_X1 U7219 ( .A1(n6303), .A2(n6268), .B1(n6302), .B2(n6269), .ZN(n6250)
         );
  AOI22_X1 U7220 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6272), .B1(n6248), 
        .B2(n6270), .ZN(n6249) );
  OAI211_X1 U7221 ( .C1(n6251), .C2(n6341), .A(n6250), .B(n6249), .ZN(U3134)
         );
  AOI22_X1 U7222 ( .A1(n6309), .A2(n6268), .B1(n6308), .B2(n6269), .ZN(n6254)
         );
  AOI22_X1 U7223 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6272), .B1(n6252), 
        .B2(n6270), .ZN(n6253) );
  OAI211_X1 U7224 ( .C1(n6255), .C2(n6341), .A(n6254), .B(n6253), .ZN(U3135)
         );
  AOI22_X1 U7225 ( .A1(n6315), .A2(n6268), .B1(n6314), .B2(n6269), .ZN(n6258)
         );
  AOI22_X1 U7226 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6272), .B1(n6256), 
        .B2(n6270), .ZN(n6257) );
  OAI211_X1 U7227 ( .C1(n6259), .C2(n6341), .A(n6258), .B(n6257), .ZN(U3136)
         );
  AOI22_X1 U7228 ( .A1(n6321), .A2(n6268), .B1(n6320), .B2(n6269), .ZN(n6262)
         );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6272), .B1(n6260), 
        .B2(n6270), .ZN(n6261) );
  OAI211_X1 U7230 ( .C1(n6263), .C2(n6341), .A(n6262), .B(n6261), .ZN(U3137)
         );
  AOI22_X1 U7231 ( .A1(n6327), .A2(n6268), .B1(n6326), .B2(n6269), .ZN(n6266)
         );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6272), .B1(n6264), 
        .B2(n6270), .ZN(n6265) );
  OAI211_X1 U7233 ( .C1(n6267), .C2(n6341), .A(n6266), .B(n6265), .ZN(U3138)
         );
  AOI22_X1 U7234 ( .A1(n6335), .A2(n6269), .B1(n6333), .B2(n6268), .ZN(n6274)
         );
  AOI22_X1 U7235 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6272), .B1(n6271), 
        .B2(n6270), .ZN(n6273) );
  OAI211_X1 U7236 ( .C1(n6275), .C2(n6341), .A(n6274), .B(n6273), .ZN(U3139)
         );
  AOI21_X1 U7237 ( .B1(n6277), .B2(n6276), .A(n6332), .ZN(n6285) );
  OAI22_X1 U7238 ( .A1(n6285), .A2(n6278), .B1(n6281), .B2(n3391), .ZN(n6334)
         );
  AOI22_X1 U7239 ( .A1(n6280), .A2(n6332), .B1(n6279), .B2(n6334), .ZN(n6294)
         );
  INV_X1 U7240 ( .A(n6281), .ZN(n6291) );
  AOI21_X1 U7241 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(n6287) );
  OAI21_X1 U7242 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(n6288) );
  OAI211_X1 U7243 ( .C1(n6291), .C2(n6290), .A(n6289), .B(n6288), .ZN(n6338)
         );
  AOI22_X1 U7244 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6338), .B1(n6292), 
        .B2(n6336), .ZN(n6293) );
  OAI211_X1 U7245 ( .C1(n6295), .C2(n6341), .A(n6294), .B(n6293), .ZN(U3140)
         );
  AOI22_X1 U7246 ( .A1(n6297), .A2(n6332), .B1(n6296), .B2(n6334), .ZN(n6300)
         );
  AOI22_X1 U7247 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6338), .B1(n6298), 
        .B2(n6336), .ZN(n6299) );
  OAI211_X1 U7248 ( .C1(n6301), .C2(n6341), .A(n6300), .B(n6299), .ZN(U3141)
         );
  AOI22_X1 U7249 ( .A1(n6303), .A2(n6332), .B1(n6302), .B2(n6334), .ZN(n6306)
         );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6338), .B1(n6304), 
        .B2(n6336), .ZN(n6305) );
  OAI211_X1 U7251 ( .C1(n6307), .C2(n6341), .A(n6306), .B(n6305), .ZN(U3142)
         );
  AOI22_X1 U7252 ( .A1(n6309), .A2(n6332), .B1(n6308), .B2(n6334), .ZN(n6312)
         );
  AOI22_X1 U7253 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6338), .B1(n6310), 
        .B2(n6336), .ZN(n6311) );
  OAI211_X1 U7254 ( .C1(n6313), .C2(n6341), .A(n6312), .B(n6311), .ZN(U3143)
         );
  AOI22_X1 U7255 ( .A1(n6315), .A2(n6332), .B1(n6314), .B2(n6334), .ZN(n6318)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6338), .B1(n6316), 
        .B2(n6336), .ZN(n6317) );
  OAI211_X1 U7257 ( .C1(n6319), .C2(n6341), .A(n6318), .B(n6317), .ZN(U3144)
         );
  AOI22_X1 U7258 ( .A1(n6321), .A2(n6332), .B1(n6320), .B2(n6334), .ZN(n6324)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6338), .B1(n6322), 
        .B2(n6336), .ZN(n6323) );
  OAI211_X1 U7260 ( .C1(n6325), .C2(n6341), .A(n6324), .B(n6323), .ZN(U3145)
         );
  AOI22_X1 U7261 ( .A1(n6327), .A2(n6332), .B1(n6326), .B2(n6334), .ZN(n6330)
         );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6338), .B1(n6328), 
        .B2(n6336), .ZN(n6329) );
  OAI211_X1 U7263 ( .C1(n6331), .C2(n6341), .A(n6330), .B(n6329), .ZN(U3146)
         );
  AOI22_X1 U7264 ( .A1(n6335), .A2(n6334), .B1(n6333), .B2(n6332), .ZN(n6340)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6338), .B1(n6337), 
        .B2(n6336), .ZN(n6339) );
  OAI211_X1 U7266 ( .C1(n6342), .C2(n6341), .A(n6340), .B(n6339), .ZN(U3147)
         );
  OAI22_X1 U7267 ( .A1(n6345), .A2(n6344), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6343), .ZN(n6467) );
  NAND2_X1 U7268 ( .A1(n6346), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6475) );
  INV_X1 U7269 ( .A(n6475), .ZN(n6348) );
  NOR3_X1 U7270 ( .A1(n6467), .A2(n6348), .A3(n6347), .ZN(n6352) );
  INV_X1 U7271 ( .A(n6352), .ZN(n6355) );
  INV_X1 U7272 ( .A(n6349), .ZN(n6350) );
  OAI22_X1 U7273 ( .A1(n6352), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6351), .B2(n6350), .ZN(n6353) );
  OAI21_X1 U7274 ( .B1(n6355), .B2(n6354), .A(n6353), .ZN(n6356) );
  AOI222_X1 U7275 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6357), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6356), .C1(n6357), .C2(n6356), 
        .ZN(n6359) );
  AOI222_X1 U7276 ( .A1(n6360), .A2(n6359), .B1(n6360), .B2(n6358), .C1(n6359), 
        .C2(n6358), .ZN(n6363) );
  OAI21_X1 U7277 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6361), 
        .ZN(n6362) );
  OAI21_X1 U7278 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6363), .A(n6362), 
        .ZN(n6368) );
  NOR2_X1 U7279 ( .A1(n6364), .A2(n2999), .ZN(n6365) );
  NAND2_X1 U7280 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  NOR2_X1 U7281 ( .A1(n6368), .A2(n6367), .ZN(n6383) );
  OR2_X1 U7282 ( .A1(n6370), .A2(n6369), .ZN(n6374) );
  AOI21_X1 U7283 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6371) );
  INV_X1 U7284 ( .A(n6371), .ZN(n6372) );
  AND2_X1 U7285 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6372), .ZN(n6373) );
  AND2_X1 U7286 ( .A1(n6374), .A2(n6373), .ZN(n6377) );
  OAI221_X1 U7287 ( .B1(n6634), .B2(n6383), .C1(n6634), .C2(n6468), .A(n6377), 
        .ZN(n6465) );
  OAI21_X1 U7288 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6486), .A(n6465), .ZN(
        n6384) );
  AOI221_X1 U7289 ( .B1(n6376), .B2(STATE2_REG_0__SCAN_IN), .C1(n6384), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6375), .ZN(n6382) );
  INV_X1 U7290 ( .A(n6377), .ZN(n6378) );
  OAI211_X1 U7291 ( .C1(n6380), .C2(n6379), .A(n6634), .B(n6378), .ZN(n6381)
         );
  OAI211_X1 U7292 ( .C1(n6383), .C2(n6385), .A(n6382), .B(n6381), .ZN(U3148)
         );
  NAND3_X1 U7293 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6391), .A3(n6384), .ZN(
        n6390) );
  OAI21_X1 U7294 ( .B1(READY_N), .B2(n6386), .A(n6385), .ZN(n6388) );
  AOI21_X1 U7295 ( .B1(n6388), .B2(n6465), .A(n6387), .ZN(n6389) );
  NAND2_X1 U7296 ( .A1(n6390), .A2(n6389), .ZN(U3149) );
  OAI211_X1 U7297 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6486), .A(n6463), .B(
        n6391), .ZN(n6393) );
  OAI21_X1 U7298 ( .B1(n6489), .B2(n6393), .A(n6392), .ZN(U3150) );
  AND2_X1 U7299 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6458), .ZN(U3151) );
  AND2_X1 U7300 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6458), .ZN(U3152) );
  AND2_X1 U7301 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6458), .ZN(U3153) );
  AND2_X1 U7302 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6458), .ZN(U3154) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6458), .ZN(U3155) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6458), .ZN(U3156) );
  INV_X1 U7305 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U7306 ( .A1(n6462), .A2(n6501), .ZN(U3157) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6458), .ZN(U3158) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6458), .ZN(U3159) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6458), .ZN(U3160) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6458), .ZN(U3161) );
  AND2_X1 U7311 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6458), .ZN(U3162) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6458), .ZN(U3163) );
  AND2_X1 U7313 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6458), .ZN(U3164) );
  INV_X1 U7314 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6571) );
  NOR2_X1 U7315 ( .A1(n6462), .A2(n6571), .ZN(U3165) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6458), .ZN(U3166) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6458), .ZN(U3167) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6458), .ZN(U3168) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6458), .ZN(U3169) );
  AND2_X1 U7320 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6458), .ZN(U3170) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6458), .ZN(U3171) );
  AND2_X1 U7322 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6458), .ZN(U3172) );
  AND2_X1 U7323 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6458), .ZN(U3173) );
  INV_X1 U7324 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6541) );
  NOR2_X1 U7325 ( .A1(n6462), .A2(n6541), .ZN(U3174) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6458), .ZN(U3175) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6458), .ZN(U3176) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6458), .ZN(U3177) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6458), .ZN(U3178) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6458), .ZN(U3179) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6458), .ZN(U3180) );
  INV_X1 U7332 ( .A(n6411), .ZN(n6407) );
  NOR2_X1 U7333 ( .A1(n6486), .A2(n6563), .ZN(n6408) );
  AOI21_X1 U7334 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6408), .ZN(n6412)
         );
  OAI21_X1 U7335 ( .B1(NA_N), .B2(n6403), .A(n6405), .ZN(n6406) );
  INV_X1 U7336 ( .A(HOLD), .ZN(n6402) );
  NOR2_X1 U7337 ( .A1(n6563), .A2(n6402), .ZN(n6396) );
  INV_X1 U7338 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6394) );
  OAI21_X1 U7339 ( .B1(n6396), .B2(n6394), .A(n6483), .ZN(n6395) );
  OAI221_X1 U7340 ( .B1(n6407), .B2(n6412), .C1(n6407), .C2(n6406), .A(n6395), 
        .ZN(U3181) );
  NOR2_X1 U7341 ( .A1(n6403), .A2(n6402), .ZN(n6400) );
  AOI21_X1 U7342 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6396), .ZN(n6399) );
  INV_X1 U7343 ( .A(n6408), .ZN(n6397) );
  OAI211_X1 U7344 ( .C1(n6400), .C2(n6399), .A(n6398), .B(n6397), .ZN(U3182)
         );
  INV_X1 U7345 ( .A(NA_N), .ZN(n6515) );
  AOI21_X1 U7346 ( .B1(READY_N), .B2(n6515), .A(n6563), .ZN(n6401) );
  AOI211_X1 U7347 ( .C1(n6403), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6402), 
        .B(n6401), .ZN(n6404) );
  OAI22_X1 U7348 ( .A1(n6407), .A2(n6406), .B1(n6405), .B2(n6404), .ZN(n6410)
         );
  NAND4_X1 U7349 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .A3(n6408), .A4(n6515), .ZN(n6409) );
  OAI211_X1 U7350 ( .C1(n6412), .C2(n6411), .A(n6410), .B(n6409), .ZN(U3183)
         );
  AND2_X1 U7351 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6494), .ZN(n6445) );
  NOR2_X2 U7352 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6483), .ZN(n6450) );
  AOI22_X1 U7353 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6483), .ZN(n6413) );
  OAI21_X1 U7354 ( .B1(n5615), .B2(n6453), .A(n6413), .ZN(U3184) );
  AOI22_X1 U7355 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6483), .ZN(n6414) );
  OAI21_X1 U7356 ( .B1(n6415), .B2(n6453), .A(n6414), .ZN(U3185) );
  INV_X1 U7357 ( .A(n6450), .ZN(n6456) );
  AOI22_X1 U7358 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6483), .ZN(n6416) );
  OAI21_X1 U7359 ( .B1(n6418), .B2(n6456), .A(n6416), .ZN(U3186) );
  AOI22_X1 U7360 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6483), .ZN(n6417) );
  OAI21_X1 U7361 ( .B1(n6418), .B2(n6453), .A(n6417), .ZN(U3187) );
  INV_X1 U7362 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6601) );
  INV_X1 U7363 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6608) );
  OAI222_X1 U7364 ( .A1(n6453), .A2(n6601), .B1(n6608), .B2(n6494), .C1(n6419), 
        .C2(n6456), .ZN(U3188) );
  INV_X1 U7365 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6524) );
  OAI222_X1 U7366 ( .A1(n6456), .A2(n6421), .B1(n6524), .B2(n6494), .C1(n6419), 
        .C2(n6453), .ZN(U3189) );
  AOI22_X1 U7367 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6483), .ZN(n6420) );
  OAI21_X1 U7368 ( .B1(n6421), .B2(n6453), .A(n6420), .ZN(U3190) );
  AOI22_X1 U7369 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6483), .ZN(n6422) );
  OAI21_X1 U7370 ( .B1(n6424), .B2(n6456), .A(n6422), .ZN(U3191) );
  AOI22_X1 U7371 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6483), .ZN(n6423) );
  OAI21_X1 U7372 ( .B1(n6424), .B2(n6453), .A(n6423), .ZN(U3192) );
  AOI22_X1 U7373 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6483), .ZN(n6425) );
  OAI21_X1 U7374 ( .B1(n4729), .B2(n6453), .A(n6425), .ZN(U3193) );
  AOI22_X1 U7375 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6483), .ZN(n6426) );
  OAI21_X1 U7376 ( .B1(n6517), .B2(n6456), .A(n6426), .ZN(U3194) );
  AOI22_X1 U7377 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6483), .ZN(n6427) );
  OAI21_X1 U7378 ( .B1(n6517), .B2(n6453), .A(n6427), .ZN(U3195) );
  AOI22_X1 U7379 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6483), .ZN(n6428) );
  OAI21_X1 U7380 ( .B1(n6561), .B2(n6453), .A(n6428), .ZN(U3196) );
  AOI22_X1 U7381 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6483), .ZN(n6429) );
  OAI21_X1 U7382 ( .B1(n6430), .B2(n6456), .A(n6429), .ZN(U3197) );
  INV_X1 U7383 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U7384 ( .A1(n6453), .A2(n6430), .B1(n6591), .B2(n6494), .C1(n5192), 
        .C2(n6456), .ZN(U3198) );
  AOI22_X1 U7385 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6483), .ZN(n6431) );
  OAI21_X1 U7386 ( .B1(n5192), .B2(n6453), .A(n6431), .ZN(U3199) );
  INV_X1 U7387 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6587) );
  OAI222_X1 U7388 ( .A1(n6456), .A2(n6434), .B1(n6587), .B2(n6494), .C1(n6432), 
        .C2(n6453), .ZN(U3200) );
  AOI22_X1 U7389 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6483), .ZN(n6433) );
  OAI21_X1 U7390 ( .B1(n6434), .B2(n6453), .A(n6433), .ZN(U3201) );
  INV_X1 U7391 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6581) );
  OAI222_X1 U7392 ( .A1(n6453), .A2(n6435), .B1(n6581), .B2(n6494), .C1(n6437), 
        .C2(n6456), .ZN(U3202) );
  AOI22_X1 U7393 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6483), .ZN(n6436) );
  OAI21_X1 U7394 ( .B1(n6437), .B2(n6453), .A(n6436), .ZN(U3203) );
  INV_X1 U7395 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6532) );
  OAI222_X1 U7396 ( .A1(n6453), .A2(n6438), .B1(n6532), .B2(n6494), .C1(n6440), 
        .C2(n6456), .ZN(U3204) );
  AOI22_X1 U7397 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6483), .ZN(n6439) );
  OAI21_X1 U7398 ( .B1(n6440), .B2(n6453), .A(n6439), .ZN(U3205) );
  AOI22_X1 U7399 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6483), .ZN(n6441) );
  OAI21_X1 U7400 ( .B1(n6442), .B2(n6453), .A(n6441), .ZN(U3206) );
  AOI22_X1 U7401 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6483), .ZN(n6443) );
  OAI21_X1 U7402 ( .B1(n5130), .B2(n6456), .A(n6443), .ZN(U3207) );
  AOI22_X1 U7403 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6483), .ZN(n6444) );
  OAI21_X1 U7404 ( .B1(n5130), .B2(n6453), .A(n6444), .ZN(U3208) );
  AOI22_X1 U7405 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6445), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6483), .ZN(n6446) );
  OAI21_X1 U7406 ( .B1(n6448), .B2(n6456), .A(n6446), .ZN(U3209) );
  AOI22_X1 U7407 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6483), .ZN(n6447) );
  OAI21_X1 U7408 ( .B1(n6448), .B2(n6453), .A(n6447), .ZN(U3210) );
  INV_X1 U7409 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6594) );
  OAI222_X1 U7410 ( .A1(n6453), .A2(n6449), .B1(n6594), .B2(n6494), .C1(n6452), 
        .C2(n6456), .ZN(U3211) );
  AOI22_X1 U7411 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6450), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6483), .ZN(n6451) );
  OAI21_X1 U7412 ( .B1(n6452), .B2(n6453), .A(n6451), .ZN(U3212) );
  INV_X1 U7413 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6455) );
  INV_X1 U7414 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6547) );
  OAI222_X1 U7415 ( .A1(n6456), .A2(n6455), .B1(n6547), .B2(n6494), .C1(n6454), 
        .C2(n6453), .ZN(U3213) );
  MUX2_X1 U7416 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6494), .Z(U3445) );
  MUX2_X1 U7417 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6494), .Z(U3446) );
  MUX2_X1 U7418 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6494), .Z(U3447) );
  MUX2_X1 U7419 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6494), .Z(U3448) );
  INV_X1 U7420 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6459) );
  INV_X1 U7421 ( .A(n6460), .ZN(n6457) );
  AOI21_X1 U7422 ( .B1(n6459), .B2(n6458), .A(n6457), .ZN(U3451) );
  OAI21_X1 U7423 ( .B1(n6462), .B2(n6461), .A(n6460), .ZN(U3452) );
  OAI211_X1 U7424 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n6463), .ZN(U3453)
         );
  INV_X1 U7425 ( .A(n6467), .ZN(n6469) );
  OAI22_X1 U7426 ( .A1(n6469), .A2(n6474), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6468), .ZN(n6471) );
  OAI22_X1 U7427 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6472), .B1(n6471), .B2(n6470), .ZN(n6473) );
  OAI21_X1 U7428 ( .B1(n6475), .B2(n6474), .A(n6473), .ZN(U3461) );
  AOI21_X1 U7429 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6476) );
  AOI22_X1 U7430 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6476), .B2(n5615), .ZN(n6478) );
  INV_X1 U7431 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U7432 ( .A1(n6479), .A2(n6478), .B1(n6477), .B2(n6481), .ZN(U3468)
         );
  INV_X1 U7433 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6482) );
  NOR2_X1 U7434 ( .A1(n6481), .A2(REIP_REG_1__SCAN_IN), .ZN(n6480) );
  AOI22_X1 U7435 ( .A1(n6482), .A2(n6481), .B1(n6527), .B2(n6480), .ZN(U3469)
         );
  INV_X1 U7436 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6542) );
  AOI22_X1 U7437 ( .A1(n6494), .A2(READREQUEST_REG_SCAN_IN), .B1(n6542), .B2(
        n6483), .ZN(U3470) );
  AOI211_X1 U7438 ( .C1(n5663), .C2(n6486), .A(n6485), .B(n6484), .ZN(n6493)
         );
  OAI211_X1 U7439 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6488), .A(n6487), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6490) );
  AOI21_X1 U7440 ( .B1(n6490), .B2(STATE2_REG_0__SCAN_IN), .A(n6489), .ZN(
        n6492) );
  NAND2_X1 U7441 ( .A1(n6493), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6491) );
  OAI21_X1 U7442 ( .B1(n6493), .B2(n6492), .A(n6491), .ZN(U3472) );
  MUX2_X1 U7443 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6494), .Z(U3473) );
  AOI22_X1 U7444 ( .A1(n6621), .A2(keyinput49), .B1(n6496), .B2(keyinput14), 
        .ZN(n6495) );
  OAI221_X1 U7445 ( .B1(n6621), .B2(keyinput49), .C1(n6496), .C2(keyinput14), 
        .A(n6495), .ZN(n6508) );
  AOI22_X1 U7446 ( .A1(n6499), .A2(keyinput0), .B1(n6498), .B2(keyinput34), 
        .ZN(n6497) );
  OAI221_X1 U7447 ( .B1(n6499), .B2(keyinput0), .C1(n6498), .C2(keyinput34), 
        .A(n6497), .ZN(n6507) );
  INV_X1 U7448 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6502) );
  AOI22_X1 U7449 ( .A1(n6502), .A2(keyinput60), .B1(n6501), .B2(keyinput11), 
        .ZN(n6500) );
  OAI221_X1 U7450 ( .B1(n6502), .B2(keyinput60), .C1(n6501), .C2(keyinput11), 
        .A(n6500), .ZN(n6506) );
  INV_X1 U7451 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U7452 ( .A1(n6504), .A2(keyinput21), .B1(n6629), .B2(keyinput26), 
        .ZN(n6503) );
  OAI221_X1 U7453 ( .B1(n6504), .B2(keyinput21), .C1(n6629), .C2(keyinput26), 
        .A(n6503), .ZN(n6505) );
  NOR4_X1 U7454 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n6555)
         );
  INV_X1 U7455 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6510) );
  AOI22_X1 U7456 ( .A1(n6511), .A2(keyinput23), .B1(n6510), .B2(keyinput62), 
        .ZN(n6509) );
  OAI221_X1 U7457 ( .B1(n6511), .B2(keyinput23), .C1(n6510), .C2(keyinput62), 
        .A(n6509), .ZN(n6522) );
  AOI22_X1 U7458 ( .A1(n6652), .A2(keyinput4), .B1(keyinput51), .B2(n6513), 
        .ZN(n6512) );
  OAI221_X1 U7459 ( .B1(n6652), .B2(keyinput4), .C1(n6513), .C2(keyinput51), 
        .A(n6512), .ZN(n6521) );
  INV_X1 U7460 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U7461 ( .A1(n6631), .A2(keyinput24), .B1(keyinput7), .B2(n6515), 
        .ZN(n6514) );
  OAI221_X1 U7462 ( .B1(n6631), .B2(keyinput24), .C1(n6515), .C2(keyinput7), 
        .A(n6514), .ZN(n6520) );
  AOI22_X1 U7463 ( .A1(n6518), .A2(keyinput41), .B1(n6517), .B2(keyinput32), 
        .ZN(n6516) );
  OAI221_X1 U7464 ( .B1(n6518), .B2(keyinput41), .C1(n6517), .C2(keyinput32), 
        .A(n6516), .ZN(n6519) );
  NOR4_X1 U7465 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n6554)
         );
  AOI22_X1 U7466 ( .A1(n6524), .A2(keyinput38), .B1(n5255), .B2(keyinput27), 
        .ZN(n6523) );
  OAI221_X1 U7467 ( .B1(n6524), .B2(keyinput38), .C1(n5255), .C2(keyinput27), 
        .A(n6523), .ZN(n6536) );
  AOI22_X1 U7468 ( .A1(n6527), .A2(keyinput52), .B1(n6526), .B2(keyinput18), 
        .ZN(n6525) );
  OAI221_X1 U7469 ( .B1(n6527), .B2(keyinput52), .C1(n6526), .C2(keyinput18), 
        .A(n6525), .ZN(n6535) );
  INV_X1 U7470 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6529) );
  AOI22_X1 U7471 ( .A1(n6529), .A2(keyinput31), .B1(n3836), .B2(keyinput35), 
        .ZN(n6528) );
  OAI221_X1 U7472 ( .B1(n6529), .B2(keyinput31), .C1(n3836), .C2(keyinput35), 
        .A(n6528), .ZN(n6534) );
  INV_X1 U7473 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7474 ( .A1(n6532), .A2(keyinput10), .B1(n6531), .B2(keyinput28), 
        .ZN(n6530) );
  OAI221_X1 U7475 ( .B1(n6532), .B2(keyinput10), .C1(n6531), .C2(keyinput28), 
        .A(n6530), .ZN(n6533) );
  NOR4_X1 U7476 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .ZN(n6553)
         );
  AOI22_X1 U7477 ( .A1(n6539), .A2(keyinput59), .B1(keyinput54), .B2(n6538), 
        .ZN(n6537) );
  OAI221_X1 U7478 ( .B1(n6539), .B2(keyinput59), .C1(n6538), .C2(keyinput54), 
        .A(n6537), .ZN(n6551) );
  AOI22_X1 U7479 ( .A1(n6542), .A2(keyinput42), .B1(n6541), .B2(keyinput2), 
        .ZN(n6540) );
  OAI221_X1 U7480 ( .B1(n6542), .B2(keyinput42), .C1(n6541), .C2(keyinput2), 
        .A(n6540), .ZN(n6550) );
  AOI22_X1 U7481 ( .A1(n6545), .A2(keyinput57), .B1(n6544), .B2(keyinput29), 
        .ZN(n6543) );
  OAI221_X1 U7482 ( .B1(n6545), .B2(keyinput57), .C1(n6544), .C2(keyinput29), 
        .A(n6543), .ZN(n6549) );
  AOI22_X1 U7483 ( .A1(n6547), .A2(keyinput37), .B1(n6632), .B2(keyinput22), 
        .ZN(n6546) );
  OAI221_X1 U7484 ( .B1(n6547), .B2(keyinput37), .C1(n6632), .C2(keyinput22), 
        .A(n6546), .ZN(n6548) );
  NOR4_X1 U7485 ( .A1(n6551), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(n6552)
         );
  NAND4_X1 U7486 ( .A1(n6555), .A2(n6554), .A3(n6553), .A4(n6552), .ZN(n6620)
         );
  INV_X1 U7487 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7488 ( .A1(n6558), .A2(keyinput12), .B1(keyinput8), .B2(n6557), 
        .ZN(n6556) );
  OAI221_X1 U7489 ( .B1(n6558), .B2(keyinput12), .C1(n6557), .C2(keyinput8), 
        .A(n6556), .ZN(n6569) );
  INV_X1 U7490 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6560) );
  AOI22_X1 U7491 ( .A1(n6561), .A2(keyinput17), .B1(n6560), .B2(keyinput43), 
        .ZN(n6559) );
  OAI221_X1 U7492 ( .B1(n6561), .B2(keyinput17), .C1(n6560), .C2(keyinput43), 
        .A(n6559), .ZN(n6568) );
  INV_X1 U7493 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6630) );
  AOI22_X1 U7494 ( .A1(n6630), .A2(keyinput63), .B1(keyinput6), .B2(n6563), 
        .ZN(n6562) );
  OAI221_X1 U7495 ( .B1(n6630), .B2(keyinput63), .C1(n6563), .C2(keyinput6), 
        .A(n6562), .ZN(n6567) );
  AOI22_X1 U7496 ( .A1(n4153), .A2(keyinput5), .B1(keyinput45), .B2(n6565), 
        .ZN(n6564) );
  OAI221_X1 U7497 ( .B1(n4153), .B2(keyinput5), .C1(n6565), .C2(keyinput45), 
        .A(n6564), .ZN(n6566) );
  NOR4_X1 U7498 ( .A1(n6569), .A2(n6568), .A3(n6567), .A4(n6566), .ZN(n6618)
         );
  INV_X1 U7499 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7500 ( .A1(n6575), .A2(keyinput39), .B1(keyinput1), .B2(n6574), 
        .ZN(n6573) );
  OAI221_X1 U7501 ( .B1(n6575), .B2(keyinput39), .C1(n6574), .C2(keyinput1), 
        .A(n6573), .ZN(n6584) );
  INV_X1 U7502 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U7503 ( .A1(n6578), .A2(keyinput3), .B1(keyinput56), .B2(n6577), 
        .ZN(n6576) );
  OAI221_X1 U7504 ( .B1(n6578), .B2(keyinput3), .C1(n6577), .C2(keyinput56), 
        .A(n6576), .ZN(n6583) );
  INV_X1 U7505 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6580) );
  AOI22_X1 U7506 ( .A1(n6581), .A2(keyinput16), .B1(n6580), .B2(keyinput25), 
        .ZN(n6579) );
  OAI221_X1 U7507 ( .B1(n6581), .B2(keyinput16), .C1(n6580), .C2(keyinput25), 
        .A(n6579), .ZN(n6582) );
  NOR4_X1 U7508 ( .A1(n6585), .A2(n6584), .A3(n6583), .A4(n6582), .ZN(n6617)
         );
  AOI22_X1 U7509 ( .A1(n6587), .A2(keyinput44), .B1(n6633), .B2(keyinput15), 
        .ZN(n6586) );
  OAI221_X1 U7510 ( .B1(n6587), .B2(keyinput44), .C1(n6633), .C2(keyinput15), 
        .A(n6586), .ZN(n6599) );
  AOI22_X1 U7511 ( .A1(n6589), .A2(keyinput40), .B1(keyinput19), .B2(n5615), 
        .ZN(n6588) );
  OAI221_X1 U7512 ( .B1(n6589), .B2(keyinput40), .C1(n5615), .C2(keyinput19), 
        .A(n6588), .ZN(n6598) );
  AOI22_X1 U7513 ( .A1(n6592), .A2(keyinput47), .B1(keyinput13), .B2(n6591), 
        .ZN(n6590) );
  OAI221_X1 U7514 ( .B1(n6592), .B2(keyinput47), .C1(n6591), .C2(keyinput13), 
        .A(n6590), .ZN(n6597) );
  INV_X1 U7515 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7516 ( .A1(n6595), .A2(keyinput58), .B1(keyinput9), .B2(n6594), 
        .ZN(n6593) );
  OAI221_X1 U7517 ( .B1(n6595), .B2(keyinput58), .C1(n6594), .C2(keyinput9), 
        .A(n6593), .ZN(n6596) );
  NOR4_X1 U7518 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n6616)
         );
  AOI22_X1 U7519 ( .A1(n6602), .A2(keyinput50), .B1(keyinput48), .B2(n6601), 
        .ZN(n6600) );
  OAI221_X1 U7520 ( .B1(n6602), .B2(keyinput50), .C1(n6601), .C2(keyinput48), 
        .A(n6600), .ZN(n6614) );
  INV_X1 U7521 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6604) );
  AOI22_X1 U7522 ( .A1(n6608), .A2(keyinput33), .B1(n6607), .B2(keyinput30), 
        .ZN(n6606) );
  OAI221_X1 U7523 ( .B1(n6608), .B2(keyinput33), .C1(n6607), .C2(keyinput30), 
        .A(n6606), .ZN(n6612) );
  AOI22_X1 U7524 ( .A1(n6610), .A2(keyinput61), .B1(n6634), .B2(keyinput55), 
        .ZN(n6609) );
  OAI221_X1 U7525 ( .B1(n6610), .B2(keyinput61), .C1(n6634), .C2(keyinput55), 
        .A(n6609), .ZN(n6611) );
  NOR4_X1 U7526 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n6615)
         );
  NAND4_X1 U7527 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n6619)
         );
  NOR2_X1 U7528 ( .A1(n6620), .A2(n6619), .ZN(n6657) );
  NOR4_X1 U7529 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .A3(REIP_REG_12__SCAN_IN), .A4(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6648) );
  NAND3_X1 U7530 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n4153), .A3(n6621), .ZN(
        n6624) );
  NAND4_X1 U7531 ( .A1(ADDRESS_REG_4__SCAN_IN), .A2(ADDRESS_REG_14__SCAN_IN), 
        .A3(ADDRESS_REG_16__SCAN_IN), .A4(ADDRESS_REG_29__SCAN_IN), .ZN(n6623)
         );
  NAND4_X1 U7532 ( .A1(W_R_N_REG_SCAN_IN), .A2(ADDRESS_REG_20__SCAN_IN), .A3(
        ADDRESS_REG_27__SCAN_IN), .A4(ADDRESS_REG_18__SCAN_IN), .ZN(n6622) );
  NOR4_X1 U7533 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6624), .A3(n6623), .A4(n6622), 
        .ZN(n6647) );
  NAND4_X1 U7534 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(LWORD_REG_14__SCAN_IN), .A4(
        LWORD_REG_0__SCAN_IN), .ZN(n6628) );
  NAND4_X1 U7535 ( .A1(EBX_REG_18__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        UWORD_REG_4__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n6627) );
  NAND4_X1 U7536 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .A3(PHYADDRPOINTER_REG_16__SCAN_IN), 
        .A4(REIP_REG_0__SCAN_IN), .ZN(n6626) );
  NAND4_X1 U7537 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .A3(DATAI_23_), .A4(DATAI_21_), .ZN(
        n6625) );
  NOR4_X1 U7538 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n6646)
         );
  NAND4_X1 U7539 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(
        INSTQUEUE_REG_14__6__SCAN_IN), .A3(n6630), .A4(n6629), .ZN(n6644) );
  NAND4_X1 U7540 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(
        INSTQUEUE_REG_7__7__SCAN_IN), .A3(n6632), .A4(n6631), .ZN(n6643) );
  NOR2_X1 U7541 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6636) );
  NOR4_X1 U7542 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUE_REG_15__3__SCAN_IN), .A3(n6634), .A4(n6633), .ZN(n6635) );
  NAND4_X1 U7543 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(
        INSTQUEUE_REG_14__3__SCAN_IN), .A3(n6636), .A4(n6635), .ZN(n6642) );
  NOR4_X1 U7544 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(ADDRESS_REG_5__SCAN_IN), 
        .A3(MEMORYFETCH_REG_SCAN_IN), .A4(n6652), .ZN(n6640) );
  NOR4_X1 U7545 ( .A1(STATE_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(EAX_REG_6__SCAN_IN), .A4(NA_N), 
        .ZN(n6639) );
  NOR4_X1 U7546 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        LWORD_REG_3__SCAN_IN), .A3(DATAO_REG_8__SCAN_IN), .A4(
        UWORD_REG_6__SCAN_IN), .ZN(n6638) );
  NOR4_X1 U7547 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        DATAI_18_), .A4(UWORD_REG_8__SCAN_IN), .ZN(n6637) );
  NAND4_X1 U7548 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6641)
         );
  NOR4_X1 U7549 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6645)
         );
  NAND4_X1 U7550 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6655)
         );
  AOI22_X1 U7551 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6650), .B1(n6649), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6651) );
  OAI21_X1 U7552 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6654) );
  XOR2_X1 U7553 ( .A(n6655), .B(n6654), .Z(n6656) );
  XNOR2_X1 U7554 ( .A(n6657), .B(n6656), .ZN(U2950) );
  CLKBUF_X1 U3405 ( .A(n3151), .Z(n3505) );
  CLKBUF_X1 U3418 ( .A(n3186), .Z(n3195) );
  INV_X1 U3433 ( .A(n3206), .ZN(n3385) );
  CLKBUF_X1 U34590 ( .A(n3887), .Z(n2978) );
  CLKBUF_X1 U3513 ( .A(n4083), .Z(n2979) );
endmodule

