

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361;

  CLKBUF_X1 U4918 ( .A(n5183), .Z(n6922) );
  INV_X1 U4919 ( .A(n7739), .ZN(n7738) );
  BUF_X2 U4920 ( .A(n5217), .Z(n7538) );
  XNOR2_X1 U4921 ( .A(n5074), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5077) );
  OR2_X1 U4923 ( .A1(n6484), .A2(n6224), .ZN(n6482) );
  NAND2_X1 U4924 ( .A1(n4510), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6850) );
  OR2_X1 U4925 ( .A1(n5378), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U4926 ( .A1(n5692), .A2(n7607), .ZN(n5690) );
  INV_X1 U4927 ( .A(n9000), .ZN(n6034) );
  NOR2_X2 U4928 ( .A1(n7902), .A2(n7901), .ZN(n7998) );
  INV_X1 U4929 ( .A(n6926), .ZN(n5211) );
  INV_X1 U4930 ( .A(n7538), .ZN(n5488) );
  OR2_X1 U4931 ( .A1(n5076), .A2(n5073), .ZN(n5074) );
  OR2_X1 U4932 ( .A1(n6830), .A2(n6831), .ZN(n7170) );
  INV_X1 U4933 ( .A(n6340), .ZN(n6125) );
  INV_X1 U4934 ( .A(n5873), .ZN(n6329) );
  INV_X1 U4935 ( .A(n8805), .ZN(n6975) );
  OAI21_X1 U4936 ( .B1(n6151), .B2(n4754), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6181) );
  NAND2_X1 U4937 ( .A1(n8058), .A2(n7882), .ZN(n7970) );
  OR3_X1 U4938 ( .A1(n7457), .A2(n7451), .A3(n7437), .ZN(n6520) );
  INV_X1 U4939 ( .A(n5830), .ZN(n4415) );
  INV_X1 U4940 ( .A(n6579), .ZN(n5197) );
  XNOR2_X1 U4941 ( .A(n5255), .B(n10177), .ZN(n6708) );
  AND4_X1 U4942 ( .A1(n6007), .A2(n6180), .A3(n5792), .A4(n5766), .ZN(n4412)
         );
  OR2_X1 U4943 ( .A1(n8123), .A2(n8138), .ZN(n4413) );
  INV_X1 U4944 ( .A(n6903), .ZN(n6630) );
  AOI21_X1 U4945 ( .B1(n8908), .B2(n8905), .A(n9065), .ZN(n4634) );
  MUX2_X2 U4946 ( .A(n8909), .B(n8903), .S(n9049), .Z(n8908) );
  INV_X1 U4947 ( .A(n6342), .ZN(n5811) );
  OAI21_X2 U4948 ( .B1(n5277), .B2(n4963), .A(n4960), .ZN(n5309) );
  NAND2_X2 U4949 ( .A1(n5275), .A2(n5274), .ZN(n5277) );
  NOR2_X2 U4950 ( .A1(n5801), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U4951 ( .A1(n6288), .A2(n9139), .ZN(n6507) );
  BUF_X8 U4952 ( .A(n6630), .Z(n4414) );
  OAI21_X2 U4953 ( .B1(n6998), .B2(n7003), .A(n6997), .ZN(n7076) );
  NOR2_X2 U4954 ( .A1(n9459), .A2(n6044), .ZN(n6045) );
  OAI22_X4 U4955 ( .A1(n5421), .A2(n4689), .B1(SI_15_), .B2(n5419), .ZN(n5441)
         );
  NAND2_X2 U4956 ( .A1(n5155), .A2(n4930), .ZN(n5421) );
  INV_X1 U4957 ( .A(n9341), .ZN(n9664) );
  NAND2_X4 U4958 ( .A1(n5680), .A2(n5681), .ZN(n5189) );
  XNOR2_X2 U4959 ( .A(n4756), .B(n5007), .ZN(n5681) );
  XNOR2_X2 U4960 ( .A(n5188), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9858) );
  AND2_X1 U4961 ( .A1(n8046), .A2(n4900), .ZN(n7943) );
  NAND2_X1 U4962 ( .A1(n6116), .A2(n6115), .ZN(n9341) );
  NAND2_X1 U4963 ( .A1(n5782), .A2(n5781), .ZN(n9375) );
  AOI21_X1 U4964 ( .B1(n6841), .B2(n6840), .A(n6839), .ZN(n6843) );
  AOI21_X1 U4965 ( .B1(n6699), .B2(n6708), .A(n6698), .ZN(n6700) );
  NOR2_X1 U4966 ( .A1(n8084), .A2(n7980), .ZN(n7014) );
  NAND2_X1 U4967 ( .A1(n8909), .A2(n8904), .ZN(n9015) );
  NAND2_X1 U4968 ( .A1(n6162), .A2(n9061), .ZN(n9014) );
  INV_X1 U4969 ( .A(n6875), .ZN(n6884) );
  NAND2_X2 U4970 ( .A1(n5227), .A2(n5226), .ZN(n7611) );
  NAND2_X2 U4971 ( .A1(n5197), .A2(n5196), .ZN(n5692) );
  INV_X2 U4972 ( .A(n9908), .ZN(n5246) );
  INV_X1 U4973 ( .A(n9169), .ZN(n6755) );
  INV_X2 U4974 ( .A(n9918), .ZN(n5196) );
  INV_X2 U4975 ( .A(n5846), .ZN(n5848) );
  INV_X1 U4976 ( .A(n5226), .ZN(n9923) );
  AND4_X1 U4977 ( .A1(n5826), .A2(n4453), .A3(n5825), .A4(n5824), .ZN(n6591)
         );
  OR2_X1 U4978 ( .A1(n5210), .A2(n6983), .ZN(n5184) );
  NAND2_X1 U4980 ( .A1(n5091), .A2(n7519), .ZN(n6926) );
  NAND2_X4 U4981 ( .A1(n5189), .A2(n7533), .ZN(n5222) );
  NAND2_X1 U4983 ( .A1(n6247), .A2(n6481), .ZN(n6251) );
  AND2_X1 U4984 ( .A1(n5072), .A2(n5005), .ZN(n5076) );
  NAND2_X1 U4985 ( .A1(n5001), .A2(n5000), .ZN(n5463) );
  NAND2_X1 U4986 ( .A1(n6789), .A2(n5097), .ZN(n4928) );
  NAND2_X1 U4987 ( .A1(n4825), .A2(n4423), .ZN(n9322) );
  NOR2_X1 U4988 ( .A1(n8197), .A2(n4620), .ZN(n4619) );
  AND2_X1 U4989 ( .A1(n8165), .A2(n8164), .ZN(n8173) );
  OAI21_X1 U4990 ( .B1(n8271), .B2(n5583), .A(n5582), .ZN(n8262) );
  OAI21_X1 U4991 ( .B1(n8329), .B2(n5706), .A(n7707), .ZN(n8322) );
  NAND2_X2 U4992 ( .A1(n6123), .A2(n6122), .ZN(n9574) );
  NAND2_X1 U4993 ( .A1(n8348), .A2(n7702), .ZN(n8329) );
  XNOR2_X1 U4994 ( .A(n7536), .B(n7535), .ZN(n8994) );
  NAND2_X1 U4995 ( .A1(n5009), .A2(n5008), .ZN(n8348) );
  OR2_X1 U4996 ( .A1(n8360), .A2(n5704), .ZN(n5009) );
  NAND2_X1 U4997 ( .A1(n4496), .A2(n6105), .ZN(n9585) );
  OR2_X1 U4998 ( .A1(n9375), .A2(n9393), .ZN(n4511) );
  NAND2_X1 U4999 ( .A1(n4974), .A2(n4972), .ZN(n8372) );
  AND2_X2 U5000 ( .A1(n5572), .A2(n5571), .ZN(n8537) );
  NAND2_X1 U5001 ( .A1(n7284), .A2(n7283), .ZN(n7413) );
  NAND2_X1 U5002 ( .A1(n6091), .A2(n6090), .ZN(n9595) );
  NAND2_X1 U5003 ( .A1(n8426), .A2(n7671), .ZN(n8417) );
  NAND2_X1 U5004 ( .A1(n6079), .A2(n6078), .ZN(n9407) );
  AOI21_X1 U5005 ( .B1(n4850), .B2(n4848), .A(n4462), .ZN(n4847) );
  NAND2_X1 U5006 ( .A1(n5541), .A2(n5540), .ZN(n8026) );
  NAND2_X1 U5007 ( .A1(n8796), .A2(n6828), .ZN(n7173) );
  NAND2_X1 U5008 ( .A1(n6036), .A2(n6035), .ZN(n9625) );
  AND2_X1 U5009 ( .A1(n4519), .A2(n6830), .ZN(n8796) );
  NAND2_X1 U5010 ( .A1(n4809), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U5011 ( .A1(n4810), .A2(n7079), .ZN(n7007) );
  NAND2_X1 U5012 ( .A1(n5360), .A2(n5359), .ZN(n7362) );
  NAND2_X1 U5013 ( .A1(n5341), .A2(n5340), .ZN(n7341) );
  NAND2_X2 U5014 ( .A1(n6613), .A2(n9898), .ZN(n9913) );
  OAI21_X1 U5015 ( .B1(n5324), .B2(n5323), .A(n5136), .ZN(n5333) );
  INV_X2 U5016 ( .A(n6355), .ZN(n6463) );
  NAND2_X1 U5017 ( .A1(n5883), .A2(n5882), .ZN(n8805) );
  NAND2_X1 U5018 ( .A1(n5311), .A2(n5132), .ZN(n5324) );
  OAI211_X1 U5019 ( .C1(n5873), .C2(n9215), .A(n5872), .B(n5871), .ZN(n6875)
         );
  CLKBUF_X1 U5020 ( .A(n6532), .Z(n8680) );
  NAND4_X1 U5021 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n6987)
         );
  NAND4_X1 U5022 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n9169)
         );
  INV_X1 U5023 ( .A(n6591), .ZN(n4416) );
  NAND4_X2 U5024 ( .A1(n5815), .A2(n5813), .A3(n5816), .A4(n5814), .ZN(n9057)
         );
  AND2_X2 U5025 ( .A1(n6521), .A2(n6221), .ZN(P1_U3973) );
  NAND2_X1 U5026 ( .A1(n5715), .A2(n5716), .ZN(n7424) );
  OR2_X1 U5027 ( .A1(n5841), .A2(n5812), .ZN(n5813) );
  CLKBUF_X2 U5028 ( .A(n6926), .Z(n4417) );
  CLKBUF_X3 U5029 ( .A(n5841), .Z(n6343) );
  INV_X1 U5030 ( .A(n5077), .ZN(n7519) );
  INV_X1 U5031 ( .A(n5772), .ZN(n9701) );
  XNOR2_X1 U5032 ( .A(n5486), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U5033 ( .A1(n5195), .A2(n5194), .ZN(n5819) );
  NAND2_X2 U5034 ( .A1(n5771), .A2(n5773), .ZN(n6342) );
  INV_X1 U5035 ( .A(n5771), .ZN(n7851) );
  XNOR2_X1 U5036 ( .A(n4757), .B(n5159), .ZN(n5680) );
  NAND2_X1 U5037 ( .A1(n4758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4756) );
  OAI21_X1 U5038 ( .B1(n4758), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4757) );
  OR2_X1 U5039 ( .A1(n5317), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U5040 ( .A1(n5072), .A2(n5071), .ZN(n4758) );
  INV_X1 U5041 ( .A(n5463), .ZN(n5069) );
  OAI21_X1 U5042 ( .B1(n5780), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4569) );
  OR2_X2 U5043 ( .A1(n5133), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9709) );
  NAND2_X1 U5044 ( .A1(n6188), .A2(n4424), .ZN(n9697) );
  OR2_X1 U5045 ( .A1(n5281), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5301) );
  AND4_X1 U5046 ( .A1(n4744), .A2(n4745), .A3(n4747), .A4(n4475), .ZN(n5798)
         );
  AND3_X1 U5047 ( .A1(n5003), .A2(n5002), .A3(n4760), .ZN(n4759) );
  AND2_X1 U5048 ( .A1(n4746), .A2(n4747), .ZN(n5980) );
  AND2_X1 U5049 ( .A1(n5004), .A2(n5673), .ZN(n5003) );
  NOR2_X1 U5050 ( .A1(n5015), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4744) );
  NAND2_X2 U5051 ( .A1(n4929), .A2(n4928), .ZN(n5160) );
  NOR2_X1 U5052 ( .A1(n5014), .A2(n5015), .ZN(n4746) );
  AND2_X1 U5053 ( .A1(n5068), .A2(n5676), .ZN(n5004) );
  AND2_X1 U5054 ( .A1(n5067), .A2(n5066), .ZN(n5000) );
  NAND2_X1 U5055 ( .A1(n6790), .A2(n5096), .ZN(n4929) );
  AND2_X1 U5056 ( .A1(n4908), .A2(n6257), .ZN(n5254) );
  INV_X1 U5057 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10053) );
  AND2_X1 U5058 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6789) );
  INV_X1 U5059 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5911) );
  NOR2_X2 U5060 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6790) );
  INV_X1 U5061 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6180) );
  INV_X1 U5062 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5792) );
  INV_X1 U5063 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5794) );
  INV_X1 U5064 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5016) );
  NOR2_X1 U5065 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5012) );
  INV_X1 U5066 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5869) );
  INV_X1 U5067 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5097) );
  INV_X1 U5068 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5337) );
  INV_X1 U5069 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5673) );
  INV_X1 U5070 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5325) );
  INV_X1 U5071 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5293) );
  INV_X1 U5072 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5066) );
  NOR2_X1 U5073 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5058) );
  NOR2_X1 U5074 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5059) );
  NOR2_X1 U5075 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4908) );
  NOR2_X1 U5076 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5060) );
  NOR2_X1 U5077 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5061) );
  NOR2_X2 U5078 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5068) );
  INV_X4 U5079 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI22_X2 U5080 ( .A1(n9543), .A2(n9544), .B1(n8892), .B2(n9561), .ZN(n9522)
         );
  NAND2_X2 U5081 ( .A1(n7346), .A2(n5994), .ZN(n9543) );
  XNOR2_X2 U5082 ( .A(n6150), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6288) );
  OAI21_X2 U5083 ( .B1(n8407), .B2(n7673), .A(n7677), .ZN(n8394) );
  INV_X4 U5084 ( .A(n6226), .ZN(n8208) );
  AOI22_X2 U5085 ( .A1(n9414), .A2(n6077), .B1(n8650), .B2(n9420), .ZN(n9398)
         );
  NAND2_X1 U5086 ( .A1(n4836), .A2(n4837), .ZN(n9414) );
  OR2_X1 U5087 ( .A1(n6343), .A2(n5850), .ZN(n5855) );
  NOR2_X1 U5088 ( .A1(n5156), .A2(n5157), .ZN(n4689) );
  INV_X1 U5089 ( .A(n5200), .ZN(n5208) );
  AND2_X1 U5090 ( .A1(n7519), .A2(n7859), .ZN(n5200) );
  AND2_X1 U5091 ( .A1(n4479), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U5092 ( .A1(n8930), .A2(n4675), .ZN(n4674) );
  OAI21_X1 U5093 ( .B1(n4668), .B2(n8936), .A(n4484), .ZN(n4666) );
  AOI21_X1 U5094 ( .B1(n4672), .B2(n4670), .A(n4669), .ZN(n4668) );
  INV_X1 U5095 ( .A(n8934), .ZN(n4669) );
  INV_X1 U5096 ( .A(n4673), .ZN(n4670) );
  NAND2_X1 U5097 ( .A1(n4471), .A2(n4691), .ZN(n4690) );
  INV_X1 U5098 ( .A(n4693), .ZN(n4692) );
  AND2_X1 U5099 ( .A1(n4660), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U5100 ( .A1(n4653), .A2(n8974), .ZN(n4652) );
  NOR2_X1 U5101 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5102 ( .A1(n9092), .A2(n4658), .ZN(n4657) );
  NOR2_X1 U5103 ( .A1(n7729), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U5104 ( .A1(n4712), .A2(n4711), .ZN(n4710) );
  INV_X1 U5105 ( .A(n7728), .ZN(n4711) );
  NAND2_X1 U5106 ( .A1(n4593), .A2(n4592), .ZN(n7258) );
  NAND2_X1 U5107 ( .A1(n4914), .A2(n7087), .ZN(n4592) );
  OAI21_X1 U5108 ( .B1(n7086), .B2(n4596), .A(n7102), .ZN(n4594) );
  OR2_X1 U5109 ( .A1(n8323), .A2(n8334), .ZN(n7589) );
  INV_X1 U5110 ( .A(n4800), .ZN(n4798) );
  AND2_X1 U5111 ( .A1(n9971), .A2(n8079), .ZN(n4808) );
  INV_X1 U5112 ( .A(n5047), .ZN(n4804) );
  OR2_X1 U5113 ( .A1(n9971), .A2(n8429), .ZN(n7665) );
  NOR2_X1 U5114 ( .A1(n7545), .A2(n7649), .ZN(n4980) );
  AND2_X1 U5115 ( .A1(n8526), .A2(n8264), .ZN(n7722) );
  OR2_X1 U5116 ( .A1(n8526), .A2(n8264), .ZN(n7721) );
  OR2_X1 U5117 ( .A1(n5530), .A2(n8320), .ZN(n7590) );
  NAND2_X1 U5118 ( .A1(n8532), .A2(n8273), .ZN(n7717) );
  OR2_X1 U5119 ( .A1(n5708), .A2(n8284), .ZN(n7713) );
  NOR2_X1 U5120 ( .A1(n5476), .A2(n5056), .ZN(n8330) );
  OR2_X1 U5121 ( .A1(n8043), .A2(n8335), .ZN(n7702) );
  OR2_X1 U5122 ( .A1(n8559), .A2(n8347), .ZN(n7703) );
  OR2_X1 U5123 ( .A1(n8570), .A2(n8346), .ZN(n7690) );
  NOR2_X1 U5124 ( .A1(n8593), .A2(n8395), .ZN(n7673) );
  INV_X1 U5125 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5067) );
  OR2_X1 U5126 ( .A1(n9574), .A2(n9341), .ZN(n4590) );
  INV_X1 U5127 ( .A(n6114), .ZN(n4828) );
  NAND2_X1 U5128 ( .A1(n9341), .A2(n8980), .ZN(n9112) );
  OR2_X1 U5129 ( .A1(n9341), .A2(n8980), .ZN(n9098) );
  OR2_X1 U5130 ( .A1(n9585), .A2(n8776), .ZN(n9108) );
  NAND2_X1 U5131 ( .A1(n9585), .A2(n8776), .ZN(n9099) );
  OR2_X1 U5132 ( .A1(n8843), .A2(n5993), .ZN(n8937) );
  INV_X1 U5133 ( .A(n9032), .ZN(n4554) );
  OR2_X1 U5134 ( .A1(n8862), .A2(n8764), .ZN(n8933) );
  XNOR2_X1 U5135 ( .A(n9057), .B(n4415), .ZN(n9017) );
  INV_X1 U5136 ( .A(n6696), .ZN(n5829) );
  OR2_X1 U5137 ( .A1(n6797), .A2(n6961), .ZN(n7029) );
  XNOR2_X1 U5138 ( .A(n7521), .B(n7520), .ZN(n7524) );
  NAND2_X1 U5139 ( .A1(n4940), .A2(n4938), .ZN(n5515) );
  AND2_X1 U5140 ( .A1(n4939), .A2(n5499), .ZN(n4938) );
  NAND2_X1 U5141 ( .A1(n5441), .A2(n4442), .ZN(n4940) );
  XNOR2_X1 U5142 ( .A(n5145), .B(SI_11_), .ZN(n5370) );
  AND2_X1 U5143 ( .A1(n5351), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U5144 ( .A1(n5135), .A2(n10113), .ZN(n5136) );
  XNOR2_X1 U5145 ( .A(n5137), .B(SI_9_), .ZN(n5332) );
  NAND2_X1 U5146 ( .A1(n5123), .A2(SI_6_), .ZN(n5127) );
  AND2_X1 U5147 ( .A1(n7864), .A2(n7199), .ZN(n4909) );
  OR2_X1 U5148 ( .A1(n5542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5556) );
  INV_X1 U5149 ( .A(n5210), .ZN(n5665) );
  AND4_X1 U5150 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n7877)
         );
  NAND2_X1 U5151 ( .A1(n4609), .A2(n4608), .ZN(n4607) );
  INV_X1 U5152 ( .A(n7261), .ZN(n4608) );
  INV_X1 U5153 ( .A(n4926), .ZN(n4609) );
  NAND2_X1 U5154 ( .A1(n4787), .A2(n4790), .ZN(n7844) );
  NAND2_X1 U5155 ( .A1(n5633), .A2(n5632), .ZN(n7875) );
  AOI21_X1 U5156 ( .B1(n8296), .B2(n8299), .A(n5547), .ZN(n8282) );
  NOR2_X1 U5157 ( .A1(n8026), .A2(n8076), .ZN(n5547) );
  NAND2_X1 U5158 ( .A1(n8323), .A2(n8334), .ZN(n8309) );
  OR2_X1 U5159 ( .A1(n7940), .A2(n8347), .ZN(n5049) );
  INV_X1 U5160 ( .A(n8395), .ZN(n8430) );
  INV_X1 U5161 ( .A(n8080), .ZN(n8440) );
  NOR2_X1 U5162 ( .A1(n5350), .A2(n4807), .ZN(n4806) );
  INV_X1 U5163 ( .A(n5331), .ZN(n4807) );
  INV_X1 U5164 ( .A(n7427), .ZN(n7361) );
  OAI21_X1 U5165 ( .B1(n5262), .B2(n4768), .A(n4765), .ZN(n7141) );
  AOI21_X1 U5166 ( .B1(n4767), .B2(n4766), .A(n4440), .ZN(n4765) );
  INV_X1 U5167 ( .A(n4772), .ZN(n4766) );
  NAND2_X1 U5168 ( .A1(n5189), .A2(n5133), .ZN(n5217) );
  OR2_X1 U5169 ( .A1(n8262), .A2(n4786), .ZN(n4782) );
  AOI21_X1 U5170 ( .B1(n8384), .B2(n7557), .A(n7559), .ZN(n8374) );
  INV_X1 U5171 ( .A(n5222), .ZN(n7537) );
  INV_X1 U5172 ( .A(n5189), .ZN(n5487) );
  NOR2_X1 U5173 ( .A1(n8423), .A2(n4999), .ZN(n4998) );
  INV_X1 U5174 ( .A(n7666), .ZN(n4999) );
  INV_X1 U5175 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5223) );
  AND2_X1 U5176 ( .A1(n8671), .A2(n8669), .ZN(n8819) );
  XNOR2_X1 U5177 ( .A(n6554), .B(n8678), .ZN(n6813) );
  NAND2_X1 U5178 ( .A1(n8773), .A2(n4741), .ZN(n4740) );
  AND2_X1 U5180 ( .A1(n9098), .A2(n9112), .ZN(n9339) );
  NOR2_X1 U5181 ( .A1(n9375), .A2(n9384), .ZN(n9374) );
  NAND2_X1 U5182 ( .A1(n9614), .A2(n9464), .ZN(n6055) );
  AND2_X1 U5183 ( .A1(n9470), .A2(n9453), .ZN(n6044) );
  OR2_X1 U5184 ( .A1(n9535), .A2(n9159), .ZN(n4856) );
  OR2_X1 U5185 ( .A1(n7294), .A2(n9164), .ZN(n5934) );
  NAND2_X1 U5186 ( .A1(n6727), .A2(n4684), .ZN(n4683) );
  INV_X1 U5187 ( .A(n9016), .ZN(n4684) );
  NAND2_X1 U5188 ( .A1(n5873), .A2(n5133), .ZN(n5837) );
  NAND2_X1 U5189 ( .A1(n5873), .A2(n7533), .ZN(n5857) );
  INV_X2 U5190 ( .A(n5979), .ZN(n8998) );
  OAI21_X1 U5191 ( .B1(n5441), .B2(n5440), .A(n5439), .ZN(n5461) );
  AND2_X1 U5192 ( .A1(n4959), .A2(n4435), .ZN(n4955) );
  INV_X1 U5193 ( .A(n5172), .ZN(n4959) );
  NAND2_X1 U5194 ( .A1(n5355), .A2(n4957), .ZN(n4956) );
  XNOR2_X1 U5195 ( .A(n5371), .B(n5370), .ZN(n6350) );
  NAND2_X1 U5196 ( .A1(n5355), .A2(n5144), .ZN(n5371) );
  NAND2_X1 U5197 ( .A1(n5118), .A2(SI_5_), .ZN(n5122) );
  INV_X1 U5198 ( .A(n6684), .ZN(n6681) );
  NAND4_X1 U5199 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8081)
         );
  OR2_X1 U5200 ( .A1(n5208), .A2(n5316), .ZN(n5321) );
  OR2_X1 U5201 ( .A1(n6407), .A2(n6406), .ZN(n4725) );
  NOR2_X1 U5202 ( .A1(n8913), .A2(n9049), .ZN(n4632) );
  NAND2_X1 U5203 ( .A1(n6157), .A2(n8910), .ZN(n4633) );
  AOI21_X1 U5204 ( .B1(n8908), .B2(n9061), .A(n4638), .ZN(n4637) );
  NAND2_X1 U5205 ( .A1(n8910), .A2(n8909), .ZN(n4638) );
  NOR2_X1 U5206 ( .A1(n8914), .A2(n9004), .ZN(n4636) );
  AOI21_X1 U5207 ( .B1(n4688), .B2(n7738), .A(n4687), .ZN(n4686) );
  NOR2_X1 U5208 ( .A1(n7596), .A2(n7738), .ZN(n4687) );
  NAND2_X1 U5209 ( .A1(n7689), .A2(n7595), .ZN(n4688) );
  INV_X1 U5210 ( .A(n7698), .ZN(n4695) );
  OAI21_X1 U5211 ( .B1(n4666), .B2(n4667), .A(n4451), .ZN(n4665) );
  NOR2_X1 U5212 ( .A1(n4671), .A2(n8936), .ZN(n4667) );
  INV_X1 U5213 ( .A(n4672), .ZN(n4671) );
  INV_X1 U5214 ( .A(n4666), .ZN(n4663) );
  NAND2_X1 U5215 ( .A1(n4682), .A2(n4680), .ZN(n4679) );
  NOR2_X1 U5216 ( .A1(n4875), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U5217 ( .A1(n8957), .A2(n9082), .ZN(n4682) );
  OR2_X1 U5218 ( .A1(n9097), .A2(n9049), .ZN(n4681) );
  NOR2_X1 U5219 ( .A1(n4678), .A2(n8958), .ZN(n4677) );
  AND2_X1 U5220 ( .A1(n8955), .A2(n9049), .ZN(n4678) );
  NAND2_X1 U5221 ( .A1(n7716), .A2(n7738), .ZN(n4517) );
  INV_X1 U5222 ( .A(n4655), .ZN(n4650) );
  INV_X1 U5223 ( .A(n4651), .ZN(n4648) );
  NAND2_X1 U5224 ( .A1(n4651), .A2(n4647), .ZN(n4646) );
  INV_X1 U5225 ( .A(n4653), .ZN(n4647) );
  AND2_X1 U5226 ( .A1(n9098), .A2(n9004), .ZN(n4659) );
  INV_X1 U5227 ( .A(n4968), .ZN(n4967) );
  OAI21_X1 U5228 ( .B1(n5644), .B2(n4969), .A(n5658), .ZN(n4968) );
  INV_X1 U5229 ( .A(n5646), .ZN(n4969) );
  NOR2_X1 U5230 ( .A1(n4896), .A2(n5053), .ZN(n4895) );
  INV_X1 U5231 ( .A(n7953), .ZN(n4896) );
  INV_X1 U5232 ( .A(n4897), .ZN(n4893) );
  NAND2_X1 U5233 ( .A1(n6257), .A2(n5223), .ZN(n4599) );
  AOI21_X1 U5234 ( .B1(n5073), .B2(n5223), .A(n9915), .ZN(n4600) );
  INV_X1 U5235 ( .A(n7298), .ZN(n5031) );
  NOR2_X1 U5236 ( .A1(n5031), .A2(n4530), .ZN(n4526) );
  INV_X1 U5237 ( .A(n4526), .ZN(n4525) );
  INV_X1 U5238 ( .A(n7440), .ZN(n4906) );
  AND2_X1 U5239 ( .A1(n4705), .A2(n4706), .ZN(n7742) );
  OAI21_X1 U5240 ( .B1(n4709), .B2(n4708), .A(n4707), .ZN(n4706) );
  INV_X1 U5241 ( .A(n7733), .ZN(n4707) );
  NAND2_X1 U5242 ( .A1(n9877), .A2(n6261), .ZN(n6262) );
  OR2_X1 U5243 ( .A1(n6705), .A2(n6840), .ZN(n4910) );
  AND2_X1 U5244 ( .A1(n4920), .A2(n4919), .ZN(n7490) );
  NAND2_X1 U5245 ( .A1(n7495), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4919) );
  OR2_X1 U5246 ( .A1(n8110), .A2(n4913), .ZN(n4912) );
  AND2_X1 U5247 ( .A1(n8111), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4913) );
  INV_X1 U5248 ( .A(n4777), .ZN(n4776) );
  OAI21_X1 U5249 ( .B1(n4779), .B2(n4778), .A(n7543), .ZN(n4777) );
  INV_X1 U5250 ( .A(n5512), .ZN(n4778) );
  NAND2_X1 U5251 ( .A1(n5492), .A2(n5491), .ZN(n5505) );
  INV_X1 U5252 ( .A(n5493), .ZN(n5492) );
  OR2_X1 U5253 ( .A1(n8082), .A2(n9946), .ZN(n7650) );
  NAND2_X1 U5254 ( .A1(n4790), .A2(n4430), .ZN(n4786) );
  NOR2_X1 U5255 ( .A1(n7875), .A2(n8236), .ZN(n7727) );
  NAND2_X1 U5256 ( .A1(n4994), .A2(n8299), .ZN(n4991) );
  OR2_X1 U5257 ( .A1(n8469), .A2(n8298), .ZN(n7710) );
  NOR2_X1 U5258 ( .A1(n4448), .A2(n4977), .ZN(n4976) );
  INV_X1 U5259 ( .A(n7595), .ZN(n4977) );
  INV_X1 U5260 ( .A(n7682), .ZN(n4978) );
  INV_X1 U5261 ( .A(n7596), .ZN(n4973) );
  NAND2_X1 U5262 ( .A1(n8576), .A2(n8064), .ZN(n7689) );
  OR2_X1 U5263 ( .A1(n8576), .A2(n8064), .ZN(n7687) );
  NOR2_X1 U5264 ( .A1(n8581), .A2(n8396), .ZN(n7559) );
  INV_X1 U5265 ( .A(n6520), .ZN(n6510) );
  NAND2_X1 U5266 ( .A1(n8754), .A2(n8644), .ZN(n8648) );
  NAND2_X1 U5267 ( .A1(n6503), .A2(n6520), .ZN(n6532) );
  NAND2_X1 U5268 ( .A1(n4735), .A2(n4520), .ZN(n8783) );
  NAND2_X1 U5269 ( .A1(n8711), .A2(n7796), .ZN(n4735) );
  NAND2_X1 U5270 ( .A1(n4521), .A2(n8709), .ZN(n4520) );
  OR2_X1 U5271 ( .A1(n9375), .A2(n8880), .ZN(n8976) );
  NAND2_X1 U5272 ( .A1(n9399), .A2(n4872), .ZN(n4871) );
  OR2_X1 U5273 ( .A1(n9595), .A2(n8777), .ZN(n9089) );
  OR2_X1 U5274 ( .A1(n9407), .A2(n8850), .ZN(n8971) );
  INV_X1 U5275 ( .A(n6055), .ZN(n4839) );
  NOR2_X1 U5276 ( .A1(n4583), .A2(n8961), .ZN(n6065) );
  OR2_X1 U5277 ( .A1(n9637), .A2(n8889), .ZN(n8947) );
  OR2_X1 U5278 ( .A1(n9647), .A2(n8892), .ZN(n8939) );
  NOR2_X1 U5279 ( .A1(n8862), .A2(n7194), .ZN(n4578) );
  AND2_X1 U5280 ( .A1(n5954), .A2(n9827), .ZN(n4579) );
  AND2_X1 U5281 ( .A1(n9055), .A2(n4541), .ZN(n4866) );
  INV_X1 U5282 ( .A(n9029), .ZN(n4541) );
  OR2_X1 U5283 ( .A1(n8731), .A2(n5953), .ZN(n9054) );
  OAI21_X1 U5284 ( .B1(n6738), .B2(n8906), .A(n8911), .ZN(n9062) );
  NOR2_X1 U5285 ( .A1(n7029), .A2(n9804), .ZN(n7028) );
  OAI21_X1 U5286 ( .B1(n7524), .B2(n7523), .A(n7522), .ZN(n7536) );
  XNOR2_X1 U5287 ( .A(n5770), .B(n10296), .ZN(n5773) );
  NAND2_X1 U5288 ( .A1(n5608), .A2(n5607), .ZN(n5625) );
  NAND2_X1 U5289 ( .A1(n5606), .A2(n5605), .ZN(n5608) );
  NAND2_X1 U5290 ( .A1(n5587), .A2(n5586), .ZN(n5606) );
  NAND2_X1 U5291 ( .A1(n5585), .A2(n5584), .ZN(n5587) );
  AND3_X1 U5292 ( .A1(n10053), .A2(n5789), .A3(n5794), .ZN(n5769) );
  NAND2_X1 U5293 ( .A1(n5391), .A2(n5154), .ZN(n5405) );
  NOR2_X1 U5294 ( .A1(n4954), .A2(n4701), .ZN(n4700) );
  INV_X1 U5295 ( .A(n4955), .ZN(n4954) );
  INV_X1 U5296 ( .A(n4702), .ZN(n4701) );
  INV_X1 U5297 ( .A(n4957), .ZN(n4953) );
  INV_X1 U5298 ( .A(n5150), .ZN(n4952) );
  NAND2_X1 U5299 ( .A1(n4700), .A2(n4698), .ZN(n4697) );
  INV_X1 U5300 ( .A(n5332), .ZN(n4698) );
  NAND2_X1 U5301 ( .A1(n5151), .A2(SI_13_), .ZN(n5154) );
  NOR2_X1 U5302 ( .A1(n5370), .A2(n4958), .ZN(n4957) );
  INV_X1 U5303 ( .A(n5144), .ZN(n4958) );
  XNOR2_X1 U5304 ( .A(n5134), .B(SI_8_), .ZN(n5323) );
  NAND2_X1 U5305 ( .A1(n5113), .A2(SI_4_), .ZN(n5117) );
  INV_X1 U5306 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5765) );
  INV_X1 U5307 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5308 ( .A1(n7753), .A2(n7598), .ZN(n7739) );
  OR2_X1 U5309 ( .A1(n5505), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U5310 ( .A1(n5089), .A2(n5088), .ZN(n5430) );
  INV_X1 U5311 ( .A(n5428), .ZN(n5089) );
  OR2_X1 U5312 ( .A1(n5430), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5451) );
  INV_X1 U5313 ( .A(n7988), .ZN(n4890) );
  INV_X1 U5314 ( .A(n7987), .ZN(n4887) );
  NAND2_X1 U5315 ( .A1(n7952), .A2(n7953), .ZN(n7951) );
  XNOR2_X1 U5316 ( .A(n6903), .B(n5196), .ZN(n6631) );
  AND4_X1 U5317 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n7198)
         );
  OR2_X1 U5318 ( .A1(n5208), .A2(n5280), .ZN(n5286) );
  NAND2_X1 U5319 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  INV_X1 U5320 ( .A(n6262), .ZN(n4614) );
  NAND2_X1 U5321 ( .A1(n6262), .A2(n6481), .ZN(n6265) );
  NOR2_X1 U5322 ( .A1(n6233), .A2(n6234), .ZN(n6698) );
  NOR2_X1 U5323 ( .A1(n6700), .A2(n6701), .ZN(n6839) );
  INV_X1 U5324 ( .A(n6994), .ZN(n4918) );
  AND2_X1 U5325 ( .A1(n4915), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U5326 ( .A1(n6995), .A2(n6994), .ZN(n4916) );
  OAI21_X1 U5327 ( .B1(n7110), .B2(n7259), .A(n7109), .ZN(n7111) );
  NAND2_X1 U5328 ( .A1(n7110), .A2(n7259), .ZN(n7109) );
  NAND2_X1 U5329 ( .A1(n7258), .A2(n7259), .ZN(n4926) );
  AND2_X1 U5330 ( .A1(n7380), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4822) );
  NOR2_X1 U5331 ( .A1(n7469), .A2(n7470), .ZN(n7473) );
  OR2_X1 U5332 ( .A1(n7473), .A2(n7472), .ZN(n4920) );
  XNOR2_X1 U5333 ( .A(n7490), .B(n8097), .ZN(n8093) );
  XNOR2_X1 U5334 ( .A(n4912), .B(n4911), .ZN(n8113) );
  INV_X1 U5335 ( .A(n8138), .ZN(n4911) );
  NOR2_X1 U5336 ( .A1(n8113), .A2(n8112), .ZN(n8139) );
  AOI21_X1 U5337 ( .B1(n4413), .B2(n10199), .A(n8127), .ZN(n4820) );
  AOI21_X1 U5338 ( .B1(n8207), .B2(n8206), .A(n8205), .ZN(n8211) );
  NAND2_X1 U5339 ( .A1(n5635), .A2(n5634), .ZN(n5649) );
  INV_X1 U5340 ( .A(n5636), .ZN(n5635) );
  NAND2_X1 U5341 ( .A1(n8072), .A2(n8410), .ZN(n7846) );
  AND2_X1 U5342 ( .A1(n5621), .A2(n5620), .ZN(n8264) );
  NAND2_X1 U5343 ( .A1(n5595), .A2(n5594), .ZN(n5615) );
  INV_X1 U5344 ( .A(n5596), .ZN(n5595) );
  OR2_X1 U5345 ( .A1(n5556), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5575) );
  NOR2_X1 U5346 ( .A1(n8321), .A2(n4780), .ZN(n4779) );
  INV_X1 U5347 ( .A(n5049), .ZN(n4780) );
  AND2_X1 U5348 ( .A1(n7589), .A2(n8309), .ZN(n8321) );
  OR2_X1 U5349 ( .A1(n5469), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5493) );
  OR2_X1 U5350 ( .A1(n5457), .A2(n8346), .ZN(n5048) );
  AND4_X1 U5351 ( .A1(n5498), .A2(n5497), .A3(n5496), .A4(n5495), .ZN(n8347)
         );
  AND2_X1 U5352 ( .A1(n5705), .A2(n7700), .ZN(n5008) );
  NAND2_X1 U5353 ( .A1(n5087), .A2(n10200), .ZN(n5411) );
  INV_X1 U5354 ( .A(n5397), .ZN(n5087) );
  AND2_X1 U5355 ( .A1(n5182), .A2(n5181), .ZN(n7670) );
  AND4_X1 U5356 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n8441)
         );
  AOI21_X1 U5357 ( .B1(n4803), .B2(n4801), .A(n4470), .ZN(n4800) );
  INV_X1 U5358 ( .A(n4806), .ZN(n4801) );
  AND4_X1 U5359 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n8429)
         );
  NAND2_X1 U5360 ( .A1(n7216), .A2(n5057), .ZN(n7214) );
  OR2_X1 U5361 ( .A1(n8082), .A2(n7868), .ZN(n7215) );
  NAND2_X1 U5362 ( .A1(n5083), .A2(n7000), .ZN(n5317) );
  INV_X1 U5363 ( .A(n5301), .ZN(n5083) );
  NAND2_X1 U5364 ( .A1(n7139), .A2(n7628), .ZN(n4997) );
  NAND2_X1 U5365 ( .A1(n7650), .A2(n7211), .ZN(n7642) );
  NAND2_X1 U5366 ( .A1(n7161), .A2(n7642), .ZN(n7216) );
  NAND2_X1 U5367 ( .A1(n5082), .A2(n5081), .ZN(n5281) );
  INV_X1 U5368 ( .A(n5264), .ZN(n5082) );
  NAND2_X1 U5369 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  NAND2_X1 U5370 ( .A1(n7611), .A2(n7612), .ZN(n9901) );
  NAND2_X1 U5371 ( .A1(n5819), .A2(n7533), .ZN(n4882) );
  AND2_X1 U5372 ( .A1(n7534), .A2(n5189), .ZN(n7579) );
  NAND2_X1 U5373 ( .A1(n5663), .A2(n5662), .ZN(n5750) );
  AND2_X1 U5374 ( .A1(n5648), .A2(n5647), .ZN(n7565) );
  NAND2_X1 U5375 ( .A1(n4785), .A2(n4430), .ZN(n4784) );
  INV_X1 U5376 ( .A(n4788), .ZN(n4785) );
  AOI21_X1 U5377 ( .B1(n4789), .B2(n4790), .A(n4459), .ZN(n4788) );
  XNOR2_X1 U5378 ( .A(n7565), .B(n7916), .ZN(n8234) );
  OR2_X1 U5379 ( .A1(n7727), .A2(n7726), .ZN(n7843) );
  NOR2_X1 U5380 ( .A1(n8537), .A2(n8284), .ZN(n5583) );
  NAND2_X1 U5381 ( .A1(n4986), .A2(n7718), .ZN(n4985) );
  INV_X1 U5382 ( .A(n4983), .ZN(n4982) );
  INV_X1 U5383 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U5384 ( .A1(n4988), .A2(n7713), .ZN(n4987) );
  NAND2_X1 U5385 ( .A1(n4989), .A2(n4992), .ZN(n4988) );
  INV_X1 U5386 ( .A(n4994), .ZN(n4992) );
  NAND2_X1 U5387 ( .A1(n7718), .A2(n7717), .ZN(n8267) );
  AND2_X1 U5388 ( .A1(n7710), .A2(n4995), .ZN(n4994) );
  AND2_X1 U5389 ( .A1(n7710), .A2(n7709), .ZN(n8285) );
  NAND2_X1 U5390 ( .A1(n8300), .A2(n8295), .ZN(n4996) );
  NAND2_X1 U5391 ( .A1(n7305), .A2(n7537), .ZN(n5541) );
  NAND2_X1 U5392 ( .A1(n8330), .A2(n8331), .ZN(n8337) );
  OR2_X1 U5393 ( .A1(n6652), .A2(n7739), .ZN(n9910) );
  OAI22_X1 U5394 ( .A1(n8394), .A2(n5418), .B1(n8411), .B2(n8587), .ZN(n8384)
         );
  NAND2_X1 U5395 ( .A1(n5702), .A2(n5701), .ZN(n8403) );
  INV_X1 U5396 ( .A(n9910), .ZN(n8408) );
  AND3_X1 U5397 ( .A1(n5244), .A2(n5243), .A3(n5242), .ZN(n9927) );
  AND2_X1 U5398 ( .A1(n5070), .A2(n5000), .ZN(n4760) );
  NAND2_X1 U5399 ( .A1(n5712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5714) );
  INV_X1 U5400 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n10177) );
  OAI21_X1 U5401 ( .B1(n6257), .B2(n5073), .A(n5223), .ZN(n4818) );
  NAND2_X1 U5402 ( .A1(n4817), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U5403 ( .A1(n5073), .A2(n5223), .ZN(n4816) );
  NAND2_X1 U5404 ( .A1(n7793), .A2(n4736), .ZN(n8711) );
  OR2_X1 U5405 ( .A1(n7828), .A2(n7827), .ZN(n8628) );
  OR2_X1 U5406 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  NAND2_X1 U5407 ( .A1(n8614), .A2(n7181), .ZN(n7184) );
  AND3_X1 U5408 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U5409 ( .A1(n4527), .A2(n4529), .ZN(n7295) );
  NAND3_X1 U5410 ( .A1(n7185), .A2(n4748), .A3(n7295), .ZN(n7296) );
  INV_X1 U5411 ( .A(n7188), .ZN(n4748) );
  NOR2_X1 U5412 ( .A1(n5033), .A2(n8831), .ZN(n5032) );
  INV_X1 U5413 ( .A(n8632), .ZN(n5033) );
  AND2_X1 U5414 ( .A1(n5021), .A2(n4537), .ZN(n4536) );
  AND2_X1 U5415 ( .A1(n8762), .A2(n5022), .ZN(n5021) );
  NAND2_X1 U5416 ( .A1(n8856), .A2(n5023), .ZN(n5022) );
  INV_X1 U5417 ( .A(n8857), .ZN(n5023) );
  INV_X1 U5418 ( .A(n8856), .ZN(n5024) );
  OR2_X1 U5419 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U5420 ( .A1(n8648), .A2(n8647), .ZN(n8719) );
  INV_X1 U5421 ( .A(n6507), .ZN(n4532) );
  NAND2_X1 U5422 ( .A1(n8726), .A2(n4538), .ZN(n4537) );
  INV_X1 U5423 ( .A(n7773), .ZN(n4538) );
  NAND2_X1 U5424 ( .A1(n6815), .A2(n4452), .ZN(n6830) );
  AND2_X1 U5425 ( .A1(n7169), .A2(n6826), .ZN(n6829) );
  OAI21_X1 U5426 ( .B1(n8670), .B2(n4741), .A(n4533), .ZN(n8771) );
  INV_X1 U5427 ( .A(n4534), .ZN(n4533) );
  OAI21_X1 U5428 ( .B1(n8819), .B2(n4741), .A(n8773), .ZN(n4534) );
  OR2_X1 U5429 ( .A1(n6131), .A2(n6833), .ZN(n5888) );
  OR2_X1 U5430 ( .A1(n6125), .A2(n6385), .ZN(n5878) );
  NAND2_X1 U5431 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U5432 ( .A1(n7851), .A2(n9701), .ZN(n5841) );
  NAND2_X1 U5433 ( .A1(n6340), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5816) );
  OR2_X1 U5434 ( .A1(n9762), .A2(n9761), .ZN(n4721) );
  AND2_X1 U5435 ( .A1(n4721), .A2(n4720), .ZN(n9781) );
  NAND2_X1 U5436 ( .A1(n9248), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4720) );
  OR2_X1 U5437 ( .A1(n9781), .A2(n9780), .ZN(n4719) );
  NOR2_X1 U5438 ( .A1(n9314), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5439 ( .A1(n4588), .A2(n9356), .ZN(n4587) );
  INV_X1 U5440 ( .A(n4590), .ZN(n4588) );
  AOI21_X1 U5441 ( .B1(n9382), .B2(n6102), .A(n6101), .ZN(n9365) );
  NAND2_X1 U5442 ( .A1(n9407), .A2(n8850), .ZN(n9390) );
  NOR2_X1 U5443 ( .A1(n9415), .A2(n9407), .ZN(n9383) );
  INV_X1 U5444 ( .A(n4436), .ZN(n4844) );
  OR2_X1 U5445 ( .A1(n9625), .A2(n9492), .ZN(n6042) );
  AND2_X1 U5446 ( .A1(n4879), .A2(n8952), .ZN(n4878) );
  INV_X1 U5447 ( .A(n9485), .ZN(n4879) );
  NAND2_X1 U5448 ( .A1(n9490), .A2(n9495), .ZN(n4880) );
  AND2_X1 U5449 ( .A1(n8947), .A2(n9076), .ZN(n9511) );
  AND2_X1 U5450 ( .A1(n9525), .A2(n8926), .ZN(n4861) );
  AND2_X1 U5451 ( .A1(n9548), .A2(n8926), .ZN(n9526) );
  NAND2_X1 U5452 ( .A1(n4549), .A2(n4548), .ZN(n9545) );
  INV_X1 U5453 ( .A(n4550), .ZN(n4548) );
  OAI21_X1 U5454 ( .B1(n4554), .B2(n4551), .A(n8937), .ZN(n4550) );
  NAND2_X1 U5455 ( .A1(n4863), .A2(n4862), .ZN(n9548) );
  INV_X1 U5456 ( .A(n9545), .ZN(n4863) );
  NAND2_X1 U5457 ( .A1(n4555), .A2(n4554), .ZN(n7224) );
  INV_X1 U5458 ( .A(n7226), .ZN(n4555) );
  AND2_X1 U5459 ( .A1(n9029), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5460 ( .A1(n4834), .A2(n5934), .ZN(n4833) );
  INV_X1 U5461 ( .A(n6937), .ZN(n4834) );
  INV_X1 U5462 ( .A(n5934), .ZN(n4835) );
  NAND2_X1 U5463 ( .A1(n9054), .A2(n8930), .ZN(n9029) );
  NAND2_X1 U5464 ( .A1(n5925), .A2(n5924), .ZN(n7294) );
  NAND2_X1 U5465 ( .A1(n6946), .A2(n5921), .ZN(n6938) );
  NAND2_X1 U5466 ( .A1(n6938), .A2(n6937), .ZN(n6936) );
  NAND2_X1 U5467 ( .A1(n6947), .A2(n6948), .ZN(n6946) );
  NAND2_X1 U5468 ( .A1(n6552), .A2(n6807), .ZN(n5861) );
  NAND2_X1 U5469 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U5470 ( .A1(n6160), .A2(n6159), .ZN(n6727) );
  NAND2_X1 U5471 ( .A1(n6276), .A2(n5831), .ZN(n6724) );
  OR2_X1 U5472 ( .A1(n9057), .A2(n6890), .ZN(n5831) );
  NAND2_X1 U5473 ( .A1(n6724), .A2(n9016), .ZN(n6723) );
  OR2_X1 U5474 ( .A1(n6498), .A2(n6208), .ZN(n6284) );
  OR2_X1 U5475 ( .A1(n9049), .A2(n9137), .ZN(n9651) );
  NAND2_X1 U5476 ( .A1(n6278), .A2(n9651), .ZN(n9836) );
  NOR2_X1 U5477 ( .A1(n4425), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5038) );
  INV_X1 U5478 ( .A(n5773), .ZN(n5772) );
  NAND2_X1 U5479 ( .A1(n5627), .A2(n5626), .ZN(n5645) );
  NAND2_X1 U5480 ( .A1(n5625), .A2(n5624), .ZN(n5627) );
  XNOR2_X1 U5481 ( .A(n5645), .B(n5644), .ZN(n7458) );
  XNOR2_X1 U5482 ( .A(n5625), .B(n5624), .ZN(n7452) );
  NAND2_X1 U5483 ( .A1(n6185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U5484 ( .A1(n6188), .A2(n6190), .ZN(n6185) );
  XNOR2_X1 U5485 ( .A(n5606), .B(n5605), .ZN(n7446) );
  XNOR2_X1 U5486 ( .A(n5585), .B(n5584), .ZN(n7422) );
  OAI21_X1 U5487 ( .B1(n5441), .B2(n4945), .A(n4942), .ZN(n5501) );
  NAND2_X1 U5488 ( .A1(n4946), .A2(n4947), .ZN(n5480) );
  NAND2_X1 U5489 ( .A1(n5441), .A2(n4949), .ZN(n4946) );
  XNOR2_X1 U5490 ( .A(n5441), .B(n5158), .ZN(n6599) );
  NAND2_X1 U5491 ( .A1(n5150), .A2(n5149), .ZN(n5172) );
  INV_X1 U5492 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4566) );
  INV_X1 U5493 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4565) );
  INV_X1 U5494 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5495 ( .A1(n4622), .A2(n5869), .ZN(n5015) );
  NOR2_X1 U5496 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4622) );
  NOR2_X2 U5497 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5936) );
  NAND2_X1 U5498 ( .A1(n4704), .A2(n4702), .ZN(n5355) );
  NAND2_X1 U5499 ( .A1(n4558), .A2(n4561), .ZN(n4704) );
  AND2_X1 U5500 ( .A1(n5127), .A2(n5126), .ZN(n5288) );
  NAND2_X1 U5501 ( .A1(n5259), .A2(n5117), .ZN(n5275) );
  AND2_X1 U5502 ( .A1(n5122), .A2(n5121), .ZN(n5274) );
  AND3_X1 U5503 ( .A1(n5017), .A2(n5765), .A3(n5016), .ZN(n5868) );
  NOR2_X1 U5504 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4717) );
  AND3_X1 U5505 ( .A1(n5546), .A2(n5545), .A3(n5544), .ZN(n8308) );
  NAND2_X1 U5506 ( .A1(n4497), .A2(n6679), .ZN(n6680) );
  AND4_X1 U5507 ( .A1(n5511), .A2(n5510), .A3(n5509), .A4(n5508), .ZN(n8334)
         );
  NAND2_X1 U5508 ( .A1(n5504), .A2(n5503), .ZN(n8323) );
  INV_X1 U5509 ( .A(n8256), .ZN(n8236) );
  OR2_X1 U5510 ( .A1(n6653), .A2(n6654), .ZN(n8063) );
  AND2_X1 U5511 ( .A1(n6924), .A2(n5669), .ZN(n8237) );
  INV_X1 U5512 ( .A(n8334), .ZN(n8077) );
  NAND4_X1 U5513 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n8080)
         );
  AND4_X1 U5514 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n7427)
         );
  OR2_X1 U5515 ( .A1(n5210), .A2(n7339), .ZN(n5347) );
  INV_X1 U5516 ( .A(n7198), .ZN(n8083) );
  OR2_X1 U5517 ( .A1(n5199), .A2(n6227), .ZN(n5202) );
  OR2_X1 U5518 ( .A1(n5210), .A2(n5198), .ZN(n5203) );
  NAND2_X1 U5519 ( .A1(n9890), .A2(n9891), .ZN(n9889) );
  NAND2_X1 U5520 ( .A1(n7103), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7257) );
  OR2_X1 U5521 ( .A1(n8104), .A2(n10199), .ZN(n4821) );
  NOR2_X1 U5522 ( .A1(n4621), .A2(n8194), .ZN(n4620) );
  INV_X1 U5523 ( .A(n8198), .ZN(n4621) );
  INV_X1 U5524 ( .A(n7670), .ZN(n8509) );
  NAND2_X1 U5525 ( .A1(n5377), .A2(n5376), .ZN(n9971) );
  NAND2_X1 U5526 ( .A1(n5695), .A2(n7648), .ZN(n7332) );
  AND3_X1 U5527 ( .A1(n5297), .A2(n5296), .A3(n5295), .ZN(n9942) );
  NAND2_X1 U5528 ( .A1(n4763), .A2(n4420), .ZN(n4764) );
  INV_X1 U5529 ( .A(n5750), .ZN(n7855) );
  NAND2_X1 U5530 ( .A1(n5069), .A2(n5068), .ZN(n5675) );
  AOI21_X1 U5531 ( .B1(n8820), .B2(n4428), .A(n4738), .ZN(n8744) );
  NAND2_X1 U5532 ( .A1(n8701), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5533 ( .A1(n4428), .A2(n4742), .ZN(n4739) );
  OR2_X1 U5534 ( .A1(n8749), .A2(n5035), .ZN(n5034) );
  NAND2_X1 U5535 ( .A1(n5037), .A2(n5036), .ZN(n5035) );
  INV_X1 U5536 ( .A(n8748), .ZN(n5037) );
  NOR2_X1 U5537 ( .A1(n8696), .A2(n8695), .ZN(n8748) );
  NAND2_X1 U5538 ( .A1(n9704), .A2(n8998), .ZN(n6123) );
  NAND2_X1 U5539 ( .A1(n6024), .A2(n6023), .ZN(n9498) );
  NAND2_X1 U5540 ( .A1(n6558), .A2(n6559), .ZN(n6815) );
  AND2_X1 U5541 ( .A1(n6560), .A2(n6561), .ZN(n6558) );
  NAND2_X1 U5542 ( .A1(n6048), .A2(n6047), .ZN(n9614) );
  INV_X1 U5543 ( .A(n9529), .ZN(n8892) );
  NAND2_X1 U5544 ( .A1(n6012), .A2(n6011), .ZN(n9535) );
  AND2_X1 U5545 ( .A1(n9218), .A2(n4726), .ZN(n6407) );
  NAND2_X1 U5546 ( .A1(n6371), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U5547 ( .A1(n9292), .A2(n4732), .ZN(n4731) );
  INV_X1 U5548 ( .A(n4733), .ZN(n4732) );
  OAI21_X1 U5549 ( .B1(n9293), .B2(n10319), .A(n9769), .ZN(n4733) );
  OAI22_X1 U5550 ( .A1(n9295), .A2(n10323), .B1(n10319), .B2(n9294), .ZN(n4729) );
  AOI21_X1 U5551 ( .B1(n6176), .B2(n9523), .A(n6175), .ZN(n9321) );
  XNOR2_X1 U5552 ( .A(n4540), .B(n8992), .ZN(n6176) );
  AND2_X1 U5553 ( .A1(n4507), .A2(n4505), .ZN(n9576) );
  AOI21_X1 U5554 ( .B1(n9330), .B2(n9528), .A(n4506), .ZN(n4505) );
  NAND2_X1 U5555 ( .A1(n9331), .A2(n9523), .ZN(n4507) );
  AND2_X1 U5556 ( .A1(n9360), .A2(n9530), .ZN(n4506) );
  OAI21_X1 U5557 ( .B1(n4431), .B2(n4824), .A(n9322), .ZN(n9577) );
  NAND2_X1 U5558 ( .A1(n4829), .A2(n6114), .ZN(n9340) );
  NAND2_X1 U5559 ( .A1(n9349), .A2(n9348), .ZN(n4829) );
  AND2_X1 U5560 ( .A1(n9342), .A2(n4439), .ZN(n9580) );
  NAND2_X1 U5561 ( .A1(n5970), .A2(n5969), .ZN(n8768) );
  OR2_X1 U5562 ( .A1(n6366), .A2(n5979), .ZN(n5970) );
  NAND2_X1 U5563 ( .A1(n5893), .A2(n5892), .ZN(n6961) );
  NAND2_X1 U5564 ( .A1(n5793), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5795) );
  OAI21_X1 U5565 ( .B1(n5690), .B2(n7601), .A(n7606), .ZN(n7602) );
  NAND2_X1 U5566 ( .A1(n4635), .A2(n4631), .ZN(n8916) );
  OAI21_X1 U5567 ( .B1(n4637), .B2(n4466), .A(n4636), .ZN(n4635) );
  OAI21_X1 U5568 ( .B1(n4634), .B2(n4633), .A(n4632), .ZN(n4631) );
  AND2_X1 U5569 ( .A1(n7687), .A2(n4686), .ZN(n4685) );
  AOI21_X1 U5570 ( .B1(n4673), .B2(n8925), .A(n4472), .ZN(n4672) );
  OAI22_X1 U5571 ( .A1(n7699), .A2(n7739), .B1(n7738), .B2(n4694), .ZN(n4693)
         );
  AOI21_X1 U5572 ( .B1(n7708), .B2(n4695), .A(n4468), .ZN(n4694) );
  NOR2_X1 U5573 ( .A1(n7593), .A2(n7738), .ZN(n4691) );
  INV_X1 U5574 ( .A(n4665), .ZN(n4664) );
  NOR2_X1 U5575 ( .A1(n4661), .A2(n4654), .ZN(n4653) );
  NOR2_X1 U5576 ( .A1(n8959), .A2(n4676), .ZN(n8966) );
  NAND2_X1 U5577 ( .A1(n4679), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5578 ( .A1(n4518), .A2(n4517), .ZN(n7720) );
  NAND2_X1 U5579 ( .A1(n7731), .A2(n7739), .ZN(n4502) );
  NAND2_X1 U5580 ( .A1(n7730), .A2(n7738), .ZN(n4503) );
  AND2_X1 U5581 ( .A1(n4712), .A2(n7735), .ZN(n4708) );
  INV_X1 U5582 ( .A(n8537), .ZN(n5708) );
  AND2_X1 U5583 ( .A1(n4736), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U5584 ( .A1(n4644), .A2(n4648), .ZN(n4641) );
  NAND2_X1 U5585 ( .A1(n4427), .A2(n4650), .ZN(n4640) );
  NAND2_X1 U5586 ( .A1(n4645), .A2(n4643), .ZN(n4642) );
  INV_X1 U5587 ( .A(n4427), .ZN(n4643) );
  NAND2_X1 U5588 ( .A1(n4870), .A2(n9089), .ZN(n4869) );
  AOI21_X1 U5589 ( .B1(n4967), .B2(n4969), .A(n4493), .ZN(n4964) );
  INV_X1 U5590 ( .A(n5500), .ZN(n4941) );
  INV_X1 U5591 ( .A(SI_14_), .ZN(n4932) );
  INV_X1 U5592 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5096) );
  NAND2_X1 U5593 ( .A1(n4893), .A2(n4899), .ZN(n4892) );
  NAND2_X1 U5594 ( .A1(n4602), .A2(n4601), .ZN(n9879) );
  NAND2_X1 U5595 ( .A1(n4815), .A2(n4598), .ZN(n4602) );
  AND2_X1 U5596 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U5597 ( .A1(n9878), .A2(n9879), .ZN(n9877) );
  NAND2_X1 U5598 ( .A1(n4612), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5599 ( .A1(n4910), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4604) );
  AND3_X1 U5600 ( .A1(n4606), .A2(n4607), .A3(n4491), .ZN(n7467) );
  OR2_X1 U5601 ( .A1(n5750), .A2(n8237), .ZN(n7540) );
  NOR2_X1 U5602 ( .A1(n5622), .A2(n4792), .ZN(n4791) );
  INV_X1 U5603 ( .A(n8267), .ZN(n4792) );
  NAND2_X1 U5604 ( .A1(n5084), .A2(n7112), .ZN(n5362) );
  INV_X1 U5605 ( .A(n5343), .ZN(n5084) );
  AND2_X1 U5606 ( .A1(n7048), .A2(n7633), .ZN(n7621) );
  NAND2_X1 U5607 ( .A1(n6901), .A2(n9934), .ZN(n4771) );
  NAND2_X1 U5608 ( .A1(n8085), .A2(n8011), .ZN(n4772) );
  OR2_X1 U5609 ( .A1(n5246), .A2(n9927), .ZN(n7626) );
  INV_X1 U5610 ( .A(n4791), .ZN(n4789) );
  OAI21_X1 U5611 ( .B1(n4987), .B2(n4984), .A(n7717), .ZN(n4983) );
  NAND2_X1 U5612 ( .A1(n4990), .A2(n7718), .ZN(n4984) );
  NAND4_X1 U5613 ( .A1(n5325), .A2(n5293), .A3(n5337), .A4(n5062), .ZN(n5063)
         );
  NAND2_X1 U5614 ( .A1(n4737), .A2(n7792), .ZN(n4736) );
  INV_X1 U5615 ( .A(n7794), .ZN(n4737) );
  AND2_X1 U5616 ( .A1(n6532), .A2(n6530), .ZN(n6527) );
  INV_X1 U5617 ( .A(n5030), .ZN(n5029) );
  OAI21_X1 U5618 ( .B1(n4528), .B2(n4525), .A(n4524), .ZN(n5030) );
  AOI21_X1 U5619 ( .B1(n4526), .B2(n4531), .A(n4456), .ZN(n4524) );
  AND2_X1 U5620 ( .A1(n7307), .A2(n9143), .ZN(n9004) );
  OR2_X1 U5621 ( .A1(n9574), .A2(n8979), .ZN(n9114) );
  NAND2_X1 U5622 ( .A1(n5885), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5900) );
  AND2_X1 U5623 ( .A1(n4719), .A2(n4718), .ZN(n9251) );
  NAND2_X1 U5624 ( .A1(n9784), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5625 ( .A1(n9574), .A2(n8979), .ZN(n9111) );
  NAND2_X1 U5626 ( .A1(n9335), .A2(n9112), .ZN(n9328) );
  NAND2_X1 U5627 ( .A1(n9328), .A2(n9329), .ZN(n9327) );
  NOR2_X1 U5628 ( .A1(n4869), .A2(n4547), .ZN(n4546) );
  INV_X1 U5629 ( .A(n9401), .ZN(n4547) );
  INV_X1 U5630 ( .A(n8967), .ZN(n4544) );
  INV_X1 U5631 ( .A(n4869), .ZN(n4868) );
  AND2_X1 U5632 ( .A1(n4584), .A2(n4583), .ZN(n4582) );
  NOR2_X1 U5633 ( .A1(n9614), .A2(n9470), .ZN(n4584) );
  OR2_X1 U5634 ( .A1(n9614), .A2(n7838), .ZN(n8964) );
  NOR2_X1 U5635 ( .A1(n4852), .A2(n4855), .ZN(n4848) );
  NAND2_X1 U5636 ( .A1(n4850), .A2(n6032), .ZN(n4849) );
  NOR2_X1 U5637 ( .A1(n9535), .A2(n9647), .ZN(n4574) );
  NOR2_X1 U5638 ( .A1(n5999), .A2(n5998), .ZN(n6013) );
  INV_X1 U5639 ( .A(n9070), .ZN(n4553) );
  OR2_X1 U5640 ( .A1(n5986), .A2(n5985), .ZN(n5999) );
  OR2_X1 U5641 ( .A1(n5946), .A2(n8727), .ZN(n5960) );
  NOR2_X1 U5642 ( .A1(n5900), .A2(n5899), .ZN(n5915) );
  NOR2_X1 U5643 ( .A1(n6761), .A2(n6875), .ZN(n6736) );
  NAND2_X1 U5644 ( .A1(n6736), .A2(n6975), .ZN(n6797) );
  AOI21_X1 U5645 ( .B1(n4944), .B2(n4943), .A(n4489), .ZN(n4942) );
  INV_X1 U5646 ( .A(n4949), .ZN(n4943) );
  NOR2_X1 U5647 ( .A1(n5460), .A2(n4950), .ZN(n4949) );
  INV_X1 U5648 ( .A(n5439), .ZN(n4950) );
  AOI21_X1 U5649 ( .B1(n4949), .B2(n5440), .A(n4948), .ZN(n4947) );
  INV_X1 U5650 ( .A(n5459), .ZN(n4948) );
  INV_X1 U5651 ( .A(n5122), .ZN(n4962) );
  OAI21_X1 U5652 ( .B1(n5133), .B2(n4509), .A(n4508), .ZN(n5123) );
  NAND2_X1 U5653 ( .A1(n5133), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4508) );
  OR2_X1 U5654 ( .A1(n5880), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U5655 ( .B1(n5160), .B2(n5099), .A(n5098), .ZN(n5100) );
  NAND2_X1 U5656 ( .A1(n5160), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U5657 ( .A1(n5100), .A2(SI_3_), .ZN(n5112) );
  INV_X1 U5658 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7000) );
  AND2_X1 U5659 ( .A1(n7959), .A2(n7905), .ZN(n7997) );
  AND2_X1 U5660 ( .A1(n7863), .A2(n7203), .ZN(n7270) );
  NOR2_X1 U5661 ( .A1(n8027), .A2(n4898), .ZN(n4897) );
  INV_X1 U5662 ( .A(n7897), .ZN(n4898) );
  NAND2_X1 U5663 ( .A1(n5524), .A2(n5523), .ZN(n5542) );
  XNOR2_X1 U5664 ( .A(n6630), .B(n9923), .ZN(n6677) );
  AOI21_X1 U5665 ( .B1(n4905), .B2(n4904), .A(n4465), .ZN(n4903) );
  INV_X1 U5666 ( .A(n7438), .ZN(n4904) );
  OR2_X1 U5667 ( .A1(n6610), .A2(n5745), .ZN(n6646) );
  INV_X1 U5668 ( .A(n7741), .ZN(n4936) );
  AND4_X1 U5669 ( .A1(n5095), .A2(n5094), .A3(n5093), .A4(n5092), .ZN(n8064)
         );
  NAND4_X1 U5670 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n6579)
         );
  NAND2_X1 U5671 ( .A1(n9851), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U5672 ( .A1(n4610), .A2(n6265), .ZN(n6488) );
  INV_X1 U5673 ( .A(n4611), .ZN(n4610) );
  NAND2_X1 U5674 ( .A1(n4910), .A2(n6854), .ZN(n6707) );
  NAND2_X1 U5675 ( .A1(n4605), .A2(n6853), .ZN(n6995) );
  NAND2_X1 U5676 ( .A1(n4604), .A2(n6854), .ZN(n4605) );
  NAND2_X1 U5677 ( .A1(n4603), .A2(n6854), .ZN(n6856) );
  INV_X1 U5678 ( .A(n4604), .ZN(n4603) );
  NAND2_X1 U5679 ( .A1(n4500), .A2(n4499), .ZN(n4810) );
  INV_X1 U5680 ( .A(n4811), .ZN(n4500) );
  NOR2_X1 U5681 ( .A1(n7494), .A2(n4823), .ZN(n7496) );
  AND2_X1 U5682 ( .A1(n7495), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4823) );
  NOR2_X1 U5683 ( .A1(n8093), .A2(n5396), .ZN(n8092) );
  AOI21_X1 U5684 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8111), .A(n8103), .ZN(
        n8123) );
  INV_X1 U5685 ( .A(n4912), .ZN(n8137) );
  AND2_X1 U5686 ( .A1(n8152), .A2(n8151), .ZN(n8190) );
  INV_X1 U5687 ( .A(n5664), .ZN(n7853) );
  AOI21_X1 U5688 ( .B1(n4784), .B2(n4786), .A(n4455), .ZN(n4783) );
  OR2_X1 U5689 ( .A1(n5649), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5664) );
  OR2_X1 U5690 ( .A1(n5615), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U5691 ( .A1(n5574), .A2(n5573), .ZN(n5596) );
  INV_X1 U5692 ( .A(n5575), .ZN(n5574) );
  NAND2_X1 U5693 ( .A1(n4774), .A2(n4773), .ZN(n8296) );
  AOI21_X1 U5694 ( .B1(n4776), .B2(n4778), .A(n4454), .ZN(n4773) );
  NAND2_X1 U5695 ( .A1(n5450), .A2(n5449), .ZN(n5469) );
  INV_X1 U5696 ( .A(n5451), .ZN(n5450) );
  AND4_X1 U5697 ( .A1(n5456), .A2(n5455), .A3(n5454), .A4(n5453), .ZN(n8346)
         );
  NAND2_X1 U5698 ( .A1(n5086), .A2(n5085), .ZN(n5397) );
  INV_X1 U5699 ( .A(n5380), .ZN(n5086) );
  INV_X1 U5700 ( .A(n4795), .ZN(n8427) );
  NAND2_X1 U5701 ( .A1(n8438), .A2(n4803), .ZN(n4799) );
  AOI21_X1 U5702 ( .B1(n4798), .B2(n8438), .A(n4808), .ZN(n4797) );
  NAND2_X1 U5703 ( .A1(n7331), .A2(n5697), .ZN(n7429) );
  NAND2_X1 U5704 ( .A1(n7648), .A2(n7637), .ZN(n7550) );
  AOI21_X1 U5705 ( .B1(n7141), .B2(n5299), .A(n5298), .ZN(n7161) );
  NAND2_X1 U5706 ( .A1(n6772), .A2(n5080), .ZN(n5264) );
  INV_X1 U5707 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5708 ( .A1(n4770), .A2(n4771), .ZN(n7015) );
  NAND2_X1 U5709 ( .A1(n5262), .A2(n4772), .ZN(n4770) );
  AND2_X1 U5710 ( .A1(n7626), .A2(n7620), .ZN(n7546) );
  NOR2_X1 U5711 ( .A1(n5690), .A2(n6985), .ZN(n6986) );
  NAND2_X1 U5712 ( .A1(n4970), .A2(n7539), .ZN(n7577) );
  NAND2_X1 U5713 ( .A1(n8994), .A2(n7537), .ZN(n4970) );
  AND2_X1 U5714 ( .A1(n7721), .A2(n7542), .ZN(n8253) );
  INV_X1 U5715 ( .A(n8253), .ZN(n8251) );
  AND2_X1 U5716 ( .A1(n5603), .A2(n5602), .ZN(n8273) );
  NAND2_X1 U5717 ( .A1(n5555), .A2(n5554), .ZN(n8469) );
  AND4_X1 U5718 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n8335)
         );
  NAND2_X1 U5719 ( .A1(n7690), .A2(n7700), .ZN(n8359) );
  AOI21_X1 U5720 ( .B1(n4976), .B2(n4979), .A(n4973), .ZN(n4972) );
  NAND2_X1 U5721 ( .A1(n8403), .A2(n4976), .ZN(n4974) );
  INV_X1 U5722 ( .A(n7681), .ZN(n4979) );
  INV_X1 U5723 ( .A(n9909), .ZN(n8410) );
  INV_X1 U5724 ( .A(n7341), .ZN(n9955) );
  AND2_X1 U5725 ( .A1(n5329), .A2(n5328), .ZN(n9951) );
  NAND2_X1 U5726 ( .A1(n5003), .A2(n5002), .ZN(n4761) );
  NOR2_X1 U5727 ( .A1(n5006), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U5728 ( .A1(n5159), .A2(n5007), .ZN(n5006) );
  OR2_X1 U5729 ( .A1(n5271), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5292) );
  OR2_X1 U5730 ( .A1(n7774), .A2(n7773), .ZN(n4749) );
  NAND2_X1 U5731 ( .A1(n7774), .A2(n7773), .ZN(n7776) );
  OR2_X1 U5732 ( .A1(n6534), .A2(n6533), .ZN(n6549) );
  INV_X1 U5733 ( .A(n9371), .ZN(n8776) );
  OR2_X1 U5734 ( .A1(n5928), .A2(n5927), .ZN(n5946) );
  AOI21_X1 U5735 ( .B1(n4416), .B2(n8740), .A(n6506), .ZN(n6512) );
  NAND2_X1 U5736 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  NAND2_X1 U5737 ( .A1(n5829), .A2(n8736), .ZN(n6505) );
  NOR2_X1 U5738 ( .A1(n5040), .A2(n5039), .ZN(n8632) );
  NOR2_X1 U5739 ( .A1(n8629), .A2(n8628), .ZN(n5040) );
  AND2_X1 U5740 ( .A1(n8626), .A2(n8625), .ZN(n8627) );
  NAND2_X1 U5741 ( .A1(n6058), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6068) );
  OR2_X1 U5742 ( .A1(n6068), .A2(n8849), .ZN(n6081) );
  NAND2_X1 U5743 ( .A1(n5027), .A2(n5026), .ZN(n8718) );
  INV_X1 U5744 ( .A(n8848), .ZN(n5026) );
  INV_X1 U5745 ( .A(n8847), .ZN(n5027) );
  NAND2_X1 U5746 ( .A1(n4751), .A2(n4750), .ZN(n6540) );
  AOI21_X1 U5747 ( .B1(n6815), .B2(n6814), .A(n4434), .ZN(n4743) );
  INV_X1 U5748 ( .A(n6107), .ZN(n6108) );
  INV_X1 U5749 ( .A(n8773), .ZN(n4742) );
  CLKBUF_X1 U5750 ( .A(n8783), .Z(n8785) );
  NAND2_X1 U5751 ( .A1(n6149), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U5752 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n4755) );
  XNOR2_X1 U5753 ( .A(n6152), .B(n10053), .ZN(n9139) );
  INV_X1 U5754 ( .A(n6342), .ZN(n6095) );
  INV_X1 U5755 ( .A(n6343), .ZN(n6124) );
  NAND2_X1 U5756 ( .A1(n9173), .A2(n9185), .ZN(n9172) );
  OR2_X1 U5757 ( .A1(n6396), .A2(n6397), .ZN(n9233) );
  NOR2_X1 U5758 ( .A1(n9246), .A2(n4715), .ZN(n9716) );
  INV_X1 U5759 ( .A(n9714), .ZN(n4715) );
  NOR2_X1 U5760 ( .A1(n9716), .A2(n4714), .ZN(n9737) );
  AND2_X1 U5761 ( .A1(n9717), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5762 ( .A1(n9737), .A2(n9736), .ZN(n9735) );
  NOR2_X1 U5763 ( .A1(n9735), .A2(n4713), .ZN(n9748) );
  AND2_X1 U5764 ( .A1(n9743), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4713) );
  AND2_X1 U5765 ( .A1(n9264), .A2(n9263), .ZN(n9267) );
  NAND2_X1 U5766 ( .A1(n9327), .A2(n9111), .ZN(n4540) );
  INV_X1 U5767 ( .A(n9337), .ZN(n8979) );
  AOI21_X1 U5768 ( .B1(n4827), .B2(n9359), .A(n4469), .ZN(n4826) );
  NAND2_X1 U5769 ( .A1(n4512), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U5770 ( .A1(n9357), .A2(n9099), .ZN(n9336) );
  NAND2_X1 U5771 ( .A1(n9336), .A2(n9339), .ZN(n9335) );
  OAI211_X1 U5772 ( .C1(n4545), .C2(n9421), .A(n4867), .B(n4543), .ZN(n9358)
         );
  NAND2_X1 U5773 ( .A1(n4546), .A2(n4544), .ZN(n4543) );
  INV_X1 U5774 ( .A(n4546), .ZN(n4545) );
  AOI21_X1 U5775 ( .B1(n4868), .B2(n4873), .A(n4661), .ZN(n4867) );
  NAND2_X1 U5776 ( .A1(n9358), .A2(n9359), .ZN(n9357) );
  NAND2_X1 U5777 ( .A1(n4871), .A2(n9089), .ZN(n9367) );
  NAND2_X1 U5778 ( .A1(n4871), .A2(n4868), .ZN(n9369) );
  NAND2_X1 U5779 ( .A1(n9383), .A2(n9389), .ZN(n9384) );
  AND2_X1 U5780 ( .A1(n9089), .A2(n9104), .ZN(n9391) );
  NAND2_X1 U5781 ( .A1(n9400), .A2(n9401), .ZN(n9399) );
  NAND2_X1 U5782 ( .A1(n9421), .A2(n8967), .ZN(n9400) );
  AND2_X1 U5783 ( .A1(n8971), .A2(n9390), .ZN(n9401) );
  NAND2_X1 U5784 ( .A1(n9467), .A2(n4580), .ZN(n9415) );
  NOR2_X1 U5785 ( .A1(n9605), .A2(n4581), .ZN(n4580) );
  INV_X1 U5786 ( .A(n4582), .ZN(n4581) );
  AOI21_X1 U5787 ( .B1(n4842), .B2(n4838), .A(n4426), .ZN(n4837) );
  INV_X1 U5788 ( .A(n4542), .ZN(n9431) );
  OAI21_X1 U5789 ( .B1(n9451), .B2(n9452), .A(n8964), .ZN(n4542) );
  NAND2_X1 U5790 ( .A1(n9460), .A2(n8954), .ZN(n9451) );
  NAND2_X1 U5791 ( .A1(n9467), .A2(n6177), .ZN(n9468) );
  NAND2_X1 U5792 ( .A1(n9467), .A2(n4584), .ZN(n9445) );
  AOI21_X1 U5793 ( .B1(n4878), .B2(n4876), .A(n4875), .ZN(n4874) );
  INV_X1 U5794 ( .A(n4878), .ZN(n4877) );
  NAND2_X1 U5795 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
  AND2_X1 U5796 ( .A1(n9083), .A2(n8954), .ZN(n9462) );
  OR2_X1 U5797 ( .A1(n6026), .A2(n6025), .ZN(n6038) );
  NAND2_X1 U5798 ( .A1(n9637), .A2(n9527), .ZN(n4850) );
  NAND2_X1 U5799 ( .A1(n7350), .A2(n4570), .ZN(n9496) );
  NOR2_X1 U5800 ( .A1(n9498), .A2(n4572), .ZN(n4570) );
  NAND2_X1 U5801 ( .A1(n7350), .A2(n4574), .ZN(n9533) );
  NOR2_X1 U5802 ( .A1(n9511), .A2(n4853), .ZN(n4852) );
  INV_X1 U5803 ( .A(n4856), .ZN(n4853) );
  NAND2_X1 U5804 ( .A1(n4858), .A2(n4859), .ZN(n9508) );
  AOI21_X1 U5805 ( .B1(n4861), .B2(n9544), .A(n4860), .ZN(n4859) );
  INV_X1 U5806 ( .A(n8940), .ZN(n4860) );
  NAND2_X1 U5807 ( .A1(n7350), .A2(n9561), .ZN(n9555) );
  NAND2_X1 U5808 ( .A1(n7228), .A2(n5978), .ZN(n7347) );
  NAND2_X1 U5809 ( .A1(n4864), .A2(n8933), .ZN(n7226) );
  NAND4_X1 U5810 ( .A1(n5977), .A2(n4578), .A3(n4579), .A4(n7028), .ZN(n7351)
         );
  NOR2_X1 U5811 ( .A1(n4576), .A2(n4577), .ZN(n7230) );
  INV_X1 U5812 ( .A(n4579), .ZN(n4576) );
  NAND2_X1 U5813 ( .A1(n4579), .A2(n6954), .ZN(n7130) );
  AND2_X1 U5814 ( .A1(n7028), .A2(n9821), .ZN(n6954) );
  NAND2_X1 U5815 ( .A1(n6793), .A2(n5055), .ZN(n7027) );
  OAI21_X1 U5816 ( .B1(n8905), .B2(n6163), .A(n8909), .ZN(n6738) );
  NAND2_X1 U5817 ( .A1(n8902), .A2(n9061), .ZN(n8905) );
  NAND2_X1 U5818 ( .A1(n4567), .A2(n6807), .ZN(n6761) );
  INV_X1 U5819 ( .A(n6751), .ZN(n4567) );
  CLKBUF_X1 U5820 ( .A(n9017), .Z(n4514) );
  NAND2_X1 U5821 ( .A1(n8997), .A2(n8996), .ZN(n9305) );
  NAND2_X1 U5822 ( .A1(n7446), .A2(n8998), .ZN(n5782) );
  OR2_X1 U5823 ( .A1(n6284), .A2(n6210), .ZN(n6217) );
  XNOR2_X1 U5824 ( .A(n7532), .B(n7531), .ZN(n8999) );
  OAI21_X1 U5825 ( .B1(n7536), .B2(n7535), .A(n7529), .ZN(n7532) );
  XNOR2_X1 U5826 ( .A(n7524), .B(SI_29_), .ZN(n7518) );
  XNOR2_X1 U5827 ( .A(n4569), .B(n5779), .ZN(n6170) );
  XNOR2_X1 U5828 ( .A(n5550), .B(n5549), .ZN(n7305) );
  NAND2_X1 U5829 ( .A1(n5791), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6033) );
  INV_X1 U5830 ( .A(n4700), .ZN(n4699) );
  AND2_X1 U5831 ( .A1(n4697), .A2(n4951), .ZN(n4696) );
  AOI21_X1 U5832 ( .B1(n4953), .B2(n4955), .A(n4952), .ZN(n4951) );
  AND2_X1 U5833 ( .A1(n5154), .A2(n5153), .ZN(n5388) );
  AOI21_X1 U5834 ( .B1(n4561), .B2(n4560), .A(n5139), .ZN(n4559) );
  INV_X1 U5835 ( .A(n5136), .ZN(n4560) );
  NAND2_X1 U5836 ( .A1(n5323), .A2(n5136), .ZN(n4563) );
  AND2_X1 U5837 ( .A1(n5144), .A2(n5143), .ZN(n5351) );
  INV_X1 U5838 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5940) );
  INV_X1 U5839 ( .A(n5288), .ZN(n4963) );
  AOI21_X1 U5840 ( .B1(n5288), .B2(n4962), .A(n4961), .ZN(n4960) );
  INV_X1 U5841 ( .A(n5127), .ZN(n4961) );
  AND2_X1 U5842 ( .A1(n5132), .A2(n5131), .ZN(n5308) );
  OR2_X1 U5843 ( .A1(n5938), .A2(n5833), .ZN(n5910) );
  AND2_X1 U5844 ( .A1(n5117), .A2(n5116), .ZN(n5256) );
  INV_X1 U5845 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10285) );
  AND2_X1 U5846 ( .A1(n5112), .A2(n5101), .ZN(n5235) );
  OR2_X1 U5847 ( .A1(n5100), .A2(SI_3_), .ZN(n5101) );
  INV_X1 U5848 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5833) );
  AND2_X1 U5849 ( .A1(n7200), .A2(n7199), .ZN(n7865) );
  NAND2_X1 U5850 ( .A1(n4907), .A2(n7440), .ZN(n7880) );
  NAND2_X1 U5851 ( .A1(n7439), .A2(n7438), .ZN(n4907) );
  AND2_X1 U5852 ( .A1(n7941), .A2(n8256), .ZN(n7942) );
  AND3_X1 U5853 ( .A1(n5560), .A2(n5559), .A3(n5558), .ZN(n8298) );
  AND2_X1 U5854 ( .A1(n6655), .A2(n6654), .ZN(n8061) );
  AND2_X1 U5855 ( .A1(n6898), .A2(n6897), .ZN(n8008) );
  INV_X1 U5856 ( .A(n4889), .ZN(n4888) );
  AOI21_X1 U5857 ( .B1(n4889), .B2(n4887), .A(n4458), .ZN(n4886) );
  NOR2_X1 U5858 ( .A1(n7891), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U5859 ( .A1(n7951), .A2(n7897), .ZN(n8028) );
  AND4_X1 U5860 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), .ZN(n9908)
         );
  OR2_X1 U5861 ( .A1(n5210), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U5862 ( .A1(n4891), .A2(n7988), .ZN(n8036) );
  NAND2_X1 U5863 ( .A1(n7989), .A2(n7987), .ZN(n4891) );
  AND2_X1 U5864 ( .A1(n5614), .A2(n5613), .ZN(n8054) );
  INV_X1 U5865 ( .A(n8273), .ZN(n8255) );
  INV_X1 U5866 ( .A(n8298), .ZN(n8075) );
  INV_X1 U5867 ( .A(n8308), .ZN(n8076) );
  NAND4_X1 U5868 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n8396)
         );
  INV_X1 U5869 ( .A(n7877), .ZN(n8411) );
  NAND4_X1 U5870 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n8395)
         );
  INV_X1 U5871 ( .A(n8429), .ZN(n8079) );
  NAND4_X1 U5872 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n8082)
         );
  OR2_X1 U5873 ( .A1(n5208), .A2(n5300), .ZN(n5306) );
  NAND4_X1 U5874 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n8084)
         );
  OR2_X1 U5875 ( .A1(n5210), .A2(n7981), .ZN(n5268) );
  NAND2_X1 U5876 ( .A1(n5183), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5214) );
  OR2_X1 U5877 ( .A1(n5208), .A2(n5207), .ZN(n5216) );
  CLKBUF_X1 U5878 ( .A(n6579), .Z(n8086) );
  OR2_X1 U5879 ( .A1(n6238), .A2(P2_U3151), .ZN(n8185) );
  OAI21_X1 U5880 ( .B1(n8208), .B2(P2_REG2_REG_0__SCAN_IN), .A(n4498), .ZN(
        n9851) );
  NAND2_X1 U5881 ( .A1(n8208), .A2(n6227), .ZN(n4498) );
  OR2_X1 U5882 ( .A1(n4815), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5883 ( .A1(n6265), .A2(n4612), .ZN(n6486) );
  NAND2_X1 U5884 ( .A1(n7086), .A2(n4915), .ZN(n6996) );
  INV_X1 U5885 ( .A(n4914), .ZN(n4597) );
  INV_X1 U5886 ( .A(n7109), .ZN(n4812) );
  AND2_X1 U5887 ( .A1(n7257), .A2(n4926), .ZN(n7262) );
  INV_X1 U5888 ( .A(n4920), .ZN(n7489) );
  OAI21_X1 U5889 ( .B1(n8093), .B2(n4616), .A(n4615), .ZN(n8110) );
  NAND2_X1 U5890 ( .A1(n4617), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4616) );
  INV_X1 U5891 ( .A(n7493), .ZN(n4617) );
  NOR2_X1 U5892 ( .A1(n8174), .A2(n4501), .ZN(n8167) );
  AND2_X1 U5893 ( .A1(n8166), .A2(n8492), .ZN(n4501) );
  INV_X1 U5894 ( .A(n8222), .ZN(n4923) );
  NAND2_X1 U5895 ( .A1(n8223), .A2(n9872), .ZN(n4924) );
  XNOR2_X1 U5896 ( .A(n8219), .B(n8220), .ZN(n4925) );
  INV_X1 U5897 ( .A(n5688), .ZN(n4762) );
  NAND2_X1 U5898 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U5899 ( .A1(n8073), .A2(n8408), .ZN(n7845) );
  NAND2_X1 U5900 ( .A1(n4775), .A2(n5512), .ZN(n8306) );
  NAND2_X1 U5901 ( .A1(n8337), .A2(n4779), .ZN(n4775) );
  NAND2_X1 U5902 ( .A1(n8337), .A2(n5049), .ZN(n8318) );
  AND2_X1 U5903 ( .A1(n5410), .A2(n5409), .ZN(n8399) );
  OR2_X1 U5904 ( .A1(n7214), .A2(n4802), .ZN(n4796) );
  INV_X1 U5905 ( .A(n7362), .ZN(n9962) );
  NAND2_X1 U5906 ( .A1(n4805), .A2(n5047), .ZN(n7425) );
  NAND2_X1 U5907 ( .A1(n7214), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5908 ( .A1(n7214), .A2(n5331), .ZN(n7333) );
  INV_X1 U5909 ( .A(n9951), .ZN(n5330) );
  AND3_X1 U5910 ( .A1(n5315), .A2(n5314), .A3(n5313), .ZN(n9946) );
  NAND2_X1 U5911 ( .A1(n4997), .A2(n7631), .ZN(n7159) );
  NAND2_X1 U5912 ( .A1(n5690), .A2(n6629), .ZN(n6981) );
  OAI21_X1 U5913 ( .B1(n5189), .B2(n4883), .A(n4881), .ZN(n4884) );
  OR2_X1 U5914 ( .A1(n5217), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U5915 ( .A1(n5189), .A2(n4882), .ZN(n4881) );
  OR2_X1 U5916 ( .A1(n6645), .A2(n6602), .ZN(n9898) );
  INV_X1 U5917 ( .A(n8352), .ZN(n8445) );
  INV_X1 U5918 ( .A(n7579), .ZN(n8515) );
  INV_X1 U5919 ( .A(n7565), .ZN(n8520) );
  AOI21_X1 U5920 ( .B1(n8239), .B2(n8413), .A(n8238), .ZN(n8519) );
  NAND2_X1 U5921 ( .A1(n4782), .A2(n4784), .ZN(n8235) );
  INV_X1 U5922 ( .A(n8054), .ZN(n8526) );
  NAND2_X1 U5923 ( .A1(n5593), .A2(n5592), .ZN(n8532) );
  NAND2_X1 U5924 ( .A1(n7446), .A2(n7537), .ZN(n5593) );
  XNOR2_X1 U5925 ( .A(n8266), .B(n8267), .ZN(n8533) );
  AOI21_X1 U5926 ( .B1(n8300), .B2(n4989), .A(n4987), .ZN(n4981) );
  XOR2_X1 U5927 ( .A(n8278), .B(n8277), .Z(n8538) );
  NOR2_X1 U5928 ( .A1(n4993), .A2(n7591), .ZN(n8287) );
  INV_X1 U5929 ( .A(n4996), .ZN(n4993) );
  NAND2_X1 U5930 ( .A1(n5490), .A2(n5489), .ZN(n8559) );
  AND2_X1 U5931 ( .A1(n5468), .A2(n5467), .ZN(n8567) );
  NAND2_X1 U5932 ( .A1(n5448), .A2(n5447), .ZN(n8570) );
  NAND2_X1 U5933 ( .A1(n5166), .A2(n5165), .ZN(n8576) );
  NAND2_X1 U5934 ( .A1(n5427), .A2(n5426), .ZN(n8581) );
  NAND2_X1 U5935 ( .A1(n4975), .A2(n7681), .ZN(n8383) );
  NAND2_X1 U5936 ( .A1(n8403), .A2(n7682), .ZN(n4975) );
  INV_X1 U5937 ( .A(n8399), .ZN(n8587) );
  NAND2_X1 U5938 ( .A1(n5395), .A2(n5394), .ZN(n8593) );
  NAND2_X1 U5939 ( .A1(n5698), .A2(n7666), .ZN(n8424) );
  XNOR2_X1 U5940 ( .A(n5079), .B(n5078), .ZN(n7859) );
  XNOR2_X1 U5941 ( .A(n5718), .B(n5717), .ZN(n7448) );
  XNOR2_X1 U5942 ( .A(n5273), .B(n5272), .ZN(n6840) );
  INV_X1 U5943 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5099) );
  AND2_X1 U5944 ( .A1(n6257), .A2(n5223), .ZN(n5239) );
  NAND2_X1 U5945 ( .A1(n4815), .A2(n4818), .ZN(n6306) );
  NAND2_X1 U5946 ( .A1(n7458), .A2(n8998), .ZN(n6116) );
  NAND2_X1 U5947 ( .A1(n7776), .A2(n4749), .ZN(n8725) );
  NAND2_X1 U5948 ( .A1(n5945), .A2(n5944), .ZN(n8731) );
  OR2_X1 U5949 ( .A1(n6334), .A2(n5979), .ZN(n5945) );
  NAND2_X1 U5950 ( .A1(n7185), .A2(n7295), .ZN(n7187) );
  NAND2_X1 U5951 ( .A1(n5020), .A2(n8856), .ZN(n8763) );
  NAND2_X1 U5952 ( .A1(n8855), .A2(n8857), .ZN(n5020) );
  NAND2_X1 U5953 ( .A1(n8820), .A2(n8671), .ZN(n8772) );
  NAND2_X1 U5954 ( .A1(n5028), .A2(n4734), .ZN(n8717) );
  AOI21_X1 U5955 ( .B1(n8719), .B2(n8848), .A(n4486), .ZN(n4734) );
  NAND2_X1 U5956 ( .A1(n7422), .A2(n8998), .ZN(n6091) );
  XNOR2_X1 U5957 ( .A(n6813), .B(n6811), .ZN(n6560) );
  INV_X1 U5958 ( .A(n9165), .ZN(n8619) );
  NAND2_X1 U5959 ( .A1(n7297), .A2(n7298), .ZN(n7771) );
  NAND2_X1 U5960 ( .A1(n8633), .A2(n8632), .ZN(n8830) );
  AOI21_X1 U5961 ( .B1(n5021), .B2(n5024), .A(n4457), .ZN(n5018) );
  NAND2_X1 U5962 ( .A1(n8649), .A2(n8719), .ZN(n8847) );
  INV_X1 U5963 ( .A(n6830), .ZN(n6827) );
  NAND2_X1 U5964 ( .A1(n7452), .A2(n8998), .ZN(n4496) );
  INV_X1 U5965 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U5966 ( .B1(n9146), .B2(n6153), .A(n9051), .ZN(n4624) );
  INV_X1 U5967 ( .A(n9053), .ZN(n9330) );
  NAND4_X1 U5968 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n9168)
         );
  NAND2_X1 U5969 ( .A1(n5855), .A2(n5854), .ZN(n9170) );
  INV_X1 U5970 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5102) );
  OR2_X1 U5971 ( .A1(n6070), .A2(n6287), .ZN(n5815) );
  NAND2_X1 U5972 ( .A1(n5811), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5814) );
  AND2_X1 U5973 ( .A1(n4725), .A2(n4724), .ZN(n6419) );
  NAND2_X1 U5974 ( .A1(n6386), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4724) );
  NOR2_X1 U5975 ( .A1(n6417), .A2(n4723), .ZN(n6446) );
  AND2_X1 U5976 ( .A1(n6424), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5977 ( .A1(n6446), .A2(n6445), .ZN(n6444) );
  NOR2_X1 U5978 ( .A1(n6444), .A2(n4722), .ZN(n6434) );
  AND2_X1 U5979 ( .A1(n6391), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4722) );
  NOR2_X1 U5980 ( .A1(n6434), .A2(n6433), .ZN(n6432) );
  INV_X1 U5981 ( .A(n4721), .ZN(n9760) );
  INV_X1 U5982 ( .A(n4719), .ZN(n9779) );
  OR2_X1 U5983 ( .A1(n9255), .A2(n9254), .ZN(n9264) );
  NAND2_X1 U5984 ( .A1(n4841), .A2(n4843), .ZN(n4840) );
  INV_X1 U5985 ( .A(n6045), .ZN(n4841) );
  NAND2_X1 U5986 ( .A1(n4880), .A2(n8952), .ZN(n9484) );
  NAND2_X1 U5987 ( .A1(n4854), .A2(n4856), .ZN(n9512) );
  NAND2_X1 U5988 ( .A1(n9548), .A2(n4861), .ZN(n9524) );
  NAND2_X1 U5989 ( .A1(n7224), .A2(n9070), .ZN(n7348) );
  NAND2_X1 U5990 ( .A1(n6166), .A2(n9055), .ZN(n7059) );
  OAI21_X1 U5991 ( .B1(n6938), .B2(n4835), .A(n4832), .ZN(n7056) );
  NAND2_X1 U5992 ( .A1(n6936), .A2(n5934), .ZN(n7057) );
  CLKBUF_X1 U5993 ( .A(n6793), .Z(n6794) );
  NAND2_X1 U5994 ( .A1(n4683), .A2(n6161), .ZN(n6753) );
  CLKBUF_X1 U5995 ( .A(n6748), .Z(n6749) );
  NAND2_X1 U5996 ( .A1(n4557), .A2(n9321), .ZN(n6218) );
  AOI21_X1 U5997 ( .B1(n9309), .B2(n9836), .A(n4513), .ZN(n4557) );
  INV_X1 U5998 ( .A(n9317), .ZN(n4513) );
  NAND2_X1 U5999 ( .A1(n4556), .A2(n9839), .ZN(n6215) );
  INV_X1 U6000 ( .A(n6218), .ZN(n4556) );
  AOI211_X1 U6001 ( .C1(n9581), .C2(n9836), .A(n9580), .B(n9579), .ZN(n9662)
         );
  AOI211_X1 U6002 ( .C1(n9591), .C2(n9836), .A(n9590), .B(n9589), .ZN(n9666)
         );
  INV_X1 U6003 ( .A(n9407), .ZN(n9673) );
  INV_X1 U6004 ( .A(n9535), .ZN(n9690) );
  NAND2_X1 U6005 ( .A1(n5983), .A2(n5982), .ZN(n8843) );
  OR2_X1 U6006 ( .A1(n6456), .A2(n5979), .ZN(n5983) );
  NAND2_X1 U6007 ( .A1(n5958), .A2(n5957), .ZN(n8862) );
  NAND2_X1 U6008 ( .A1(n5898), .A2(n5897), .ZN(n9804) );
  XNOR2_X1 U6009 ( .A(n5659), .B(n5658), .ZN(n9704) );
  NAND2_X1 U6010 ( .A1(n4966), .A2(n5646), .ZN(n5659) );
  NAND2_X1 U6011 ( .A1(n5645), .A2(n5644), .ZN(n4966) );
  CLKBUF_X1 U6012 ( .A(n6170), .Z(n9705) );
  NAND2_X1 U6013 ( .A1(n5780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4568) );
  XNOR2_X1 U6014 ( .A(n6187), .B(n10047), .ZN(n7457) );
  NAND2_X1 U6015 ( .A1(n4956), .A2(n4955), .ZN(n5174) );
  NAND2_X1 U6016 ( .A1(n4956), .A2(n4435), .ZN(n5173) );
  NOR2_X1 U6017 ( .A1(n5014), .A2(n5015), .ZN(n5013) );
  NAND2_X1 U6018 ( .A1(n5288), .A2(n5289), .ZN(n5291) );
  NAND2_X1 U6019 ( .A1(n5277), .A2(n5122), .ZN(n5289) );
  NAND2_X1 U6020 ( .A1(n4716), .A2(n5818), .ZN(n6378) );
  AOI21_X1 U6021 ( .B1(n4467), .B2(P1_IR_REG_1__SCAN_IN), .A(n4717), .ZN(n4716) );
  OAI211_X1 U6022 ( .C1(n7914), .C2(n4432), .A(n8048), .B(n7913), .ZN(n7919)
         );
  AOI21_X1 U6023 ( .B1(n7749), .B2(n7748), .A(n7747), .ZN(n7756) );
  AND2_X1 U6024 ( .A1(n4821), .A2(n4413), .ZN(n8128) );
  OAI211_X1 U6025 ( .C1(n8199), .C2(n8224), .A(n4619), .B(n4618), .ZN(P2_U3200) );
  OAI21_X1 U6026 ( .B1(n8218), .B2(n4449), .A(n9883), .ZN(n4618) );
  NAND2_X1 U6027 ( .A1(n4764), .A2(n5761), .ZN(n5762) );
  OR2_X1 U6028 ( .A1(n8744), .A2(n5034), .ZN(n8753) );
  INV_X1 U6029 ( .A(n4725), .ZN(n6405) );
  AOI21_X1 U6030 ( .B1(n9731), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9296), .ZN(
        n4727) );
  NAND2_X1 U6031 ( .A1(n4729), .A2(n6153), .ZN(n4728) );
  NAND2_X1 U6032 ( .A1(n4731), .A2(n9143), .ZN(n4730) );
  CLKBUF_X1 U6033 ( .A(n9309), .Z(n9319) );
  NOR2_X1 U6034 ( .A1(n9576), .A2(n9521), .ZN(n9332) );
  NOR2_X1 U6035 ( .A1(n8532), .A2(n8255), .ZN(n5604) );
  OR2_X1 U6036 ( .A1(n8532), .A2(n8273), .ZN(n7718) );
  AND2_X1 U6037 ( .A1(n5711), .A2(n4762), .ZN(n4419) );
  AND2_X1 U6038 ( .A1(n4419), .A2(n9992), .ZN(n4420) );
  NAND2_X1 U6039 ( .A1(n5520), .A2(n5519), .ZN(n5530) );
  AND4_X1 U6040 ( .A1(n9111), .A2(n9049), .A3(n9099), .A4(n9112), .ZN(n4421)
         );
  INV_X1 U6041 ( .A(n8953), .ZN(n4875) );
  NAND2_X1 U6042 ( .A1(n9108), .A2(n9099), .ZN(n9348) );
  OR2_X1 U6043 ( .A1(n8081), .A2(n9951), .ZN(n7648) );
  OR2_X1 U6044 ( .A1(n9132), .A2(n9049), .ZN(n4422) );
  INV_X1 U6045 ( .A(n9498), .ZN(n9685) );
  AND2_X1 U6046 ( .A1(n4826), .A2(n4824), .ZN(n4423) );
  AND2_X1 U6047 ( .A1(n5038), .A2(n4450), .ZN(n4424) );
  NOR2_X1 U6048 ( .A1(n9350), .A2(n4590), .ZN(n4589) );
  INV_X1 U6049 ( .A(n7181), .ZN(n4531) );
  INV_X1 U6050 ( .A(n5604), .ZN(n4794) );
  OR2_X1 U6051 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4425) );
  NOR2_X1 U6052 ( .A1(n9437), .A2(n9454), .ZN(n4426) );
  INV_X1 U6053 ( .A(n8973), .ZN(n4654) );
  NAND2_X1 U6054 ( .A1(n4473), .A2(n4793), .ZN(n4790) );
  CLKBUF_X3 U6055 ( .A(n6903), .Z(n6674) );
  AND2_X1 U6056 ( .A1(n4464), .A2(n4844), .ZN(n4843) );
  NAND2_X1 U6057 ( .A1(n5001), .A2(n5066), .ZN(n5163) );
  OR2_X1 U6058 ( .A1(n6217), .A2(n9694), .ZN(n9838) );
  INV_X1 U6059 ( .A(n7796), .ZN(n4523) );
  NAND2_X2 U6060 ( .A1(n5077), .A2(n5091), .ZN(n5210) );
  AND3_X1 U6061 ( .A1(n4649), .A2(n4659), .A3(n9114), .ZN(n4427) );
  INV_X1 U6062 ( .A(n9360), .ZN(n8980) );
  AND2_X1 U6063 ( .A1(n8685), .A2(n4740), .ZN(n4428) );
  INV_X1 U6064 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5007) );
  INV_X1 U6065 ( .A(n4981), .ZN(n8266) );
  BUF_X1 U6066 ( .A(n6070), .Z(n6131) );
  AND2_X1 U6067 ( .A1(n5017), .A2(n5016), .ZN(n5817) );
  AND4_X1 U6068 ( .A1(n4412), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n4429)
         );
  OR2_X1 U6069 ( .A1(n7875), .A2(n8256), .ZN(n4430) );
  AND2_X1 U6070 ( .A1(n4825), .A2(n4826), .ZN(n4431) );
  AND2_X1 U6071 ( .A1(n8046), .A2(n7911), .ZN(n4432) );
  OR2_X1 U6072 ( .A1(n5463), .A2(n4761), .ZN(n4433) );
  XNOR2_X1 U6073 ( .A(n8674), .B(n6816), .ZN(n4434) );
  OR2_X1 U6074 ( .A1(n5145), .A2(SI_11_), .ZN(n4435) );
  NAND2_X1 U6075 ( .A1(n5797), .A2(n5796), .ZN(n9470) );
  AND2_X1 U6076 ( .A1(n6177), .A2(n9487), .ZN(n4436) );
  INV_X1 U6077 ( .A(n9171), .ZN(n5847) );
  AND2_X1 U6078 ( .A1(n4840), .A2(n6055), .ZN(n4437) );
  INV_X1 U6079 ( .A(n4945), .ZN(n4944) );
  NAND2_X1 U6080 ( .A1(n4947), .A2(n5477), .ZN(n4945) );
  INV_X1 U6081 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6082 ( .A1(n5997), .A2(n5996), .ZN(n9647) );
  INV_X1 U6083 ( .A(n8992), .ZN(n9046) );
  XNOR2_X1 U6084 ( .A(n9314), .B(n9330), .ZN(n8992) );
  AND2_X1 U6085 ( .A1(n7887), .A2(n8078), .ZN(n4438) );
  NAND2_X2 U6086 ( .A1(n5077), .A2(n7859), .ZN(n5199) );
  INV_X1 U6087 ( .A(n8423), .ZN(n5699) );
  INV_X1 U6088 ( .A(n8299), .ZN(n8295) );
  XNOR2_X1 U6089 ( .A(n8026), .B(n8308), .ZN(n8299) );
  OR2_X1 U6090 ( .A1(n9350), .A2(n9341), .ZN(n4439) );
  AND2_X1 U6091 ( .A1(n8084), .A2(n7980), .ZN(n4440) );
  AND2_X1 U6092 ( .A1(n8007), .A2(n6897), .ZN(n4441) );
  AND2_X1 U6093 ( .A1(n4942), .A2(n4941), .ZN(n4442) );
  AND2_X1 U6094 ( .A1(n4996), .A2(n4994), .ZN(n4443) );
  AND3_X1 U6095 ( .A1(n4641), .A2(n8989), .A3(n4640), .ZN(n4444) );
  NAND2_X1 U6096 ( .A1(n5069), .A2(n5003), .ZN(n5671) );
  NAND2_X1 U6097 ( .A1(n4885), .A2(n4884), .ZN(n9918) );
  INV_X1 U6098 ( .A(n9605), .ZN(n9420) );
  NAND2_X1 U6099 ( .A1(n6067), .A2(n6066), .ZN(n9605) );
  NOR2_X1 U6100 ( .A1(n8318), .A2(n8321), .ZN(n4445) );
  INV_X1 U6101 ( .A(n7087), .ZN(n4596) );
  AND2_X1 U6102 ( .A1(n9114), .A2(n9111), .ZN(n9329) );
  INV_X1 U6103 ( .A(n9329), .ZN(n4824) );
  OR2_X1 U6104 ( .A1(n7294), .A2(n8728), .ZN(n9026) );
  INV_X1 U6105 ( .A(n9026), .ZN(n4675) );
  OR2_X1 U6106 ( .A1(n9479), .A2(n8812), .ZN(n4446) );
  NOR2_X1 U6107 ( .A1(n6342), .A2(n6370), .ZN(n4447) );
  AND2_X1 U6108 ( .A1(n4978), .A2(n7681), .ZN(n4448) );
  INV_X1 U6109 ( .A(n4803), .ZN(n4802) );
  NOR2_X1 U6110 ( .A1(n5369), .A2(n4804), .ZN(n4803) );
  AND2_X1 U6111 ( .A1(n8196), .A2(n8195), .ZN(n4449) );
  INV_X1 U6112 ( .A(n4873), .ZN(n4872) );
  AND2_X1 U6113 ( .A1(n10046), .A2(n5779), .ZN(n4450) );
  NOR2_X1 U6114 ( .A1(n9339), .A2(n4828), .ZN(n4827) );
  INV_X1 U6115 ( .A(n4589), .ZN(n4591) );
  AND2_X1 U6116 ( .A1(n9076), .A2(n9073), .ZN(n4451) );
  AND2_X1 U6117 ( .A1(n4434), .A2(n6814), .ZN(n4452) );
  OR2_X1 U6118 ( .A1(n6342), .A2(n10051), .ZN(n4453) );
  AND2_X1 U6119 ( .A1(n8552), .A2(n8320), .ZN(n4454) );
  INV_X1 U6120 ( .A(n6032), .ZN(n4855) );
  INV_X1 U6121 ( .A(n5622), .ZN(n4793) );
  NOR2_X1 U6122 ( .A1(n8054), .A2(n8264), .ZN(n5622) );
  NAND2_X1 U6123 ( .A1(n6139), .A2(n6138), .ZN(n9314) );
  AND2_X1 U6124 ( .A1(n7565), .A2(n7916), .ZN(n4455) );
  NOR2_X1 U6125 ( .A1(n7770), .A2(n7769), .ZN(n4456) );
  NOR2_X1 U6126 ( .A1(n7791), .A2(n7790), .ZN(n4457) );
  NOR2_X1 U6127 ( .A1(n4438), .A2(n7931), .ZN(n4458) );
  INV_X1 U6128 ( .A(n4530), .ZN(n4529) );
  OAI21_X1 U6129 ( .B1(n8616), .B2(n4531), .A(n7183), .ZN(n4530) );
  AND2_X1 U6130 ( .A1(n7875), .A2(n8256), .ZN(n4459) );
  NOR2_X1 U6131 ( .A1(n8026), .A2(n8308), .ZN(n7591) );
  INV_X1 U6132 ( .A(n7591), .ZN(n4995) );
  NAND2_X1 U6133 ( .A1(n9375), .A2(n8880), .ZN(n8987) );
  INV_X1 U6134 ( .A(n8987), .ZN(n4661) );
  AND2_X1 U6135 ( .A1(n5954), .A2(n5953), .ZN(n4460) );
  AND2_X1 U6136 ( .A1(n7711), .A2(n7709), .ZN(n4461) );
  INV_X1 U6137 ( .A(n5053), .ZN(n4899) );
  AND2_X1 U6138 ( .A1(n9685), .A2(n9510), .ZN(n4462) );
  NAND2_X1 U6139 ( .A1(n7540), .A2(n7571), .ZN(n7732) );
  INV_X1 U6140 ( .A(n7732), .ZN(n4712) );
  NAND2_X1 U6141 ( .A1(n5069), .A2(n5004), .ZN(n4463) );
  NAND2_X1 U6142 ( .A1(n9450), .A2(n7838), .ZN(n4464) );
  INV_X1 U6143 ( .A(n4572), .ZN(n4571) );
  NAND2_X1 U6144 ( .A1(n4573), .A2(n4574), .ZN(n4572) );
  AND2_X1 U6145 ( .A1(n7878), .A2(n7877), .ZN(n4465) );
  OR2_X1 U6146 ( .A1(n8913), .A2(n8912), .ZN(n4466) );
  INV_X1 U6147 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5789) );
  INV_X1 U6148 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6190) );
  AND2_X1 U6149 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4467) );
  AND2_X1 U6150 ( .A1(n8026), .A2(n8308), .ZN(n4468) );
  INV_X1 U6151 ( .A(n6901), .ZN(n8085) );
  AND4_X1 U6152 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n6901)
         );
  INV_X1 U6153 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5071) );
  INV_X1 U6154 ( .A(n4768), .ZN(n4767) );
  NAND2_X1 U6155 ( .A1(n4771), .A2(n4769), .ZN(n4768) );
  INV_X1 U6156 ( .A(n5139), .ZN(n4703) );
  NOR2_X1 U6157 ( .A1(n5138), .A2(SI_9_), .ZN(n5139) );
  AND2_X1 U6158 ( .A1(n9664), .A2(n8980), .ZN(n4469) );
  NOR2_X1 U6159 ( .A1(n9962), .A2(n8440), .ZN(n4470) );
  INV_X1 U6160 ( .A(n4843), .ZN(n4842) );
  NAND2_X1 U6161 ( .A1(n7697), .A2(n7696), .ZN(n4471) );
  NAND2_X1 U6162 ( .A1(n9070), .A2(n8931), .ZN(n4472) );
  INV_X1 U6163 ( .A(n4990), .ZN(n4989) );
  NAND2_X1 U6164 ( .A1(n4461), .A2(n4991), .ZN(n4990) );
  INV_X1 U6165 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U6166 ( .A1(n4421), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U6167 ( .A1(n5623), .A2(n4794), .ZN(n4473) );
  NAND2_X1 U6168 ( .A1(n6057), .A2(n6056), .ZN(n9437) );
  INV_X1 U6169 ( .A(n9437), .ZN(n4583) );
  AND2_X1 U6170 ( .A1(n7269), .A2(n7203), .ZN(n4474) );
  NOR2_X1 U6171 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4475) );
  NOR2_X1 U6172 ( .A1(n7261), .A2(n5345), .ZN(n4476) );
  OR2_X1 U6173 ( .A1(n4818), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4477) );
  INV_X1 U6174 ( .A(n6571), .ZN(n5010) );
  AOI22_X1 U6175 ( .A1(n8740), .A2(n9057), .B1(n8736), .B2(n6890), .ZN(n6571)
         );
  OR2_X1 U6176 ( .A1(n9092), .A2(n4654), .ZN(n4478) );
  INV_X1 U6177 ( .A(n9009), .ZN(n9656) );
  AND2_X1 U6178 ( .A1(n8933), .A2(n9054), .ZN(n4479) );
  AND2_X1 U6179 ( .A1(n5694), .A2(n7631), .ZN(n4480) );
  NOR2_X1 U6180 ( .A1(n6065), .A2(n4839), .ZN(n4838) );
  NOR2_X1 U6181 ( .A1(n7879), .A2(n4906), .ZN(n4905) );
  AND2_X1 U6182 ( .A1(n5154), .A2(n4932), .ZN(n4481) );
  INV_X1 U6183 ( .A(n4552), .ZN(n4551) );
  NOR2_X1 U6184 ( .A1(n4553), .A2(n8936), .ZN(n4552) );
  INV_X1 U6185 ( .A(n4562), .ZN(n4561) );
  NAND2_X1 U6186 ( .A1(n4563), .A2(n5332), .ZN(n4562) );
  NAND2_X1 U6187 ( .A1(n7773), .A2(n7775), .ZN(n4482) );
  INV_X1 U6188 ( .A(n9495), .ZN(n4876) );
  INV_X1 U6189 ( .A(n8671), .ZN(n4741) );
  INV_X1 U6190 ( .A(n5419), .ZN(n5156) );
  INV_X1 U6191 ( .A(n7577), .ZN(n8518) );
  AND2_X1 U6192 ( .A1(n4539), .A2(n4537), .ZN(n8855) );
  AND2_X1 U6193 ( .A1(n4851), .A2(n4850), .ZN(n4483) );
  INV_X1 U6194 ( .A(n5011), .ZN(n4747) );
  NOR2_X1 U6195 ( .A1(n9496), .A2(n9625), .ZN(n9467) );
  NAND2_X1 U6196 ( .A1(n8939), .A2(n8926), .ZN(n9544) );
  INV_X1 U6197 ( .A(n9544), .ZN(n4862) );
  INV_X1 U6198 ( .A(n9393), .ZN(n8880) );
  AND2_X1 U6199 ( .A1(n8937), .A2(n8939), .ZN(n4484) );
  AND3_X1 U6200 ( .A1(n4749), .A2(n7775), .A3(n7776), .ZN(n4485) );
  NAND2_X1 U6201 ( .A1(n9467), .A2(n4582), .ZN(n4585) );
  NAND2_X1 U6202 ( .A1(n7350), .A2(n4571), .ZN(n4575) );
  NAND2_X1 U6203 ( .A1(n8817), .A2(n8660), .ZN(n4486) );
  AND2_X1 U6204 ( .A1(n4880), .A2(n4878), .ZN(n4487) );
  NAND2_X1 U6205 ( .A1(n7951), .A2(n4897), .ZN(n4488) );
  INV_X1 U6206 ( .A(n9858), .ZN(n4883) );
  AND2_X1 U6207 ( .A1(n5479), .A2(SI_18_), .ZN(n4489) );
  INV_X1 U6208 ( .A(n4851), .ZN(n9640) );
  NAND2_X1 U6209 ( .A1(n4854), .A2(n4852), .ZN(n4851) );
  NOR2_X1 U6210 ( .A1(n8092), .A2(n7491), .ZN(n4490) );
  OR2_X1 U6211 ( .A1(n7254), .A2(n5364), .ZN(n4491) );
  INV_X1 U6212 ( .A(n8899), .ZN(n5036) );
  INV_X1 U6213 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4509) );
  INV_X1 U6214 ( .A(n5262), .ZN(n7050) );
  NAND2_X1 U6215 ( .A1(n4433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6216 ( .A1(n4796), .A2(n4800), .ZN(n8437) );
  NAND2_X1 U6217 ( .A1(n5804), .A2(n5803), .ZN(n9637) );
  INV_X1 U6218 ( .A(n9637), .ZN(n4573) );
  NOR2_X1 U6219 ( .A1(n7351), .A2(n8843), .ZN(n7350) );
  NAND2_X1 U6220 ( .A1(n7173), .A2(n7170), .ZN(n4492) );
  AND2_X1 U6221 ( .A1(n5661), .A2(n5660), .ZN(n4493) );
  AND2_X1 U6222 ( .A1(n4914), .A2(n7086), .ZN(n4494) );
  NOR2_X1 U6223 ( .A1(n6538), .A2(n6537), .ZN(n6570) );
  AND2_X1 U6224 ( .A1(n4595), .A2(n7087), .ZN(n4495) );
  INV_X2 U6225 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U6226 ( .A1(n4811), .A2(n7006), .ZN(n7079) );
  INV_X1 U6227 ( .A(n7006), .ZN(n4499) );
  NOR2_X1 U6228 ( .A1(n4918), .A2(n7006), .ZN(n4917) );
  NAND2_X1 U6229 ( .A1(n4916), .A2(n7006), .ZN(n7086) );
  AOI21_X1 U6230 ( .B1(n8180), .B2(n8191), .A(n8179), .ZN(n8182) );
  NAND2_X1 U6231 ( .A1(n5405), .A2(SI_14_), .ZN(n5155) );
  NAND2_X1 U6232 ( .A1(n4965), .A2(n4964), .ZN(n7521) );
  NAND2_X1 U6233 ( .A1(n4503), .A2(n4502), .ZN(n7734) );
  NAND2_X1 U6234 ( .A1(n7578), .A2(n7540), .ZN(n7730) );
  NAND2_X1 U6235 ( .A1(n5389), .A2(n5388), .ZN(n5391) );
  NAND2_X1 U6236 ( .A1(n5517), .A2(n5516), .ZN(n5535) );
  INV_X1 U6237 ( .A(n9366), .ZN(n4870) );
  NAND2_X1 U6238 ( .A1(n5238), .A2(n5112), .ZN(n5257) );
  INV_X1 U6239 ( .A(n8988), .ZN(n4656) );
  NAND2_X1 U6240 ( .A1(n4627), .A2(n4626), .ZN(n9048) );
  MUX2_X1 U6241 ( .A(n9006), .B(n9049), .S(n9305), .Z(n9003) );
  NAND2_X1 U6242 ( .A1(n4655), .A2(n4478), .ZN(n4649) );
  NAND2_X1 U6243 ( .A1(n4931), .A2(n5403), .ZN(n4930) );
  INV_X1 U6244 ( .A(n5072), .ZN(n5720) );
  AND2_X2 U6245 ( .A1(n4759), .A2(n5001), .ZN(n5072) );
  NAND2_X1 U6246 ( .A1(n6675), .A2(n6676), .ZN(n4497) );
  NAND2_X2 U6247 ( .A1(n6627), .A2(n6626), .ZN(n6903) );
  AOI21_X1 U6248 ( .B1(n4925), .B2(n9883), .A(n4922), .ZN(n4921) );
  AOI21_X1 U6249 ( .B1(n6230), .B2(n6306), .A(n9876), .ZN(n6479) );
  OAI21_X2 U6250 ( .B1(n7413), .B2(n8409), .A(n7412), .ZN(n7415) );
  OAI22_X1 U6251 ( .A1(n7098), .A2(n7097), .B1(n7096), .B2(n7095), .ZN(n7100)
         );
  NOR2_X1 U6252 ( .A1(n7503), .A2(n7502), .ZN(n8090) );
  AOI21_X2 U6253 ( .B1(n7996), .B2(n7959), .A(n7960), .ZN(n7962) );
  OAI21_X2 U6254 ( .B1(n7989), .B2(n4888), .A(n4886), .ZN(n8020) );
  NAND2_X1 U6255 ( .A1(n5190), .A2(n5191), .ZN(n5195) );
  AND2_X1 U6256 ( .A1(n5104), .A2(n5106), .ZN(n5190) );
  NAND2_X1 U6257 ( .A1(n5309), .A2(n5308), .ZN(n5311) );
  AOI21_X2 U6258 ( .B1(n8273), .B2(n7907), .A(n7962), .ZN(n7910) );
  NAND2_X1 U6259 ( .A1(n5257), .A2(n5256), .ZN(n5259) );
  NOR2_X2 U6260 ( .A1(n7920), .A2(n8075), .ZN(n7999) );
  INV_X1 U6261 ( .A(n9349), .ZN(n4512) );
  NAND2_X1 U6262 ( .A1(n9365), .A2(n4511), .ZN(n6104) );
  OAI21_X1 U6263 ( .B1(n6218), .B2(n9843), .A(n6219), .ZN(n6220) );
  NOR2_X1 U6264 ( .A1(n8492), .A2(n8166), .ZN(n8174) );
  NAND2_X1 U6265 ( .A1(n7077), .A2(n7078), .ZN(n7108) );
  NOR2_X1 U6266 ( .A1(n5342), .A2(n7111), .ZN(n7245) );
  NOR2_X1 U6267 ( .A1(n7372), .A2(n5381), .ZN(n7462) );
  NOR2_X1 U6268 ( .A1(n7248), .A2(n7247), .ZN(n7371) );
  NOR2_X1 U6269 ( .A1(n7462), .A2(n7463), .ZN(n7466) );
  NOR2_X1 U6270 ( .A1(n8087), .A2(n7497), .ZN(n7500) );
  XNOR2_X1 U6271 ( .A(n7496), .B(n8097), .ZN(n8088) );
  OR2_X1 U6272 ( .A1(n9867), .A2(n10182), .ZN(n9866) );
  INV_X1 U6273 ( .A(n7007), .ZN(n4809) );
  NOR2_X1 U6274 ( .A1(n8088), .A2(n8503), .ZN(n8087) );
  NAND2_X1 U6275 ( .A1(n7005), .A2(n7004), .ZN(n4811) );
  XNOR2_X1 U6276 ( .A(n7461), .B(n7468), .ZN(n7372) );
  NOR2_X1 U6277 ( .A1(n7466), .A2(n7465), .ZN(n7494) );
  NAND2_X1 U6278 ( .A1(n4924), .A2(n4923), .ZN(n4922) );
  NOR2_X2 U6279 ( .A1(n8182), .A2(n8181), .ZN(n8205) );
  AOI21_X1 U6280 ( .B1(n7742), .B2(n7739), .A(n7572), .ZN(n4504) );
  NAND2_X1 U6281 ( .A1(n5515), .A2(n10235), .ZN(n5516) );
  NAND2_X1 U6282 ( .A1(n5221), .A2(n5111), .ZN(n5236) );
  OAI21_X1 U6283 ( .B1(n5333), .B2(n4699), .A(n4696), .ZN(n5389) );
  OAI21_X1 U6284 ( .B1(n5102), .B2(n5160), .A(n4927), .ZN(n5103) );
  OAI21_X1 U6285 ( .B1(n5535), .B2(n5534), .A(n5533), .ZN(n5550) );
  NAND2_X1 U6286 ( .A1(n4515), .A2(n4504), .ZN(n4935) );
  NAND2_X1 U6287 ( .A1(n5567), .A2(n5566), .ZN(n5585) );
  OR2_X1 U6288 ( .A1(n5103), .A2(SI_1_), .ZN(n5104) );
  OAI21_X1 U6289 ( .B1(n5515), .B2(n10235), .A(n5514), .ZN(n5517) );
  NAND2_X1 U6290 ( .A1(n5565), .A2(n5564), .ZN(n5567) );
  OAI21_X2 U6291 ( .B1(n7999), .B2(n7998), .A(n7997), .ZN(n7996) );
  NOR2_X2 U6292 ( .A1(n7943), .A2(n7942), .ZN(n7945) );
  NAND2_X1 U6293 ( .A1(n4894), .A2(n4892), .ZN(n7899) );
  NAND2_X1 U6294 ( .A1(n8006), .A2(n6902), .ZN(n7978) );
  NAND2_X1 U6295 ( .A1(n7978), .A2(n7977), .ZN(n6907) );
  NAND2_X1 U6296 ( .A1(n6850), .A2(n6846), .ZN(n6848) );
  INV_X1 U6297 ( .A(n6712), .ZN(n4510) );
  NAND2_X1 U6298 ( .A1(n4820), .A2(n4819), .ZN(n8165) );
  OAI21_X1 U6299 ( .B1(n8225), .B2(n8224), .A(n4921), .ZN(P2_U3201) );
  NOR2_X1 U6300 ( .A1(n7371), .A2(n4822), .ZN(n7461) );
  NOR2_X1 U6301 ( .A1(n7245), .A2(n4812), .ZN(n7248) );
  XNOR2_X2 U6302 ( .A(n5241), .B(n5240), .ZN(n6481) );
  INV_X1 U6303 ( .A(n4845), .ZN(n9477) );
  NAND2_X1 U6304 ( .A1(n4937), .A2(n4936), .ZN(n4515) );
  NAND3_X1 U6305 ( .A1(n4690), .A2(n4516), .A3(n4692), .ZN(n7715) );
  NAND4_X1 U6306 ( .A1(n4471), .A2(n7706), .A3(n7707), .A4(n7708), .ZN(n4516)
         );
  NAND2_X1 U6307 ( .A1(n7685), .A2(n4685), .ZN(n7686) );
  AOI21_X1 U6308 ( .B1(n4709), .B2(n7735), .A(n7734), .ZN(n4705) );
  NAND3_X1 U6309 ( .A1(n7712), .A2(n7711), .A3(n7739), .ZN(n4518) );
  INV_X1 U6310 ( .A(n4743), .ZN(n4519) );
  NAND2_X1 U6311 ( .A1(n7793), .A2(n4522), .ZN(n4521) );
  NAND2_X2 U6312 ( .A1(n8783), .A2(n7807), .ZN(n8867) );
  INV_X1 U6313 ( .A(n8615), .ZN(n4528) );
  NAND2_X1 U6314 ( .A1(n8615), .A2(n8616), .ZN(n8614) );
  OR2_X1 U6315 ( .A1(n8615), .A2(n4531), .ZN(n4527) );
  NAND2_X2 U6316 ( .A1(n4532), .A2(n6520), .ZN(n8651) );
  NAND2_X1 U6317 ( .A1(n8670), .A2(n8819), .ZN(n8820) );
  INV_X1 U6318 ( .A(n8771), .ZN(n8878) );
  INV_X1 U6319 ( .A(n7774), .ZN(n4535) );
  NAND2_X1 U6320 ( .A1(n4535), .A2(n4482), .ZN(n4539) );
  NAND2_X1 U6321 ( .A1(n4539), .A2(n4536), .ZN(n5019) );
  AND2_X2 U6322 ( .A1(n5980), .A2(n4429), .ZN(n6188) );
  NAND2_X1 U6323 ( .A1(n7226), .A2(n4552), .ZN(n4549) );
  NAND2_X1 U6324 ( .A1(n9545), .A2(n4861), .ZN(n4858) );
  NAND2_X1 U6325 ( .A1(n5324), .A2(n5136), .ZN(n4558) );
  OAI21_X1 U6326 ( .B1(n5324), .B2(n4562), .A(n4559), .ZN(n5353) );
  NAND4_X1 U6327 ( .A1(n5911), .A2(n4566), .A3(n4565), .A4(n4564), .ZN(n5014)
         );
  NAND2_X2 U6328 ( .A1(n6170), .A2(n9183), .ZN(n5873) );
  XNOR2_X2 U6329 ( .A(n4568), .B(n10046), .ZN(n9183) );
  INV_X1 U6330 ( .A(n4575), .ZN(n9514) );
  NAND2_X1 U6331 ( .A1(n4578), .A2(n7028), .ZN(n4577) );
  INV_X1 U6332 ( .A(n4585), .ZN(n9436) );
  NAND2_X1 U6333 ( .A1(n9374), .A2(n4586), .ZN(n9304) );
  NAND2_X1 U6334 ( .A1(n9374), .A2(n9356), .ZN(n9350) );
  INV_X1 U6335 ( .A(n4594), .ZN(n4593) );
  NAND2_X1 U6336 ( .A1(n4597), .A2(n7086), .ZN(n4595) );
  NAND2_X1 U6337 ( .A1(n6306), .A2(n9915), .ZN(n4601) );
  NAND2_X1 U6338 ( .A1(n7103), .A2(n4476), .ZN(n4606) );
  NAND2_X1 U6339 ( .A1(n4606), .A2(n4607), .ZN(n7379) );
  NAND2_X1 U6340 ( .A1(n4611), .A2(n6265), .ZN(n6263) );
  INV_X1 U6341 ( .A(n6481), .ZN(n4613) );
  NAND2_X1 U6342 ( .A1(n7491), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U6343 ( .A1(n4625), .A2(n4623), .ZN(n9154) );
  NAND2_X1 U6344 ( .A1(n9048), .A2(n4422), .ZN(n4625) );
  NAND2_X1 U6345 ( .A1(n9008), .A2(n9126), .ZN(n4626) );
  NAND2_X1 U6346 ( .A1(n4628), .A2(n9009), .ZN(n4627) );
  NAND2_X1 U6347 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  INV_X1 U6348 ( .A(n9007), .ZN(n4629) );
  NAND2_X1 U6349 ( .A1(n9008), .A2(n9011), .ZN(n4630) );
  NAND2_X1 U6350 ( .A1(n4639), .A2(n4444), .ZN(n8993) );
  NAND2_X1 U6351 ( .A1(n8975), .A2(n4642), .ZN(n4639) );
  NAND2_X1 U6352 ( .A1(n8974), .A2(n8973), .ZN(n4658) );
  INV_X1 U6353 ( .A(n9092), .ZN(n4660) );
  NAND2_X1 U6354 ( .A1(n8929), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U6355 ( .A1(n4664), .A2(n4662), .ZN(n8927) );
  OAI21_X2 U6356 ( .B1(n8951), .B2(n8950), .A(n9495), .ZN(n8957) );
  NAND3_X1 U6357 ( .A1(n4683), .A2(n6161), .A3(n6162), .ZN(n8902) );
  MUX2_X1 U6358 ( .A(n6368), .B(P1_REG2_REG_1__SCAN_IN), .S(n6378), .Z(n9173)
         );
  NAND3_X1 U6359 ( .A1(n4730), .A2(n4728), .A3(n4727), .ZN(P1_U3262) );
  OAI21_X2 U6360 ( .B1(n8820), .B2(n4742), .A(n4428), .ZN(n8702) );
  INV_X1 U6361 ( .A(n5014), .ZN(n4745) );
  NAND3_X1 U6362 ( .A1(n4744), .A2(n4745), .A3(n4747), .ZN(n5995) );
  NAND2_X1 U6363 ( .A1(n6571), .A2(n6572), .ZN(n4750) );
  NAND2_X1 U6364 ( .A1(n6570), .A2(n4752), .ZN(n4751) );
  NAND2_X1 U6365 ( .A1(n4753), .A2(n5010), .ZN(n4752) );
  INV_X1 U6366 ( .A(n6572), .ZN(n4753) );
  XNOR2_X1 U6367 ( .A(n6181), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6154) );
  OAI21_X2 U6368 ( .B1(n6151), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6150) );
  OAI211_X1 U6369 ( .C1(n6306), .C2(n5189), .A(n5224), .B(n5225), .ZN(n5226)
         );
  INV_X2 U6370 ( .A(n5161), .ZN(n5001) );
  NAND2_X1 U6371 ( .A1(n5689), .A2(n8413), .ZN(n4763) );
  NAND2_X1 U6372 ( .A1(n4763), .A2(n4419), .ZN(n5760) );
  AND2_X1 U6373 ( .A1(n4763), .A2(n4762), .ZN(n7852) );
  INV_X1 U6374 ( .A(n7014), .ZN(n4769) );
  NAND2_X1 U6375 ( .A1(n8337), .A2(n4776), .ZN(n4774) );
  NAND2_X1 U6376 ( .A1(n4781), .A2(n4783), .ZN(n5657) );
  NAND2_X1 U6377 ( .A1(n8262), .A2(n4784), .ZN(n4781) );
  NAND2_X1 U6378 ( .A1(n8262), .A2(n4791), .ZN(n4787) );
  AOI21_X1 U6379 ( .B1(n8262), .B2(n8267), .A(n5604), .ZN(n8254) );
  OAI21_X1 U6380 ( .B1(n7214), .B2(n4799), .A(n4797), .ZN(n4795) );
  NAND2_X1 U6381 ( .A1(n9900), .A2(n5230), .ZN(n6767) );
  NAND2_X1 U6382 ( .A1(n5563), .A2(n5562), .ZN(n8271) );
  NAND2_X1 U6383 ( .A1(n6540), .A2(n5044), .ZN(n6550) );
  NAND2_X1 U6384 ( .A1(n5019), .A2(n5018), .ZN(n8837) );
  NAND2_X1 U6385 ( .A1(n8828), .A2(n8637), .ZN(n8755) );
  NOR2_X1 U6386 ( .A1(n8344), .A2(n5475), .ZN(n5476) );
  NAND2_X1 U6387 ( .A1(n5228), .A2(n9901), .ZN(n9900) );
  OR2_X1 U6388 ( .A1(n5222), .A2(n6305), .ZN(n5224) );
  MUX2_X1 U6389 ( .A(n7694), .B(n7693), .S(n7739), .Z(n7705) );
  OAI21_X1 U6390 ( .B1(n7720), .B2(n8267), .A(n7719), .ZN(n7725) );
  NAND2_X1 U6391 ( .A1(n5236), .A2(n5235), .ZN(n5238) );
  NOR2_X4 U6392 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6257) );
  NAND3_X1 U6393 ( .A1(n4814), .A2(n4477), .A3(n4813), .ZN(n9891) );
  NAND3_X1 U6394 ( .A1(n4818), .A2(n4815), .A3(P2_REG1_REG_2__SCAN_IN), .ZN(
        n4814) );
  INV_X1 U6395 ( .A(n6257), .ZN(n4817) );
  NAND2_X1 U6396 ( .A1(n4413), .A2(n8104), .ZN(n4819) );
  XNOR2_X1 U6397 ( .A(n8123), .B(n8138), .ZN(n8104) );
  INV_X1 U6398 ( .A(n4821), .ZN(n8124) );
  NAND2_X1 U6399 ( .A1(n6938), .A2(n4832), .ZN(n4830) );
  NAND2_X1 U6400 ( .A1(n4830), .A2(n4831), .ZN(n7129) );
  AOI21_X1 U6401 ( .B1(n4832), .B2(n4835), .A(n4460), .ZN(n4831) );
  NAND2_X1 U6402 ( .A1(n6045), .A2(n4838), .ZN(n4836) );
  NOR2_X1 U6403 ( .A1(n6045), .A2(n4436), .ZN(n9444) );
  INV_X1 U6404 ( .A(n4514), .ZN(n6158) );
  NAND2_X1 U6405 ( .A1(n6277), .A2(n9017), .ZN(n6276) );
  OAI21_X1 U6406 ( .B1(n9522), .B2(n4846), .A(n4847), .ZN(n4845) );
  OR2_X1 U6407 ( .A1(n9522), .A2(n6021), .ZN(n4854) );
  OR2_X1 U6408 ( .A1(n4849), .A2(n6021), .ZN(n4846) );
  XNOR2_X2 U6409 ( .A(n4857), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5771) );
  OAI21_X2 U6410 ( .B1(n9697), .B2(P1_IR_REG_29__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U6411 ( .A1(n4865), .A2(n6167), .ZN(n4864) );
  NAND2_X1 U6412 ( .A1(n6166), .A2(n4866), .ZN(n4865) );
  NAND2_X1 U6413 ( .A1(n7124), .A2(n6167), .ZN(n7122) );
  NAND2_X1 U6414 ( .A1(n6166), .A2(n4866), .ZN(n7124) );
  NAND2_X1 U6415 ( .A1(n9391), .A2(n9390), .ZN(n4873) );
  OAI21_X1 U6416 ( .B1(n9490), .B2(n4877), .A(n4874), .ZN(n9461) );
  NAND3_X1 U6417 ( .A1(n5980), .A2(n5038), .A3(n4429), .ZN(n5780) );
  NAND2_X1 U6418 ( .A1(n7883), .A2(n7884), .ZN(n7989) );
  NAND2_X1 U6419 ( .A1(n6898), .A2(n4441), .ZN(n8006) );
  NAND2_X1 U6420 ( .A1(n7952), .A2(n4895), .ZN(n4894) );
  INV_X1 U6421 ( .A(n7911), .ZN(n4901) );
  NOR2_X1 U6422 ( .A1(n4901), .A2(n7912), .ZN(n4900) );
  NAND2_X1 U6423 ( .A1(n4902), .A2(n4903), .ZN(n8055) );
  NAND3_X1 U6424 ( .A1(n7415), .A2(n7414), .A3(n4905), .ZN(n4902) );
  NAND2_X1 U6425 ( .A1(n7415), .A2(n7414), .ZN(n7439) );
  NAND2_X1 U6426 ( .A1(n5065), .A2(n5254), .ZN(n5161) );
  NAND2_X1 U6427 ( .A1(n7200), .A2(n4909), .ZN(n7863) );
  NAND2_X1 U6428 ( .A1(n7863), .A2(n4474), .ZN(n7276) );
  NAND2_X1 U6429 ( .A1(n6705), .A2(n6840), .ZN(n6854) );
  NAND2_X1 U6430 ( .A1(n6995), .A2(n4917), .ZN(n4915) );
  NAND2_X1 U6431 ( .A1(n5160), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U6432 ( .A1(n5391), .A2(n4481), .ZN(n4931) );
  OAI21_X1 U6433 ( .B1(n4934), .B2(n7746), .A(n4933), .ZN(n7747) );
  NAND2_X1 U6434 ( .A1(n4934), .A2(n7745), .ZN(n4933) );
  NAND2_X1 U6435 ( .A1(n4935), .A2(n7743), .ZN(n4934) );
  INV_X1 U6436 ( .A(n7742), .ZN(n4937) );
  NAND3_X1 U6437 ( .A1(n4942), .A2(n4945), .A3(n4941), .ZN(n4939) );
  NAND2_X1 U6438 ( .A1(n5645), .A2(n4967), .ZN(n4965) );
  NAND2_X1 U6439 ( .A1(n6982), .A2(n5692), .ZN(n4971) );
  NAND2_X1 U6440 ( .A1(n4971), .A2(n9897), .ZN(n9896) );
  OAI21_X1 U6441 ( .B1(n9897), .B2(n4971), .A(n9896), .ZN(n9926) );
  NAND3_X1 U6442 ( .A1(n7519), .A2(n5091), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n5187) );
  XNOR2_X2 U6443 ( .A(n5079), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6444 ( .A1(n5695), .A2(n4980), .ZN(n7331) );
  OAI21_X2 U6445 ( .B1(n8300), .B2(n4985), .A(n4982), .ZN(n8252) );
  NAND2_X1 U6446 ( .A1(n4997), .A2(n4480), .ZN(n7212) );
  NAND2_X1 U6447 ( .A1(n5698), .A2(n4998), .ZN(n8426) );
  INV_X1 U6448 ( .A(n5690), .ZN(n7547) );
  NAND2_X1 U6449 ( .A1(n5009), .A2(n7700), .ZN(n8350) );
  NAND4_X1 U6450 ( .A1(n5936), .A2(n5016), .A3(n5765), .A4(n5012), .ZN(n5011)
         );
  NAND3_X1 U6451 ( .A1(n5013), .A2(n5868), .A3(n5936), .ZN(n5967) );
  INV_X1 U6452 ( .A(n8649), .ZN(n5025) );
  NAND2_X1 U6453 ( .A1(n5025), .A2(n8719), .ZN(n5028) );
  OAI21_X2 U6454 ( .B1(n7296), .B2(n5031), .A(n5029), .ZN(n7774) );
  NAND2_X1 U6455 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  NAND2_X1 U6456 ( .A1(n8633), .A2(n5032), .ZN(n8828) );
  NOR2_X1 U6457 ( .A1(n8674), .A2(n6536), .ZN(n6537) );
  XNOR2_X1 U6458 ( .A(n9340), .B(n9339), .ZN(n9581) );
  INV_X1 U6459 ( .A(n9902), .ZN(n5206) );
  AOI22_X2 U6460 ( .A1(n9398), .A2(n6089), .B1(n9424), .B2(n9407), .ZN(n9382)
         );
  NAND2_X1 U6461 ( .A1(n5211), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5204) );
  CLKBUF_X1 U6462 ( .A(n6559), .Z(n6583) );
  NAND2_X1 U6463 ( .A1(n9697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6464 ( .A1(n5183), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6465 ( .A1(n4418), .A2(n7101), .ZN(n5319) );
  AND2_X1 U6466 ( .A1(n8631), .A2(n8630), .ZN(n5039) );
  INV_X1 U6467 ( .A(n9992), .ZN(n9990) );
  AND2_X1 U6468 ( .A1(n5747), .A2(n5746), .ZN(n9975) );
  OR2_X1 U6469 ( .A1(n5246), .A2(n5245), .ZN(n5041) );
  OR2_X1 U6470 ( .A1(n8805), .A2(n9168), .ZN(n5042) );
  INV_X1 U6471 ( .A(n8731), .ZN(n5954) );
  AND2_X1 U6472 ( .A1(n8788), .A2(n7809), .ZN(n5043) );
  AND2_X1 U6473 ( .A1(n6549), .A2(n6535), .ZN(n5044) );
  INV_X1 U6474 ( .A(n9170), .ZN(n6552) );
  OR2_X1 U6475 ( .A1(n7855), .A2(n8566), .ZN(n5045) );
  OR2_X1 U6476 ( .A1(n6178), .A2(n9689), .ZN(n5046) );
  OR2_X1 U6477 ( .A1(n7361), .A2(n7341), .ZN(n5047) );
  OR2_X1 U6478 ( .A1(n9169), .A2(n6875), .ZN(n5050) );
  OR2_X1 U6479 ( .A1(n6178), .A2(n9645), .ZN(n5051) );
  OR2_X1 U6480 ( .A1(n7855), .A2(n8491), .ZN(n5052) );
  INV_X1 U6481 ( .A(n7545), .ZN(n5696) );
  INV_X1 U6482 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5078) );
  AND2_X1 U6483 ( .A1(n7898), .A2(n8076), .ZN(n5053) );
  AND2_X1 U6484 ( .A1(n5960), .A2(n5959), .ZN(n5054) );
  INV_X1 U6485 ( .A(n8768), .ZN(n5977) );
  INV_X1 U6486 ( .A(n8081), .ZN(n7334) );
  INV_X4 U6487 ( .A(n7533), .ZN(n5133) );
  INV_X1 U6488 ( .A(n5160), .ZN(n7533) );
  OR2_X1 U6489 ( .A1(n6961), .A2(n9167), .ZN(n5055) );
  INV_X1 U6490 ( .A(n9383), .ZN(n9406) );
  AND2_X1 U6491 ( .A1(n8567), .A2(n8335), .ZN(n5056) );
  NAND2_X1 U6492 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  INV_X1 U6493 ( .A(n7642), .ZN(n5694) );
  AND2_X1 U6494 ( .A1(n7550), .A2(n7215), .ZN(n5057) );
  NAND2_X1 U6495 ( .A1(n5798), .A2(n5790), .ZN(n5801) );
  OAI211_X1 U6496 ( .C1(n7593), .C2(n7592), .A(n7710), .B(n4995), .ZN(n7594)
         );
  INV_X1 U6497 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5062) );
  INV_X1 U6498 ( .A(n9927), .ZN(n5245) );
  INV_X1 U6499 ( .A(n6811), .ZN(n6812) );
  NAND2_X1 U6500 ( .A1(n8520), .A2(n8072), .ZN(n5656) );
  OR2_X1 U6501 ( .A1(n8323), .A2(n8077), .ZN(n5512) );
  AND2_X1 U6502 ( .A1(n8083), .A2(n6916), .ZN(n5298) );
  NAND2_X1 U6503 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U6504 ( .A1(n8537), .A2(n8284), .ZN(n5582) );
  AND2_X1 U6505 ( .A1(n7625), .A2(n7138), .ZN(n7628) );
  INV_X1 U6506 ( .A(n8351), .ZN(n5705) );
  OR2_X1 U6507 ( .A1(n8509), .A2(n8409), .ZN(n5386) );
  OR2_X1 U6508 ( .A1(n5229), .A2(n5226), .ZN(n5230) );
  NOR2_X1 U6509 ( .A1(n8786), .A2(n8784), .ZN(n7806) );
  NAND2_X1 U6510 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  NAND2_X1 U6511 ( .A1(n6153), .A2(n9139), .ZN(n6501) );
  INV_X1 U6512 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5899) );
  INV_X1 U6513 ( .A(n9160), .ZN(n5993) );
  INV_X1 U6514 ( .A(n9163), .ZN(n5953) );
  INV_X1 U6515 ( .A(n6866), .ZN(n5860) );
  INV_X1 U6516 ( .A(SI_15_), .ZN(n5157) );
  INV_X1 U6517 ( .A(n7899), .ZN(n7902) );
  INV_X1 U6518 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6519 ( .A1(n8559), .A2(n8347), .ZN(n7707) );
  OR2_X1 U6520 ( .A1(n7538), .A2(n5099), .ZN(n5244) );
  NOR2_X1 U6521 ( .A1(n5043), .A2(n7806), .ZN(n7807) );
  OAI22_X1 U6522 ( .A1(n6527), .A2(n6696), .B1(n6591), .B2(n8651), .ZN(n6536)
         );
  BUF_X4 U6523 ( .A(n8736), .Z(n8741) );
  AND2_X1 U6524 ( .A1(n6013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U6525 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6108), .ZN(n6127) );
  OR2_X1 U6526 ( .A1(n6081), .A2(n6080), .ZN(n6092) );
  NAND2_X1 U6527 ( .A1(n6015), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6026) );
  INV_X1 U6528 ( .A(n9314), .ZN(n6178) );
  INV_X1 U6529 ( .A(n9470), .ZN(n6177) );
  NOR2_X1 U6530 ( .A1(n5960), .A2(n5959), .ZN(n5971) );
  NAND2_X1 U6531 ( .A1(n6552), .A2(n6866), .ZN(n6162) );
  NAND2_X1 U6532 ( .A1(n5146), .A2(SI_12_), .ZN(n5150) );
  NAND2_X1 U6533 ( .A1(n5128), .A2(SI_7_), .ZN(n5132) );
  OAI21_X1 U6534 ( .B1(n7970), .B2(n7968), .A(n8386), .ZN(n7883) );
  OR2_X1 U6535 ( .A1(n5210), .A2(n8442), .ZN(n5383) );
  OR2_X1 U6536 ( .A1(n4417), .A2(n6225), .ZN(n5231) );
  OR2_X1 U6537 ( .A1(n6606), .A2(n5726), .ZN(n5758) );
  NOR2_X1 U6538 ( .A1(n4443), .A2(n8276), .ZN(n8277) );
  NAND2_X1 U6539 ( .A1(n7703), .A2(n7707), .ZN(n8331) );
  NOR2_X1 U6540 ( .A1(n6092), .A2(n8823), .ZN(n6093) );
  AND2_X1 U6541 ( .A1(n6049), .A2(n5763), .ZN(n6058) );
  NOR2_X1 U6542 ( .A1(n6038), .A2(n6037), .ZN(n6049) );
  NAND2_X1 U6543 ( .A1(n8976), .A2(n8987), .ZN(n9366) );
  INV_X1 U6544 ( .A(n7350), .ZN(n9558) );
  NAND2_X1 U6545 ( .A1(n6748), .A2(n5861), .ZN(n6759) );
  INV_X2 U6546 ( .A(n9004), .ZN(n9049) );
  INV_X1 U6547 ( .A(n9164), .ZN(n8728) );
  NAND2_X1 U6548 ( .A1(n7026), .A2(n5908), .ZN(n6947) );
  AND2_X1 U6549 ( .A1(n5111), .A2(n5110), .ZN(n5218) );
  NAND2_X1 U6550 ( .A1(n7422), .A2(n7537), .ZN(n5572) );
  AND2_X1 U6551 ( .A1(n5655), .A2(n5654), .ZN(n7916) );
  AND2_X1 U6552 ( .A1(n5581), .A2(n5580), .ZN(n8284) );
  OR2_X1 U6553 ( .A1(n5210), .A2(n7869), .ZN(n5305) );
  XNOR2_X1 U6554 ( .A(n7844), .B(n7843), .ZN(n7848) );
  AND2_X1 U6555 ( .A1(n9913), .A2(n9912), .ZN(n8419) );
  OR2_X1 U6556 ( .A1(n9992), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5761) );
  AND2_X1 U6557 ( .A1(n5758), .A2(n5757), .ZN(n6612) );
  OR2_X1 U6558 ( .A1(n9973), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5748) );
  AND2_X1 U6559 ( .A1(n5725), .A2(n5724), .ZN(n6610) );
  OR2_X1 U6560 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  INV_X1 U6561 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5240) );
  AND4_X1 U6562 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n9053)
         );
  OR2_X1 U6563 ( .A1(n6070), .A2(n9190), .ZN(n5844) );
  AOI211_X1 U6564 ( .C1(n9574), .C2(n4439), .A(n9557), .B(n4589), .ZN(n9573)
         );
  AND2_X1 U6565 ( .A1(n8962), .A2(n8967), .ZN(n9423) );
  INV_X1 U6566 ( .A(n9521), .ZN(n9502) );
  INV_X1 U6567 ( .A(n8469), .ZN(n8290) );
  AND2_X1 U6568 ( .A1(n6621), .A2(n6620), .ZN(n8056) );
  INV_X1 U6569 ( .A(n7916), .ZN(n8072) );
  AND3_X1 U6570 ( .A1(n5529), .A2(n5528), .A3(n5527), .ZN(n8320) );
  INV_X1 U6571 ( .A(n8441), .ZN(n8409) );
  OR2_X1 U6572 ( .A1(P2_U3150), .A2(n6235), .ZN(n9887) );
  INV_X1 U6573 ( .A(n8419), .ZN(n8448) );
  XNOR2_X1 U6574 ( .A(n8233), .B(n8232), .ZN(n8523) );
  INV_X1 U6575 ( .A(n5530), .ZN(n8552) );
  OR2_X1 U6576 ( .A1(n6514), .A2(n6513), .ZN(n8899) );
  INV_X1 U6577 ( .A(n9313), .ZN(n9811) );
  INV_X1 U6578 ( .A(n9513), .ZN(n9541) );
  OR2_X1 U6579 ( .A1(n6217), .A2(n6497), .ZN(n9843) );
  INV_X1 U6580 ( .A(n9375), .ZN(n9669) );
  INV_X1 U6581 ( .A(n9838), .ZN(n9839) );
  INV_X1 U6582 ( .A(n9838), .ZN(n9691) );
  AND2_X1 U6583 ( .A1(n6521), .A2(n6194), .ZN(n9693) );
  NAND4_X1 U6584 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n5064)
         );
  NOR2_X1 U6585 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NOR3_X1 U6586 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5070) );
  INV_X1 U6587 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5159) );
  INV_X1 U6588 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  INV_X1 U6589 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6590 ( .A1(n5076), .A2(n5075), .ZN(n8604) );
  NAND2_X2 U6591 ( .A1(n8604), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6592 ( .A1(n6922), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5095) );
  INV_X1 U6593 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8575) );
  OR2_X1 U6594 ( .A1(n5208), .A2(n8575), .ZN(n5094) );
  INV_X2 U6595 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6772) );
  INV_X1 U6596 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7112) );
  INV_X1 U6598 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5085) );
  INV_X1 U6599 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10200) );
  OR2_X2 U6600 ( .A1(n5411), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5428) );
  INV_X1 U6601 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6602 ( .A1(n5430), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5090) );
  AND2_X1 U6603 ( .A1(n5451), .A2(n5090), .ZN(n8378) );
  OR2_X1 U6604 ( .A1(n5210), .A2(n8378), .ZN(n5093) );
  INV_X1 U6605 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8377) );
  OR2_X1 U6606 ( .A1(n4417), .A2(n8377), .ZN(n5092) );
  NAND2_X1 U6607 ( .A1(n5103), .A2(SI_1_), .ZN(n5106) );
  MUX2_X1 U6608 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5160), .Z(n5105) );
  AND2_X1 U6609 ( .A1(n5105), .A2(SI_0_), .ZN(n5191) );
  NAND2_X1 U6610 ( .A1(n5195), .A2(n5106), .ZN(n5219) );
  MUX2_X1 U6611 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5160), .Z(n5107) );
  NAND2_X1 U6612 ( .A1(n5107), .A2(SI_2_), .ZN(n5111) );
  INV_X1 U6613 ( .A(n5107), .ZN(n5109) );
  INV_X1 U6614 ( .A(SI_2_), .ZN(n5108) );
  NAND2_X1 U6615 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  NAND2_X1 U6616 ( .A1(n5219), .A2(n5218), .ZN(n5221) );
  MUX2_X1 U6617 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5160), .Z(n5113) );
  INV_X1 U6618 ( .A(n5113), .ZN(n5115) );
  INV_X1 U6619 ( .A(SI_4_), .ZN(n5114) );
  NAND2_X1 U6620 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  MUX2_X1 U6621 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5133), .Z(n5118) );
  INV_X1 U6622 ( .A(n5118), .ZN(n5120) );
  INV_X1 U6623 ( .A(SI_5_), .ZN(n5119) );
  NAND2_X1 U6624 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  INV_X1 U6625 ( .A(n5123), .ZN(n5125) );
  INV_X1 U6626 ( .A(SI_6_), .ZN(n5124) );
  NAND2_X1 U6627 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  MUX2_X1 U6628 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5133), .Z(n5128) );
  INV_X1 U6629 ( .A(n5128), .ZN(n5130) );
  INV_X1 U6630 ( .A(SI_7_), .ZN(n5129) );
  NAND2_X1 U6631 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  MUX2_X1 U6632 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5133), .Z(n5134) );
  INV_X1 U6633 ( .A(n5134), .ZN(n5135) );
  INV_X1 U6634 ( .A(SI_8_), .ZN(n10113) );
  INV_X1 U6635 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6331) );
  INV_X1 U6636 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6458) );
  MUX2_X1 U6637 ( .A(n6331), .B(n6458), .S(n5133), .Z(n5137) );
  INV_X1 U6638 ( .A(n5137), .ZN(n5138) );
  MUX2_X1 U6639 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5133), .Z(n5140) );
  NAND2_X1 U6640 ( .A1(n5140), .A2(SI_10_), .ZN(n5144) );
  INV_X1 U6641 ( .A(n5140), .ZN(n5142) );
  INV_X1 U6642 ( .A(SI_10_), .ZN(n5141) );
  NAND2_X1 U6643 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  MUX2_X1 U6644 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5133), .Z(n5145) );
  MUX2_X1 U6645 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5133), .Z(n5146) );
  INV_X1 U6646 ( .A(n5146), .ZN(n5148) );
  INV_X1 U6647 ( .A(SI_12_), .ZN(n5147) );
  NAND2_X1 U6648 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  MUX2_X1 U6649 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5133), .Z(n5151) );
  INV_X1 U6650 ( .A(n5151), .ZN(n5152) );
  INV_X1 U6651 ( .A(SI_13_), .ZN(n10094) );
  NAND2_X1 U6652 ( .A1(n5152), .A2(n10094), .ZN(n5153) );
  MUX2_X1 U6653 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5133), .Z(n5403) );
  MUX2_X1 U6654 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5133), .Z(n5419) );
  INV_X1 U6655 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6600) );
  INV_X1 U6656 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10228) );
  MUX2_X1 U6657 ( .A(n6600), .B(n10228), .S(n5133), .Z(n5437) );
  XNOR2_X1 U6658 ( .A(n5437), .B(SI_16_), .ZN(n5158) );
  NAND2_X1 U6659 ( .A1(n6599), .A2(n7537), .ZN(n5166) );
  NAND2_X1 U6660 ( .A1(n5161), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6661 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5162), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5164) );
  AND2_X1 U6662 ( .A1(n5164), .A2(n5163), .ZN(n8141) );
  AOI22_X1 U6663 ( .A1(n5488), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5487), .B2(
        n8141), .ZN(n5165) );
  INV_X1 U6664 ( .A(n8576), .ZN(n5436) );
  CLKBUF_X3 U6665 ( .A(n5200), .Z(n6921) );
  NAND2_X1 U6666 ( .A1(n6921), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5171) );
  INV_X1 U6667 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8432) );
  OR2_X1 U6668 ( .A1(n4418), .A2(n8432), .ZN(n5170) );
  NAND2_X1 U6669 ( .A1(n5380), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5167) );
  AND2_X1 U6670 ( .A1(n5397), .A2(n5167), .ZN(n8431) );
  OR2_X1 U6671 ( .A1(n5210), .A2(n8431), .ZN(n5169) );
  INV_X1 U6672 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8510) );
  OR2_X1 U6673 ( .A1(n5199), .A2(n8510), .ZN(n5168) );
  NAND2_X1 U6674 ( .A1(n5173), .A2(n5172), .ZN(n5175) );
  NAND2_X1 U6675 ( .A1(n5175), .A2(n5174), .ZN(n6366) );
  OR2_X1 U6676 ( .A1(n6366), .A2(n5222), .ZN(n5182) );
  NAND2_X1 U6677 ( .A1(n5254), .A2(n10177), .ZN(n5271) );
  NOR2_X1 U6678 ( .A1(n5292), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5312) );
  INV_X1 U6679 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5176) );
  INV_X1 U6680 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5357) );
  AND4_X1 U6681 ( .A1(n5325), .A2(n5337), .A3(n5176), .A4(n5357), .ZN(n5177)
         );
  AND2_X1 U6682 ( .A1(n5312), .A2(n5177), .ZN(n5372) );
  INV_X1 U6683 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6684 ( .A1(n5372), .A2(n5178), .ZN(n5392) );
  NAND2_X1 U6685 ( .A1(n5392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5180) );
  INV_X1 U6686 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6687 ( .A(n5180), .B(n5179), .ZN(n7495) );
  INV_X1 U6688 ( .A(n7495), .ZN(n7479) );
  AOI22_X1 U6689 ( .A1(n5488), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5487), .B2(
        n7479), .ZN(n5181) );
  INV_X1 U6690 ( .A(n5199), .ZN(n5183) );
  NAND2_X1 U6691 ( .A1(n5200), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5185) );
  INV_X1 U6692 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U6693 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5188) );
  INV_X1 U6694 ( .A(n5190), .ZN(n5193) );
  INV_X1 U6695 ( .A(n5191), .ZN(n5192) );
  NAND2_X1 U6696 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  NOR2_X1 U6697 ( .A1(n6579), .A2(n5196), .ZN(n9902) );
  NAND2_X1 U6698 ( .A1(n6579), .A2(n9918), .ZN(n7607) );
  INV_X1 U6699 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5198) );
  INV_X1 U6700 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U6701 ( .A1(n5200), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6702 ( .A1(n7533), .A2(SI_0_), .ZN(n5205) );
  XNOR2_X1 U6703 ( .A(n5205), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8613) );
  MUX2_X1 U6704 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8613), .S(n5189), .Z(n7758) );
  NAND2_X1 U6705 ( .A1(n6987), .A2(n7758), .ZN(n6985) );
  NAND2_X1 U6706 ( .A1(n5690), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U6707 ( .A1(n5206), .A2(n6984), .ZN(n5228) );
  INV_X1 U6708 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5207) );
  INV_X1 U6709 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6710 ( .A1(n5210), .A2(n5209), .ZN(n5213) );
  NAND2_X1 U6711 ( .A1(n5211), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5212) );
  AND2_X1 U6712 ( .A1(n5213), .A2(n5212), .ZN(n5215) );
  NAND3_X2 U6713 ( .A1(n5216), .A2(n5215), .A3(n5214), .ZN(n5229) );
  INV_X1 U6714 ( .A(n5229), .ZN(n5227) );
  INV_X1 U6715 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6307) );
  OR2_X1 U6716 ( .A1(n5217), .A2(n6307), .ZN(n5225) );
  OR2_X1 U6717 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  NAND2_X1 U6718 ( .A1(n5221), .A2(n5220), .ZN(n6305) );
  NAND2_X1 U6719 ( .A1(n5229), .A2(n9923), .ZN(n7612) );
  NAND2_X1 U6720 ( .A1(n6921), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5234) );
  INV_X1 U6721 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6224) );
  OR2_X1 U6722 ( .A1(n5199), .A2(n6224), .ZN(n5233) );
  INV_X1 U6723 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6225) );
  OR2_X1 U6724 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  NAND2_X1 U6725 ( .A1(n5238), .A2(n5237), .ZN(n6308) );
  OR2_X1 U6726 ( .A1(n5222), .A2(n6308), .ZN(n5243) );
  OR2_X1 U6727 ( .A1(n5239), .A2(n5073), .ZN(n5241) );
  OR2_X1 U6728 ( .A1(n5189), .A2(n6481), .ZN(n5242) );
  NAND2_X1 U6729 ( .A1(n6767), .A2(n5247), .ZN(n5248) );
  NAND2_X1 U6730 ( .A1(n5248), .A2(n5041), .ZN(n5262) );
  NAND2_X1 U6731 ( .A1(n6921), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5253) );
  INV_X1 U6732 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7052) );
  OR2_X1 U6733 ( .A1(n4418), .A2(n7052), .ZN(n5252) );
  NAND2_X1 U6734 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5249) );
  AND2_X1 U6735 ( .A1(n5264), .A2(n5249), .ZN(n7053) );
  OR2_X1 U6736 ( .A1(n5210), .A2(n7053), .ZN(n5251) );
  INV_X1 U6737 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6248) );
  OR2_X1 U6738 ( .A1(n5199), .A2(n6248), .ZN(n5250) );
  OR2_X1 U6739 ( .A1(n5254), .A2(n5073), .ZN(n5255) );
  INV_X1 U6740 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6310) );
  OR2_X1 U6741 ( .A1(n7538), .A2(n6310), .ZN(n5261) );
  OR2_X1 U6742 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6743 ( .A1(n5259), .A2(n5258), .ZN(n6309) );
  OR2_X1 U6744 ( .A1(n5222), .A2(n6309), .ZN(n5260) );
  OAI211_X1 U6745 ( .C1(n5189), .C2(n6708), .A(n5261), .B(n5260), .ZN(n8011)
         );
  NAND2_X1 U6746 ( .A1(n6921), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5270) );
  INV_X1 U6747 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5263) );
  OR2_X1 U6748 ( .A1(n5199), .A2(n5263), .ZN(n5269) );
  NAND2_X1 U6749 ( .A1(n5264), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6750 ( .A1(n5281), .A2(n5265), .ZN(n7981) );
  INV_X1 U6751 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6752 ( .A1(n4417), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U6753 ( .A1(n5271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  INV_X1 U6754 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5272) );
  INV_X1 U6755 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6304) );
  OR2_X1 U6756 ( .A1(n7538), .A2(n6304), .ZN(n5279) );
  OR2_X1 U6757 ( .A1(n5275), .A2(n5274), .ZN(n5276) );
  NAND2_X1 U6758 ( .A1(n5277), .A2(n5276), .ZN(n6303) );
  OR2_X1 U6759 ( .A1(n5222), .A2(n6303), .ZN(n5278) );
  OAI211_X1 U6760 ( .C1(n5189), .C2(n6840), .A(n5279), .B(n5278), .ZN(n7980)
         );
  NAND2_X1 U6761 ( .A1(n6922), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5287) );
  INV_X1 U6762 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6763 ( .A1(n5281), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5282) );
  AND2_X1 U6764 ( .A1(n5301), .A2(n5282), .ZN(n7145) );
  OR2_X1 U6765 ( .A1(n5210), .A2(n7145), .ZN(n5285) );
  INV_X1 U6766 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5283) );
  OR2_X1 U6767 ( .A1(n4417), .A2(n5283), .ZN(n5284) );
  OR2_X1 U6768 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6769 ( .A1(n5291), .A2(n5290), .ZN(n6302) );
  OR2_X1 U6770 ( .A1(n5222), .A2(n6302), .ZN(n5297) );
  OR2_X1 U6771 ( .A1(n7538), .A2(n4509), .ZN(n5296) );
  NAND2_X1 U6772 ( .A1(n5292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6773 ( .A(n5294), .B(n5293), .ZN(n7003) );
  OR2_X1 U6774 ( .A1(n5189), .A2(n7003), .ZN(n5295) );
  NAND2_X1 U6775 ( .A1(n7198), .A2(n9942), .ZN(n5299) );
  INV_X1 U6776 ( .A(n9942), .ZN(n6916) );
  NAND2_X1 U6777 ( .A1(n6922), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5307) );
  INV_X1 U6778 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6779 ( .A1(n5301), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5302) );
  AND2_X1 U6780 ( .A1(n5317), .A2(n5302), .ZN(n7869) );
  INV_X1 U6781 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5303) );
  OR2_X1 U6782 ( .A1(n4418), .A2(n5303), .ZN(n5304) );
  OR2_X1 U6783 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U6784 ( .A1(n5311), .A2(n5310), .ZN(n6312) );
  OR2_X1 U6785 ( .A1(n5222), .A2(n6312), .ZN(n5315) );
  INV_X1 U6786 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6311) );
  OR2_X1 U6787 ( .A1(n7538), .A2(n6311), .ZN(n5314) );
  OR2_X1 U6788 ( .A1(n5312), .A2(n5073), .ZN(n5335) );
  XNOR2_X1 U6789 ( .A(n5335), .B(n5325), .ZN(n7006) );
  OR2_X1 U6790 ( .A1(n5189), .A2(n7006), .ZN(n5313) );
  NAND2_X1 U6791 ( .A1(n8082), .A2(n9946), .ZN(n7211) );
  NAND2_X1 U6792 ( .A1(n6922), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5322) );
  INV_X1 U6793 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6794 ( .A1(n5317), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5318) );
  AND2_X1 U6795 ( .A1(n5343), .A2(n5318), .ZN(n7220) );
  OR2_X1 U6796 ( .A1(n5210), .A2(n7220), .ZN(n5320) );
  INV_X1 U6797 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7101) );
  XNOR2_X1 U6798 ( .A(n5324), .B(n5323), .ZN(n6314) );
  NAND2_X1 U6799 ( .A1(n6314), .A2(n7537), .ZN(n5329) );
  NAND2_X1 U6800 ( .A1(n5335), .A2(n5325), .ZN(n5326) );
  NAND2_X1 U6801 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5327) );
  XNOR2_X1 U6802 ( .A(n5327), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7106) );
  AOI22_X1 U6803 ( .A1(n5488), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5487), .B2(
        n7106), .ZN(n5328) );
  NAND2_X1 U6804 ( .A1(n8081), .A2(n9951), .ZN(n7637) );
  INV_X1 U6805 ( .A(n9946), .ZN(n7868) );
  NAND2_X1 U6806 ( .A1(n8081), .A2(n5330), .ZN(n5331) );
  XNOR2_X1 U6807 ( .A(n5333), .B(n5332), .ZN(n6324) );
  NAND2_X1 U6808 ( .A1(n6324), .A2(n7537), .ZN(n5341) );
  OAI21_X1 U6809 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5334) );
  AND2_X1 U6810 ( .A1(n5335), .A2(n5334), .ZN(n5338) );
  INV_X1 U6811 ( .A(n5338), .ZN(n5336) );
  NAND2_X1 U6812 ( .A1(n5336), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6813 ( .A1(n5338), .A2(n5337), .ZN(n5356) );
  AND2_X1 U6814 ( .A1(n5339), .A2(n5356), .ZN(n7113) );
  AOI22_X1 U6815 ( .A1(n5488), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5487), .B2(
        n7113), .ZN(n5340) );
  NAND2_X1 U6816 ( .A1(n6921), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5349) );
  INV_X1 U6817 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6818 ( .A1(n5199), .A2(n5342), .ZN(n5348) );
  NAND2_X1 U6819 ( .A1(n5343), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5344) );
  AND2_X1 U6820 ( .A1(n5362), .A2(n5344), .ZN(n7339) );
  INV_X1 U6821 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6822 ( .A1(n4417), .A2(n5345), .ZN(n5346) );
  NOR2_X1 U6823 ( .A1(n9955), .A2(n7427), .ZN(n5350) );
  INV_X1 U6824 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6825 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U6826 ( .A1(n5355), .A2(n5354), .ZN(n6334) );
  OR2_X1 U6827 ( .A1(n6334), .A2(n5222), .ZN(n5360) );
  NAND2_X1 U6828 ( .A1(n5356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6829 ( .A(n5358), .B(n5357), .ZN(n7380) );
  INV_X1 U6830 ( .A(n7380), .ZN(n7254) );
  AOI22_X1 U6831 ( .A1(n5488), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5487), .B2(
        n7254), .ZN(n5359) );
  NAND2_X1 U6832 ( .A1(n6921), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5368) );
  INV_X1 U6833 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6834 ( .A1(n5199), .A2(n5361), .ZN(n5367) );
  NAND2_X1 U6835 ( .A1(n5362), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5363) );
  AND2_X1 U6836 ( .A1(n5378), .A2(n5363), .ZN(n7363) );
  OR2_X1 U6837 ( .A1(n5210), .A2(n7363), .ZN(n5366) );
  INV_X1 U6838 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5364) );
  OR2_X1 U6839 ( .A1(n4417), .A2(n5364), .ZN(n5365) );
  NOR2_X1 U6840 ( .A1(n7362), .A2(n8080), .ZN(n5369) );
  NAND2_X1 U6841 ( .A1(n6350), .A2(n7537), .ZN(n5377) );
  NOR2_X1 U6842 ( .A1(n5372), .A2(n5073), .ZN(n5373) );
  MUX2_X1 U6843 ( .A(n5073), .B(n5373), .S(P2_IR_REG_11__SCAN_IN), .Z(n5375)
         );
  INV_X1 U6844 ( .A(n5392), .ZN(n5374) );
  OR2_X1 U6845 ( .A1(n5375), .A2(n5374), .ZN(n7476) );
  INV_X1 U6846 ( .A(n7476), .ZN(n7468) );
  AOI22_X1 U6847 ( .A1(n5488), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5487), .B2(
        n7468), .ZN(n5376) );
  NAND2_X1 U6848 ( .A1(n6921), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5385) );
  INV_X1 U6849 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8443) );
  OR2_X1 U6850 ( .A1(n4418), .A2(n8443), .ZN(n5384) );
  NAND2_X1 U6851 ( .A1(n5378), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5379) );
  AND2_X1 U6852 ( .A1(n5380), .A2(n5379), .ZN(n8442) );
  INV_X1 U6853 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5381) );
  OR2_X1 U6854 ( .A1(n5199), .A2(n5381), .ZN(n5382) );
  NAND2_X1 U6855 ( .A1(n9971), .A2(n8429), .ZN(n7666) );
  NAND2_X2 U6856 ( .A1(n7665), .A2(n7666), .ZN(n8438) );
  OAI21_X1 U6857 ( .B1(n8441), .B2(n7670), .A(n8427), .ZN(n5387) );
  NAND2_X1 U6858 ( .A1(n5387), .A2(n5386), .ZN(n8407) );
  OR2_X1 U6859 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  NAND2_X1 U6860 ( .A1(n5391), .A2(n5390), .ZN(n6456) );
  OR2_X1 U6861 ( .A1(n6456), .A2(n5222), .ZN(n5395) );
  OR2_X1 U6862 ( .A1(n5392), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6863 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U6864 ( .A(n5407), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8097) );
  AOI22_X1 U6865 ( .A1(n5488), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5487), .B2(
        n8097), .ZN(n5394) );
  NAND2_X1 U6866 ( .A1(n6921), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5402) );
  INV_X1 U6867 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6868 ( .A1(n4418), .A2(n5396), .ZN(n5401) );
  NAND2_X1 U6869 ( .A1(n5397), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5398) );
  AND2_X1 U6870 ( .A1(n5411), .A2(n5398), .ZN(n8406) );
  OR2_X1 U6871 ( .A1(n5210), .A2(n8406), .ZN(n5400) );
  INV_X1 U6872 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8503) );
  OR2_X1 U6873 ( .A1(n5199), .A2(n8503), .ZN(n5399) );
  NAND2_X1 U6874 ( .A1(n8593), .A2(n8395), .ZN(n7677) );
  XNOR2_X1 U6875 ( .A(n5403), .B(SI_14_), .ZN(n5404) );
  XNOR2_X1 U6876 ( .A(n5405), .B(n5404), .ZN(n6461) );
  NAND2_X1 U6877 ( .A1(n6461), .A2(n7537), .ZN(n5410) );
  INV_X1 U6878 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6879 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  NAND2_X1 U6880 ( .A1(n5408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5423) );
  INV_X1 U6881 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5422) );
  XNOR2_X1 U6882 ( .A(n5423), .B(n5422), .ZN(n8111) );
  INV_X1 U6883 ( .A(n8111), .ZN(n7506) );
  AOI22_X1 U6884 ( .A1(n5488), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5487), .B2(
        n7506), .ZN(n5409) );
  NAND2_X1 U6885 ( .A1(n6921), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5417) );
  INV_X1 U6886 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8500) );
  OR2_X1 U6887 ( .A1(n5199), .A2(n8500), .ZN(n5416) );
  NAND2_X1 U6888 ( .A1(n5411), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5412) );
  AND2_X1 U6889 ( .A1(n5428), .A2(n5412), .ZN(n8398) );
  OR2_X1 U6890 ( .A1(n5210), .A2(n8398), .ZN(n5415) );
  INV_X1 U6891 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6892 ( .A1(n4417), .A2(n5413), .ZN(n5414) );
  NOR2_X1 U6893 ( .A1(n8399), .A2(n7877), .ZN(n5418) );
  XNOR2_X1 U6894 ( .A(n5419), .B(SI_15_), .ZN(n5420) );
  XNOR2_X1 U6895 ( .A(n5421), .B(n5420), .ZN(n6545) );
  NAND2_X1 U6896 ( .A1(n6545), .A2(n7537), .ZN(n5427) );
  NAND2_X1 U6897 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6898 ( .A1(n5424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6899 ( .A(n5425), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8138) );
  AOI22_X1 U6900 ( .A1(n5488), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5487), .B2(
        n8138), .ZN(n5426) );
  NAND2_X1 U6901 ( .A1(n5211), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5434) );
  INV_X1 U6902 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10199) );
  OR2_X1 U6903 ( .A1(n5199), .A2(n10199), .ZN(n5433) );
  INV_X1 U6904 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10096) );
  OR2_X1 U6905 ( .A1(n5208), .A2(n10096), .ZN(n5432) );
  NAND2_X1 U6906 ( .A1(n5428), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5429) );
  AND2_X1 U6907 ( .A1(n5430), .A2(n5429), .ZN(n8060) );
  OR2_X1 U6908 ( .A1(n5210), .A2(n8060), .ZN(n5431) );
  NAND2_X1 U6909 ( .A1(n8581), .A2(n8396), .ZN(n7557) );
  NAND2_X1 U6910 ( .A1(n7687), .A2(n7689), .ZN(n8371) );
  NAND2_X1 U6911 ( .A1(n8374), .A2(n8371), .ZN(n5435) );
  OAI21_X1 U6912 ( .B1(n8064), .B2(n5436), .A(n5435), .ZN(n8362) );
  INV_X1 U6913 ( .A(n5437), .ZN(n5438) );
  NOR2_X1 U6914 ( .A1(n5438), .A2(SI_16_), .ZN(n5440) );
  NAND2_X1 U6915 ( .A1(n5438), .A2(SI_16_), .ZN(n5439) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6673) );
  INV_X1 U6917 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6671) );
  MUX2_X1 U6918 ( .A(n6673), .B(n6671), .S(n5133), .Z(n5443) );
  INV_X1 U6919 ( .A(SI_17_), .ZN(n5442) );
  NAND2_X1 U6920 ( .A1(n5443), .A2(n5442), .ZN(n5459) );
  INV_X1 U6921 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6922 ( .A1(n5444), .A2(SI_17_), .ZN(n5445) );
  NAND2_X1 U6923 ( .A1(n5459), .A2(n5445), .ZN(n5460) );
  XNOR2_X1 U6924 ( .A(n5461), .B(n5460), .ZN(n6670) );
  NAND2_X1 U6925 ( .A1(n6670), .A2(n7537), .ZN(n5448) );
  NAND2_X1 U6926 ( .A1(n5163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6927 ( .A(n5446), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8191) );
  AOI22_X1 U6928 ( .A1(n5488), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5487), .B2(
        n8191), .ZN(n5447) );
  NAND2_X1 U6929 ( .A1(n6921), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5456) );
  INV_X1 U6930 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8492) );
  OR2_X1 U6931 ( .A1(n5199), .A2(n8492), .ZN(n5455) );
  INV_X1 U6932 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6933 ( .A1(n5451), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5452) );
  AND2_X1 U6934 ( .A1(n5469), .A2(n5452), .ZN(n8366) );
  OR2_X1 U6935 ( .A1(n5210), .A2(n8366), .ZN(n5454) );
  INV_X1 U6936 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8365) );
  OR2_X1 U6937 ( .A1(n4418), .A2(n8365), .ZN(n5453) );
  NAND2_X1 U6938 ( .A1(n8570), .A2(n8346), .ZN(n7700) );
  NAND2_X1 U6939 ( .A1(n8362), .A2(n8359), .ZN(n5458) );
  INV_X1 U6940 ( .A(n8570), .ZN(n5457) );
  NAND2_X1 U6941 ( .A1(n5458), .A2(n5048), .ZN(n8344) );
  INV_X1 U6942 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10128) );
  INV_X1 U6943 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5462) );
  MUX2_X1 U6944 ( .A(n10128), .B(n5462), .S(n5133), .Z(n5478) );
  XNOR2_X1 U6945 ( .A(n5478), .B(SI_18_), .ZN(n5477) );
  XNOR2_X1 U6946 ( .A(n5480), .B(n5477), .ZN(n6801) );
  NAND2_X1 U6947 ( .A1(n6801), .A2(n7537), .ZN(n5468) );
  NAND2_X1 U6948 ( .A1(n5463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5465) );
  INV_X1 U6949 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6950 ( .A1(n5465), .A2(n5464), .ZN(n5485) );
  OR2_X1 U6951 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  AND2_X1 U6952 ( .A1(n5485), .A2(n5466), .ZN(n8207) );
  AOI22_X1 U6953 ( .A1(n5488), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5487), .B2(
        n8207), .ZN(n5467) );
  NAND2_X1 U6954 ( .A1(n6922), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5474) );
  INV_X1 U6955 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8564) );
  OR2_X1 U6956 ( .A1(n5208), .A2(n8564), .ZN(n5473) );
  NAND2_X1 U6957 ( .A1(n5469), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5470) );
  AND2_X1 U6958 ( .A1(n5493), .A2(n5470), .ZN(n8353) );
  OR2_X1 U6959 ( .A1(n5210), .A2(n8353), .ZN(n5472) );
  INV_X1 U6960 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8354) );
  OR2_X1 U6961 ( .A1(n4418), .A2(n8354), .ZN(n5471) );
  NOR2_X1 U6962 ( .A1(n8567), .A2(n8335), .ZN(n5475) );
  INV_X1 U6963 ( .A(n5478), .ZN(n5479) );
  INV_X1 U6964 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6929) );
  INV_X1 U6965 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7517) );
  MUX2_X1 U6966 ( .A(n6929), .B(n7517), .S(n5133), .Z(n5482) );
  INV_X1 U6967 ( .A(SI_19_), .ZN(n5481) );
  NAND2_X1 U6968 ( .A1(n5482), .A2(n5481), .ZN(n5499) );
  INV_X1 U6969 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U6970 ( .A1(n5483), .A2(SI_19_), .ZN(n5484) );
  NAND2_X1 U6971 ( .A1(n5499), .A2(n5484), .ZN(n5500) );
  XNOR2_X1 U6972 ( .A(n5501), .B(n5500), .ZN(n6928) );
  NAND2_X1 U6973 ( .A1(n6928), .A2(n7537), .ZN(n5490) );
  NAND2_X1 U6974 ( .A1(n5485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5486) );
  AOI22_X1 U6975 ( .A1(n5488), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8212), .B2(
        n5487), .ZN(n5489) );
  NAND2_X1 U6976 ( .A1(n6921), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5498) );
  INV_X1 U6977 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8484) );
  OR2_X1 U6978 ( .A1(n5199), .A2(n8484), .ZN(n5497) );
  INV_X1 U6979 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6980 ( .A1(n5493), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5494) );
  AND2_X1 U6981 ( .A1(n5505), .A2(n5494), .ZN(n7935) );
  OR2_X1 U6982 ( .A1(n5210), .A2(n7935), .ZN(n5496) );
  INV_X1 U6983 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8339) );
  OR2_X1 U6984 ( .A1(n4417), .A2(n8339), .ZN(n5495) );
  INV_X1 U6985 ( .A(n8559), .ZN(n7940) );
  MUX2_X1 U6986 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5133), .Z(n5513) );
  INV_X1 U6987 ( .A(SI_20_), .ZN(n10235) );
  XNOR2_X1 U6988 ( .A(n5513), .B(n10235), .ZN(n5502) );
  XNOR2_X1 U6989 ( .A(n5515), .B(n5502), .ZN(n7069) );
  NAND2_X1 U6990 ( .A1(n7069), .A2(n7537), .ZN(n5504) );
  INV_X1 U6991 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7092) );
  OR2_X1 U6992 ( .A1(n7538), .A2(n7092), .ZN(n5503) );
  NAND2_X1 U6993 ( .A1(n5505), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U6994 ( .A1(n5525), .A2(n5506), .ZN(n8324) );
  NAND2_X1 U6995 ( .A1(n5665), .A2(n8324), .ZN(n5511) );
  INV_X1 U6996 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8554) );
  OR2_X1 U6997 ( .A1(n5208), .A2(n8554), .ZN(n5510) );
  INV_X1 U6998 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8482) );
  OR2_X1 U6999 ( .A1(n5199), .A2(n8482), .ZN(n5509) );
  INV_X1 U7000 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5507) );
  OR2_X1 U7001 ( .A1(n4418), .A2(n5507), .ZN(n5508) );
  INV_X1 U7002 ( .A(n5513), .ZN(n5514) );
  INV_X1 U7003 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7150) );
  INV_X1 U7004 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10284) );
  MUX2_X1 U7005 ( .A(n7150), .B(n10284), .S(n5133), .Z(n5531) );
  XNOR2_X1 U7006 ( .A(n5531), .B(SI_21_), .ZN(n5518) );
  XNOR2_X1 U7007 ( .A(n5535), .B(n5518), .ZN(n7149) );
  NAND2_X1 U7008 ( .A1(n7149), .A2(n7537), .ZN(n5520) );
  OR2_X1 U7009 ( .A1(n7538), .A2(n7150), .ZN(n5519) );
  INV_X1 U7010 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8550) );
  OR2_X1 U7011 ( .A1(n5208), .A2(n8550), .ZN(n5522) );
  INV_X1 U7012 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10226) );
  OR2_X1 U7013 ( .A1(n5199), .A2(n10226), .ZN(n5521) );
  AND2_X1 U7014 ( .A1(n5522), .A2(n5521), .ZN(n5529) );
  INV_X1 U7015 ( .A(n5525), .ZN(n5524) );
  INV_X1 U7016 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7017 ( .A1(n5525), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7018 ( .A1(n5542), .A2(n5526), .ZN(n8313) );
  NAND2_X1 U7019 ( .A1(n8313), .A2(n5665), .ZN(n5528) );
  NAND2_X1 U7020 ( .A1(n5211), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7021 ( .A1(n5530), .A2(n8320), .ZN(n7586) );
  NAND2_X1 U7022 ( .A1(n7590), .A2(n7586), .ZN(n7543) );
  INV_X1 U7023 ( .A(n5531), .ZN(n5532) );
  NOR2_X1 U7024 ( .A1(n5532), .A2(SI_21_), .ZN(n5534) );
  NAND2_X1 U7025 ( .A1(n5532), .A2(SI_21_), .ZN(n5533) );
  INV_X1 U7026 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7306) );
  INV_X1 U7027 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7309) );
  MUX2_X1 U7028 ( .A(n7306), .B(n7309), .S(n5133), .Z(n5537) );
  INV_X1 U7029 ( .A(SI_22_), .ZN(n5536) );
  NAND2_X1 U7030 ( .A1(n5537), .A2(n5536), .ZN(n5548) );
  INV_X1 U7031 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U7032 ( .A1(n5538), .A2(SI_22_), .ZN(n5539) );
  NAND2_X1 U7033 ( .A1(n5548), .A2(n5539), .ZN(n5549) );
  OR2_X1 U7034 ( .A1(n7538), .A2(n7306), .ZN(n5540) );
  NAND2_X1 U7035 ( .A1(n5542), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7036 ( .A1(n5556), .A2(n5543), .ZN(n8301) );
  NAND2_X1 U7037 ( .A1(n8301), .A2(n5665), .ZN(n5546) );
  AOI22_X1 U7038 ( .A1(n6922), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6921), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7039 ( .A1(n5211), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5544) );
  OAI21_X1 U7040 ( .B1(n5550), .B2(n5549), .A(n5548), .ZN(n5565) );
  INV_X1 U7041 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7330) );
  INV_X1 U7042 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7326) );
  MUX2_X1 U7043 ( .A(n7330), .B(n7326), .S(n5133), .Z(n5551) );
  INV_X1 U7044 ( .A(SI_23_), .ZN(n10258) );
  NAND2_X1 U7045 ( .A1(n5551), .A2(n10258), .ZN(n5566) );
  INV_X1 U7046 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U7047 ( .A1(n5552), .A2(SI_23_), .ZN(n5553) );
  AND2_X1 U7048 ( .A1(n5566), .A2(n5553), .ZN(n5564) );
  XNOR2_X1 U7049 ( .A(n5565), .B(n5564), .ZN(n7327) );
  NAND2_X1 U7050 ( .A1(n7327), .A2(n7537), .ZN(n5555) );
  OR2_X1 U7051 ( .A1(n7538), .A2(n7330), .ZN(n5554) );
  NAND2_X1 U7052 ( .A1(n5556), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7053 ( .A1(n5575), .A2(n5557), .ZN(n8288) );
  NAND2_X1 U7054 ( .A1(n8288), .A2(n5665), .ZN(n5560) );
  AOI22_X1 U7055 ( .A1(n6922), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6921), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7056 ( .A1(n5211), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7057 ( .A1(n8290), .A2(n8298), .ZN(n5561) );
  NAND2_X1 U7058 ( .A1(n8282), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U7059 ( .A1(n8469), .A2(n8075), .ZN(n5562) );
  INV_X1 U7060 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7423) );
  INV_X1 U7061 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U7062 ( .A(n7423), .B(n10079), .S(n5133), .Z(n5568) );
  INV_X1 U7063 ( .A(SI_24_), .ZN(n10283) );
  NAND2_X1 U7064 ( .A1(n5568), .A2(n10283), .ZN(n5586) );
  INV_X1 U7065 ( .A(n5568), .ZN(n5569) );
  NAND2_X1 U7066 ( .A1(n5569), .A2(SI_24_), .ZN(n5570) );
  AND2_X1 U7067 ( .A1(n5586), .A2(n5570), .ZN(n5584) );
  OR2_X1 U7068 ( .A1(n7538), .A2(n7423), .ZN(n5571) );
  INV_X1 U7069 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7070 ( .A1(n5575), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7071 ( .A1(n5596), .A2(n5576), .ZN(n8275) );
  NAND2_X1 U7072 ( .A1(n8275), .A2(n5665), .ZN(n5581) );
  INV_X1 U7073 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U7074 ( .A1(n6922), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7075 ( .A1(n5211), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U7076 ( .C1(n5208), .C2(n10125), .A(n5578), .B(n5577), .ZN(n5579)
         );
  INV_X1 U7077 ( .A(n5579), .ZN(n5580) );
  INV_X1 U7078 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7447) );
  INV_X1 U7079 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7449) );
  MUX2_X1 U7080 ( .A(n7447), .B(n7449), .S(n5133), .Z(n5589) );
  INV_X1 U7081 ( .A(SI_25_), .ZN(n5588) );
  NAND2_X1 U7082 ( .A1(n5589), .A2(n5588), .ZN(n5607) );
  INV_X1 U7083 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7084 ( .A1(n5590), .A2(SI_25_), .ZN(n5591) );
  AND2_X1 U7085 ( .A1(n5607), .A2(n5591), .ZN(n5605) );
  OR2_X1 U7086 ( .A1(n7538), .A2(n7447), .ZN(n5592) );
  INV_X1 U7087 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7088 ( .A1(n5596), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7089 ( .A1(n5615), .A2(n5597), .ZN(n8265) );
  NAND2_X1 U7090 ( .A1(n8265), .A2(n5665), .ZN(n5603) );
  INV_X1 U7091 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7092 ( .A1(n6922), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7093 ( .A1(n6921), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U7094 ( .C1(n5600), .C2(n4417), .A(n5599), .B(n5598), .ZN(n5601)
         );
  INV_X1 U7095 ( .A(n5601), .ZN(n5602) );
  INV_X1 U7096 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7453) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7455) );
  MUX2_X1 U7098 ( .A(n7453), .B(n7455), .S(n5133), .Z(n5610) );
  INV_X1 U7099 ( .A(SI_26_), .ZN(n5609) );
  NAND2_X1 U7100 ( .A1(n5610), .A2(n5609), .ZN(n5626) );
  INV_X1 U7101 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7102 ( .A1(n5611), .A2(SI_26_), .ZN(n5612) );
  AND2_X1 U7103 ( .A1(n5626), .A2(n5612), .ZN(n5624) );
  NAND2_X1 U7104 ( .A1(n7452), .A2(n7537), .ZN(n5614) );
  OR2_X1 U7105 ( .A1(n7538), .A2(n7453), .ZN(n5613) );
  NAND2_X1 U7106 ( .A1(n5615), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7107 ( .A1(n5636), .A2(n5616), .ZN(n8259) );
  NAND2_X1 U7108 ( .A1(n8259), .A2(n5665), .ZN(n5621) );
  INV_X1 U7109 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U7110 ( .A1(n6922), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7111 ( .A1(n6921), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U7112 ( .C1(n8258), .C2(n4418), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U7113 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7114 ( .A1(n8054), .A2(n8264), .ZN(n5623) );
  INV_X1 U7115 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5631) );
  INV_X1 U7116 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7764) );
  MUX2_X1 U7117 ( .A(n5631), .B(n7764), .S(n5133), .Z(n5628) );
  INV_X1 U7118 ( .A(SI_27_), .ZN(n10090) );
  NAND2_X1 U7119 ( .A1(n5628), .A2(n10090), .ZN(n5646) );
  INV_X1 U7120 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7121 ( .A1(n5629), .A2(SI_27_), .ZN(n5630) );
  AND2_X1 U7122 ( .A1(n5646), .A2(n5630), .ZN(n5644) );
  NAND2_X1 U7123 ( .A1(n7458), .A2(n7537), .ZN(n5633) );
  OR2_X1 U7124 ( .A1(n7538), .A2(n5631), .ZN(n5632) );
  INV_X1 U7125 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7126 ( .A1(n5636), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7127 ( .A1(n5649), .A2(n5637), .ZN(n8244) );
  NAND2_X1 U7128 ( .A1(n8244), .A2(n5665), .ZN(n5643) );
  INV_X1 U7129 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7130 ( .A1(n6922), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7131 ( .A1(n6921), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5638) );
  OAI211_X1 U7132 ( .C1(n5640), .C2(n4417), .A(n5639), .B(n5638), .ZN(n5641)
         );
  INV_X1 U7133 ( .A(n5641), .ZN(n5642) );
  NAND2_X2 U7134 ( .A1(n5643), .A2(n5642), .ZN(n8256) );
  INV_X1 U7135 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8611) );
  INV_X1 U7136 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9708) );
  MUX2_X1 U7137 ( .A(n8611), .B(n9708), .S(n5133), .Z(n5661) );
  XNOR2_X1 U7138 ( .A(n5661), .B(SI_28_), .ZN(n5658) );
  NAND2_X1 U7139 ( .A1(n9704), .A2(n7537), .ZN(n5648) );
  OR2_X1 U7140 ( .A1(n7538), .A2(n8611), .ZN(n5647) );
  NAND2_X1 U7141 ( .A1(n5649), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7142 ( .A1(n5664), .A2(n5650), .ZN(n8241) );
  NAND2_X1 U7143 ( .A1(n8241), .A2(n5665), .ZN(n5655) );
  INV_X1 U7144 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U7145 ( .A1(n6922), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7146 ( .A1(n5211), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5651) );
  OAI211_X1 U7147 ( .C1(n5208), .C2(n10129), .A(n5652), .B(n5651), .ZN(n5653)
         );
  INV_X1 U7148 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7149 ( .A1(n5657), .A2(n5656), .ZN(n5670) );
  INV_X1 U7150 ( .A(SI_28_), .ZN(n5660) );
  INV_X1 U7151 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10078) );
  INV_X1 U7152 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9703) );
  MUX2_X1 U7153 ( .A(n10078), .B(n9703), .S(n5133), .Z(n7520) );
  NAND2_X1 U7154 ( .A1(n7518), .A2(n7537), .ZN(n5663) );
  OR2_X1 U7155 ( .A1(n7538), .A2(n10078), .ZN(n5662) );
  NAND2_X1 U7156 ( .A1(n7853), .A2(n5665), .ZN(n6924) );
  INV_X1 U7157 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U7158 ( .A1(n6921), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7159 ( .A1(n6922), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5666) );
  OAI211_X1 U7160 ( .C1(n4418), .C2(n10212), .A(n5667), .B(n5666), .ZN(n5668)
         );
  INV_X1 U7161 ( .A(n5668), .ZN(n5669) );
  NAND2_X1 U7162 ( .A1(n5750), .A2(n8237), .ZN(n7571) );
  XNOR2_X1 U7163 ( .A(n5670), .B(n4712), .ZN(n5689) );
  NAND2_X1 U7164 ( .A1(n5671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U7165 ( .A(n5672), .B(n5002), .ZN(n7597) );
  INV_X1 U7166 ( .A(n7597), .ZN(n7753) );
  NAND2_X1 U7167 ( .A1(n7753), .A2(n8212), .ZN(n5679) );
  NAND2_X1 U7168 ( .A1(n4463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  XNOR2_X1 U7169 ( .A(n5674), .B(n5673), .ZN(n7151) );
  INV_X1 U7170 ( .A(n7151), .ZN(n7598) );
  NAND2_X1 U7171 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  INV_X1 U7172 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U7173 ( .A(n5677), .B(n5676), .ZN(n7093) );
  INV_X1 U7174 ( .A(n7093), .ZN(n7748) );
  NAND2_X1 U7175 ( .A1(n7598), .A2(n7748), .ZN(n5678) );
  NAND2_X1 U7176 ( .A1(n5679), .A2(n5678), .ZN(n8413) );
  INV_X1 U7177 ( .A(n5680), .ZN(n7750) );
  INV_X1 U7178 ( .A(n5681), .ZN(n6226) );
  NAND2_X1 U7179 ( .A1(n7750), .A2(n6226), .ZN(n5682) );
  NAND2_X1 U7180 ( .A1(n5189), .A2(n5682), .ZN(n6652) );
  INV_X1 U7181 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U7182 ( .A1(n5211), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7183 ( .A1(n6921), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7184 ( .C1(n5199), .C2(n10076), .A(n5684), .B(n5683), .ZN(n5685)
         );
  INV_X1 U7185 ( .A(n5685), .ZN(n5686) );
  AND2_X1 U7186 ( .A1(n6924), .A2(n5686), .ZN(n7570) );
  NAND2_X1 U7187 ( .A1(n6652), .A2(n7738), .ZN(n9909) );
  AND2_X1 U7188 ( .A1(n5189), .A2(P2_B_REG_SCAN_IN), .ZN(n5687) );
  OR2_X1 U7189 ( .A1(n9909), .A2(n5687), .ZN(n8226) );
  OAI22_X1 U7190 ( .A1(n7916), .A2(n9910), .B1(n7570), .B2(n8226), .ZN(n5688)
         );
  INV_X1 U7191 ( .A(n7758), .ZN(n6580) );
  OR2_X1 U7192 ( .A1(n6987), .A2(n6580), .ZN(n6629) );
  INV_X1 U7193 ( .A(n6629), .ZN(n5691) );
  NAND2_X1 U7194 ( .A1(n7547), .A2(n5691), .ZN(n6982) );
  INV_X1 U7195 ( .A(n9901), .ZN(n9897) );
  NAND2_X1 U7196 ( .A1(n9896), .A2(n7611), .ZN(n5693) );
  NAND2_X1 U7197 ( .A1(n5246), .A2(n9927), .ZN(n7620) );
  NAND2_X1 U7198 ( .A1(n5693), .A2(n7546), .ZN(n6771) );
  NAND2_X1 U7199 ( .A1(n6771), .A2(n7626), .ZN(n7049) );
  INV_X1 U7200 ( .A(n8011), .ZN(n9934) );
  NAND2_X1 U7201 ( .A1(n8085), .A2(n9934), .ZN(n7627) );
  NAND2_X1 U7202 ( .A1(n7049), .A2(n7627), .ZN(n7016) );
  OR2_X1 U7203 ( .A1(n8085), .A2(n9934), .ZN(n7048) );
  INV_X1 U7204 ( .A(n7980), .ZN(n9938) );
  OR2_X1 U7205 ( .A1(n8084), .A2(n9938), .ZN(n7633) );
  NAND2_X1 U7206 ( .A1(n7016), .A2(n7621), .ZN(n7139) );
  NAND2_X1 U7207 ( .A1(n8083), .A2(n9942), .ZN(n7625) );
  NAND2_X1 U7208 ( .A1(n8084), .A2(n9938), .ZN(n7138) );
  OR2_X1 U7209 ( .A1(n8083), .A2(n9942), .ZN(n7631) );
  AND2_X1 U7210 ( .A1(n7637), .A2(n7211), .ZN(n7644) );
  NAND2_X1 U7211 ( .A1(n7212), .A2(n7644), .ZN(n5695) );
  OR2_X1 U7212 ( .A1(n7427), .A2(n7341), .ZN(n7646) );
  NAND2_X1 U7213 ( .A1(n7427), .A2(n7341), .ZN(n7653) );
  NAND2_X1 U7214 ( .A1(n7646), .A2(n7653), .ZN(n7545) );
  OR2_X1 U7215 ( .A1(n7362), .A2(n8440), .ZN(n7662) );
  NAND2_X1 U7216 ( .A1(n7362), .A2(n8440), .ZN(n7661) );
  NAND2_X1 U7217 ( .A1(n7662), .A2(n7661), .ZN(n7553) );
  INV_X1 U7218 ( .A(n7646), .ZN(n7640) );
  NOR2_X1 U7219 ( .A1(n7553), .A2(n7640), .ZN(n5697) );
  NAND2_X1 U7220 ( .A1(n7429), .A2(n7661), .ZN(n8436) );
  INV_X1 U7221 ( .A(n8438), .ZN(n7555) );
  NAND2_X1 U7222 ( .A1(n8436), .A2(n7555), .ZN(n5698) );
  XNOR2_X1 U7223 ( .A(n8509), .B(n8441), .ZN(n8423) );
  OR2_X1 U7224 ( .A1(n8509), .A2(n8441), .ZN(n7671) );
  NAND2_X1 U7225 ( .A1(n8593), .A2(n8430), .ZN(n5700) );
  NAND2_X1 U7226 ( .A1(n8417), .A2(n5700), .ZN(n5702) );
  OR2_X1 U7227 ( .A1(n8593), .A2(n8430), .ZN(n5701) );
  NAND2_X1 U7228 ( .A1(n8587), .A2(n7877), .ZN(n7682) );
  OR2_X1 U7229 ( .A1(n8587), .A2(n7877), .ZN(n7681) );
  INV_X1 U7230 ( .A(n8396), .ZN(n7971) );
  NAND2_X1 U7231 ( .A1(n8581), .A2(n7971), .ZN(n7595) );
  OR2_X1 U7232 ( .A1(n8581), .A2(n7971), .ZN(n7596) );
  NAND2_X1 U7233 ( .A1(n8372), .A2(n7689), .ZN(n5703) );
  NAND2_X1 U7234 ( .A1(n5703), .A2(n7687), .ZN(n8360) );
  INV_X1 U7235 ( .A(n7690), .ZN(n5704) );
  INV_X1 U7236 ( .A(n8567), .ZN(n8043) );
  NAND2_X1 U7237 ( .A1(n8043), .A2(n8335), .ZN(n7701) );
  NAND2_X1 U7238 ( .A1(n7702), .A2(n7701), .ZN(n8351) );
  INV_X1 U7239 ( .A(n7703), .ZN(n5706) );
  NAND2_X1 U7240 ( .A1(n8322), .A2(n7589), .ZN(n8310) );
  AND2_X1 U7241 ( .A1(n7586), .A2(n8309), .ZN(n7698) );
  NAND2_X1 U7242 ( .A1(n8310), .A2(n7698), .ZN(n5707) );
  NAND2_X1 U7243 ( .A1(n5707), .A2(n7590), .ZN(n8300) );
  NAND2_X1 U7244 ( .A1(n5708), .A2(n8284), .ZN(n7711) );
  NAND2_X1 U7245 ( .A1(n8469), .A2(n8298), .ZN(n7709) );
  OAI21_X2 U7246 ( .B1(n8252), .B2(n7722), .A(n7721), .ZN(n7842) );
  NAND2_X1 U7247 ( .A1(n7875), .A2(n8236), .ZN(n7541) );
  AOI21_X2 U7248 ( .B1(n7842), .B2(n7541), .A(n7727), .ZN(n8233) );
  NOR2_X1 U7249 ( .A1(n7565), .A2(n8072), .ZN(n5709) );
  OAI22_X1 U7250 ( .A1(n8233), .A2(n5709), .B1(n7916), .B2(n8520), .ZN(n7574)
         );
  XNOR2_X1 U7251 ( .A(n7574), .B(n7732), .ZN(n7857) );
  INV_X1 U7252 ( .A(n8212), .ZN(n7584) );
  NAND2_X1 U7253 ( .A1(n7584), .A2(n7093), .ZN(n6626) );
  OR2_X1 U7254 ( .A1(n7739), .A2(n6626), .ZN(n6649) );
  NAND2_X1 U7255 ( .A1(n7597), .A2(n7151), .ZN(n9961) );
  NAND2_X1 U7256 ( .A1(n6649), .A2(n9961), .ZN(n6603) );
  NAND2_X1 U7257 ( .A1(n7753), .A2(n7584), .ZN(n5752) );
  AND2_X1 U7258 ( .A1(n5752), .A2(n6626), .ZN(n5710) );
  OR2_X1 U7259 ( .A1(n6603), .A2(n5710), .ZN(n7165) );
  AND2_X1 U7260 ( .A1(n8212), .A2(n7093), .ZN(n7744) );
  AND2_X1 U7261 ( .A1(n7597), .A2(n7744), .ZN(n9958) );
  INV_X1 U7262 ( .A(n9958), .ZN(n9947) );
  NAND2_X1 U7263 ( .A1(n7165), .A2(n9947), .ZN(n9966) );
  NAND2_X1 U7264 ( .A1(n7857), .A2(n9966), .ZN(n5711) );
  INV_X1 U7265 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7266 ( .A1(n5740), .A2(n5741), .ZN(n5712) );
  INV_X1 U7267 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7268 ( .A1(n5714), .A2(n5713), .ZN(n5716) );
  XNOR2_X1 U7269 ( .A(n7424), .B(P2_B_REG_SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7270 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U7271 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7272 ( .A1(n5719), .A2(n7448), .ZN(n5723) );
  NAND2_X1 U7273 ( .A1(n5720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5721) );
  XNOR2_X1 U7274 ( .A(n5721), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6320) );
  INV_X1 U7275 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6323) );
  AND2_X1 U7276 ( .A1(n6320), .A2(n6323), .ZN(n5722) );
  NAND2_X1 U7277 ( .A1(n5723), .A2(n5722), .ZN(n6625) );
  INV_X1 U7278 ( .A(n6320), .ZN(n7454) );
  NAND2_X1 U7279 ( .A1(n7454), .A2(n7424), .ZN(n6623) );
  NAND2_X1 U7280 ( .A1(n6625), .A2(n6623), .ZN(n6606) );
  NAND2_X1 U7281 ( .A1(n5723), .A2(n6320), .ZN(n6318) );
  OR2_X1 U7282 ( .A1(n6318), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7283 ( .A1(n7448), .A2(n7454), .ZN(n5724) );
  INV_X1 U7284 ( .A(n6610), .ZN(n5726) );
  NOR2_X1 U7285 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .ZN(
        n10045) );
  NOR4_X1 U7286 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5729) );
  NOR4_X1 U7287 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5728) );
  NOR4_X1 U7288 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5727) );
  NAND4_X1 U7289 ( .A1(n10045), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n5735)
         );
  NOR4_X1 U7290 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5733) );
  NOR4_X1 U7291 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U7292 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U7293 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5730) );
  NAND4_X1 U7294 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5734)
         );
  NOR2_X1 U7295 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  OR2_X1 U7296 ( .A1(n6318), .A2(n5736), .ZN(n5755) );
  INV_X1 U7297 ( .A(n5755), .ZN(n5737) );
  NOR2_X1 U7298 ( .A1(n5758), .A2(n5737), .ZN(n6643) );
  INV_X1 U7299 ( .A(n7448), .ZN(n5739) );
  NOR2_X1 U7300 ( .A1(n7454), .A2(n7424), .ZN(n5738) );
  NAND2_X1 U7301 ( .A1(n5739), .A2(n5738), .ZN(n6638) );
  XNOR2_X1 U7302 ( .A(n5740), .B(n5741), .ZN(n6319) );
  AND2_X1 U7303 ( .A1(n6319), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7304 ( .A1(n6638), .A2(n5742), .ZN(n6645) );
  INV_X1 U7305 ( .A(n6645), .ZN(n6328) );
  NAND2_X1 U7306 ( .A1(n6643), .A2(n6328), .ZN(n6656) );
  NAND3_X1 U7307 ( .A1(n7151), .A2(n8212), .A3(n7748), .ZN(n5743) );
  OR2_X1 U7308 ( .A1(n7597), .A2(n5743), .ZN(n6619) );
  AND2_X1 U7309 ( .A1(n6649), .A2(n6619), .ZN(n5744) );
  OR2_X1 U7310 ( .A1(n6656), .A2(n5744), .ZN(n5747) );
  NAND2_X1 U7311 ( .A1(n6606), .A2(n5755), .ZN(n5745) );
  NOR2_X1 U7312 ( .A1(n6646), .A2(n6645), .ZN(n6651) );
  NAND3_X1 U7313 ( .A1(n7739), .A2(n6619), .A3(n9961), .ZN(n6618) );
  OR2_X1 U7314 ( .A1(n9961), .A2(n7744), .ZN(n9899) );
  NAND2_X1 U7315 ( .A1(n6618), .A2(n9899), .ZN(n6635) );
  NAND2_X1 U7316 ( .A1(n6651), .A2(n6635), .ZN(n5746) );
  INV_X2 U7317 ( .A(n9975), .ZN(n9973) );
  OR2_X1 U7318 ( .A1(n5760), .A2(n9975), .ZN(n5749) );
  NAND2_X1 U7319 ( .A1(n5749), .A2(n5748), .ZN(n5751) );
  OR2_X1 U7320 ( .A1(n9975), .A2(n9961), .ZN(n8566) );
  NAND2_X1 U7321 ( .A1(n5751), .A2(n5045), .ZN(P2_U3456) );
  AND2_X1 U7322 ( .A1(n9958), .A2(n7151), .ZN(n6601) );
  NOR2_X1 U7323 ( .A1(n6606), .A2(n6601), .ZN(n5754) );
  OR2_X1 U7324 ( .A1(n5752), .A2(n7093), .ZN(n5753) );
  AND2_X1 U7325 ( .A1(n5753), .A2(n7739), .ZN(n6607) );
  MUX2_X1 U7326 ( .A(n6610), .B(n5754), .S(n6607), .Z(n5759) );
  AND2_X1 U7327 ( .A1(n7738), .A2(n6626), .ZN(n6636) );
  NOR2_X1 U7328 ( .A1(n6645), .A2(n6636), .ZN(n5756) );
  AND2_X1 U7329 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  AND2_X2 U7330 ( .A1(n5759), .A2(n6612), .ZN(n9992) );
  INV_X1 U7331 ( .A(n9961), .ZN(n9972) );
  NAND2_X1 U7332 ( .A1(n9992), .A2(n9972), .ZN(n8491) );
  NAND2_X1 U7333 ( .A1(n5762), .A2(n5052), .ZN(P2_U3488) );
  NAND2_X1 U7334 ( .A1(n5915), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5928) );
  INV_X1 U7335 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5927) );
  INV_X1 U7336 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8727) );
  INV_X1 U7337 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7338 ( .A1(n5971), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5986) );
  INV_X1 U7339 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5985) );
  INV_X1 U7340 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5998) );
  INV_X1 U7341 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6025) );
  INV_X1 U7342 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6037) );
  AND2_X1 U7343 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5763) );
  INV_X1 U7344 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8849) );
  INV_X1 U7345 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6080) );
  INV_X1 U7346 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8823) );
  OR2_X1 U7347 ( .A1(n6093), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7348 ( .A1(n6093), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6107) );
  AND2_X1 U7349 ( .A1(n5764), .A2(n6107), .ZN(n9376) );
  INV_X1 U7350 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6007) );
  INV_X1 U7351 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5766) );
  NOR2_X1 U7352 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5768) );
  NOR2_X1 U7353 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5767) );
  INV_X1 U7354 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10046) );
  INV_X1 U7355 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9695) );
  NAND2_X2 U7356 ( .A1(n5771), .A2(n5772), .ZN(n6070) );
  INV_X1 U7357 ( .A(n6070), .ZN(n6083) );
  NAND2_X1 U7358 ( .A1(n9376), .A2(n6083), .ZN(n5778) );
  AND2_X4 U7359 ( .A1(n7851), .A2(n5772), .ZN(n6340) );
  INV_X1 U7360 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U7361 ( .A1(n6124), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7362 ( .A1(n6095), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5774) );
  OAI211_X1 U7363 ( .C1(n6125), .C2(n9592), .A(n5775), .B(n5774), .ZN(n5776)
         );
  INV_X1 U7364 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7365 ( .A1(n5778), .A2(n5777), .ZN(n9393) );
  INV_X1 U7366 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7367 ( .A1(n9000), .A2(n7449), .ZN(n5781) );
  INV_X1 U7368 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5783) );
  XNOR2_X1 U7369 ( .A(n6049), .B(n5783), .ZN(n9471) );
  NAND2_X1 U7370 ( .A1(n9471), .A2(n6083), .ZN(n5788) );
  INV_X1 U7371 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U7372 ( .A1(n6340), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7373 ( .A1(n6095), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5784) );
  OAI211_X1 U7374 ( .C1(n10236), .C2(n6343), .A(n5785), .B(n5784), .ZN(n5786)
         );
  INV_X1 U7375 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U7376 ( .A1(n5788), .A2(n5787), .ZN(n9453) );
  INV_X1 U7377 ( .A(n9453), .ZN(n9487) );
  NAND2_X1 U7378 ( .A1(n6928), .A2(n8998), .ZN(n5797) );
  INV_X1 U7379 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5790) );
  INV_X1 U7380 ( .A(n6148), .ZN(n5791) );
  NAND2_X1 U7381 ( .A1(n6033), .A2(n5792), .ZN(n5793) );
  XNOR2_X2 U7382 ( .A(n5795), .B(n5794), .ZN(n6153) );
  INV_X1 U7383 ( .A(n6153), .ZN(n9143) );
  AOI22_X1 U7384 ( .A1(n6034), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6329), .B2(
        n9143), .ZN(n5796) );
  NAND2_X1 U7385 ( .A1(n6599), .A2(n8998), .ZN(n5804) );
  INV_X1 U7386 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U7387 ( .A1(n5799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  MUX2_X1 U7388 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5800), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5802) );
  NAND2_X1 U7389 ( .A1(n5802), .A2(n5801), .ZN(n9258) );
  INV_X1 U7390 ( .A(n9258), .ZN(n9270) );
  AOI22_X1 U7391 ( .A1(n6034), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6329), .B2(
        n9270), .ZN(n5803) );
  OR2_X1 U7392 ( .A1(n6015), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5805) );
  AND2_X1 U7393 ( .A1(n6026), .A2(n5805), .ZN(n9515) );
  NAND2_X1 U7394 ( .A1(n6083), .A2(n9515), .ZN(n5810) );
  INV_X1 U7395 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5806) );
  OR2_X1 U7396 ( .A1(n6343), .A2(n5806), .ZN(n5809) );
  INV_X1 U7397 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9241) );
  OR2_X1 U7398 ( .A1(n6125), .A2(n9241), .ZN(n5808) );
  INV_X1 U7399 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9253) );
  OR2_X1 U7400 ( .A1(n6342), .A2(n9253), .ZN(n5807) );
  NAND4_X1 U7401 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n9527)
         );
  INV_X1 U7402 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6287) );
  INV_X1 U7403 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5812) );
  INV_X1 U7404 ( .A(n5817), .ZN(n5818) );
  INV_X1 U7405 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6298) );
  OR2_X1 U7406 ( .A1(n5857), .A2(n6298), .ZN(n5821) );
  OR2_X1 U7407 ( .A1(n5837), .A2(n5819), .ZN(n5820) );
  OAI211_X1 U7408 ( .C1(n5873), .C2(n6378), .A(n5821), .B(n5820), .ZN(n5830)
         );
  INV_X1 U7409 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5822) );
  OR2_X1 U7410 ( .A1(n6070), .A2(n5822), .ZN(n5826) );
  INV_X1 U7411 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10051) );
  INV_X1 U7412 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7413 ( .A1(n5841), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U7414 ( .A1(n6340), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7415 ( .A1(n5133), .A2(SI_0_), .ZN(n5828) );
  INV_X1 U7416 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5827) );
  XNOR2_X1 U7417 ( .A(n5828), .B(n5827), .ZN(n6294) );
  MUX2_X1 U7418 ( .A(n5016), .B(n6294), .S(n5873), .Z(n6696) );
  NAND2_X1 U7419 ( .A1(n4416), .A2(n5829), .ZN(n6277) );
  INV_X1 U7420 ( .A(n4415), .ZN(n6890) );
  NOR2_X1 U7421 ( .A1(n5817), .A2(n5833), .ZN(n5832) );
  MUX2_X1 U7422 ( .A(n5833), .B(n5832), .S(P1_IR_REG_2__SCAN_IN), .Z(n5834) );
  INV_X1 U7423 ( .A(n5834), .ZN(n5836) );
  INV_X1 U7424 ( .A(n5868), .ZN(n5835) );
  NAND2_X1 U7425 ( .A1(n5836), .A2(n5835), .ZN(n9189) );
  INV_X1 U7426 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6299) );
  OR2_X1 U7427 ( .A1(n5857), .A2(n6299), .ZN(n5839) );
  OR2_X1 U7428 ( .A1(n5837), .A2(n6305), .ZN(n5838) );
  OAI211_X1 U7429 ( .C1(n5873), .C2(n9189), .A(n5839), .B(n5838), .ZN(n5846)
         );
  NAND2_X1 U7430 ( .A1(n6340), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5845) );
  INV_X1 U7431 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9190) );
  INV_X1 U7432 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7433 ( .A1(n6342), .A2(n6369), .ZN(n5843) );
  INV_X1 U7434 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5840) );
  OR2_X1 U7435 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  NAND4_X2 U7436 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9171)
         );
  XNOR2_X1 U7437 ( .A(n5848), .B(n9171), .ZN(n9016) );
  NAND2_X1 U7438 ( .A1(n6723), .A2(n5849), .ZN(n6750) );
  INV_X1 U7439 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5850) );
  OR2_X1 U7440 ( .A1(n6070), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7441 ( .A1(n6340), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5851) );
  INV_X1 U7442 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6370) );
  NOR2_X1 U7443 ( .A1(n5853), .A2(n4447), .ZN(n5854) );
  OR2_X1 U7444 ( .A1(n5868), .A2(n5833), .ZN(n5856) );
  XNOR2_X1 U7445 ( .A(n5856), .B(n10285), .ZN(n6381) );
  INV_X1 U7446 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6296) );
  OR2_X1 U7447 ( .A1(n5857), .A2(n6296), .ZN(n5859) );
  OR2_X1 U7448 ( .A1(n5979), .A2(n6308), .ZN(n5858) );
  OAI211_X1 U7449 ( .C1(n5873), .C2(n6381), .A(n5859), .B(n5858), .ZN(n6866)
         );
  NAND2_X1 U7450 ( .A1(n9170), .A2(n5860), .ZN(n9061) );
  NAND2_X1 U7451 ( .A1(n6750), .A2(n9014), .ZN(n6748) );
  INV_X1 U7452 ( .A(n6866), .ZN(n6807) );
  NAND2_X1 U7453 ( .A1(n6340), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5867) );
  INV_X1 U7454 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5862) );
  OR2_X1 U7455 ( .A1(n6342), .A2(n5862), .ZN(n5866) );
  XNOR2_X1 U7456 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6564) );
  OR2_X1 U7457 ( .A1(n6131), .A2(n6564), .ZN(n5865) );
  INV_X1 U7458 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7459 ( .A1(n6343), .A2(n5863), .ZN(n5864) );
  NAND2_X1 U7460 ( .A1(n5868), .A2(n10285), .ZN(n5880) );
  NAND2_X1 U7461 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U7462 ( .A(n5870), .B(n5869), .ZN(n9215) );
  OR2_X1 U7463 ( .A1(n5979), .A2(n6309), .ZN(n5872) );
  INV_X1 U7464 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6297) );
  OR2_X1 U7465 ( .A1(n9000), .A2(n6297), .ZN(n5871) );
  NAND2_X1 U7466 ( .A1(n6755), .A2(n6875), .ZN(n8909) );
  NAND2_X1 U7467 ( .A1(n9169), .A2(n6884), .ZN(n8904) );
  NAND2_X1 U7468 ( .A1(n6759), .A2(n9015), .ZN(n6758) );
  NAND2_X1 U7469 ( .A1(n6758), .A2(n5050), .ZN(n6735) );
  AOI21_X1 U7470 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5874) );
  NOR2_X1 U7471 ( .A1(n5874), .A2(n5885), .ZN(n8799) );
  NAND2_X1 U7472 ( .A1(n6083), .A2(n8799), .ZN(n5879) );
  INV_X1 U7473 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6385) );
  INV_X1 U7474 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10052) );
  OR2_X1 U7475 ( .A1(n6342), .A2(n10052), .ZN(n5877) );
  INV_X1 U7476 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5875) );
  OR2_X1 U7477 ( .A1(n6343), .A2(n5875), .ZN(n5876) );
  INV_X1 U7478 ( .A(n9168), .ZN(n6799) );
  OR2_X1 U7479 ( .A1(n6303), .A2(n5979), .ZN(n5883) );
  NAND2_X1 U7480 ( .A1(n5891), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7481 ( .A(n5881), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U7482 ( .A1(n6034), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6329), .B2(
        n6386), .ZN(n5882) );
  NAND2_X1 U7483 ( .A1(n6799), .A2(n8805), .ZN(n8910) );
  NAND2_X1 U7484 ( .A1(n6975), .A2(n9168), .ZN(n8911) );
  NAND2_X1 U7485 ( .A1(n8910), .A2(n8911), .ZN(n9013) );
  NAND2_X1 U7486 ( .A1(n6735), .A2(n9013), .ZN(n6734) );
  NAND2_X1 U7487 ( .A1(n6734), .A2(n5042), .ZN(n6795) );
  NAND2_X1 U7488 ( .A1(n6340), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5890) );
  INV_X1 U7489 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5884) );
  OR2_X1 U7490 ( .A1(n6343), .A2(n5884), .ZN(n5889) );
  OAI21_X1 U7491 ( .B1(n5885), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5900), .ZN(
        n6833) );
  INV_X1 U7492 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7493 ( .A1(n6342), .A2(n5886), .ZN(n5887) );
  NAND4_X1 U7494 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n9167)
         );
  INV_X1 U7495 ( .A(n9167), .ZN(n8803) );
  OR2_X1 U7496 ( .A1(n6302), .A2(n5979), .ZN(n5893) );
  NOR2_X1 U7497 ( .A1(n5891), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7498 ( .A(n5910), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6424) );
  AOI22_X1 U7499 ( .A1(n6034), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6329), .B2(
        n6424), .ZN(n5892) );
  OR2_X1 U7500 ( .A1(n8803), .A2(n6961), .ZN(n8907) );
  NAND2_X1 U7501 ( .A1(n6961), .A2(n8803), .ZN(n6157) );
  NAND2_X1 U7502 ( .A1(n8907), .A2(n6157), .ZN(n9022) );
  NAND2_X1 U7503 ( .A1(n6795), .A2(n9022), .ZN(n6793) );
  OR2_X1 U7504 ( .A1(n6312), .A2(n5979), .ZN(n5898) );
  INV_X1 U7505 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7506 ( .A1(n5910), .A2(n5894), .ZN(n5895) );
  NAND2_X1 U7507 ( .A1(n5895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  XNOR2_X1 U7508 ( .A(n5896), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6391) );
  AOI22_X1 U7509 ( .A1(n6034), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6329), .B2(
        n6391), .ZN(n5897) );
  NAND2_X1 U7510 ( .A1(n6340), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5907) );
  AND2_X1 U7511 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  OR2_X1 U7512 ( .A1(n5901), .A2(n5915), .ZN(n8618) );
  OR2_X1 U7513 ( .A1(n6070), .A2(n8618), .ZN(n5906) );
  INV_X1 U7514 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5902) );
  OR2_X1 U7515 ( .A1(n6342), .A2(n5902), .ZN(n5905) );
  INV_X1 U7516 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5903) );
  OR2_X1 U7517 ( .A1(n6343), .A2(n5903), .ZN(n5904) );
  NAND4_X1 U7518 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n9166)
         );
  INV_X1 U7519 ( .A(n9166), .ZN(n7190) );
  OR2_X1 U7520 ( .A1(n9804), .A2(n7190), .ZN(n6164) );
  NAND2_X1 U7521 ( .A1(n9804), .A2(n7190), .ZN(n6931) );
  NAND2_X1 U7522 ( .A1(n6164), .A2(n6931), .ZN(n8915) );
  NAND2_X1 U7523 ( .A1(n7027), .A2(n8915), .ZN(n7026) );
  NAND2_X1 U7524 ( .A1(n9812), .A2(n7190), .ZN(n5908) );
  NAND2_X1 U7525 ( .A1(n6314), .A2(n8998), .ZN(n5913) );
  OAI21_X1 U7526 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7527 ( .A1(n5910), .A2(n5909), .ZN(n5922) );
  XNOR2_X1 U7528 ( .A(n5922), .B(n5911), .ZN(n6393) );
  AOI22_X1 U7529 ( .A1(n6034), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6329), .B2(
        n6393), .ZN(n5912) );
  NAND2_X1 U7530 ( .A1(n5913), .A2(n5912), .ZN(n7194) );
  NAND2_X1 U7531 ( .A1(n6340), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5920) );
  INV_X1 U7532 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7533 ( .A1(n6343), .A2(n5914), .ZN(n5919) );
  OR2_X1 U7534 ( .A1(n5915), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7535 ( .A1(n5928), .A2(n5916), .ZN(n7191) );
  OR2_X1 U7536 ( .A1(n6131), .A2(n7191), .ZN(n5918) );
  INV_X1 U7537 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6953) );
  OR2_X1 U7538 ( .A1(n6342), .A2(n6953), .ZN(n5917) );
  NAND4_X1 U7539 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n9165)
         );
  OR2_X1 U7540 ( .A1(n7194), .A2(n8619), .ZN(n8918) );
  NAND2_X1 U7541 ( .A1(n7194), .A2(n8619), .ZN(n8901) );
  NAND2_X1 U7542 ( .A1(n8918), .A2(n8901), .ZN(n6948) );
  OR2_X1 U7543 ( .A1(n7194), .A2(n9165), .ZN(n5921) );
  NAND2_X1 U7544 ( .A1(n6324), .A2(n8998), .ZN(n5925) );
  OAI21_X1 U7545 ( .B1(n5922), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U7546 ( .A(n5923), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9245) );
  AOI22_X1 U7547 ( .A1(n6034), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6329), .B2(
        n9245), .ZN(n5924) );
  NAND2_X1 U7548 ( .A1(n6124), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5933) );
  INV_X1 U7549 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7550 ( .A1(n6125), .A2(n5926), .ZN(n5932) );
  NAND2_X1 U7551 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7552 ( .A1(n5946), .A2(n5929), .ZN(n7300) );
  OR2_X1 U7553 ( .A1(n6070), .A2(n7300), .ZN(n5931) );
  INV_X1 U7554 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6940) );
  OR2_X1 U7555 ( .A1(n6342), .A2(n6940), .ZN(n5930) );
  NAND4_X1 U7556 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n9164)
         );
  NAND2_X1 U7557 ( .A1(n7294), .A2(n8728), .ZN(n8928) );
  NAND2_X1 U7558 ( .A1(n9026), .A2(n8928), .ZN(n6937) );
  NOR2_X1 U7559 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5935) );
  AND2_X1 U7560 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  AND2_X1 U7561 ( .A1(n5938), .A2(n5937), .ZN(n5941) );
  NOR2_X1 U7562 ( .A1(n5941), .A2(n5833), .ZN(n5939) );
  MUX2_X1 U7563 ( .A(n5833), .B(n5939), .S(P1_IR_REG_10__SCAN_IN), .Z(n5943)
         );
  NAND2_X1 U7564 ( .A1(n5941), .A2(n5940), .ZN(n5955) );
  INV_X1 U7565 ( .A(n5955), .ZN(n5942) );
  NOR2_X1 U7566 ( .A1(n5943), .A2(n5942), .ZN(n9717) );
  AOI22_X1 U7567 ( .A1(n6034), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6329), .B2(
        n9717), .ZN(n5944) );
  NAND2_X1 U7568 ( .A1(n6340), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5952) );
  INV_X1 U7569 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9243) );
  OR2_X1 U7570 ( .A1(n6342), .A2(n9243), .ZN(n5951) );
  NAND2_X1 U7571 ( .A1(n5946), .A2(n8727), .ZN(n5947) );
  NAND2_X1 U7572 ( .A1(n5960), .A2(n5947), .ZN(n8729) );
  OR2_X1 U7573 ( .A1(n6131), .A2(n8729), .ZN(n5950) );
  INV_X1 U7574 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7575 ( .A1(n6343), .A2(n5948), .ZN(n5949) );
  NAND4_X1 U7576 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n9163)
         );
  NAND2_X1 U7577 ( .A1(n8731), .A2(n5953), .ZN(n8930) );
  NAND2_X1 U7578 ( .A1(n6350), .A2(n8998), .ZN(n5958) );
  NAND2_X1 U7579 ( .A1(n5955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7580 ( .A(n5956), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U7581 ( .A1(n6034), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6329), .B2(
        n9743), .ZN(n5957) );
  NAND2_X1 U7582 ( .A1(n6340), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5965) );
  INV_X1 U7583 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7132) );
  OR2_X1 U7584 ( .A1(n6342), .A2(n7132), .ZN(n5964) );
  OR2_X1 U7585 ( .A1(n5054), .A2(n5971), .ZN(n8859) );
  OR2_X1 U7586 ( .A1(n6070), .A2(n8859), .ZN(n5963) );
  INV_X1 U7587 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5961) );
  OR2_X1 U7588 ( .A1(n6343), .A2(n5961), .ZN(n5962) );
  NAND4_X1 U7589 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n9162)
         );
  INV_X1 U7590 ( .A(n9162), .ZN(n8764) );
  NAND2_X1 U7591 ( .A1(n8862), .A2(n8764), .ZN(n8931) );
  NAND2_X1 U7592 ( .A1(n8933), .A2(n8931), .ZN(n9031) );
  NAND2_X1 U7593 ( .A1(n7129), .A2(n9031), .ZN(n7128) );
  NAND2_X1 U7594 ( .A1(n7131), .A2(n8764), .ZN(n5966) );
  NAND2_X1 U7595 ( .A1(n7128), .A2(n5966), .ZN(n7229) );
  NAND2_X1 U7596 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7597 ( .A(n5968), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U7598 ( .A1(n6034), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6329), .B2(
        n9754), .ZN(n5969) );
  NAND2_X1 U7599 ( .A1(n6124), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5976) );
  INV_X1 U7600 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9236) );
  OR2_X1 U7601 ( .A1(n6125), .A2(n9236), .ZN(n5975) );
  OR2_X1 U7602 ( .A1(n5971), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7603 ( .A1(n5986), .A2(n5972), .ZN(n8765) );
  OR2_X1 U7604 ( .A1(n6070), .A2(n8765), .ZN(n5974) );
  INV_X1 U7605 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7233) );
  OR2_X1 U7606 ( .A1(n6342), .A2(n7233), .ZN(n5973) );
  NAND4_X1 U7607 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n9161)
         );
  INV_X1 U7608 ( .A(n9161), .ZN(n8839) );
  OR2_X1 U7609 ( .A1(n8768), .A2(n8839), .ZN(n8934) );
  NAND2_X1 U7610 ( .A1(n8768), .A2(n8839), .ZN(n9070) );
  NAND2_X1 U7611 ( .A1(n8934), .A2(n9070), .ZN(n9032) );
  NAND2_X1 U7612 ( .A1(n7229), .A2(n9032), .ZN(n7228) );
  NAND2_X1 U7613 ( .A1(n5977), .A2(n8839), .ZN(n5978) );
  OR2_X1 U7614 ( .A1(n5980), .A2(n5833), .ZN(n5981) );
  XNOR2_X1 U7615 ( .A(n5981), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9248) );
  AOI22_X1 U7616 ( .A1(n6034), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6329), .B2(
        n9248), .ZN(n5982) );
  NAND2_X1 U7617 ( .A1(n6340), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5992) );
  INV_X1 U7618 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7619 ( .A1(n6342), .A2(n5984), .ZN(n5991) );
  NAND2_X1 U7620 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7621 ( .A1(n5999), .A2(n5987), .ZN(n8840) );
  OR2_X1 U7622 ( .A1(n6131), .A2(n8840), .ZN(n5990) );
  INV_X1 U7623 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7624 ( .A1(n6343), .A2(n5988), .ZN(n5989) );
  NAND4_X1 U7625 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n9160)
         );
  NAND2_X1 U7626 ( .A1(n8843), .A2(n5993), .ZN(n9069) );
  NAND2_X1 U7627 ( .A1(n8937), .A2(n9069), .ZN(n9034) );
  NAND2_X1 U7628 ( .A1(n7347), .A2(n9034), .ZN(n7346) );
  NAND2_X1 U7629 ( .A1(n7355), .A2(n5993), .ZN(n5994) );
  NAND2_X1 U7630 ( .A1(n6461), .A2(n8998), .ZN(n5997) );
  NAND2_X1 U7631 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7632 ( .A(n6008), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U7633 ( .A1(n6034), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6329), .B2(
        n9784), .ZN(n5996) );
  AND2_X1 U7634 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NOR2_X1 U7635 ( .A1(n6013), .A2(n6000), .ZN(n9559) );
  NAND2_X1 U7636 ( .A1(n6083), .A2(n9559), .ZN(n6006) );
  INV_X1 U7637 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7638 ( .A1(n6343), .A2(n6001), .ZN(n6005) );
  INV_X1 U7639 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9228) );
  OR2_X1 U7640 ( .A1(n6125), .A2(n9228), .ZN(n6004) );
  INV_X1 U7641 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7642 ( .A1(n6342), .A2(n6002), .ZN(n6003) );
  NAND4_X1 U7643 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n9529)
         );
  NAND2_X1 U7644 ( .A1(n9647), .A2(n8892), .ZN(n8926) );
  INV_X1 U7645 ( .A(n9647), .ZN(n9561) );
  NAND2_X1 U7646 ( .A1(n6545), .A2(n8998), .ZN(n6012) );
  NAND2_X1 U7647 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7648 ( .A1(n6009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7649 ( .A(n6010), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U7650 ( .A1(n6034), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6329), .B2(
        n10328), .ZN(n6011) );
  NOR2_X1 U7651 ( .A1(n6013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7652 ( .A1(n6015), .A2(n6014), .ZN(n8893) );
  INV_X1 U7653 ( .A(n8893), .ZN(n9536) );
  NAND2_X1 U7654 ( .A1(n6083), .A2(n9536), .ZN(n6020) );
  INV_X1 U7655 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10321) );
  OR2_X1 U7656 ( .A1(n6125), .A2(n10321), .ZN(n6019) );
  INV_X1 U7657 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10223) );
  OR2_X1 U7658 ( .A1(n6343), .A2(n10223), .ZN(n6018) );
  INV_X1 U7659 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7660 ( .A1(n6342), .A2(n6016), .ZN(n6017) );
  NAND4_X1 U7661 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n9159)
         );
  INV_X1 U7662 ( .A(n9159), .ZN(n9550) );
  NOR2_X1 U7663 ( .A1(n9690), .A2(n9550), .ZN(n6021) );
  INV_X1 U7664 ( .A(n9527), .ZN(n8889) );
  NAND2_X1 U7665 ( .A1(n9637), .A2(n8889), .ZN(n9076) );
  NAND2_X1 U7666 ( .A1(n6670), .A2(n8998), .ZN(n6024) );
  NAND2_X1 U7667 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7668 ( .A(n6022), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9288) );
  AOI22_X1 U7669 ( .A1(n6034), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6329), .B2(
        n9288), .ZN(n6023) );
  NAND2_X1 U7670 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7671 ( .A1(n6038), .A2(n6027), .ZN(n9500) );
  INV_X1 U7672 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9632) );
  OR2_X1 U7673 ( .A1(n6125), .A2(n9632), .ZN(n6029) );
  INV_X1 U7674 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9501) );
  OR2_X1 U7675 ( .A1(n6342), .A2(n9501), .ZN(n6028) );
  AND2_X1 U7676 ( .A1(n6029), .A2(n6028), .ZN(n6031) );
  NAND2_X1 U7677 ( .A1(n6124), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6030) );
  OAI211_X1 U7678 ( .C1(n9500), .C2(n6131), .A(n6031), .B(n6030), .ZN(n9158)
         );
  NAND2_X1 U7679 ( .A1(n9498), .A2(n9158), .ZN(n6032) );
  INV_X1 U7680 ( .A(n9158), .ZN(n9510) );
  NAND2_X1 U7681 ( .A1(n6801), .A2(n8998), .ZN(n6036) );
  XNOR2_X1 U7682 ( .A(n6033), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U7683 ( .A1(n6034), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6329), .B2(
        n9799), .ZN(n6035) );
  AND2_X1 U7684 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  OR2_X1 U7685 ( .A1(n6039), .A2(n6049), .ZN(n9480) );
  AOI22_X1 U7686 ( .A1(n6340), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6124), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7687 ( .A1(n6095), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6040) );
  OAI211_X1 U7688 ( .C1(n9480), .C2(n6070), .A(n6041), .B(n6040), .ZN(n9492)
         );
  NAND2_X1 U7689 ( .A1(n9477), .A2(n6042), .ZN(n6043) );
  INV_X1 U7690 ( .A(n9625), .ZN(n9479) );
  INV_X1 U7691 ( .A(n9492), .ZN(n8812) );
  NAND2_X1 U7692 ( .A1(n6043), .A2(n4446), .ZN(n9459) );
  NAND2_X1 U7693 ( .A1(n7069), .A2(n8998), .ZN(n6048) );
  INV_X1 U7694 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7695 ( .A1(n9000), .A2(n6046), .ZN(n6047) );
  INV_X1 U7696 ( .A(n9614), .ZN(n9450) );
  AOI21_X1 U7697 ( .B1(n6049), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7698 ( .A1(n6058), .A2(n6050), .ZN(n9447) );
  INV_X1 U7699 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U7700 ( .A1(n6340), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7701 ( .A1(n6095), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7702 ( .C1(n10272), .C2(n6343), .A(n6052), .B(n6051), .ZN(n6053)
         );
  INV_X1 U7703 ( .A(n6053), .ZN(n6054) );
  OAI21_X1 U7704 ( .B1(n9447), .B2(n6070), .A(n6054), .ZN(n9464) );
  INV_X1 U7705 ( .A(n9464), .ZN(n7838) );
  NAND2_X1 U7706 ( .A1(n7149), .A2(n8998), .ZN(n6057) );
  OR2_X1 U7707 ( .A1(n9000), .A2(n10284), .ZN(n6056) );
  OR2_X1 U7708 ( .A1(n6058), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6059) );
  AND2_X1 U7709 ( .A1(n6068), .A2(n6059), .ZN(n9438) );
  NAND2_X1 U7710 ( .A1(n9438), .A2(n6083), .ZN(n6064) );
  INV_X1 U7711 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U7712 ( .A1(n6095), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7713 ( .A1(n6124), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6060) );
  OAI211_X1 U7714 ( .C1(n6125), .C2(n10123), .A(n6061), .B(n6060), .ZN(n6062)
         );
  INV_X1 U7715 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7716 ( .A1(n6064), .A2(n6063), .ZN(n9454) );
  INV_X1 U7717 ( .A(n9454), .ZN(n8961) );
  NAND2_X1 U7718 ( .A1(n7305), .A2(n8998), .ZN(n6067) );
  OR2_X1 U7719 ( .A1(n9000), .A2(n7309), .ZN(n6066) );
  NAND2_X1 U7720 ( .A1(n6068), .A2(n8849), .ZN(n6069) );
  NAND2_X1 U7721 ( .A1(n6081), .A2(n6069), .ZN(n9417) );
  OR2_X1 U7722 ( .A1(n9417), .A2(n6070), .ZN(n6076) );
  INV_X1 U7723 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7724 ( .A1(n6095), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7725 ( .A1(n6124), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6071) );
  OAI211_X1 U7726 ( .C1(n6125), .C2(n6073), .A(n6072), .B(n6071), .ZN(n6074)
         );
  INV_X1 U7727 ( .A(n6074), .ZN(n6075) );
  NAND2_X1 U7728 ( .A1(n6076), .A2(n6075), .ZN(n9433) );
  NAND2_X1 U7729 ( .A1(n9605), .A2(n9433), .ZN(n6077) );
  INV_X1 U7730 ( .A(n9433), .ZN(n8650) );
  NAND2_X1 U7731 ( .A1(n7327), .A2(n8998), .ZN(n6079) );
  OR2_X1 U7732 ( .A1(n9000), .A2(n7326), .ZN(n6078) );
  NAND2_X1 U7733 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  AND2_X1 U7734 ( .A1(n6092), .A2(n6082), .ZN(n9408) );
  NAND2_X1 U7735 ( .A1(n9408), .A2(n6083), .ZN(n6088) );
  INV_X1 U7736 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U7737 ( .A1(n6340), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7738 ( .A1(n6095), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6084) );
  OAI211_X1 U7739 ( .C1(n6343), .C2(n10165), .A(n6085), .B(n6084), .ZN(n6086)
         );
  INV_X1 U7740 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7741 ( .A1(n6088), .A2(n6087), .ZN(n9424) );
  INV_X1 U7742 ( .A(n9424), .ZN(n8850) );
  NAND2_X1 U7743 ( .A1(n9673), .A2(n8850), .ZN(n6089) );
  OR2_X1 U7744 ( .A1(n9000), .A2(n10079), .ZN(n6090) );
  AND2_X1 U7745 ( .A1(n6092), .A2(n8823), .ZN(n6094) );
  OR2_X1 U7746 ( .A1(n6094), .A2(n6093), .ZN(n9386) );
  INV_X1 U7747 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7748 ( .A1(n6095), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7749 ( .A1(n6124), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7750 ( .C1(n6125), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6099)
         );
  INV_X1 U7751 ( .A(n6099), .ZN(n6100) );
  OAI21_X1 U7752 ( .B1(n9386), .B2(n6131), .A(n6100), .ZN(n9403) );
  NAND2_X1 U7753 ( .A1(n9595), .A2(n9403), .ZN(n6102) );
  NOR2_X1 U7754 ( .A1(n9595), .A2(n9403), .ZN(n6101) );
  NAND2_X1 U7755 ( .A1(n9375), .A2(n9393), .ZN(n6103) );
  NAND2_X1 U7756 ( .A1(n6104), .A2(n6103), .ZN(n9349) );
  OR2_X1 U7757 ( .A1(n9000), .A2(n7455), .ZN(n6105) );
  NAND2_X1 U7758 ( .A1(n6340), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6113) );
  INV_X1 U7759 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7760 ( .A1(n6343), .A2(n6106), .ZN(n6112) );
  OAI21_X1 U7761 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6108), .A(n6127), .ZN(
        n9353) );
  OR2_X1 U7762 ( .A1(n6131), .A2(n9353), .ZN(n6111) );
  INV_X1 U7763 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7764 ( .A1(n6342), .A2(n6109), .ZN(n6110) );
  NAND4_X1 U7765 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n9371)
         );
  NAND2_X1 U7766 ( .A1(n9585), .A2(n9371), .ZN(n6114) );
  OR2_X1 U7767 ( .A1(n9000), .A2(n7764), .ZN(n6115) );
  NAND2_X1 U7768 ( .A1(n6340), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6121) );
  INV_X1 U7769 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10098) );
  OR2_X1 U7770 ( .A1(n6343), .A2(n10098), .ZN(n6120) );
  INV_X1 U7771 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6126) );
  XNOR2_X1 U7772 ( .A(n6127), .B(n6126), .ZN(n8704) );
  OR2_X1 U7773 ( .A1(n6131), .A2(n8704), .ZN(n6119) );
  INV_X1 U7774 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7775 ( .A1(n6342), .A2(n6117), .ZN(n6118) );
  NAND4_X1 U7776 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n9360)
         );
  OR2_X1 U7777 ( .A1(n9000), .A2(n9708), .ZN(n6122) );
  NAND2_X1 U7778 ( .A1(n6124), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6136) );
  INV_X1 U7779 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10099) );
  OR2_X1 U7780 ( .A1(n6125), .A2(n10099), .ZN(n6135) );
  INV_X1 U7781 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8745) );
  OAI21_X1 U7782 ( .B1(n6127), .B2(n6126), .A(n8745), .ZN(n6130) );
  INV_X1 U7783 ( .A(n6127), .ZN(n6129) );
  AND2_X1 U7784 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6128) );
  NAND2_X1 U7785 ( .A1(n6129), .A2(n6128), .ZN(n9311) );
  NAND2_X1 U7786 ( .A1(n6130), .A2(n9311), .ZN(n9323) );
  OR2_X1 U7787 ( .A1(n6131), .A2(n9323), .ZN(n6134) );
  INV_X1 U7788 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6132) );
  OR2_X1 U7789 ( .A1(n6342), .A2(n6132), .ZN(n6133) );
  NAND4_X1 U7790 ( .A1(n6136), .A2(n6135), .A3(n6134), .A4(n6133), .ZN(n9337)
         );
  NAND2_X1 U7791 ( .A1(n9574), .A2(n9337), .ZN(n6137) );
  NAND2_X1 U7792 ( .A1(n9322), .A2(n6137), .ZN(n6146) );
  NAND2_X1 U7793 ( .A1(n7518), .A2(n8998), .ZN(n6139) );
  OR2_X1 U7794 ( .A1(n9000), .A2(n9703), .ZN(n6138) );
  NAND2_X1 U7795 ( .A1(n6340), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6145) );
  INV_X1 U7796 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7797 ( .A1(n6343), .A2(n6140), .ZN(n6144) );
  OR2_X1 U7798 ( .A1(n6131), .A2(n9311), .ZN(n6143) );
  INV_X1 U7799 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7800 ( .A1(n6342), .A2(n6141), .ZN(n6142) );
  XNOR2_X1 U7801 ( .A(n6146), .B(n8992), .ZN(n9309) );
  NOR2_X1 U7802 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6147) );
  NAND2_X1 U7803 ( .A1(n6148), .A2(n6147), .ZN(n6151) );
  INV_X1 U7804 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7805 ( .A1(n6154), .A2(n6288), .ZN(n6729) );
  INV_X1 U7806 ( .A(n6729), .ZN(n9133) );
  NAND2_X1 U7807 ( .A1(n6151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6152) );
  INV_X1 U7808 ( .A(n6501), .ZN(n9147) );
  AND2_X1 U7809 ( .A1(n9133), .A2(n9147), .ZN(n6689) );
  INV_X1 U7810 ( .A(n6154), .ZN(n7307) );
  INV_X1 U7811 ( .A(n6288), .ZN(n9056) );
  NAND2_X1 U7812 ( .A1(n7307), .A2(n9056), .ZN(n6597) );
  INV_X1 U7813 ( .A(n6597), .ZN(n6690) );
  NAND2_X1 U7814 ( .A1(n6154), .A2(n6153), .ZN(n6509) );
  AND2_X1 U7815 ( .A1(n6501), .A2(n6509), .ZN(n6155) );
  OR3_X1 U7816 ( .A1(n6689), .A2(n6690), .A3(n6155), .ZN(n6278) );
  INV_X1 U7817 ( .A(n9139), .ZN(n9137) );
  INV_X1 U7818 ( .A(n9403), .ZN(n8777) );
  NAND2_X1 U7819 ( .A1(n9595), .A2(n8777), .ZN(n9104) );
  NAND2_X1 U7820 ( .A1(n8901), .A2(n6931), .ZN(n8917) );
  AND2_X1 U7821 ( .A1(n8917), .A2(n8918), .ZN(n6932) );
  NAND2_X1 U7822 ( .A1(n6932), .A2(n9026), .ZN(n6156) );
  NAND2_X1 U7823 ( .A1(n6156), .A2(n8928), .ZN(n9028) );
  INV_X1 U7824 ( .A(n6157), .ZN(n8914) );
  NOR2_X1 U7825 ( .A1(n9028), .A2(n8914), .ZN(n9063) );
  AND2_X1 U7826 ( .A1(n6591), .A2(n5829), .ZN(n6593) );
  NAND2_X1 U7827 ( .A1(n6158), .A2(n6593), .ZN(n6160) );
  INV_X1 U7828 ( .A(n9057), .ZN(n6594) );
  NAND2_X1 U7829 ( .A1(n6594), .A2(n6890), .ZN(n6159) );
  NAND2_X1 U7830 ( .A1(n5847), .A2(n5846), .ZN(n6161) );
  INV_X1 U7831 ( .A(n8904), .ZN(n6163) );
  INV_X1 U7832 ( .A(n8910), .ZN(n8906) );
  NAND2_X1 U7833 ( .A1(n9063), .A2(n9062), .ZN(n6166) );
  AND2_X1 U7834 ( .A1(n8918), .A2(n6164), .ZN(n9025) );
  AND3_X1 U7835 ( .A1(n9026), .A2(n9025), .A3(n8907), .ZN(n6165) );
  OR2_X1 U7836 ( .A1(n9028), .A2(n6165), .ZN(n9055) );
  INV_X1 U7837 ( .A(n8930), .ZN(n8925) );
  NOR2_X1 U7838 ( .A1(n9031), .A2(n8925), .ZN(n6167) );
  INV_X1 U7839 ( .A(n9069), .ZN(n8936) );
  XNOR2_X1 U7840 ( .A(n9535), .B(n9159), .ZN(n9525) );
  OR2_X1 U7841 ( .A1(n9535), .A2(n9550), .ZN(n8940) );
  NAND2_X1 U7842 ( .A1(n9508), .A2(n9511), .ZN(n6168) );
  NAND2_X1 U7843 ( .A1(n6168), .A2(n8947), .ZN(n9490) );
  XNOR2_X1 U7844 ( .A(n9498), .B(n9158), .ZN(n9495) );
  OR2_X1 U7845 ( .A1(n9498), .A2(n9510), .ZN(n8952) );
  OR2_X1 U7846 ( .A1(n9625), .A2(n8812), .ZN(n9084) );
  NAND2_X1 U7847 ( .A1(n9625), .A2(n8812), .ZN(n8953) );
  NAND2_X1 U7848 ( .A1(n9084), .A2(n8953), .ZN(n9485) );
  OR2_X1 U7849 ( .A1(n9470), .A2(n9487), .ZN(n9083) );
  NAND2_X1 U7850 ( .A1(n9470), .A2(n9487), .ZN(n8954) );
  NAND2_X1 U7851 ( .A1(n9614), .A2(n7838), .ZN(n8960) );
  NAND2_X1 U7852 ( .A1(n8964), .A2(n8960), .ZN(n9452) );
  XNOR2_X1 U7853 ( .A(n9437), .B(n9454), .ZN(n9430) );
  NAND2_X1 U7854 ( .A1(n9431), .A2(n9430), .ZN(n9429) );
  NAND2_X1 U7855 ( .A1(n9437), .A2(n8961), .ZN(n8965) );
  NAND2_X1 U7856 ( .A1(n9429), .A2(n8965), .ZN(n9422) );
  OR2_X1 U7857 ( .A1(n9605), .A2(n8650), .ZN(n8962) );
  NAND2_X1 U7858 ( .A1(n9605), .A2(n8650), .ZN(n8967) );
  NAND2_X1 U7859 ( .A1(n9422), .A2(n9423), .ZN(n9421) );
  INV_X1 U7860 ( .A(n9348), .ZN(n9359) );
  NAND2_X1 U7861 ( .A1(n6154), .A2(n9143), .ZN(n6169) );
  NAND2_X1 U7862 ( .A1(n6288), .A2(n9137), .ZN(n9050) );
  NAND2_X1 U7863 ( .A1(n6169), .A2(n9050), .ZN(n9523) );
  OR2_X1 U7864 ( .A1(n6729), .A2(n9705), .ZN(n9551) );
  INV_X1 U7865 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7866 ( .A1(n6340), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6172) );
  INV_X1 U7867 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9658) );
  OR2_X1 U7868 ( .A1(n6343), .A2(n9658), .ZN(n6171) );
  OAI211_X1 U7869 ( .C1(n6342), .C2(n6173), .A(n6172), .B(n6171), .ZN(n9157)
         );
  INV_X1 U7870 ( .A(n9183), .ZN(n9729) );
  NAND2_X1 U7871 ( .A1(n9729), .A2(P1_B_REG_SCAN_IN), .ZN(n9298) );
  NAND2_X1 U7872 ( .A1(n9157), .A2(n9298), .ZN(n6174) );
  INV_X1 U7873 ( .A(n9705), .ZN(n9186) );
  OR2_X1 U7874 ( .A1(n6729), .A2(n9186), .ZN(n9549) );
  OAI22_X1 U7875 ( .A1(n8979), .A2(n9551), .B1(n6174), .B2(n9549), .ZN(n6175)
         );
  INV_X1 U7876 ( .A(n9585), .ZN(n9356) );
  NAND2_X1 U7877 ( .A1(n4415), .A2(n6696), .ZN(n6725) );
  OR2_X1 U7878 ( .A1(n6725), .A2(n5846), .ZN(n6751) );
  INV_X1 U7879 ( .A(n7194), .ZN(n9821) );
  INV_X1 U7880 ( .A(n7294), .ZN(n9827) );
  OR2_X2 U7881 ( .A1(n6597), .A2(n9137), .ZN(n9557) );
  AOI21_X1 U7882 ( .B1(n9314), .B2(n4591), .A(n9557), .ZN(n6179) );
  NAND2_X1 U7883 ( .A1(n6179), .A2(n9304), .ZN(n9317) );
  NAND2_X1 U7884 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  NAND2_X1 U7885 ( .A1(n6182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6184) );
  INV_X1 U7886 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6183) );
  XNOR2_X1 U7887 ( .A(n6184), .B(n6183), .ZN(n6521) );
  INV_X1 U7888 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7889 ( .A1(n6193), .A2(n6192), .ZN(n6186) );
  NAND2_X1 U7890 ( .A1(n6186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6187) );
  INV_X1 U7891 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10047) );
  INV_X1 U7892 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7893 ( .A1(n6189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7894 ( .A(n6191), .B(n6190), .ZN(n7437) );
  XNOR2_X1 U7895 ( .A(n6193), .B(n6192), .ZN(n7451) );
  AND2_X1 U7896 ( .A1(n6520), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7897 ( .A1(n7451), .A2(P1_B_REG_SCAN_IN), .ZN(n6195) );
  MUX2_X1 U7898 ( .A(P1_B_REG_SCAN_IN), .B(n6195), .S(n7437), .Z(n6197) );
  INV_X1 U7899 ( .A(n7457), .ZN(n6196) );
  NAND2_X1 U7900 ( .A1(n6197), .A2(n6196), .ZN(n6335) );
  NOR4_X1 U7901 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6199) );
  NOR4_X1 U7902 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6198) );
  AND2_X1 U7903 ( .A1(n6199), .A2(n6198), .ZN(n10043) );
  NOR4_X1 U7904 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6200) );
  INV_X1 U7905 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10161) );
  INV_X1 U7906 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10206) );
  NAND4_X1 U7907 ( .A1(n10043), .A2(n6200), .A3(n10161), .A4(n10206), .ZN(
        n6206) );
  NOR4_X1 U7908 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6204) );
  NOR4_X1 U7909 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6203) );
  NOR4_X1 U7910 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6202) );
  NOR4_X1 U7911 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6201) );
  NAND4_X1 U7912 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n6205)
         );
  NOR2_X1 U7913 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  OR2_X1 U7914 ( .A1(n6335), .A2(n6207), .ZN(n6515) );
  NAND2_X1 U7915 ( .A1(n9693), .A2(n6515), .ZN(n6498) );
  OR2_X1 U7916 ( .A1(n6729), .A2(n9147), .ZN(n6522) );
  INV_X1 U7917 ( .A(n6522), .ZN(n6208) );
  NOR2_X1 U7918 ( .A1(n9651), .A2(n6288), .ZN(n6285) );
  INV_X1 U7919 ( .A(n6335), .ZN(n6211) );
  INV_X1 U7920 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7921 ( .A1(n6211), .A2(n6338), .ZN(n6209) );
  NAND2_X1 U7922 ( .A1(n7457), .A2(n7451), .ZN(n6336) );
  NAND2_X1 U7923 ( .A1(n6209), .A2(n6336), .ZN(n6496) );
  INV_X1 U7924 ( .A(n6496), .ZN(n6282) );
  OR2_X1 U7925 ( .A1(n6285), .A2(n6282), .ZN(n6210) );
  INV_X1 U7926 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U7927 ( .A1(n6211), .A2(n10083), .ZN(n6213) );
  NAND2_X1 U7928 ( .A1(n7457), .A2(n7437), .ZN(n6212) );
  NAND2_X1 U7929 ( .A1(n6213), .A2(n6212), .ZN(n6497) );
  INV_X1 U7930 ( .A(n6497), .ZN(n9694) );
  OR2_X1 U7931 ( .A1(n9839), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7932 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  OR2_X1 U7933 ( .A1(n6597), .A2(n9147), .ZN(n9833) );
  INV_X1 U7934 ( .A(n9833), .ZN(n9648) );
  NAND2_X1 U7935 ( .A1(n9691), .A2(n9648), .ZN(n9689) );
  NAND2_X1 U7936 ( .A1(n6216), .A2(n5046), .ZN(P1_U3519) );
  OR2_X1 U7937 ( .A1(n9845), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6219) );
  INV_X2 U7938 ( .A(n9843), .ZN(n9845) );
  NAND2_X1 U7939 ( .A1(n9845), .A2(n9648), .ZN(n9645) );
  NAND2_X1 U7940 ( .A1(n6220), .A2(n5051), .ZN(P1_U3551) );
  INV_X1 U7941 ( .A(n6319), .ZN(n7328) );
  OR2_X1 U7942 ( .A1(n6638), .A2(n7328), .ZN(n6238) );
  INV_X2 U7943 ( .A(n8185), .ZN(P2_U3893) );
  NOR2_X1 U7944 ( .A1(n6520), .A2(P1_U3086), .ZN(n6221) );
  NAND2_X1 U7945 ( .A1(n6638), .A2(n7739), .ZN(n6222) );
  NAND2_X1 U7946 ( .A1(n6222), .A2(n6319), .ZN(n9847) );
  NAND2_X1 U7947 ( .A1(n9847), .A2(n5189), .ZN(n6223) );
  NAND2_X1 U7948 ( .A1(n6223), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U7949 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8208), .Z(n6699) );
  XNOR2_X1 U7950 ( .A(n6699), .B(n6708), .ZN(n6234) );
  MUX2_X1 U7951 ( .A(n6225), .B(n6224), .S(n8208), .Z(n6231) );
  INV_X1 U7952 ( .A(n6231), .ZN(n6232) );
  MUX2_X1 U7953 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8208), .Z(n6230) );
  MUX2_X1 U7954 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5681), .Z(n6228) );
  XNOR2_X1 U7955 ( .A(n9858), .B(n6228), .ZN(n9862) );
  NAND2_X1 U7956 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  NAND2_X1 U7957 ( .A1(n6228), .A2(n4883), .ZN(n6229) );
  NAND2_X1 U7958 ( .A1(n9860), .A2(n6229), .ZN(n9874) );
  INV_X1 U7959 ( .A(n6306), .ZN(n9880) );
  XNOR2_X1 U7960 ( .A(n6230), .B(n9880), .ZN(n9873) );
  AND2_X1 U7961 ( .A1(n9874), .A2(n9873), .ZN(n9876) );
  XNOR2_X1 U7962 ( .A(n6231), .B(n6481), .ZN(n6478) );
  NAND2_X1 U7963 ( .A1(n6479), .A2(n6478), .ZN(n6477) );
  OAI21_X1 U7964 ( .B1(n6232), .B2(n6481), .A(n6477), .ZN(n6233) );
  NOR2_X2 U7965 ( .A1(n8185), .A2(n7750), .ZN(n9872) );
  INV_X1 U7966 ( .A(n9872), .ZN(n9848) );
  AOI211_X1 U7967 ( .C1(n6234), .C2(n6233), .A(n9848), .B(n6698), .ZN(n6275)
         );
  INV_X1 U7968 ( .A(n6238), .ZN(n6235) );
  INV_X1 U7969 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6236) );
  NOR2_X1 U7970 ( .A1(n9887), .A2(n6236), .ZN(n6274) );
  NOR2_X1 U7971 ( .A1(n8208), .A2(P2_U3151), .ZN(n7459) );
  AND2_X1 U7972 ( .A1(n7459), .A2(n5680), .ZN(n6237) );
  NAND2_X1 U7973 ( .A1(n9847), .A2(n6237), .ZN(n6240) );
  OR2_X1 U7974 ( .A1(n5680), .A2(P2_U3151), .ZN(n9849) );
  OR2_X1 U7975 ( .A1(n6238), .A2(n9849), .ZN(n6239) );
  NAND2_X1 U7976 ( .A1(n6240), .A2(n6239), .ZN(n9881) );
  INV_X1 U7977 ( .A(n6708), .ZN(n6241) );
  AND2_X1 U7978 ( .A1(n9881), .A2(n6241), .ZN(n6273) );
  NOR2_X1 U7979 ( .A1(n9849), .A2(n6226), .ZN(n6242) );
  NAND2_X1 U7980 ( .A1(n6242), .A2(n9847), .ZN(n8224) );
  INV_X1 U7981 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9977) );
  INV_X1 U7982 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7983 ( .A1(n6255), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7984 ( .A1(n9858), .A2(n6243), .ZN(n6244) );
  NAND2_X1 U7985 ( .A1(n6257), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7986 ( .A1(n6244), .A2(n6245), .ZN(n9867) );
  INV_X1 U7987 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U7988 ( .A1(n9866), .A2(n6245), .ZN(n9890) );
  NAND2_X1 U7989 ( .A1(n6306), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7990 ( .A1(n9889), .A2(n6246), .ZN(n6247) );
  OAI21_X1 U7991 ( .B1(n6247), .B2(n6481), .A(n6251), .ZN(n6484) );
  NAND2_X1 U7992 ( .A1(n6482), .A2(n6251), .ZN(n6249) );
  XNOR2_X1 U7993 ( .A(n6708), .B(n6248), .ZN(n6250) );
  NAND2_X1 U7994 ( .A1(n6249), .A2(n6250), .ZN(n6710) );
  INV_X1 U7995 ( .A(n6250), .ZN(n6252) );
  NAND3_X1 U7996 ( .A1(n6482), .A2(n6252), .A3(n6251), .ZN(n6253) );
  AND2_X1 U7997 ( .A1(n6710), .A2(n6253), .ZN(n6271) );
  NOR2_X1 U7998 ( .A1(n9849), .A2(n8208), .ZN(n6254) );
  NAND2_X1 U7999 ( .A1(n6254), .A2(n9847), .ZN(n8221) );
  INV_X1 U8000 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U8001 ( .A1(n6255), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U8002 ( .A1(n9858), .A2(n6256), .ZN(n6258) );
  NAND2_X1 U8003 ( .A1(n6257), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U8004 ( .A1(n6258), .A2(n6259), .ZN(n9857) );
  INV_X1 U8005 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9856) );
  OR2_X1 U8006 ( .A1(n9857), .A2(n9856), .ZN(n6260) );
  NAND2_X1 U8007 ( .A1(n6260), .A2(n6259), .ZN(n9878) );
  NAND2_X1 U8008 ( .A1(n6306), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6261) );
  XNOR2_X1 U8009 ( .A(n6708), .B(n7052), .ZN(n6264) );
  NAND2_X1 U8010 ( .A1(n6263), .A2(n6264), .ZN(n6704) );
  INV_X1 U8011 ( .A(n6264), .ZN(n6266) );
  NAND3_X1 U8012 ( .A1(n6488), .A2(n6266), .A3(n6265), .ZN(n6267) );
  AND2_X1 U8013 ( .A1(n6704), .A2(n6267), .ZN(n6268) );
  OR2_X1 U8014 ( .A1(n8221), .A2(n6268), .ZN(n6270) );
  AND2_X1 U8015 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8010) );
  INV_X1 U8016 ( .A(n8010), .ZN(n6269) );
  OAI211_X1 U8017 ( .C1(n8224), .C2(n6271), .A(n6270), .B(n6269), .ZN(n6272)
         );
  OR4_X1 U8018 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(P2_U3186)
         );
  XNOR2_X1 U8019 ( .A(n4514), .B(n6593), .ZN(n6281) );
  INV_X1 U8020 ( .A(n9523), .ZN(n9546) );
  OAI21_X1 U8021 ( .B1(n4514), .B2(n6277), .A(n6276), .ZN(n6745) );
  INV_X1 U8022 ( .A(n6278), .ZN(n9554) );
  NAND2_X1 U8023 ( .A1(n6745), .A2(n9554), .ZN(n6280) );
  INV_X1 U8024 ( .A(n9551), .ZN(n9530) );
  INV_X1 U8025 ( .A(n9549), .ZN(n9528) );
  AOI22_X1 U8026 ( .A1(n4416), .A2(n9530), .B1(n9528), .B2(n9171), .ZN(n6279)
         );
  OAI211_X1 U8027 ( .C1(n6281), .C2(n9546), .A(n6280), .B(n6279), .ZN(n6743)
         );
  NAND2_X1 U8028 ( .A1(n6282), .A2(n6497), .ZN(n6283) );
  OR2_X1 U8029 ( .A1(n6284), .A2(n6283), .ZN(n6286) );
  NAND2_X1 U8030 ( .A1(n6285), .A2(n9693), .ZN(n9499) );
  AND2_X2 U8031 ( .A1(n6286), .A2(n9499), .ZN(n9521) );
  MUX2_X1 U8032 ( .A(n6743), .B(P1_REG2_REG_1__SCAN_IN), .S(n9521), .Z(n6293)
         );
  OR2_X1 U8033 ( .A1(n6597), .A2(n9139), .ZN(n6499) );
  NOR2_X1 U8034 ( .A1(n9521), .A2(n6499), .ZN(n9313) );
  OAI22_X1 U8035 ( .A1(n9811), .A2(n4415), .B1(n9499), .B2(n6287), .ZN(n6292)
         );
  INV_X1 U8036 ( .A(n6745), .ZN(n6290) );
  NOR2_X1 U8037 ( .A1(n6507), .A2(n6153), .ZN(n6289) );
  NAND2_X1 U8038 ( .A1(n9502), .A2(n6289), .ZN(n9803) );
  NAND2_X1 U8039 ( .A1(n9502), .A2(n6153), .ZN(n9316) );
  INV_X1 U8040 ( .A(n9557), .ZN(n7062) );
  OAI211_X1 U8041 ( .C1(n4415), .C2(n6696), .A(n7062), .B(n6725), .ZN(n6742)
         );
  OAI22_X1 U8042 ( .A1(n6290), .A2(n9803), .B1(n9316), .B2(n6742), .ZN(n6291)
         );
  OR3_X1 U8043 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(P1_U3292) );
  XNOR2_X1 U8044 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8045 ( .A(n6294), .B(n5016), .S(P1_STATE_REG_SCAN_IN), .Z(n6295) );
  INV_X1 U8046 ( .A(n6295), .ZN(P1_U3355) );
  AND2_X1 U8047 ( .A1(n5133), .A2(P1_U3086), .ZN(n7324) );
  INV_X2 U8048 ( .A(n7324), .ZN(n9707) );
  OAI222_X1 U8049 ( .A1(P1_U3086), .A2(n6381), .B1(n9707), .B2(n6308), .C1(
        n6296), .C2(n9709), .ZN(P1_U3352) );
  OAI222_X1 U8050 ( .A1(n9709), .A2(n6297), .B1(n9707), .B2(n6309), .C1(n9215), 
        .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U8051 ( .A1(P1_U3086), .A2(n6378), .B1(n9707), .B2(n5819), .C1(
        n6298), .C2(n9709), .ZN(P1_U3354) );
  OAI222_X1 U8052 ( .A1(P1_U3086), .A2(n9189), .B1(n9707), .B2(n6305), .C1(
        n6299), .C2(n9709), .ZN(P1_U3353) );
  OR2_X1 U8053 ( .A1(n5133), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8608) );
  AND2_X1 U8054 ( .A1(n5133), .A2(P2_U3151), .ZN(n8606) );
  INV_X2 U8055 ( .A(n8606), .ZN(n8612) );
  OAI222_X1 U8056 ( .A1(n8608), .A2(n5819), .B1(n8612), .B2(n5102), .C1(
        P2_U3151), .C2(n4883), .ZN(P2_U3294) );
  INV_X1 U8057 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6300) );
  INV_X1 U8058 ( .A(n6386), .ZN(n6414) );
  OAI222_X1 U8059 ( .A1(n9709), .A2(n6300), .B1(n9707), .B2(n6303), .C1(n6414), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U8060 ( .A(n9709), .ZN(n7071) );
  AOI22_X1 U8061 ( .A1(n6424), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7071), .ZN(n6301) );
  OAI21_X1 U8062 ( .B1(n6302), .B2(n9707), .A(n6301), .ZN(P1_U3349) );
  INV_X1 U8063 ( .A(n8608), .ZN(n8609) );
  INV_X1 U8064 ( .A(n8609), .ZN(n7861) );
  OAI222_X1 U8065 ( .A1(n7861), .A2(n6302), .B1(n7003), .B2(P2_U3151), .C1(
        n4509), .C2(n8612), .ZN(P2_U3289) );
  OAI222_X1 U8066 ( .A1(n8612), .A2(n6304), .B1(n6840), .B2(P2_U3151), .C1(
        n7861), .C2(n6303), .ZN(P2_U3290) );
  OAI222_X1 U8067 ( .A1(n8612), .A2(n6307), .B1(n6306), .B2(P2_U3151), .C1(
        n7861), .C2(n6305), .ZN(P2_U3293) );
  OAI222_X1 U8068 ( .A1(n8612), .A2(n5099), .B1(n6481), .B2(P2_U3151), .C1(
        n7861), .C2(n6308), .ZN(P2_U3292) );
  OAI222_X1 U8069 ( .A1(n8612), .A2(n6310), .B1(n6708), .B2(P2_U3151), .C1(
        n7861), .C2(n6309), .ZN(P2_U3291) );
  OAI222_X1 U8070 ( .A1(n8608), .A2(n6312), .B1(n7006), .B2(P2_U3151), .C1(
        n6311), .C2(n8612), .ZN(P2_U3288) );
  INV_X1 U8071 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6313) );
  INV_X1 U8072 ( .A(n6391), .ZN(n6452) );
  OAI222_X1 U8073 ( .A1(n9709), .A2(n6313), .B1(n9707), .B2(n6312), .C1(n6452), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8074 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6315) );
  INV_X1 U8075 ( .A(n6314), .ZN(n6316) );
  INV_X1 U8076 ( .A(n7106), .ZN(n7095) );
  OAI222_X1 U8077 ( .A1(n8612), .A2(n6315), .B1(n8608), .B2(n6316), .C1(
        P2_U3151), .C2(n7095), .ZN(P2_U3287) );
  INV_X1 U8078 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6317) );
  INV_X1 U8079 ( .A(n6393), .ZN(n6441) );
  OAI222_X1 U8080 ( .A1(n6317), .A2(n9709), .B1(P1_U3086), .B2(n6441), .C1(
        n9707), .C2(n6316), .ZN(P1_U3347) );
  NAND2_X1 U8081 ( .A1(n6328), .A2(n6318), .ZN(n6355) );
  NAND3_X1 U8082 ( .A1(n7424), .A2(P2_STATE_REG_SCAN_IN), .A3(n6319), .ZN(
        n6321) );
  NOR2_X1 U8083 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  AOI21_X1 U8084 ( .B1(n6355), .B2(n6323), .A(n6322), .ZN(P2_U3376) );
  INV_X1 U8085 ( .A(n6324), .ZN(n6332) );
  AOI22_X1 U8086 ( .A1(n9245), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7071), .ZN(n6325) );
  OAI21_X1 U8087 ( .B1(n6332), .B2(n9707), .A(n6325), .ZN(P1_U3346) );
  INV_X1 U8088 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U8089 ( .A1(n6610), .A2(n6328), .ZN(n6326) );
  OAI21_X1 U8090 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(P2_U3377) );
  INV_X1 U8091 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10220) );
  OAI222_X1 U8092 ( .A1(n8608), .A2(n6334), .B1(n7380), .B2(P2_U3151), .C1(
        n10220), .C2(n8612), .ZN(P2_U3285) );
  AOI21_X1 U8093 ( .B1(n9133), .B2(n6521), .A(n6329), .ZN(n6374) );
  INV_X1 U8094 ( .A(n6374), .ZN(n6330) );
  OR2_X1 U8095 ( .A1(n6521), .A2(P1_U3086), .ZN(n9142) );
  INV_X1 U8096 ( .A(n9142), .ZN(n9140) );
  OR2_X1 U8097 ( .A1(n9140), .A2(n9693), .ZN(n6375) );
  AND2_X1 U8098 ( .A1(n6330), .A2(n6375), .ZN(n9731) );
  NOR2_X1 U8099 ( .A1(n9731), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8100 ( .A(n7113), .ZN(n7259) );
  OAI222_X1 U8101 ( .A1(n8608), .A2(n6332), .B1(n7259), .B2(P2_U3151), .C1(
        n6331), .C2(n8612), .ZN(P2_U3286) );
  INV_X1 U8102 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10257) );
  INV_X1 U8103 ( .A(n9717), .ZN(n6333) );
  OAI222_X1 U8104 ( .A1(n9709), .A2(n10257), .B1(n9707), .B2(n6334), .C1(n6333), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8105 ( .A1(n9693), .A2(n6335), .ZN(n9818) );
  INV_X1 U8106 ( .A(n9818), .ZN(n9819) );
  OAI21_X1 U8107 ( .B1(n9819), .B2(P1_D_REG_1__SCAN_IN), .A(n6336), .ZN(n6337)
         );
  OAI21_X1 U8108 ( .B1(n9693), .B2(n6338), .A(n6337), .ZN(P1_U3440) );
  INV_X1 U8109 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U8110 ( .A1(n4416), .A2(P1_U3973), .ZN(n6339) );
  OAI21_X1 U8111 ( .B1(P1_U3973), .B2(n10222), .A(n6339), .ZN(P1_U3554) );
  INV_X1 U8112 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8113 ( .A1(n6340), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6346) );
  INV_X1 U8114 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6341) );
  OR2_X1 U8115 ( .A1(n6342), .A2(n6341), .ZN(n6345) );
  INV_X1 U8116 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9654) );
  OR2_X1 U8117 ( .A1(n6343), .A2(n9654), .ZN(n6344) );
  AND3_X1 U8118 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(n9126) );
  INV_X1 U8119 ( .A(n9126), .ZN(n9299) );
  NAND2_X1 U8120 ( .A1(n9299), .A2(P1_U3973), .ZN(n6347) );
  OAI21_X1 U8121 ( .B1(P1_U3973), .B2(n6348), .A(n6347), .ZN(P1_U3585) );
  NAND2_X1 U8122 ( .A1(P1_U3973), .A2(n9057), .ZN(n6349) );
  OAI21_X1 U8123 ( .B1(P1_U3973), .B2(n5102), .A(n6349), .ZN(P1_U3555) );
  INV_X1 U8124 ( .A(n6350), .ZN(n6353) );
  AOI22_X1 U8125 ( .A1(n9743), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7071), .ZN(n6351) );
  OAI21_X1 U8126 ( .B1(n6353), .B2(n9707), .A(n6351), .ZN(P1_U3344) );
  AOI22_X1 U8127 ( .A1(n9754), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7071), .ZN(n6352) );
  OAI21_X1 U8128 ( .B1(n6366), .B2(n9707), .A(n6352), .ZN(P1_U3343) );
  INV_X1 U8129 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6354) );
  OAI222_X1 U8130 ( .A1(n8612), .A2(n6354), .B1(n8608), .B2(n6353), .C1(
        P2_U3151), .C2(n7476), .ZN(P2_U3284) );
  INV_X1 U8131 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6356) );
  NOR2_X1 U8132 ( .A1(n6463), .A2(n6356), .ZN(P2_U3249) );
  INV_X1 U8133 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U8134 ( .A1(n6463), .A2(n10106), .ZN(P2_U3246) );
  INV_X1 U8135 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6357) );
  NOR2_X1 U8136 ( .A1(n6463), .A2(n6357), .ZN(P2_U3252) );
  INV_X1 U8137 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6358) );
  NOR2_X1 U8138 ( .A1(n6463), .A2(n6358), .ZN(P2_U3253) );
  INV_X1 U8139 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U8140 ( .A1(n6463), .A2(n10267), .ZN(P2_U3254) );
  INV_X1 U8141 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U8142 ( .A1(n6463), .A2(n6359), .ZN(P2_U3255) );
  INV_X1 U8143 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6360) );
  NOR2_X1 U8144 ( .A1(n6463), .A2(n6360), .ZN(P2_U3256) );
  INV_X1 U8145 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6361) );
  NOR2_X1 U8146 ( .A1(n6463), .A2(n6361), .ZN(P2_U3247) );
  INV_X1 U8147 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6362) );
  NOR2_X1 U8148 ( .A1(n6463), .A2(n6362), .ZN(P2_U3250) );
  INV_X1 U8149 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6363) );
  NOR2_X1 U8150 ( .A1(n6463), .A2(n6363), .ZN(P2_U3251) );
  INV_X1 U8151 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U8152 ( .A1(n6463), .A2(n10184), .ZN(P2_U3248) );
  INV_X1 U8153 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6364) );
  NOR2_X1 U8154 ( .A1(n6463), .A2(n6364), .ZN(P2_U3257) );
  INV_X1 U8155 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6365) );
  OAI222_X1 U8156 ( .A1(n8608), .A2(n6366), .B1(n7495), .B2(P2_U3151), .C1(
        n6365), .C2(n8612), .ZN(P2_U3283) );
  NOR2_X1 U8157 ( .A1(n9245), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6367) );
  AOI21_X1 U8158 ( .B1(n9245), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6367), .ZN(
        n6373) );
  INV_X1 U8159 ( .A(n9215), .ZN(n6371) );
  MUX2_X1 U8160 ( .A(n6369), .B(P1_REG2_REG_2__SCAN_IN), .S(n9189), .Z(n9196)
         );
  INV_X1 U8161 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6368) );
  AND2_X1 U8162 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9185) );
  OAI21_X1 U8163 ( .B1(n6368), .B2(n6378), .A(n9172), .ZN(n9195) );
  NAND2_X1 U8164 ( .A1(n9196), .A2(n9195), .ZN(n9194) );
  OAI21_X1 U8165 ( .B1(n9189), .B2(n6369), .A(n9194), .ZN(n9204) );
  XNOR2_X1 U8166 ( .A(n6381), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U8167 ( .A1(n9204), .A2(n9205), .ZN(n9203) );
  OAI21_X1 U8168 ( .B1(n6381), .B2(n6370), .A(n9203), .ZN(n9219) );
  XNOR2_X1 U8169 ( .A(n9215), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U8170 ( .A1(n9219), .A2(n9220), .ZN(n9218) );
  XNOR2_X1 U8171 ( .A(n6386), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6406) );
  XNOR2_X1 U8172 ( .A(n6424), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6418) );
  NOR2_X1 U8173 ( .A1(n6419), .A2(n6418), .ZN(n6417) );
  XNOR2_X1 U8174 ( .A(n6391), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6445) );
  XNOR2_X1 U8175 ( .A(n6393), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6433) );
  AOI21_X1 U8176 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6393), .A(n6432), .ZN(
        n6372) );
  NAND2_X1 U8177 ( .A1(n6372), .A2(n6373), .ZN(n9244) );
  OAI21_X1 U8178 ( .B1(n6373), .B2(n6372), .A(n9244), .ZN(n6402) );
  NAND2_X1 U8179 ( .A1(n6375), .A2(n6374), .ZN(n9734) );
  NOR2_X1 U8180 ( .A1(n9734), .A2(n9183), .ZN(n9291) );
  NAND2_X1 U8181 ( .A1(n9291), .A2(n9186), .ZN(n10323) );
  INV_X1 U8182 ( .A(n10323), .ZN(n9755) );
  MUX2_X1 U8183 ( .A(n5926), .B(P1_REG1_REG_9__SCAN_IN), .S(n9245), .Z(n6397)
         );
  INV_X1 U8184 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6376) );
  MUX2_X1 U8185 ( .A(n6376), .B(P1_REG1_REG_2__SCAN_IN), .S(n9189), .Z(n9199)
         );
  INV_X1 U8186 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6377) );
  MUX2_X1 U8187 ( .A(n6377), .B(P1_REG1_REG_1__SCAN_IN), .S(n6378), .Z(n9176)
         );
  AND2_X1 U8188 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9175) );
  NAND2_X1 U8189 ( .A1(n9176), .A2(n9175), .ZN(n9174) );
  INV_X1 U8190 ( .A(n6378), .ZN(n9177) );
  NAND2_X1 U8191 ( .A1(n9177), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8192 ( .A1(n9174), .A2(n6379), .ZN(n9198) );
  NAND2_X1 U8193 ( .A1(n9199), .A2(n9198), .ZN(n9197) );
  OR2_X1 U8194 ( .A1(n9189), .A2(n6376), .ZN(n6380) );
  NAND2_X1 U8195 ( .A1(n9197), .A2(n6380), .ZN(n9208) );
  XNOR2_X1 U8196 ( .A(n6381), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U8197 ( .A1(n9208), .A2(n9209), .ZN(n9207) );
  INV_X1 U8198 ( .A(n6381), .ZN(n9210) );
  NAND2_X1 U8199 ( .A1(n9210), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8200 ( .A1(n9207), .A2(n6382), .ZN(n9222) );
  XNOR2_X1 U8201 ( .A(n9215), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U8202 ( .A1(n9222), .A2(n9223), .ZN(n9221) );
  INV_X1 U8203 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6383) );
  OR2_X1 U8204 ( .A1(n9215), .A2(n6383), .ZN(n6384) );
  NAND2_X1 U8205 ( .A1(n9221), .A2(n6384), .ZN(n6409) );
  XNOR2_X1 U8206 ( .A(n6386), .B(n6385), .ZN(n6410) );
  NAND2_X1 U8207 ( .A1(n6409), .A2(n6410), .ZN(n6408) );
  NAND2_X1 U8208 ( .A1(n6386), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8209 ( .A1(n6408), .A2(n6387), .ZN(n6421) );
  INV_X1 U8210 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U8211 ( .A(n6424), .B(n6388), .ZN(n6422) );
  NAND2_X1 U8212 ( .A1(n6421), .A2(n6422), .ZN(n6420) );
  NAND2_X1 U8213 ( .A1(n6424), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8214 ( .A1(n6420), .A2(n6389), .ZN(n6448) );
  INV_X1 U8215 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6390) );
  XNOR2_X1 U8216 ( .A(n6391), .B(n6390), .ZN(n6449) );
  NAND2_X1 U8217 ( .A1(n6448), .A2(n6449), .ZN(n6447) );
  NAND2_X1 U8218 ( .A1(n6391), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8219 ( .A1(n6447), .A2(n6392), .ZN(n6436) );
  INV_X1 U8220 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9840) );
  MUX2_X1 U8221 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9840), .S(n6393), .Z(n6437)
         );
  NAND2_X1 U8222 ( .A1(n6436), .A2(n6437), .ZN(n6435) );
  NAND2_X1 U8223 ( .A1(n6393), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8224 ( .A1(n6435), .A2(n6394), .ZN(n6396) );
  INV_X1 U8225 ( .A(n9233), .ZN(n6395) );
  AOI21_X1 U8226 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6400) );
  OR2_X1 U8227 ( .A1(n9734), .A2(n9729), .ZN(n10319) );
  AND2_X1 U8228 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7302) );
  AOI21_X1 U8229 ( .B1(n9731), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7302), .ZN(
        n6399) );
  OR2_X1 U8230 ( .A1(n9734), .A2(n9186), .ZN(n9769) );
  INV_X1 U8231 ( .A(n9769), .ZN(n10329) );
  NAND2_X1 U8232 ( .A1(n10329), .A2(n9245), .ZN(n6398) );
  OAI211_X1 U8233 ( .C1(n6400), .C2(n10319), .A(n6399), .B(n6398), .ZN(n6401)
         );
  AOI21_X1 U8234 ( .B1(n6402), .B2(n9755), .A(n6401), .ZN(n6403) );
  INV_X1 U8235 ( .A(n6403), .ZN(P1_U3252) );
  NAND2_X1 U8236 ( .A1(n6987), .A2(P2_U3893), .ZN(n6404) );
  OAI21_X1 U8237 ( .B1(P2_U3893), .B2(n5827), .A(n6404), .ZN(P2_U3491) );
  AOI211_X1 U8238 ( .C1(n6407), .C2(n6406), .A(n6405), .B(n10323), .ZN(n6416)
         );
  INV_X1 U8239 ( .A(n10319), .ZN(n9764) );
  OAI211_X1 U8240 ( .C1(n6410), .C2(n6409), .A(n9764), .B(n6408), .ZN(n6413)
         );
  NAND2_X1 U8241 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n8802) );
  INV_X1 U8242 ( .A(n8802), .ZN(n6411) );
  AOI21_X1 U8243 ( .B1(n9731), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6411), .ZN(
        n6412) );
  OAI211_X1 U8244 ( .C1(n9769), .C2(n6414), .A(n6413), .B(n6412), .ZN(n6415)
         );
  OR2_X1 U8245 ( .A1(n6416), .A2(n6415), .ZN(P1_U3248) );
  AOI211_X1 U8246 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n10323), .ZN(n6430)
         );
  OAI211_X1 U8247 ( .C1(n6422), .C2(n6421), .A(n9764), .B(n6420), .ZN(n6428)
         );
  INV_X1 U8248 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6423) );
  NOR2_X1 U8249 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6423), .ZN(n6835) );
  INV_X1 U8250 ( .A(n6835), .ZN(n6427) );
  NAND2_X1 U8251 ( .A1(n10329), .A2(n6424), .ZN(n6426) );
  NAND2_X1 U8252 ( .A1(n9731), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6425) );
  NAND4_X1 U8253 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6425), .ZN(n6429)
         );
  OR2_X1 U8254 ( .A1(n6430), .A2(n6429), .ZN(P1_U3249) );
  INV_X1 U8255 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8256 ( .A1(n8395), .A2(P2_U3893), .ZN(n6431) );
  OAI21_X1 U8257 ( .B1(P2_U3893), .B2(n6457), .A(n6431), .ZN(P2_U3504) );
  AOI211_X1 U8258 ( .C1(n6434), .C2(n6433), .A(n10323), .B(n6432), .ZN(n6443)
         );
  OAI211_X1 U8259 ( .C1(n6437), .C2(n6436), .A(n9764), .B(n6435), .ZN(n6440)
         );
  NAND2_X1 U8260 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7189) );
  INV_X1 U8261 ( .A(n7189), .ZN(n6438) );
  AOI21_X1 U8262 ( .B1(n9731), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6438), .ZN(
        n6439) );
  OAI211_X1 U8263 ( .C1(n6441), .C2(n9769), .A(n6440), .B(n6439), .ZN(n6442)
         );
  OR2_X1 U8264 ( .A1(n6443), .A2(n6442), .ZN(P1_U3251) );
  AOI211_X1 U8265 ( .C1(n6446), .C2(n6445), .A(n10323), .B(n6444), .ZN(n6454)
         );
  OAI211_X1 U8266 ( .C1(n6449), .C2(n6448), .A(n9764), .B(n6447), .ZN(n6451)
         );
  AND2_X1 U8267 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8621) );
  AOI21_X1 U8268 ( .B1(n9731), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n8621), .ZN(
        n6450) );
  OAI211_X1 U8269 ( .C1(n9769), .C2(n6452), .A(n6451), .B(n6450), .ZN(n6453)
         );
  OR2_X1 U8270 ( .A1(n6454), .A2(n6453), .ZN(P1_U3250) );
  INV_X1 U8271 ( .A(n8097), .ZN(n7504) );
  INV_X1 U8272 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6455) );
  OAI222_X1 U8273 ( .A1(n8608), .A2(n6456), .B1(n7504), .B2(P2_U3151), .C1(
        n6455), .C2(n8612), .ZN(P2_U3282) );
  INV_X1 U8274 ( .A(n9248), .ZN(n9768) );
  OAI222_X1 U8275 ( .A1(P1_U3086), .A2(n9768), .B1(n9709), .B2(n6457), .C1(
        n6456), .C2(n9707), .ZN(P1_U3342) );
  MUX2_X1 U8276 ( .A(n6458), .B(n7427), .S(P2_U3893), .Z(n6459) );
  INV_X1 U8277 ( .A(n6459), .ZN(P2_U3500) );
  NAND2_X1 U8278 ( .A1(n8185), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6460) );
  OAI21_X1 U8279 ( .B1(n8320), .B2(n8185), .A(n6460), .ZN(P2_U3512) );
  INV_X1 U8280 ( .A(n6461), .ZN(n6494) );
  AOI22_X1 U8281 ( .A1(n9784), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7071), .ZN(n6462) );
  OAI21_X1 U8282 ( .B1(n6494), .B2(n9707), .A(n6462), .ZN(P1_U3341) );
  INV_X1 U8283 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U8284 ( .A1(n6463), .A2(n6464), .ZN(P2_U3260) );
  INV_X1 U8285 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U8286 ( .A1(n6463), .A2(n6465), .ZN(P2_U3258) );
  INV_X1 U8287 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U8288 ( .A1(n6463), .A2(n6466), .ZN(P2_U3234) );
  INV_X1 U8289 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U8290 ( .A1(n6463), .A2(n10207), .ZN(P2_U3263) );
  INV_X1 U8291 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6467) );
  NOR2_X1 U8292 ( .A1(n6463), .A2(n6467), .ZN(P2_U3259) );
  INV_X1 U8293 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U8294 ( .A1(n6463), .A2(n6468), .ZN(P2_U3261) );
  INV_X1 U8295 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U8296 ( .A1(n6463), .A2(n6469), .ZN(P2_U3245) );
  INV_X1 U8297 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10108) );
  NOR2_X1 U8298 ( .A1(n6463), .A2(n10108), .ZN(P2_U3243) );
  INV_X1 U8299 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U8300 ( .A1(n6463), .A2(n6470), .ZN(P2_U3242) );
  INV_X1 U8301 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U8302 ( .A1(n6463), .A2(n6471), .ZN(P2_U3241) );
  INV_X1 U8303 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U8304 ( .A1(n6463), .A2(n10110), .ZN(P2_U3262) );
  INV_X1 U8305 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U8306 ( .A1(n6463), .A2(n6472), .ZN(P2_U3239) );
  INV_X1 U8307 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10254) );
  NOR2_X1 U8308 ( .A1(n6463), .A2(n10254), .ZN(P2_U3238) );
  INV_X1 U8309 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8310 ( .A1(n6463), .A2(n6473), .ZN(P2_U3237) );
  INV_X1 U8311 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10139) );
  NOR2_X1 U8312 ( .A1(n6463), .A2(n10139), .ZN(P2_U3236) );
  INV_X1 U8313 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6474) );
  NOR2_X1 U8314 ( .A1(n6463), .A2(n6474), .ZN(P2_U3235) );
  INV_X1 U8315 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6475) );
  NOR2_X1 U8316 ( .A1(n6463), .A2(n6475), .ZN(P2_U3240) );
  INV_X1 U8317 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6476) );
  NOR2_X1 U8318 ( .A1(n6463), .A2(n6476), .ZN(P2_U3244) );
  INV_X1 U8319 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U8320 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6480) );
  NAND2_X1 U8321 ( .A1(n6480), .A2(n9872), .ZN(n6492) );
  INV_X1 U8322 ( .A(n6482), .ZN(n6483) );
  AOI21_X1 U8323 ( .B1(n6224), .B2(n6484), .A(n6483), .ZN(n6485) );
  OAI22_X1 U8324 ( .A1(n8224), .A2(n6485), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6772), .ZN(n6490) );
  NAND2_X1 U8325 ( .A1(n6486), .A2(n6225), .ZN(n6487) );
  AOI21_X1 U8326 ( .B1(n6488), .B2(n6487), .A(n8221), .ZN(n6489) );
  AOI211_X1 U8327 ( .C1(n4613), .C2(n9881), .A(n6490), .B(n6489), .ZN(n6491)
         );
  OAI211_X1 U8328 ( .C1(n9887), .C2(n6493), .A(n6492), .B(n6491), .ZN(P2_U3185) );
  INV_X1 U8329 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6495) );
  OAI222_X1 U8330 ( .A1(n8612), .A2(n6495), .B1(n8608), .B2(n6494), .C1(
        P2_U3151), .C2(n8111), .ZN(P2_U3281) );
  OR2_X1 U8331 ( .A1(n6497), .A2(n6496), .ZN(n6517) );
  OR2_X1 U8332 ( .A1(n6498), .A2(n6517), .ZN(n6514) );
  OR2_X1 U8333 ( .A1(n6514), .A2(n6499), .ZN(n6500) );
  NAND2_X1 U8334 ( .A1(n6500), .A2(n9499), .ZN(n8897) );
  INV_X1 U8335 ( .A(n8897), .ZN(n8782) );
  NAND2_X1 U8336 ( .A1(n6507), .A2(n6501), .ZN(n6502) );
  NAND2_X1 U8337 ( .A1(n6509), .A2(n6502), .ZN(n6503) );
  INV_X2 U8338 ( .A(n6532), .ZN(n8740) );
  INV_X4 U8339 ( .A(n8651), .ZN(n8736) );
  NAND2_X1 U8340 ( .A1(n6510), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6504) );
  AND2_X1 U8341 ( .A1(n6507), .A2(n6520), .ZN(n6508) );
  NAND2_X1 U8342 ( .A1(n6509), .A2(n6508), .ZN(n6530) );
  AOI21_X1 U8343 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n6510), .A(n6536), .ZN(
        n6511) );
  NOR2_X1 U8344 ( .A1(n6512), .A2(n6511), .ZN(n6538) );
  AOI21_X1 U8345 ( .B1(n6512), .B2(n6511), .A(n6538), .ZN(n9182) );
  NAND2_X1 U8346 ( .A1(n9833), .A2(n6729), .ZN(n6513) );
  NAND2_X1 U8347 ( .A1(n9182), .A2(n5036), .ZN(n6526) );
  INV_X1 U8348 ( .A(n6515), .ZN(n6516) );
  NOR2_X1 U8349 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND3_X1 U8350 ( .A1(n6689), .A2(n9693), .A3(n6518), .ZN(n6562) );
  OR2_X1 U8351 ( .A1(n6562), .A2(n9186), .ZN(n8890) );
  INV_X1 U8352 ( .A(n8890), .ZN(n8861) );
  AND2_X1 U8353 ( .A1(n9137), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7070) );
  INV_X1 U8354 ( .A(n6518), .ZN(n6519) );
  OAI21_X1 U8355 ( .B1(n9833), .B2(n7070), .A(n6519), .ZN(n6524) );
  AND3_X1 U8356 ( .A1(n6522), .A2(n6521), .A3(n6520), .ZN(n6523) );
  NAND2_X1 U8357 ( .A1(n6524), .A2(n6523), .ZN(n6563) );
  OR2_X1 U8358 ( .A1(n6563), .A2(P1_U3086), .ZN(n6576) );
  AOI22_X1 U8359 ( .A1(n8861), .A2(n9057), .B1(n6576), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6525) );
  OAI211_X1 U8360 ( .C1(n8782), .C2(n6696), .A(n6526), .B(n6525), .ZN(P1_U3232) );
  INV_X2 U8361 ( .A(n6527), .ZN(n8645) );
  NAND2_X1 U8362 ( .A1(n8645), .A2(n5846), .ZN(n6529) );
  NAND2_X1 U8363 ( .A1(n9171), .A2(n8736), .ZN(n6528) );
  NAND2_X1 U8364 ( .A1(n6529), .A2(n6528), .ZN(n6531) );
  INV_X2 U8365 ( .A(n6530), .ZN(n8678) );
  INV_X4 U8366 ( .A(n8678), .ZN(n8674) );
  XNOR2_X1 U8367 ( .A(n6531), .B(n8674), .ZN(n6534) );
  OAI22_X1 U8368 ( .A1(n5847), .A2(n8680), .B1(n5848), .B2(n8651), .ZN(n6533)
         );
  AOI22_X1 U8369 ( .A1(n8645), .A2(n6890), .B1(n8736), .B2(n9057), .ZN(n6539)
         );
  XNOR2_X1 U8370 ( .A(n6539), .B(n8674), .ZN(n6572) );
  OAI21_X1 U8371 ( .B1(n5044), .B2(n6540), .A(n6550), .ZN(n6541) );
  NAND2_X1 U8372 ( .A1(n6541), .A2(n5036), .ZN(n6544) );
  OAI22_X1 U8373 ( .A1(n6594), .A2(n9551), .B1(n6552), .B2(n9186), .ZN(n6728)
         );
  INV_X1 U8374 ( .A(n6562), .ZN(n6542) );
  AOI22_X1 U8375 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n6576), .B1(n6728), .B2(
        n6542), .ZN(n6543) );
  OAI211_X1 U8376 ( .C1(n5848), .C2(n8782), .A(n6544), .B(n6543), .ZN(P1_U3237) );
  INV_X1 U8377 ( .A(n6545), .ZN(n6547) );
  AOI22_X1 U8378 ( .A1(n8138), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8606), .ZN(n6546) );
  OAI21_X1 U8379 ( .B1(n6547), .B2(n7861), .A(n6546), .ZN(P2_U3280) );
  INV_X1 U8380 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6548) );
  INV_X1 U8381 ( .A(n10328), .ZN(n9250) );
  OAI222_X1 U8382 ( .A1(n9709), .A2(n6548), .B1(n9707), .B2(n6547), .C1(
        P1_U3086), .C2(n9250), .ZN(P1_U3340) );
  NAND2_X1 U8383 ( .A1(n6550), .A2(n6549), .ZN(n6584) );
  AOI22_X1 U8384 ( .A1(n8645), .A2(n6866), .B1(n8741), .B2(n9170), .ZN(n6551)
         );
  XNOR2_X1 U8385 ( .A(n6551), .B(n8674), .ZN(n6557) );
  OAI22_X1 U8386 ( .A1(n6552), .A2(n8680), .B1(n6807), .B2(n8651), .ZN(n6555)
         );
  XNOR2_X1 U8387 ( .A(n6557), .B(n6555), .ZN(n6585) );
  NAND2_X1 U8388 ( .A1(n6584), .A2(n6585), .ZN(n6559) );
  NOR2_X1 U8389 ( .A1(n6884), .A2(n8651), .ZN(n6553) );
  AOI21_X1 U8390 ( .B1(n8740), .B2(n9169), .A(n6553), .ZN(n6811) );
  AOI22_X1 U8391 ( .A1(n8645), .A2(n6875), .B1(n8741), .B2(n9169), .ZN(n6554)
         );
  INV_X1 U8392 ( .A(n6555), .ZN(n6556) );
  NAND2_X1 U8393 ( .A1(n6557), .A2(n6556), .ZN(n6561) );
  NAND2_X1 U8394 ( .A1(n6815), .A2(n5036), .ZN(n6569) );
  AOI21_X1 U8395 ( .B1(n6583), .B2(n6561), .A(n6560), .ZN(n6568) );
  OR2_X1 U8396 ( .A1(n6562), .A2(n9551), .ZN(n8891) );
  INV_X1 U8397 ( .A(n8891), .ZN(n8801) );
  AND2_X1 U8398 ( .A1(n6563), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8800) );
  INV_X1 U8399 ( .A(n6564), .ZN(n6876) );
  AOI22_X1 U8400 ( .A1(n8801), .A2(n9170), .B1(n8800), .B2(n6876), .ZN(n6567)
         );
  INV_X1 U8401 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U8402 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10120), .ZN(n9217) );
  NOR2_X1 U8403 ( .A1(n8890), .A2(n6799), .ZN(n6565) );
  AOI211_X1 U8404 ( .C1(n6875), .C2(n8897), .A(n9217), .B(n6565), .ZN(n6566)
         );
  OAI211_X1 U8405 ( .C1(n6569), .C2(n6568), .A(n6567), .B(n6566), .ZN(P1_U3230) );
  XNOR2_X1 U8406 ( .A(n6570), .B(n6571), .ZN(n6573) );
  XNOR2_X1 U8407 ( .A(n6573), .B(n6572), .ZN(n6578) );
  OAI22_X1 U8408 ( .A1(n5847), .A2(n8890), .B1(n8891), .B2(n6591), .ZN(n6575)
         );
  NOR2_X1 U8409 ( .A1(n8782), .A2(n4415), .ZN(n6574) );
  AOI211_X1 U8410 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6576), .A(n6575), .B(
        n6574), .ZN(n6577) );
  OAI21_X1 U8411 ( .B1(n6578), .B2(n8899), .A(n6577), .ZN(P1_U3222) );
  NOR2_X1 U8412 ( .A1(n5197), .A2(n9909), .ZN(n6605) );
  INV_X1 U8413 ( .A(n9966), .ZN(n9967) );
  INV_X1 U8414 ( .A(n8413), .ZN(n9907) );
  NAND2_X1 U8415 ( .A1(n6987), .A2(n6580), .ZN(n7600) );
  AND2_X1 U8416 ( .A1(n6629), .A2(n7600), .ZN(n7757) );
  AOI21_X1 U8417 ( .B1(n9967), .B2(n9907), .A(n7757), .ZN(n6581) );
  AOI211_X1 U8418 ( .C1(n9972), .C2(n7758), .A(n6605), .B(n6581), .ZN(n9916)
         );
  NAND2_X1 U8419 ( .A1(n9990), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6582) );
  OAI21_X1 U8420 ( .B1(n9916), .B2(n9990), .A(n6582), .ZN(P2_U3459) );
  OAI21_X1 U8421 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(n6589) );
  INV_X1 U8422 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U8423 ( .A1(n8801), .A2(n9171), .B1(n8800), .B2(n6867), .ZN(n6587)
         );
  AND2_X1 U8424 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9206) );
  AOI21_X1 U8425 ( .B1(n8861), .B2(n9169), .A(n9206), .ZN(n6586) );
  OAI211_X1 U8426 ( .C1(n6807), .C2(n8782), .A(n6587), .B(n6586), .ZN(n6588)
         );
  AOI21_X1 U8427 ( .B1(n6589), .B2(n5036), .A(n6588), .ZN(n6590) );
  INV_X1 U8428 ( .A(n6590), .ZN(P1_U3218) );
  OR2_X1 U8429 ( .A1(n6591), .A2(n5829), .ZN(n9059) );
  INV_X1 U8430 ( .A(n9059), .ZN(n6592) );
  OR2_X1 U8431 ( .A1(n6593), .A2(n6592), .ZN(n9012) );
  OAI21_X1 U8432 ( .B1(n9836), .B2(n9523), .A(n9012), .ZN(n6596) );
  NOR2_X1 U8433 ( .A1(n6594), .A2(n9549), .ZN(n6693) );
  INV_X1 U8434 ( .A(n6693), .ZN(n6595) );
  OAI211_X1 U8435 ( .C1(n6597), .C2(n6696), .A(n6596), .B(n6595), .ZN(n6668)
         );
  NAND2_X1 U8436 ( .A1(n9691), .A2(n6668), .ZN(n6598) );
  OAI21_X1 U8437 ( .B1(n9691), .B2(n5823), .A(n6598), .ZN(P1_U3453) );
  INV_X1 U8438 ( .A(n6599), .ZN(n6617) );
  INV_X1 U8439 ( .A(n8141), .ZN(n8155) );
  OAI222_X1 U8440 ( .A1(n8608), .A2(n6617), .B1(n8155), .B2(P2_U3151), .C1(
        n6600), .C2(n8612), .ZN(P2_U3279) );
  INV_X1 U8441 ( .A(n6601), .ZN(n6602) );
  INV_X1 U8442 ( .A(n9898), .ZN(n8389) );
  NOR2_X1 U8443 ( .A1(n7757), .A2(n6603), .ZN(n6604) );
  AOI211_X1 U8444 ( .C1(n8389), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6605), .B(
        n6604), .ZN(n6616) );
  INV_X1 U8445 ( .A(n6606), .ZN(n6609) );
  INV_X1 U8446 ( .A(n6607), .ZN(n6608) );
  MUX2_X1 U8447 ( .A(n6610), .B(n6609), .S(n6608), .Z(n6611) );
  NAND2_X1 U8448 ( .A1(n6612), .A2(n6611), .ZN(n6613) );
  INV_X2 U8449 ( .A(n9913), .ZN(n8421) );
  INV_X1 U8450 ( .A(n6613), .ZN(n6614) );
  INV_X1 U8451 ( .A(n9899), .ZN(n8416) );
  NAND2_X1 U8452 ( .A1(n6614), .A2(n8416), .ZN(n8352) );
  AOI22_X1 U8453 ( .A1(n8445), .A2(n7758), .B1(n8421), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6615) );
  OAI21_X1 U8454 ( .B1(n6616), .B2(n8421), .A(n6615), .ZN(P2_U3233) );
  OAI222_X1 U8455 ( .A1(P1_U3086), .A2(n9258), .B1(n9707), .B2(n6617), .C1(
        n10228), .C2(n9709), .ZN(P1_U3339) );
  OR2_X1 U8456 ( .A1(n6656), .A2(n6618), .ZN(n6621) );
  INV_X1 U8457 ( .A(n6619), .ZN(n6640) );
  NAND2_X1 U8458 ( .A1(n6651), .A2(n6640), .ZN(n6620) );
  XNOR2_X1 U8459 ( .A(n7748), .B(n7151), .ZN(n6622) );
  AND2_X1 U8460 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  NAND2_X1 U8461 ( .A1(n6625), .A2(n6624), .ZN(n6627) );
  INV_X1 U8462 ( .A(n6626), .ZN(n7745) );
  XNOR2_X1 U8463 ( .A(n6677), .B(n5229), .ZN(n6676) );
  OR2_X1 U8464 ( .A1(n7758), .A2(n6674), .ZN(n6628) );
  NAND2_X1 U8465 ( .A1(n6629), .A2(n6628), .ZN(n6662) );
  XNOR2_X1 U8466 ( .A(n6631), .B(n8086), .ZN(n6663) );
  NAND2_X1 U8467 ( .A1(n6662), .A2(n6663), .ZN(n6634) );
  INV_X1 U8468 ( .A(n6631), .ZN(n6632) );
  OR2_X1 U8469 ( .A1(n8086), .A2(n6632), .ZN(n6633) );
  NAND2_X1 U8470 ( .A1(n6634), .A2(n6633), .ZN(n6675) );
  XOR2_X1 U8471 ( .A(n6676), .B(n6675), .Z(n6661) );
  INV_X1 U8472 ( .A(n6635), .ZN(n6642) );
  NOR2_X1 U8473 ( .A1(n6636), .A2(n7328), .ZN(n6637) );
  NAND2_X1 U8474 ( .A1(n6638), .A2(n6637), .ZN(n6639) );
  AOI21_X1 U8475 ( .B1(n6646), .B2(n6640), .A(n6639), .ZN(n6641) );
  OAI21_X1 U8476 ( .B1(n6643), .B2(n6642), .A(n6641), .ZN(n6644) );
  NAND2_X1 U8477 ( .A1(n6644), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6648) );
  NOR2_X1 U8478 ( .A1(n6645), .A2(n6649), .ZN(n7751) );
  NAND2_X1 U8479 ( .A1(n6646), .A2(n7751), .ZN(n6647) );
  NAND2_X1 U8480 ( .A1(n6648), .A2(n6647), .ZN(n8066) );
  INV_X1 U8481 ( .A(n8066), .ZN(n8040) );
  NAND2_X1 U8482 ( .A1(n8040), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7760) );
  INV_X1 U8483 ( .A(n6649), .ZN(n6650) );
  AND2_X1 U8484 ( .A1(n6651), .A2(n6650), .ZN(n6655) );
  INV_X1 U8485 ( .A(n6655), .ZN(n6653) );
  INV_X1 U8486 ( .A(n6652), .ZN(n6654) );
  OR2_X1 U8487 ( .A1(n6656), .A2(n9961), .ZN(n6657) );
  NAND2_X1 U8488 ( .A1(n6657), .A2(n9898), .ZN(n8042) );
  AOI22_X1 U8489 ( .A1(n8061), .A2(n8086), .B1(n8042), .B2(n5226), .ZN(n6658)
         );
  OAI21_X1 U8490 ( .B1(n9908), .B2(n8063), .A(n6658), .ZN(n6659) );
  AOI21_X1 U8491 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7760), .A(n6659), .ZN(
        n6660) );
  OAI21_X1 U8492 ( .B1(n8056), .B2(n6661), .A(n6660), .ZN(P2_U3177) );
  XOR2_X1 U8493 ( .A(n6663), .B(n6662), .Z(n6667) );
  AOI22_X1 U8494 ( .A1(n8061), .A2(n6987), .B1(n8042), .B2(n5196), .ZN(n6664)
         );
  OAI21_X1 U8495 ( .B1(n5227), .B2(n8063), .A(n6664), .ZN(n6665) );
  AOI21_X1 U8496 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7760), .A(n6665), .ZN(
        n6666) );
  OAI21_X1 U8497 ( .B1(n8056), .B2(n6667), .A(n6666), .ZN(P2_U3162) );
  INV_X1 U8498 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U8499 ( .A1(n9845), .A2(n6668), .ZN(n6669) );
  OAI21_X1 U8500 ( .B1(n9845), .B2(n9727), .A(n6669), .ZN(P1_U3522) );
  INV_X1 U8501 ( .A(n6670), .ZN(n6672) );
  INV_X1 U8502 ( .A(n9288), .ZN(n9277) );
  OAI222_X1 U8503 ( .A1(n9709), .A2(n6671), .B1(n9707), .B2(n6672), .C1(
        P1_U3086), .C2(n9277), .ZN(P1_U3338) );
  INV_X1 U8504 ( .A(n8191), .ZN(n8154) );
  OAI222_X1 U8505 ( .A1(n8612), .A2(n6673), .B1(n8608), .B2(n6672), .C1(
        P2_U3151), .C2(n8154), .ZN(P2_U3278) );
  XNOR2_X1 U8506 ( .A(n9927), .B(n4414), .ZN(n6896) );
  XNOR2_X1 U8507 ( .A(n9908), .B(n6896), .ZN(n6684) );
  INV_X1 U8508 ( .A(n6677), .ZN(n6678) );
  OR2_X1 U8509 ( .A1(n6678), .A2(n5229), .ZN(n6679) );
  INV_X1 U8510 ( .A(n6680), .ZN(n6682) );
  NAND2_X1 U8511 ( .A1(n6682), .A2(n6681), .ZN(n6898) );
  INV_X1 U8512 ( .A(n6898), .ZN(n6683) );
  AOI211_X1 U8513 ( .C1(n6684), .C2(n6680), .A(n8056), .B(n6683), .ZN(n6688)
         );
  MUX2_X1 U8514 ( .A(P2_STATE_REG_SCAN_IN), .B(n8040), .S(n6772), .Z(n6686) );
  AOI22_X1 U8515 ( .A1(n8061), .A2(n5229), .B1(n8042), .B2(n5245), .ZN(n6685)
         );
  OAI211_X1 U8516 ( .C1(n6901), .C2(n8063), .A(n6686), .B(n6685), .ZN(n6687)
         );
  OR2_X1 U8517 ( .A1(n6688), .A2(n6687), .ZN(P2_U3158) );
  INV_X2 U8518 ( .A(n9316), .ZN(n9805) );
  AOI21_X1 U8519 ( .B1(n9805), .B2(n7062), .A(n9313), .ZN(n6697) );
  INV_X1 U8520 ( .A(n9499), .ZN(n9807) );
  INV_X1 U8521 ( .A(n9012), .ZN(n6691) );
  NOR3_X1 U8522 ( .A1(n6691), .A2(n6690), .A3(n6689), .ZN(n6692) );
  AOI211_X1 U8523 ( .C1(n9807), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6693), .B(
        n6692), .ZN(n6694) );
  MUX2_X1 U8524 ( .A(n10051), .B(n6694), .S(n9502), .Z(n6695) );
  OAI21_X1 U8525 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(P1_U3293) );
  INV_X1 U8526 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U8527 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8208), .Z(n6841) );
  XNOR2_X1 U8528 ( .A(n6841), .B(n6840), .ZN(n6701) );
  AOI211_X1 U8529 ( .C1(n6701), .C2(n6700), .A(n9848), .B(n6839), .ZN(n6702)
         );
  INV_X1 U8530 ( .A(n6702), .ZN(n6721) );
  INV_X1 U8531 ( .A(n6840), .ZN(n6719) );
  NAND2_X1 U8532 ( .A1(n6708), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8533 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  INV_X1 U8534 ( .A(n6856), .ZN(n6706) );
  AOI21_X1 U8535 ( .B1(n5266), .B2(n6707), .A(n6706), .ZN(n6717) );
  NAND2_X1 U8536 ( .A1(n6708), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8537 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  NAND2_X1 U8538 ( .A1(n6711), .A2(n6840), .ZN(n6846) );
  OAI21_X1 U8539 ( .B1(n6711), .B2(n6840), .A(n6846), .ZN(n6712) );
  INV_X1 U8540 ( .A(n6850), .ZN(n6714) );
  AND2_X1 U8541 ( .A1(n6712), .A2(n5263), .ZN(n6713) );
  INV_X1 U8542 ( .A(n8224), .ZN(n9893) );
  OAI21_X1 U8543 ( .B1(n6714), .B2(n6713), .A(n9893), .ZN(n6716) );
  NAND2_X1 U8544 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6715) );
  OAI211_X1 U8545 ( .C1(n6717), .C2(n8221), .A(n6716), .B(n6715), .ZN(n6718)
         );
  AOI21_X1 U8546 ( .B1(n6719), .B2(n9881), .A(n6718), .ZN(n6720) );
  OAI211_X1 U8547 ( .C1(n9887), .C2(n6722), .A(n6721), .B(n6720), .ZN(P2_U3187) );
  OAI21_X1 U8548 ( .B1(n6724), .B2(n9016), .A(n6723), .ZN(n7044) );
  NAND2_X1 U8549 ( .A1(n6725), .A2(n5846), .ZN(n6726) );
  AND3_X1 U8550 ( .A1(n6751), .A2(n7062), .A3(n6726), .ZN(n7043) );
  XNOR2_X1 U8551 ( .A(n6727), .B(n9016), .ZN(n6731) );
  INV_X1 U8552 ( .A(n6728), .ZN(n6730) );
  OAI22_X1 U8553 ( .A1(n6731), .A2(n9546), .B1(n6730), .B2(n6729), .ZN(n7040)
         );
  AOI211_X1 U8554 ( .C1(n9836), .C2(n7044), .A(n7043), .B(n7040), .ZN(n6920)
         );
  OAI22_X1 U8555 ( .A1(n9689), .A2(n5848), .B1(n9691), .B2(n5840), .ZN(n6732)
         );
  INV_X1 U8556 ( .A(n6732), .ZN(n6733) );
  OAI21_X1 U8557 ( .B1(n6920), .B2(n9838), .A(n6733), .ZN(P1_U3459) );
  OAI21_X1 U8558 ( .B1(n6735), .B2(n9013), .A(n6734), .ZN(n6977) );
  INV_X1 U8559 ( .A(n6736), .ZN(n6763) );
  INV_X1 U8560 ( .A(n6797), .ZN(n6737) );
  AOI211_X1 U8561 ( .C1(n8805), .C2(n6763), .A(n9557), .B(n6737), .ZN(n6972)
         );
  XNOR2_X1 U8562 ( .A(n6738), .B(n9013), .ZN(n6739) );
  OAI222_X1 U8563 ( .A1(n9549), .A2(n8803), .B1(n9551), .B2(n6755), .C1(n6739), 
        .C2(n9546), .ZN(n6971) );
  AOI211_X1 U8564 ( .C1(n9836), .C2(n6977), .A(n6972), .B(n6971), .ZN(n6805)
         );
  OAI22_X1 U8565 ( .A1(n9689), .A2(n6975), .B1(n9691), .B2(n5875), .ZN(n6740)
         );
  INV_X1 U8566 ( .A(n6740), .ZN(n6741) );
  OAI21_X1 U8567 ( .B1(n6805), .B2(n9838), .A(n6741), .ZN(P1_U3468) );
  INV_X1 U8568 ( .A(n9651), .ZN(n9825) );
  INV_X1 U8569 ( .A(n6742), .ZN(n6744) );
  AOI211_X1 U8570 ( .C1(n9825), .C2(n6745), .A(n6744), .B(n6743), .ZN(n6892)
         );
  OAI22_X1 U8571 ( .A1(n9689), .A2(n4415), .B1(n9691), .B2(n5812), .ZN(n6746)
         );
  INV_X1 U8572 ( .A(n6746), .ZN(n6747) );
  OAI21_X1 U8573 ( .B1(n6892), .B2(n9838), .A(n6747), .ZN(P1_U3456) );
  OAI21_X1 U8574 ( .B1(n6750), .B2(n9014), .A(n6749), .ZN(n6872) );
  AOI21_X1 U8575 ( .B1(n6751), .B2(n6866), .A(n9557), .ZN(n6752) );
  AND2_X1 U8576 ( .A1(n6761), .A2(n6752), .ZN(n6865) );
  XNOR2_X1 U8577 ( .A(n9014), .B(n6753), .ZN(n6754) );
  OAI222_X1 U8578 ( .A1(n9549), .A2(n6755), .B1(n9551), .B2(n5847), .C1(n6754), 
        .C2(n9546), .ZN(n6863) );
  AOI211_X1 U8579 ( .C1(n9836), .C2(n6872), .A(n6865), .B(n6863), .ZN(n6810)
         );
  OAI22_X1 U8580 ( .A1(n9689), .A2(n6807), .B1(n9691), .B2(n5850), .ZN(n6756)
         );
  INV_X1 U8581 ( .A(n6756), .ZN(n6757) );
  OAI21_X1 U8582 ( .B1(n6810), .B2(n9838), .A(n6757), .ZN(P1_U3462) );
  INV_X1 U8583 ( .A(n9836), .ZN(n9627) );
  OAI21_X1 U8584 ( .B1(n6759), .B2(n9015), .A(n6758), .ZN(n6881) );
  INV_X1 U8585 ( .A(n6881), .ZN(n6764) );
  XNOR2_X1 U8586 ( .A(n8905), .B(n9015), .ZN(n6760) );
  AOI222_X1 U8587 ( .A1(n9523), .A2(n6760), .B1(n9170), .B2(n9530), .C1(n9168), 
        .C2(n9528), .ZN(n6883) );
  AOI21_X1 U8588 ( .B1(n6761), .B2(n6875), .A(n9557), .ZN(n6762) );
  NAND2_X1 U8589 ( .A1(n6763), .A2(n6762), .ZN(n6879) );
  OAI211_X1 U8590 ( .C1(n9627), .C2(n6764), .A(n6883), .B(n6879), .ZN(n6886)
         );
  OAI22_X1 U8591 ( .A1(n9689), .A2(n6884), .B1(n9691), .B2(n5863), .ZN(n6765)
         );
  AOI21_X1 U8592 ( .B1(n6886), .B2(n9691), .A(n6765), .ZN(n6766) );
  INV_X1 U8593 ( .A(n6766), .ZN(P1_U3465) );
  XNOR2_X1 U8594 ( .A(n6767), .B(n7546), .ZN(n6768) );
  OAI222_X1 U8595 ( .A1(n9909), .A2(n6901), .B1(n9910), .B2(n5227), .C1(n9907), 
        .C2(n6768), .ZN(n9928) );
  INV_X1 U8596 ( .A(n9928), .ZN(n6776) );
  INV_X1 U8597 ( .A(n7546), .ZN(n6769) );
  NAND3_X1 U8598 ( .A1(n9896), .A2(n7611), .A3(n6769), .ZN(n6770) );
  NAND2_X1 U8599 ( .A1(n6771), .A2(n6770), .ZN(n9930) );
  NAND2_X1 U8600 ( .A1(n7598), .A2(n7744), .ZN(n6980) );
  NAND2_X1 U8601 ( .A1(n7165), .A2(n6980), .ZN(n9912) );
  AOI22_X1 U8602 ( .A1(n8445), .A2(n5245), .B1(n8389), .B2(n6772), .ZN(n6773)
         );
  OAI21_X1 U8603 ( .B1(n6225), .B2(n9913), .A(n6773), .ZN(n6774) );
  AOI21_X1 U8604 ( .B1(n9930), .B2(n8419), .A(n6774), .ZN(n6775) );
  OAI21_X1 U8605 ( .B1(n6776), .B2(n8421), .A(n6775), .ZN(P2_U3230) );
  INV_X1 U8606 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10292) );
  INV_X1 U8607 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9802) );
  INV_X1 U8608 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10238) );
  INV_X1 U8609 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8163) );
  AOI22_X1 U8610 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10238), .B2(n8163), .ZN(n10003) );
  NOR2_X1 U8611 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6777) );
  AOI21_X1 U8612 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6777), .ZN(n10006) );
  INV_X1 U8613 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10332) );
  INV_X1 U8614 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8117) );
  AOI22_X1 U8615 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n10332), .B2(n8117), .ZN(n10009) );
  NOR2_X1 U8616 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6778) );
  AOI21_X1 U8617 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6778), .ZN(n10012) );
  NOR2_X1 U8618 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6779) );
  AOI21_X1 U8619 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6779), .ZN(n10015) );
  NOR2_X1 U8620 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6780) );
  AOI21_X1 U8621 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6780), .ZN(n10018) );
  INV_X1 U8622 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10175) );
  INV_X1 U8623 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7385) );
  AOI22_X1 U8624 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n10175), .B2(n7385), .ZN(n10021) );
  NOR2_X1 U8625 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6781) );
  AOI21_X1 U8626 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6781), .ZN(n10024) );
  INV_X1 U8627 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10305) );
  INV_X1 U8628 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U8629 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(n10305), .B2(n10307), .ZN(n10346) );
  NOR2_X1 U8630 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6782) );
  AOI21_X1 U8631 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6782), .ZN(n10352) );
  INV_X1 U8632 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10105) );
  INV_X1 U8633 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U8634 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .B1(n10105), .B2(n10166), .ZN(n10349) );
  INV_X1 U8635 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10266) );
  INV_X1 U8636 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U8637 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .B1(n10266), .B2(n10122), .ZN(n10340) );
  NOR2_X1 U8638 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6783) );
  AOI21_X1 U8639 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6783), .ZN(n10343) );
  AND2_X1 U8640 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6784) );
  NOR2_X1 U8641 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6784), .ZN(n9994) );
  INV_X1 U8642 ( .A(n9994), .ZN(n9995) );
  INV_X1 U8643 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10091) );
  NAND3_X1 U8644 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U8645 ( .A1(n10091), .A2(n9996), .ZN(n9993) );
  NAND2_X1 U8646 ( .A1(n9995), .A2(n9993), .ZN(n10355) );
  NAND2_X1 U8647 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6785) );
  OAI21_X1 U8648 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6785), .ZN(n10354) );
  NOR2_X1 U8649 ( .A1(n10355), .A2(n10354), .ZN(n10353) );
  AOI21_X1 U8650 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10353), .ZN(n10358) );
  NAND2_X1 U8651 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6786) );
  OAI21_X1 U8652 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6786), .ZN(n10357) );
  NOR2_X1 U8653 ( .A1(n10358), .A2(n10357), .ZN(n10356) );
  AOI21_X1 U8654 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10356), .ZN(n10361) );
  NOR2_X1 U8655 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n6787) );
  AOI21_X1 U8656 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n6787), .ZN(n10360) );
  NAND2_X1 U8657 ( .A1(n10361), .A2(n10360), .ZN(n10359) );
  OAI21_X1 U8658 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10359), .ZN(n10342) );
  NAND2_X1 U8659 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  OAI21_X1 U8660 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10341), .ZN(n10339) );
  NAND2_X1 U8661 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  OAI21_X1 U8662 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10338), .ZN(n10348) );
  NAND2_X1 U8663 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  OAI21_X1 U8664 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10347), .ZN(n10351) );
  NAND2_X1 U8665 ( .A1(n10352), .A2(n10351), .ZN(n10350) );
  OAI21_X1 U8666 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10350), .ZN(n10345) );
  NAND2_X1 U8667 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  OAI21_X1 U8668 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10344), .ZN(n10023) );
  NAND2_X1 U8669 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U8670 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10022), .ZN(n10020) );
  NAND2_X1 U8671 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  OAI21_X1 U8672 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10019), .ZN(n10017) );
  NAND2_X1 U8673 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  OAI21_X1 U8674 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10016), .ZN(n10014) );
  NAND2_X1 U8675 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U8676 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10013), .ZN(n10011) );
  NAND2_X1 U8677 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  OAI21_X1 U8678 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10010), .ZN(n10008) );
  NAND2_X1 U8679 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  OAI21_X1 U8680 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10007), .ZN(n10005) );
  NAND2_X1 U8681 ( .A1(n10006), .A2(n10005), .ZN(n10004) );
  OAI21_X1 U8682 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10004), .ZN(n10002) );
  NAND2_X1 U8683 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  OAI21_X1 U8684 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10001), .ZN(n6788) );
  OR2_X1 U8685 ( .A1(n9802), .A2(n6788), .ZN(n10000) );
  NAND2_X1 U8686 ( .A1(n10292), .A2(n10000), .ZN(n9997) );
  NAND2_X1 U8687 ( .A1(n9802), .A2(n6788), .ZN(n9999) );
  NAND2_X1 U8688 ( .A1(n9997), .A2(n9999), .ZN(n6792) );
  NOR2_X1 U8689 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  XNOR2_X1 U8690 ( .A(n6792), .B(n6791), .ZN(ADD_1068_U4) );
  OAI21_X1 U8691 ( .B1(n6795), .B2(n9022), .A(n6794), .ZN(n6968) );
  INV_X1 U8692 ( .A(n7029), .ZN(n6796) );
  AOI211_X1 U8693 ( .C1(n6961), .C2(n6797), .A(n9557), .B(n6796), .ZN(n6962)
         );
  INV_X1 U8694 ( .A(n9062), .ZN(n6930) );
  XNOR2_X1 U8695 ( .A(n6930), .B(n9022), .ZN(n6798) );
  OAI222_X1 U8696 ( .A1(n9549), .A2(n7190), .B1(n9551), .B2(n6799), .C1(n9546), 
        .C2(n6798), .ZN(n6960) );
  AOI211_X1 U8697 ( .C1(n9836), .C2(n6968), .A(n6962), .B(n6960), .ZN(n6895)
         );
  INV_X1 U8698 ( .A(n9689), .ZN(n7405) );
  AOI22_X1 U8699 ( .A1(n7405), .A2(n6961), .B1(n9838), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U8700 ( .B1(n6895), .B2(n9838), .A(n6800), .ZN(P1_U3471) );
  INV_X1 U8701 ( .A(n6801), .ZN(n6888) );
  AOI22_X1 U8702 ( .A1(n9799), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7071), .ZN(n6802) );
  OAI21_X1 U8703 ( .B1(n6888), .B2(n9707), .A(n6802), .ZN(P1_U3337) );
  OAI22_X1 U8704 ( .A1(n9645), .A2(n6975), .B1(n9845), .B2(n6385), .ZN(n6803)
         );
  INV_X1 U8705 ( .A(n6803), .ZN(n6804) );
  OAI21_X1 U8706 ( .B1(n6805), .B2(n9843), .A(n6804), .ZN(P1_U3527) );
  INV_X1 U8707 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6806) );
  OAI22_X1 U8708 ( .A1(n9645), .A2(n6807), .B1(n9845), .B2(n6806), .ZN(n6808)
         );
  INV_X1 U8709 ( .A(n6808), .ZN(n6809) );
  OAI21_X1 U8710 ( .B1(n6810), .B2(n9843), .A(n6809), .ZN(P1_U3525) );
  AOI22_X1 U8711 ( .A1(n8645), .A2(n8805), .B1(n8741), .B2(n9168), .ZN(n6816)
         );
  NAND2_X1 U8712 ( .A1(n8645), .A2(n6961), .ZN(n6818) );
  NAND2_X1 U8713 ( .A1(n9167), .A2(n8736), .ZN(n6817) );
  NAND2_X1 U8714 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  XNOR2_X1 U8715 ( .A(n6819), .B(n8678), .ZN(n6822) );
  NAND2_X1 U8716 ( .A1(n6961), .A2(n8736), .ZN(n6821) );
  NAND2_X1 U8717 ( .A1(n8740), .A2(n9167), .ZN(n6820) );
  AND2_X1 U8718 ( .A1(n6821), .A2(n6820), .ZN(n6823) );
  NAND2_X1 U8719 ( .A1(n6822), .A2(n6823), .ZN(n7169) );
  INV_X1 U8720 ( .A(n6822), .ZN(n6825) );
  INV_X1 U8721 ( .A(n6823), .ZN(n6824) );
  NAND2_X1 U8722 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  NOR2_X1 U8723 ( .A1(n6827), .A2(n6829), .ZN(n6832) );
  AOI22_X1 U8724 ( .A1(n8740), .A2(n9168), .B1(n8741), .B2(n8805), .ZN(n8797)
         );
  NAND2_X1 U8725 ( .A1(n8796), .A2(n8797), .ZN(n8795) );
  AND2_X1 U8726 ( .A1(n8797), .A2(n6829), .ZN(n6828) );
  INV_X1 U8727 ( .A(n6829), .ZN(n6831) );
  AOI21_X1 U8728 ( .B1(n6832), .B2(n8795), .A(n4492), .ZN(n6838) );
  INV_X1 U8729 ( .A(n6833), .ZN(n6963) );
  AOI22_X1 U8730 ( .A1(n8801), .A2(n9168), .B1(n8800), .B2(n6963), .ZN(n6837)
         );
  NOR2_X1 U8731 ( .A1(n8890), .A2(n7190), .ZN(n6834) );
  AOI211_X1 U8732 ( .C1(n6961), .C2(n8897), .A(n6835), .B(n6834), .ZN(n6836)
         );
  OAI211_X1 U8733 ( .C1(n6838), .C2(n8899), .A(n6837), .B(n6836), .ZN(P1_U3239) );
  MUX2_X1 U8734 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8208), .Z(n6998) );
  XOR2_X1 U8735 ( .A(n7003), .B(n6998), .Z(n6842) );
  NAND2_X1 U8736 ( .A1(n6843), .A2(n6842), .ZN(n6997) );
  OAI21_X1 U8737 ( .B1(n6843), .B2(n6842), .A(n6997), .ZN(n6844) );
  NAND2_X1 U8738 ( .A1(n6844), .A2(n9872), .ZN(n6862) );
  INV_X1 U8739 ( .A(n7003), .ZN(n6860) );
  INV_X1 U8740 ( .A(n6846), .ZN(n6845) );
  INV_X1 U8741 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9982) );
  MUX2_X1 U8742 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9982), .S(n7003), .Z(n6847)
         );
  NOR2_X1 U8743 ( .A1(n6845), .A2(n6847), .ZN(n6851) );
  NAND2_X1 U8744 ( .A1(n6848), .A2(n6847), .ZN(n7005) );
  INV_X1 U8745 ( .A(n7005), .ZN(n6849) );
  AOI21_X1 U8746 ( .B1(n6851), .B2(n6850), .A(n6849), .ZN(n6852) );
  NAND2_X1 U8747 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6913) );
  OAI21_X1 U8748 ( .B1(n8224), .B2(n6852), .A(n6913), .ZN(n6859) );
  MUX2_X1 U8749 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5283), .S(n7003), .Z(n6853)
         );
  INV_X1 U8750 ( .A(n6853), .ZN(n6855) );
  NAND3_X1 U8751 ( .A1(n6856), .A2(n6855), .A3(n6854), .ZN(n6857) );
  AOI21_X1 U8752 ( .B1(n6995), .B2(n6857), .A(n8221), .ZN(n6858) );
  AOI211_X1 U8753 ( .C1(n6860), .C2(n9881), .A(n6859), .B(n6858), .ZN(n6861)
         );
  OAI211_X1 U8754 ( .C1(n9887), .C2(n10122), .A(n6862), .B(n6861), .ZN(
        P2_U3188) );
  INV_X1 U8755 ( .A(n6863), .ZN(n6874) );
  NAND2_X1 U8756 ( .A1(n9502), .A2(n9554), .ZN(n6864) );
  NAND2_X1 U8757 ( .A1(n9803), .A2(n6864), .ZN(n9513) );
  INV_X1 U8758 ( .A(n6865), .ZN(n6870) );
  NAND2_X1 U8759 ( .A1(n9313), .A2(n6866), .ZN(n6869) );
  AOI22_X1 U8760 ( .A1(n9521), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9807), .B2(
        n6867), .ZN(n6868) );
  OAI211_X1 U8761 ( .C1(n9316), .C2(n6870), .A(n6869), .B(n6868), .ZN(n6871)
         );
  AOI21_X1 U8762 ( .B1(n9513), .B2(n6872), .A(n6871), .ZN(n6873) );
  OAI21_X1 U8763 ( .B1(n6874), .B2(n9521), .A(n6873), .ZN(P1_U3290) );
  NAND2_X1 U8764 ( .A1(n9313), .A2(n6875), .ZN(n6878) );
  AOI22_X1 U8765 ( .A1(n9521), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6876), .B2(
        n9807), .ZN(n6877) );
  OAI211_X1 U8766 ( .C1(n9316), .C2(n6879), .A(n6878), .B(n6877), .ZN(n6880)
         );
  AOI21_X1 U8767 ( .B1(n6881), .B2(n9513), .A(n6880), .ZN(n6882) );
  OAI21_X1 U8768 ( .B1(n6883), .B2(n9521), .A(n6882), .ZN(P1_U3289) );
  OAI22_X1 U8769 ( .A1(n9645), .A2(n6884), .B1(n9845), .B2(n6383), .ZN(n6885)
         );
  AOI21_X1 U8770 ( .B1(n6886), .B2(n9845), .A(n6885), .ZN(n6887) );
  INV_X1 U8771 ( .A(n6887), .ZN(P1_U3526) );
  INV_X1 U8772 ( .A(n8207), .ZN(n8194) );
  OAI222_X1 U8773 ( .A1(n8612), .A2(n10128), .B1(n8194), .B2(P2_U3151), .C1(
        n7861), .C2(n6888), .ZN(P2_U3277) );
  NAND2_X1 U8774 ( .A1(n8185), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6889) );
  OAI21_X1 U8775 ( .B1(n8237), .B2(n8185), .A(n6889), .ZN(P2_U3520) );
  INV_X1 U8776 ( .A(n9645), .ZN(n7407) );
  AOI22_X1 U8777 ( .A1(n7407), .A2(n6890), .B1(n9843), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6891) );
  OAI21_X1 U8778 ( .B1(n6892), .B2(n9843), .A(n6891), .ZN(P1_U3523) );
  NOR2_X1 U8779 ( .A1(n9845), .A2(n6388), .ZN(n6893) );
  AOI21_X1 U8780 ( .B1(n7407), .B2(n6961), .A(n6893), .ZN(n6894) );
  OAI21_X1 U8781 ( .B1(n6895), .B2(n9843), .A(n6894), .ZN(P1_U3528) );
  OR2_X1 U8782 ( .A1(n9908), .A2(n6896), .ZN(n6897) );
  XNOR2_X1 U8783 ( .A(n8011), .B(n4414), .ZN(n6899) );
  XNOR2_X1 U8784 ( .A(n6901), .B(n6899), .ZN(n8007) );
  INV_X1 U8785 ( .A(n6899), .ZN(n6900) );
  NAND2_X1 U8786 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  XNOR2_X1 U8787 ( .A(n7980), .B(n6674), .ZN(n6904) );
  XNOR2_X1 U8788 ( .A(n6904), .B(n8084), .ZN(n7977) );
  INV_X1 U8789 ( .A(n6904), .ZN(n6905) );
  OR2_X1 U8790 ( .A1(n8084), .A2(n6905), .ZN(n6906) );
  NAND2_X1 U8791 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8792 ( .A(n9942), .B(n4414), .ZN(n7197) );
  XNOR2_X1 U8793 ( .A(n7198), .B(n7197), .ZN(n6909) );
  AOI21_X1 U8794 ( .B1(n6908), .B2(n6909), .A(n8056), .ZN(n6912) );
  INV_X1 U8795 ( .A(n6908), .ZN(n6911) );
  INV_X1 U8796 ( .A(n6909), .ZN(n6910) );
  NAND2_X1 U8797 ( .A1(n6911), .A2(n6910), .ZN(n7200) );
  NAND2_X1 U8798 ( .A1(n6912), .A2(n7200), .ZN(n6918) );
  INV_X1 U8799 ( .A(n6913), .ZN(n6915) );
  INV_X1 U8800 ( .A(n8061), .ZN(n8032) );
  INV_X1 U8801 ( .A(n8084), .ZN(n7144) );
  INV_X1 U8802 ( .A(n8082), .ZN(n7143) );
  OAI22_X1 U8803 ( .A1(n8032), .A2(n7144), .B1(n7143), .B2(n8063), .ZN(n6914)
         );
  AOI211_X1 U8804 ( .C1(n6916), .C2(n8042), .A(n6915), .B(n6914), .ZN(n6917)
         );
  OAI211_X1 U8805 ( .C1(n7145), .C2(n8040), .A(n6918), .B(n6917), .ZN(P2_U3179) );
  AOI22_X1 U8806 ( .A1(n7407), .A2(n5846), .B1(n9843), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6919) );
  OAI21_X1 U8807 ( .B1(n6920), .B2(n9843), .A(n6919), .ZN(P1_U3524) );
  INV_X1 U8808 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10195) );
  INV_X1 U8809 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U8810 ( .A1(n6922), .A2(P2_REG1_REG_31__SCAN_IN), .B1(n6921), .B2(
        P2_REG0_REG_31__SCAN_IN), .ZN(n6923) );
  OAI211_X1 U8811 ( .C1(n4417), .C2(n6925), .A(n6924), .B(n6923), .ZN(n7569)
         );
  NAND2_X1 U8812 ( .A1(n7569), .A2(P2_U3893), .ZN(n6927) );
  OAI21_X1 U8813 ( .B1(P2_U3893), .B2(n10195), .A(n6927), .ZN(P2_U3522) );
  INV_X1 U8814 ( .A(n6928), .ZN(n7516) );
  OAI222_X1 U8815 ( .A1(n8612), .A2(n6929), .B1(n8608), .B2(n7516), .C1(n7584), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  AOI21_X1 U8816 ( .B1(n6930), .B2(n8907), .A(n8914), .ZN(n7030) );
  OAI21_X1 U8817 ( .B1(n7030), .B2(n8915), .A(n6931), .ZN(n6949) );
  INV_X1 U8818 ( .A(n6948), .ZN(n6933) );
  AOI21_X1 U8819 ( .B1(n6949), .B2(n6933), .A(n6932), .ZN(n6934) );
  XOR2_X1 U8820 ( .A(n6937), .B(n6934), .Z(n6935) );
  OAI22_X1 U8821 ( .A1(n6935), .A2(n9546), .B1(n8619), .B2(n9551), .ZN(n9828)
         );
  INV_X1 U8822 ( .A(n9828), .ZN(n6945) );
  OAI21_X1 U8823 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(n9830) );
  XNOR2_X1 U8824 ( .A(n6954), .B(n7294), .ZN(n6939) );
  AOI22_X1 U8825 ( .A1(n6939), .A2(n7062), .B1(n9528), .B2(n9163), .ZN(n9826)
         );
  OAI22_X1 U8826 ( .A1(n9502), .A2(n6940), .B1(n7300), .B2(n9499), .ZN(n6941)
         );
  AOI21_X1 U8827 ( .B1(n9313), .B2(n7294), .A(n6941), .ZN(n6942) );
  OAI21_X1 U8828 ( .B1(n9826), .B2(n9316), .A(n6942), .ZN(n6943) );
  AOI21_X1 U8829 ( .B1(n9830), .B2(n9513), .A(n6943), .ZN(n6944) );
  OAI21_X1 U8830 ( .B1(n6945), .B2(n9521), .A(n6944), .ZN(P1_U3284) );
  OAI21_X1 U8831 ( .B1(n6947), .B2(n6948), .A(n6946), .ZN(n9824) );
  INV_X1 U8832 ( .A(n9824), .ZN(n6959) );
  XNOR2_X1 U8833 ( .A(n6949), .B(n6948), .ZN(n6952) );
  NAND2_X1 U8834 ( .A1(n9824), .A2(n9554), .ZN(n6951) );
  AOI22_X1 U8835 ( .A1(n9530), .A2(n9166), .B1(n9528), .B2(n9164), .ZN(n6950)
         );
  OAI211_X1 U8836 ( .C1(n9546), .C2(n6952), .A(n6951), .B(n6950), .ZN(n9822)
         );
  NAND2_X1 U8837 ( .A1(n9822), .A2(n9502), .ZN(n6958) );
  OAI22_X1 U8838 ( .A1(n9502), .A2(n6953), .B1(n7191), .B2(n9499), .ZN(n6956)
         );
  INV_X1 U8839 ( .A(n6954), .ZN(n7061) );
  OAI211_X1 U8840 ( .C1(n9821), .C2(n7028), .A(n7061), .B(n7062), .ZN(n9820)
         );
  NOR2_X1 U8841 ( .A1(n9820), .A2(n9316), .ZN(n6955) );
  AOI211_X1 U8842 ( .C1(n9313), .C2(n7194), .A(n6956), .B(n6955), .ZN(n6957)
         );
  OAI211_X1 U8843 ( .C1(n6959), .C2(n9803), .A(n6958), .B(n6957), .ZN(P1_U3285) );
  INV_X1 U8844 ( .A(n6960), .ZN(n6970) );
  INV_X1 U8845 ( .A(n6961), .ZN(n6966) );
  NAND2_X1 U8846 ( .A1(n6962), .A2(n9805), .ZN(n6965) );
  AOI22_X1 U8847 ( .A1(n9521), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6963), .B2(
        n9807), .ZN(n6964) );
  OAI211_X1 U8848 ( .C1(n6966), .C2(n9811), .A(n6965), .B(n6964), .ZN(n6967)
         );
  AOI21_X1 U8849 ( .B1(n6968), .B2(n9513), .A(n6967), .ZN(n6969) );
  OAI21_X1 U8850 ( .B1(n6970), .B2(n9521), .A(n6969), .ZN(P1_U3287) );
  INV_X1 U8851 ( .A(n6971), .ZN(n6979) );
  NAND2_X1 U8852 ( .A1(n6972), .A2(n9805), .ZN(n6974) );
  AOI22_X1 U8853 ( .A1(n9521), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8799), .B2(
        n9807), .ZN(n6973) );
  OAI211_X1 U8854 ( .C1(n6975), .C2(n9811), .A(n6974), .B(n6973), .ZN(n6976)
         );
  AOI21_X1 U8855 ( .B1(n9513), .B2(n6977), .A(n6976), .ZN(n6978) );
  OAI21_X1 U8856 ( .B1(n6979), .B2(n9521), .A(n6978), .ZN(P1_U3288) );
  OR2_X1 U8857 ( .A1(n8421), .A2(n6980), .ZN(n7344) );
  INV_X1 U8858 ( .A(n7344), .ZN(n7023) );
  NAND2_X1 U8859 ( .A1(n6982), .A2(n6981), .ZN(n9921) );
  OAI22_X1 U8860 ( .A1(n8352), .A2(n9918), .B1(n6983), .B2(n9898), .ZN(n6992)
         );
  INV_X1 U8861 ( .A(n6984), .ZN(n9903) );
  OAI21_X1 U8862 ( .B1(n9903), .B2(n6986), .A(n8413), .ZN(n6990) );
  INV_X1 U8863 ( .A(n7165), .ZN(n7336) );
  NAND2_X1 U8864 ( .A1(n9921), .A2(n7336), .ZN(n6989) );
  AOI22_X1 U8865 ( .A1(n8408), .A2(n6987), .B1(n5229), .B2(n8410), .ZN(n6988)
         );
  NAND3_X1 U8866 ( .A1(n6990), .A2(n6989), .A3(n6988), .ZN(n9919) );
  MUX2_X1 U8867 ( .A(n9919), .B(P2_REG2_REG_1__SCAN_IN), .S(n8421), .Z(n6991)
         );
  AOI211_X1 U8868 ( .C1(n7023), .C2(n9921), .A(n6992), .B(n6991), .ZN(n6993)
         );
  INV_X1 U8869 ( .A(n6993), .ZN(P2_U3232) );
  NAND2_X1 U8870 ( .A1(n7003), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6994) );
  AOI21_X1 U8871 ( .B1(n5303), .B2(n6996), .A(n4494), .ZN(n7013) );
  MUX2_X1 U8872 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8208), .Z(n7073) );
  XOR2_X1 U8873 ( .A(n7006), .B(n7073), .Z(n7075) );
  XNOR2_X1 U8874 ( .A(n7076), .B(n7075), .ZN(n6999) );
  NAND2_X1 U8875 ( .A1(n6999), .A2(n9872), .ZN(n7012) );
  INV_X1 U8876 ( .A(n9887), .ZN(n9846) );
  NAND2_X1 U8877 ( .A1(n9881), .A2(n4499), .ZN(n7002) );
  NOR2_X1 U8878 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7000), .ZN(n7867) );
  INV_X1 U8879 ( .A(n7867), .ZN(n7001) );
  NAND2_X1 U8880 ( .A1(n7002), .A2(n7001), .ZN(n7010) );
  NAND2_X1 U8881 ( .A1(n7003), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7004) );
  INV_X1 U8882 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U8883 ( .A1(n7007), .A2(n9984), .ZN(n7008) );
  AOI21_X1 U8884 ( .B1(n7081), .B2(n7008), .A(n8224), .ZN(n7009) );
  AOI211_X1 U8885 ( .C1(n9846), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7010), .B(
        n7009), .ZN(n7011) );
  OAI211_X1 U8886 ( .C1(n7013), .C2(n8221), .A(n7012), .B(n7011), .ZN(P2_U3189) );
  OR2_X1 U8887 ( .A1(n7014), .A2(n4440), .ZN(n7548) );
  XNOR2_X1 U8888 ( .A(n7015), .B(n7548), .ZN(n7020) );
  AOI22_X1 U8889 ( .A1(n8408), .A2(n8085), .B1(n8083), .B2(n8410), .ZN(n7019)
         );
  NAND2_X1 U8890 ( .A1(n7016), .A2(n7048), .ZN(n7017) );
  XNOR2_X1 U8891 ( .A(n7017), .B(n7548), .ZN(n9941) );
  NAND2_X1 U8892 ( .A1(n9941), .A2(n7336), .ZN(n7018) );
  OAI211_X1 U8893 ( .C1(n7020), .C2(n9907), .A(n7019), .B(n7018), .ZN(n9939)
         );
  INV_X1 U8894 ( .A(n9939), .ZN(n7025) );
  NOR2_X1 U8895 ( .A1(n9913), .A2(n5266), .ZN(n7022) );
  OAI22_X1 U8896 ( .A1(n8352), .A2(n9938), .B1(n7981), .B2(n9898), .ZN(n7021)
         );
  AOI211_X1 U8897 ( .C1(n9941), .C2(n7023), .A(n7022), .B(n7021), .ZN(n7024)
         );
  OAI21_X1 U8898 ( .B1(n7025), .B2(n8421), .A(n7024), .ZN(P2_U3228) );
  OAI21_X1 U8899 ( .B1(n7027), .B2(n8915), .A(n7026), .ZN(n9815) );
  AOI211_X1 U8900 ( .C1(n9804), .C2(n7029), .A(n9557), .B(n7028), .ZN(n9806)
         );
  XOR2_X1 U8901 ( .A(n8915), .B(n7030), .Z(n7032) );
  AOI22_X1 U8902 ( .A1(n9530), .A2(n9167), .B1(n9528), .B2(n9165), .ZN(n7031)
         );
  OAI21_X1 U8903 ( .B1(n7032), .B2(n9546), .A(n7031), .ZN(n7033) );
  AOI21_X1 U8904 ( .B1(n9554), .B2(n9815), .A(n7033), .ZN(n9817) );
  INV_X1 U8905 ( .A(n9817), .ZN(n7034) );
  AOI211_X1 U8906 ( .C1(n9825), .C2(n9815), .A(n9806), .B(n7034), .ZN(n7039)
         );
  NOR2_X1 U8907 ( .A1(n9691), .A2(n5903), .ZN(n7035) );
  AOI21_X1 U8908 ( .B1(n7405), .B2(n9804), .A(n7035), .ZN(n7036) );
  OAI21_X1 U8909 ( .B1(n7039), .B2(n9838), .A(n7036), .ZN(P1_U3474) );
  NOR2_X1 U8910 ( .A1(n9845), .A2(n6390), .ZN(n7037) );
  AOI21_X1 U8911 ( .B1(n7407), .B2(n9804), .A(n7037), .ZN(n7038) );
  OAI21_X1 U8912 ( .B1(n7039), .B2(n9843), .A(n7038), .ZN(P1_U3529) );
  INV_X1 U8913 ( .A(n7040), .ZN(n7047) );
  OAI22_X1 U8914 ( .A1(n9502), .A2(n6369), .B1(n9190), .B2(n9499), .ZN(n7042)
         );
  NOR2_X1 U8915 ( .A1(n9811), .A2(n5848), .ZN(n7041) );
  AOI211_X1 U8916 ( .C1(n7043), .C2(n9805), .A(n7042), .B(n7041), .ZN(n7046)
         );
  NAND2_X1 U8917 ( .A1(n9513), .A2(n7044), .ZN(n7045) );
  OAI211_X1 U8918 ( .C1(n9521), .C2(n7047), .A(n7046), .B(n7045), .ZN(P1_U3291) );
  AND2_X1 U8919 ( .A1(n7048), .A2(n7627), .ZN(n7618) );
  XOR2_X1 U8920 ( .A(n7618), .B(n7049), .Z(n9932) );
  XNOR2_X1 U8921 ( .A(n7050), .B(n7618), .ZN(n7051) );
  AOI222_X1 U8922 ( .A1(n8413), .A2(n7051), .B1(n8084), .B2(n8410), .C1(n5246), 
        .C2(n8408), .ZN(n9933) );
  MUX2_X1 U8923 ( .A(n7052), .B(n9933), .S(n9913), .Z(n7055) );
  INV_X1 U8924 ( .A(n7053), .ZN(n8012) );
  AOI22_X1 U8925 ( .A1(n8445), .A2(n8011), .B1(n8389), .B2(n8012), .ZN(n7054)
         );
  OAI211_X1 U8926 ( .C1(n8448), .C2(n9932), .A(n7055), .B(n7054), .ZN(P2_U3229) );
  OAI21_X1 U8927 ( .B1(n7057), .B2(n9029), .A(n7056), .ZN(n9837) );
  INV_X1 U8928 ( .A(n9837), .ZN(n7068) );
  INV_X1 U8929 ( .A(n7124), .ZN(n7058) );
  AOI21_X1 U8930 ( .B1(n9029), .B2(n7059), .A(n7058), .ZN(n7060) );
  OAI222_X1 U8931 ( .A1(n9549), .A2(n8764), .B1(n9551), .B2(n8728), .C1(n9546), 
        .C2(n7060), .ZN(n9834) );
  OAI21_X1 U8932 ( .B1(n7061), .B2(n7294), .A(n8731), .ZN(n7063) );
  NAND3_X1 U8933 ( .A1(n7063), .A2(n7062), .A3(n7130), .ZN(n9832) );
  OAI22_X1 U8934 ( .A1(n9502), .A2(n9243), .B1(n8729), .B2(n9499), .ZN(n7064)
         );
  AOI21_X1 U8935 ( .B1(n8731), .B2(n9313), .A(n7064), .ZN(n7065) );
  OAI21_X1 U8936 ( .B1(n9832), .B2(n9316), .A(n7065), .ZN(n7066) );
  AOI21_X1 U8937 ( .B1(n9834), .B2(n9502), .A(n7066), .ZN(n7067) );
  OAI21_X1 U8938 ( .B1(n7068), .B2(n9541), .A(n7067), .ZN(P1_U3283) );
  INV_X1 U8939 ( .A(n7069), .ZN(n7094) );
  AOI21_X1 U8940 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n7071), .A(n7070), .ZN(
        n7072) );
  OAI21_X1 U8941 ( .B1(n7094), .B2(n9707), .A(n7072), .ZN(P1_U3335) );
  MUX2_X1 U8942 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8208), .Z(n7096) );
  XOR2_X1 U8943 ( .A(n7106), .B(n7096), .Z(n7097) );
  INV_X1 U8944 ( .A(n7073), .ZN(n7074) );
  AOI22_X1 U8945 ( .A1(n7076), .A2(n7075), .B1(n4499), .B2(n7074), .ZN(n7098)
         );
  XOR2_X1 U8946 ( .A(n7097), .B(n7098), .Z(n7091) );
  INV_X1 U8947 ( .A(n9881), .ZN(n8184) );
  NAND2_X1 U8948 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7204) );
  OAI21_X1 U8949 ( .B1(n8184), .B2(n7095), .A(n7204), .ZN(n7084) );
  NAND2_X1 U8950 ( .A1(n7081), .A2(n7079), .ZN(n7077) );
  INV_X1 U8951 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9986) );
  MUX2_X1 U8952 ( .A(n9986), .B(P2_REG1_REG_8__SCAN_IN), .S(n7106), .Z(n7078)
         );
  INV_X1 U8953 ( .A(n7078), .ZN(n7080) );
  NAND3_X1 U8954 ( .A1(n7081), .A2(n7080), .A3(n7079), .ZN(n7082) );
  AOI21_X1 U8955 ( .B1(n7108), .B2(n7082), .A(n8224), .ZN(n7083) );
  AOI211_X1 U8956 ( .C1(n9846), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7084), .B(
        n7083), .ZN(n7090) );
  MUX2_X1 U8957 ( .A(n7101), .B(P2_REG2_REG_8__SCAN_IN), .S(n7106), .Z(n7087)
         );
  INV_X1 U8958 ( .A(n7086), .ZN(n7085) );
  NOR3_X1 U8959 ( .A1(n4494), .A2(n7087), .A3(n7085), .ZN(n7088) );
  INV_X1 U8960 ( .A(n8221), .ZN(n9883) );
  OAI21_X1 U8961 ( .B1(n7088), .B2(n4495), .A(n9883), .ZN(n7089) );
  OAI211_X1 U8962 ( .C1(n7091), .C2(n9848), .A(n7090), .B(n7089), .ZN(P2_U3190) );
  OAI222_X1 U8963 ( .A1(n7861), .A2(n7094), .B1(P2_U3151), .B2(n7093), .C1(
        n7092), .C2(n8612), .ZN(P2_U3275) );
  MUX2_X1 U8964 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8208), .Z(n7249) );
  XNOR2_X1 U8965 ( .A(n7249), .B(n7113), .ZN(n7099) );
  NAND2_X1 U8966 ( .A1(n7099), .A2(n7100), .ZN(n7250) );
  OAI21_X1 U8967 ( .B1(n7100), .B2(n7099), .A(n7250), .ZN(n7120) );
  OR2_X1 U8968 ( .A1(n7106), .A2(n7101), .ZN(n7102) );
  XNOR2_X1 U8969 ( .A(n7258), .B(n7113), .ZN(n7103) );
  INV_X1 U8970 ( .A(n7103), .ZN(n7104) );
  NAND2_X1 U8971 ( .A1(n7104), .A2(n5345), .ZN(n7105) );
  AOI21_X1 U8972 ( .B1(n7257), .B2(n7105), .A(n8221), .ZN(n7119) );
  OR2_X1 U8973 ( .A1(n7106), .A2(n9986), .ZN(n7107) );
  NAND2_X1 U8974 ( .A1(n7108), .A2(n7107), .ZN(n7110) );
  AOI21_X1 U8975 ( .B1(n7111), .B2(n5342), .A(n7245), .ZN(n7117) );
  NOR2_X1 U8976 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7112), .ZN(n7315) );
  AOI21_X1 U8977 ( .B1(n9881), .B2(n7113), .A(n7315), .ZN(n7114) );
  OAI21_X1 U8978 ( .B1(n9887), .B2(n10307), .A(n7114), .ZN(n7115) );
  INV_X1 U8979 ( .A(n7115), .ZN(n7116) );
  OAI21_X1 U8980 ( .B1(n7117), .B2(n8224), .A(n7116), .ZN(n7118) );
  AOI211_X1 U8981 ( .C1(n7120), .C2(n9872), .A(n7119), .B(n7118), .ZN(n7121)
         );
  INV_X1 U8982 ( .A(n7121), .ZN(P2_U3191) );
  NAND2_X1 U8983 ( .A1(n7122), .A2(n9523), .ZN(n7127) );
  INV_X1 U8984 ( .A(n9031), .ZN(n7123) );
  AOI21_X1 U8985 ( .B1(n7124), .B2(n8930), .A(n7123), .ZN(n7126) );
  AOI22_X1 U8986 ( .A1(n9530), .A2(n9163), .B1(n9528), .B2(n9161), .ZN(n7125)
         );
  OAI21_X1 U8987 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n7152) );
  INV_X1 U8988 ( .A(n7152), .ZN(n7137) );
  OAI21_X1 U8989 ( .B1(n7129), .B2(n9031), .A(n7128), .ZN(n7154) );
  NAND2_X1 U8990 ( .A1(n7154), .A2(n9513), .ZN(n7136) );
  AOI211_X1 U8991 ( .C1(n8862), .C2(n7130), .A(n9557), .B(n7230), .ZN(n7153)
         );
  INV_X1 U8992 ( .A(n8862), .ZN(n7131) );
  NOR2_X1 U8993 ( .A1(n7131), .A2(n9811), .ZN(n7134) );
  OAI22_X1 U8994 ( .A1(n9502), .A2(n7132), .B1(n8859), .B2(n9499), .ZN(n7133)
         );
  AOI211_X1 U8995 ( .C1(n7153), .C2(n9805), .A(n7134), .B(n7133), .ZN(n7135)
         );
  OAI211_X1 U8996 ( .C1(n9521), .C2(n7137), .A(n7136), .B(n7135), .ZN(P1_U3282) );
  NAND2_X1 U8997 ( .A1(n7139), .A2(n7138), .ZN(n7140) );
  AND2_X1 U8998 ( .A1(n7631), .A2(n7625), .ZN(n7549) );
  XNOR2_X1 U8999 ( .A(n7140), .B(n7549), .ZN(n9943) );
  XOR2_X1 U9000 ( .A(n7141), .B(n7549), .Z(n7142) );
  OAI222_X1 U9001 ( .A1(n9910), .A2(n7144), .B1(n9909), .B2(n7143), .C1(n7142), 
        .C2(n9907), .ZN(n9945) );
  NAND2_X1 U9002 ( .A1(n9945), .A2(n9913), .ZN(n7148) );
  OAI22_X1 U9003 ( .A1(n8352), .A2(n9942), .B1(n7145), .B2(n9898), .ZN(n7146)
         );
  AOI21_X1 U9004 ( .B1(n8421), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7146), .ZN(
        n7147) );
  OAI211_X1 U9005 ( .C1(n9943), .C2(n8448), .A(n7148), .B(n7147), .ZN(P2_U3227) );
  INV_X1 U9006 ( .A(n7149), .ZN(n7158) );
  OAI222_X1 U9007 ( .A1(n7861), .A2(n7158), .B1(P2_U3151), .B2(n7151), .C1(
        n7150), .C2(n8612), .ZN(P2_U3274) );
  AOI211_X1 U9008 ( .C1(n7154), .C2(n9836), .A(n7153), .B(n7152), .ZN(n7157)
         );
  AOI22_X1 U9009 ( .A1(n8862), .A2(n7405), .B1(n9838), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U9010 ( .B1(n7157), .B2(n9838), .A(n7155), .ZN(P1_U3486) );
  INV_X1 U9011 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9235) );
  AOI22_X1 U9012 ( .A1(n8862), .A2(n7407), .B1(n9843), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7156) );
  OAI21_X1 U9013 ( .B1(n7157), .B2(n9843), .A(n7156), .ZN(P1_U3533) );
  OAI222_X1 U9014 ( .A1(n9709), .A2(n10284), .B1(n9707), .B2(n7158), .C1(n9056), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U9015 ( .A1(n7159), .A2(n7642), .ZN(n7160) );
  NAND2_X1 U9016 ( .A1(n7212), .A2(n7160), .ZN(n9948) );
  OAI21_X1 U9017 ( .B1(n7161), .B2(n7642), .A(n7216), .ZN(n7162) );
  NAND2_X1 U9018 ( .A1(n7162), .A2(n8413), .ZN(n7164) );
  AOI22_X1 U9019 ( .A1(n8083), .A2(n8408), .B1(n8410), .B2(n8081), .ZN(n7163)
         );
  OAI211_X1 U9020 ( .C1(n7165), .C2(n9948), .A(n7164), .B(n7163), .ZN(n9950)
         );
  NAND2_X1 U9021 ( .A1(n9950), .A2(n9913), .ZN(n7168) );
  OAI22_X1 U9022 ( .A1(n8352), .A2(n9946), .B1(n7869), .B2(n9898), .ZN(n7166)
         );
  AOI21_X1 U9023 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n8421), .A(n7166), .ZN(
        n7167) );
  OAI211_X1 U9024 ( .C1(n9948), .C2(n7344), .A(n7168), .B(n7167), .ZN(P2_U3226) );
  OAI22_X1 U9025 ( .A1(n9821), .A2(n8651), .B1(n8619), .B2(n8680), .ZN(n7188)
         );
  INV_X1 U9026 ( .A(n7169), .ZN(n7172) );
  INV_X1 U9027 ( .A(n7170), .ZN(n7171) );
  NOR2_X1 U9028 ( .A1(n7172), .A2(n7171), .ZN(n7174) );
  NAND2_X1 U9029 ( .A1(n7174), .A2(n7173), .ZN(n8615) );
  NAND2_X1 U9030 ( .A1(n9804), .A2(n8735), .ZN(n7176) );
  NAND2_X1 U9031 ( .A1(n9166), .A2(n8736), .ZN(n7175) );
  NAND2_X1 U9032 ( .A1(n7176), .A2(n7175), .ZN(n7177) );
  XNOR2_X1 U9033 ( .A(n7177), .B(n8674), .ZN(n7180) );
  AOI22_X1 U9034 ( .A1(n9804), .A2(n8741), .B1(n8740), .B2(n9166), .ZN(n7178)
         );
  XNOR2_X1 U9035 ( .A(n7180), .B(n7178), .ZN(n8616) );
  INV_X1 U9036 ( .A(n7178), .ZN(n7179) );
  OR2_X1 U9037 ( .A1(n7180), .A2(n7179), .ZN(n7181) );
  AOI22_X1 U9038 ( .A1(n7194), .A2(n8645), .B1(n8741), .B2(n9165), .ZN(n7182)
         );
  XNOR2_X1 U9039 ( .A(n7182), .B(n8674), .ZN(n7183) );
  INV_X1 U9040 ( .A(n7296), .ZN(n7186) );
  AOI21_X1 U9041 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7196) );
  OAI21_X1 U9042 ( .B1(n8890), .B2(n8728), .A(n7189), .ZN(n7193) );
  INV_X1 U9043 ( .A(n8800), .ZN(n8894) );
  OAI22_X1 U9044 ( .A1(n8894), .A2(n7191), .B1(n7190), .B2(n8891), .ZN(n7192)
         );
  AOI211_X1 U9045 ( .C1(n7194), .C2(n8897), .A(n7193), .B(n7192), .ZN(n7195)
         );
  OAI21_X1 U9046 ( .B1(n7196), .B2(n8899), .A(n7195), .ZN(P1_U3221) );
  OR2_X1 U9047 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  XNOR2_X1 U9048 ( .A(n9946), .B(n4414), .ZN(n7201) );
  XNOR2_X1 U9049 ( .A(n7201), .B(n8082), .ZN(n7864) );
  INV_X1 U9050 ( .A(n7201), .ZN(n7202) );
  OR2_X1 U9051 ( .A1(n7202), .A2(n8082), .ZN(n7203) );
  XNOR2_X1 U9052 ( .A(n9951), .B(n4414), .ZN(n7271) );
  INV_X1 U9053 ( .A(n7271), .ZN(n7310) );
  XNOR2_X1 U9054 ( .A(n7270), .B(n7310), .ZN(n7311) );
  XNOR2_X1 U9055 ( .A(n7311), .B(n7334), .ZN(n7210) );
  INV_X1 U9056 ( .A(n7204), .ZN(n7206) );
  NOR2_X1 U9057 ( .A1(n8063), .A2(n7427), .ZN(n7205) );
  AOI211_X1 U9058 ( .C1(n8061), .C2(n8082), .A(n7206), .B(n7205), .ZN(n7209)
         );
  INV_X1 U9059 ( .A(n7220), .ZN(n7207) );
  AOI22_X1 U9060 ( .A1(n8066), .A2(n7207), .B1(n8042), .B2(n5330), .ZN(n7208)
         );
  OAI211_X1 U9061 ( .C1(n7210), .C2(n8056), .A(n7209), .B(n7208), .ZN(P2_U3161) );
  NAND2_X1 U9062 ( .A1(n7212), .A2(n7211), .ZN(n7213) );
  XOR2_X1 U9063 ( .A(n7550), .B(n7213), .Z(n9952) );
  NAND2_X1 U9064 ( .A1(n7214), .A2(n8413), .ZN(n7219) );
  AOI21_X1 U9065 ( .B1(n7216), .B2(n7215), .A(n7550), .ZN(n7218) );
  AOI22_X1 U9066 ( .A1(n7361), .A2(n8410), .B1(n8408), .B2(n8082), .ZN(n7217)
         );
  OAI21_X1 U9067 ( .B1(n7219), .B2(n7218), .A(n7217), .ZN(n9954) );
  NAND2_X1 U9068 ( .A1(n9954), .A2(n9913), .ZN(n7223) );
  OAI22_X1 U9069 ( .A1(n9913), .A2(n7101), .B1(n7220), .B2(n9898), .ZN(n7221)
         );
  AOI21_X1 U9070 ( .B1(n8445), .B2(n5330), .A(n7221), .ZN(n7222) );
  OAI211_X1 U9071 ( .C1(n9952), .C2(n8448), .A(n7223), .B(n7222), .ZN(P2_U3225) );
  INV_X1 U9072 ( .A(n7224), .ZN(n7225) );
  AOI21_X1 U9073 ( .B1(n9032), .B2(n7226), .A(n7225), .ZN(n7227) );
  OAI222_X1 U9074 ( .A1(n9549), .A2(n5993), .B1(n9551), .B2(n8764), .C1(n9546), 
        .C2(n7227), .ZN(n7239) );
  INV_X1 U9075 ( .A(n7239), .ZN(n7238) );
  OAI21_X1 U9076 ( .B1(n7229), .B2(n9032), .A(n7228), .ZN(n7241) );
  NAND2_X1 U9077 ( .A1(n7241), .A2(n9513), .ZN(n7237) );
  INV_X1 U9078 ( .A(n7230), .ZN(n7232) );
  INV_X1 U9079 ( .A(n7351), .ZN(n7231) );
  AOI211_X1 U9080 ( .C1(n8768), .C2(n7232), .A(n9557), .B(n7231), .ZN(n7240)
         );
  NOR2_X1 U9081 ( .A1(n5977), .A2(n9811), .ZN(n7235) );
  OAI22_X1 U9082 ( .A1(n9502), .A2(n7233), .B1(n8765), .B2(n9499), .ZN(n7234)
         );
  AOI211_X1 U9083 ( .C1(n7240), .C2(n9805), .A(n7235), .B(n7234), .ZN(n7236)
         );
  OAI211_X1 U9084 ( .C1(n9521), .C2(n7238), .A(n7237), .B(n7236), .ZN(P1_U3281) );
  AOI211_X1 U9085 ( .C1(n7241), .C2(n9836), .A(n7240), .B(n7239), .ZN(n7244)
         );
  AOI22_X1 U9086 ( .A1(n8768), .A2(n7405), .B1(n9838), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n7242) );
  OAI21_X1 U9087 ( .B1(n7244), .B2(n9838), .A(n7242), .ZN(P1_U3489) );
  AOI22_X1 U9088 ( .A1(n8768), .A2(n7407), .B1(n9843), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7243) );
  OAI21_X1 U9089 ( .B1(n7244), .B2(n9843), .A(n7243), .ZN(P1_U3534) );
  NAND2_X1 U9090 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7380), .ZN(n7246) );
  OAI21_X1 U9091 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7380), .A(n7246), .ZN(
        n7247) );
  AOI21_X1 U9092 ( .B1(n7248), .B2(n7247), .A(n7371), .ZN(n7268) );
  MUX2_X1 U9093 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8208), .Z(n7373) );
  XNOR2_X1 U9094 ( .A(n7373), .B(n7254), .ZN(n7253) );
  OR2_X1 U9095 ( .A1(n7249), .A2(n7259), .ZN(n7251) );
  NAND2_X1 U9096 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  NAND2_X1 U9097 ( .A1(n7253), .A2(n7252), .ZN(n7374) );
  OAI21_X1 U9098 ( .B1(n7253), .B2(n7252), .A(n7374), .ZN(n7266) );
  INV_X1 U9099 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7256) );
  INV_X1 U9100 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10300) );
  NOR2_X1 U9101 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10300), .ZN(n7360) );
  AOI21_X1 U9102 ( .B1(n9881), .B2(n7254), .A(n7360), .ZN(n7255) );
  OAI21_X1 U9103 ( .B1(n9887), .B2(n7256), .A(n7255), .ZN(n7265) );
  NAND2_X1 U9104 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7380), .ZN(n7260) );
  OAI21_X1 U9105 ( .B1(n7380), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7260), .ZN(
        n7261) );
  AOI21_X1 U9106 ( .B1(n7262), .B2(n7261), .A(n7379), .ZN(n7263) );
  NOR2_X1 U9107 ( .A1(n7263), .A2(n8221), .ZN(n7264) );
  AOI211_X1 U9108 ( .C1(n9872), .C2(n7266), .A(n7265), .B(n7264), .ZN(n7267)
         );
  OAI21_X1 U9109 ( .B1(n7268), .B2(n8224), .A(n7267), .ZN(P2_U3192) );
  XNOR2_X1 U9110 ( .A(n9955), .B(n4414), .ZN(n7312) );
  AOI22_X1 U9111 ( .A1(n7312), .A2(n7427), .B1(n7334), .B2(n7271), .ZN(n7269)
         );
  INV_X1 U9112 ( .A(n7312), .ZN(n7274) );
  OAI21_X1 U9113 ( .B1(n7271), .B2(n7334), .A(n7427), .ZN(n7273) );
  NOR2_X1 U9114 ( .A1(n7334), .A2(n7427), .ZN(n7272) );
  AOI22_X1 U9115 ( .A1(n7274), .A2(n7273), .B1(n7310), .B2(n7272), .ZN(n7275)
         );
  NAND2_X1 U9116 ( .A1(n7276), .A2(n7275), .ZN(n7359) );
  XNOR2_X1 U9117 ( .A(n8438), .B(n4414), .ZN(n7393) );
  XNOR2_X1 U9118 ( .A(n7362), .B(n6674), .ZN(n7391) );
  NAND2_X1 U9119 ( .A1(n7391), .A2(n8440), .ZN(n7277) );
  AND2_X1 U9120 ( .A1(n7393), .A2(n7277), .ZN(n7278) );
  NAND2_X1 U9121 ( .A1(n7359), .A2(n7278), .ZN(n7284) );
  NAND2_X1 U9122 ( .A1(n8080), .A2(n6674), .ZN(n7279) );
  OAI22_X1 U9123 ( .A1(n7362), .A2(n7279), .B1(n8429), .B2(n6674), .ZN(n7282)
         );
  NAND3_X1 U9124 ( .A1(n7362), .A2(n4414), .A3(n8080), .ZN(n7280) );
  OAI211_X1 U9125 ( .C1(n8429), .C2(n4414), .A(n8438), .B(n7280), .ZN(n7281)
         );
  OAI21_X1 U9126 ( .B1(n8438), .B2(n7282), .A(n7281), .ZN(n7283) );
  XNOR2_X1 U9127 ( .A(n7670), .B(n6674), .ZN(n7412) );
  XNOR2_X1 U9128 ( .A(n7412), .B(n8441), .ZN(n7285) );
  XNOR2_X1 U9129 ( .A(n7413), .B(n7285), .ZN(n7290) );
  AND2_X1 U9130 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7485) );
  NOR2_X1 U9131 ( .A1(n8063), .A2(n8430), .ZN(n7286) );
  AOI211_X1 U9132 ( .C1(n8061), .C2(n8079), .A(n7485), .B(n7286), .ZN(n7287)
         );
  OAI21_X1 U9133 ( .B1(n8431), .B2(n8040), .A(n7287), .ZN(n7288) );
  AOI21_X1 U9134 ( .B1(n8509), .B2(n8042), .A(n7288), .ZN(n7289) );
  OAI21_X1 U9135 ( .B1(n7290), .B2(n8056), .A(n7289), .ZN(P2_U3164) );
  NAND2_X1 U9136 ( .A1(n7294), .A2(n8735), .ZN(n7292) );
  NAND2_X1 U9137 ( .A1(n9164), .A2(n8741), .ZN(n7291) );
  NAND2_X1 U9138 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  XNOR2_X1 U9139 ( .A(n7293), .B(n8674), .ZN(n7770) );
  AOI22_X1 U9140 ( .A1(n7294), .A2(n8741), .B1(n8740), .B2(n9164), .ZN(n7768)
         );
  XNOR2_X1 U9141 ( .A(n7770), .B(n7768), .ZN(n7298) );
  OAI21_X1 U9142 ( .B1(n7298), .B2(n7297), .A(n7771), .ZN(n7299) );
  NAND2_X1 U9143 ( .A1(n7299), .A2(n5036), .ZN(n7304) );
  OAI22_X1 U9144 ( .A1(n8894), .A2(n7300), .B1(n8619), .B2(n8891), .ZN(n7301)
         );
  AOI211_X1 U9145 ( .C1(n8861), .C2(n9163), .A(n7302), .B(n7301), .ZN(n7303)
         );
  OAI211_X1 U9146 ( .C1(n9827), .C2(n8782), .A(n7304), .B(n7303), .ZN(P1_U3231) );
  INV_X1 U9147 ( .A(n7305), .ZN(n7308) );
  OAI222_X1 U9148 ( .A1(n8612), .A2(n7306), .B1(n7861), .B2(n7308), .C1(n7597), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9149 ( .A1(n9709), .A2(n7309), .B1(n9707), .B2(n7308), .C1(
        P1_U3086), .C2(n7307), .ZN(P1_U3333) );
  OAI22_X1 U9150 ( .A1(n7311), .A2(n8081), .B1(n7270), .B2(n7310), .ZN(n7314)
         );
  XNOR2_X1 U9151 ( .A(n7312), .B(n7361), .ZN(n7313) );
  XNOR2_X1 U9152 ( .A(n7314), .B(n7313), .ZN(n7322) );
  INV_X1 U9153 ( .A(n8056), .ZN(n8048) );
  AOI21_X1 U9154 ( .B1(n8061), .B2(n8081), .A(n7315), .ZN(n7320) );
  NAND2_X1 U9155 ( .A1(n8042), .A2(n7341), .ZN(n7319) );
  INV_X1 U9156 ( .A(n7339), .ZN(n7316) );
  NAND2_X1 U9157 ( .A1(n8066), .A2(n7316), .ZN(n7318) );
  INV_X1 U9158 ( .A(n8063), .ZN(n8030) );
  NAND2_X1 U9159 ( .A1(n8030), .A2(n8080), .ZN(n7317) );
  NAND4_X1 U9160 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), .ZN(n7321)
         );
  AOI21_X1 U9161 ( .B1(n7322), .B2(n8048), .A(n7321), .ZN(n7323) );
  INV_X1 U9162 ( .A(n7323), .ZN(P2_U3171) );
  NAND2_X1 U9163 ( .A1(n7327), .A2(n7324), .ZN(n7325) );
  OAI211_X1 U9164 ( .C1(n7326), .C2(n9709), .A(n7325), .B(n9142), .ZN(P1_U3332) );
  NAND2_X1 U9165 ( .A1(n7327), .A2(n8609), .ZN(n7329) );
  NAND2_X1 U9166 ( .A1(n7328), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7755) );
  OAI211_X1 U9167 ( .C1(n7330), .C2(n8612), .A(n7329), .B(n7755), .ZN(P2_U3272) );
  INV_X1 U9168 ( .A(n7331), .ZN(n7428) );
  AOI21_X1 U9169 ( .B1(n7545), .B2(n7332), .A(n7428), .ZN(n9959) );
  INV_X1 U9170 ( .A(n9959), .ZN(n7345) );
  XNOR2_X1 U9171 ( .A(n7333), .B(n7545), .ZN(n7338) );
  OAI22_X1 U9172 ( .A1(n7334), .A2(n9910), .B1(n8440), .B2(n9909), .ZN(n7335)
         );
  AOI21_X1 U9173 ( .B1(n9959), .B2(n7336), .A(n7335), .ZN(n7337) );
  OAI21_X1 U9174 ( .B1(n7338), .B2(n9907), .A(n7337), .ZN(n9956) );
  NAND2_X1 U9175 ( .A1(n9956), .A2(n9913), .ZN(n7343) );
  OAI22_X1 U9176 ( .A1(n9913), .A2(n5345), .B1(n7339), .B2(n9898), .ZN(n7340)
         );
  AOI21_X1 U9177 ( .B1(n8445), .B2(n7341), .A(n7340), .ZN(n7342) );
  OAI211_X1 U9178 ( .C1(n7345), .C2(n7344), .A(n7343), .B(n7342), .ZN(P2_U3224) );
  OAI21_X1 U9179 ( .B1(n7347), .B2(n9034), .A(n7346), .ZN(n7403) );
  INV_X1 U9180 ( .A(n7403), .ZN(n7358) );
  XNOR2_X1 U9181 ( .A(n7348), .B(n9034), .ZN(n7349) );
  OAI222_X1 U9182 ( .A1(n9551), .A2(n8839), .B1(n9549), .B2(n8892), .C1(n7349), 
        .C2(n9546), .ZN(n7401) );
  INV_X1 U9183 ( .A(n8843), .ZN(n7355) );
  AOI211_X1 U9184 ( .C1(n8843), .C2(n7351), .A(n9557), .B(n7350), .ZN(n7402)
         );
  NAND2_X1 U9185 ( .A1(n7402), .A2(n9805), .ZN(n7354) );
  INV_X1 U9186 ( .A(n8840), .ZN(n7352) );
  AOI22_X1 U9187 ( .A1(n9521), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7352), .B2(
        n9807), .ZN(n7353) );
  OAI211_X1 U9188 ( .C1(n7355), .C2(n9811), .A(n7354), .B(n7353), .ZN(n7356)
         );
  AOI21_X1 U9189 ( .B1(n7401), .B2(n9502), .A(n7356), .ZN(n7357) );
  OAI21_X1 U9190 ( .B1(n7358), .B2(n9541), .A(n7357), .ZN(P1_U3280) );
  XNOR2_X1 U9191 ( .A(n7359), .B(n8440), .ZN(n7392) );
  XNOR2_X1 U9192 ( .A(n7392), .B(n7391), .ZN(n7369) );
  AOI21_X1 U9193 ( .B1(n8061), .B2(n7361), .A(n7360), .ZN(n7367) );
  NAND2_X1 U9194 ( .A1(n7362), .A2(n8042), .ZN(n7366) );
  INV_X1 U9195 ( .A(n7363), .ZN(n7431) );
  NAND2_X1 U9196 ( .A1(n8066), .A2(n7431), .ZN(n7365) );
  NAND2_X1 U9197 ( .A1(n8030), .A2(n8079), .ZN(n7364) );
  NAND4_X1 U9198 ( .A1(n7367), .A2(n7366), .A3(n7365), .A4(n7364), .ZN(n7368)
         );
  AOI21_X1 U9199 ( .B1(n7369), .B2(n8048), .A(n7368), .ZN(n7370) );
  INV_X1 U9200 ( .A(n7370), .ZN(P2_U3157) );
  AOI21_X1 U9201 ( .B1(n5381), .B2(n7372), .A(n7462), .ZN(n7389) );
  MUX2_X1 U9202 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8208), .Z(n7477) );
  XNOR2_X1 U9203 ( .A(n7477), .B(n7468), .ZN(n7377) );
  OR2_X1 U9204 ( .A1(n7373), .A2(n7380), .ZN(n7375) );
  NAND2_X1 U9205 ( .A1(n7375), .A2(n7374), .ZN(n7376) );
  NAND2_X1 U9206 ( .A1(n7377), .A2(n7376), .ZN(n7475) );
  OAI21_X1 U9207 ( .B1(n7377), .B2(n7376), .A(n7475), .ZN(n7387) );
  INV_X1 U9208 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7378) );
  NOR2_X1 U9209 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7378), .ZN(n7396) );
  XNOR2_X1 U9210 ( .A(n7468), .B(n7467), .ZN(n7381) );
  NOR2_X1 U9211 ( .A1(n8443), .A2(n7381), .ZN(n7469) );
  AOI21_X1 U9212 ( .B1(n7381), .B2(n8443), .A(n7469), .ZN(n7382) );
  NOR2_X1 U9213 ( .A1(n8221), .A2(n7382), .ZN(n7383) );
  AOI211_X1 U9214 ( .C1(n7468), .C2(n9881), .A(n7396), .B(n7383), .ZN(n7384)
         );
  OAI21_X1 U9215 ( .B1(n7385), .B2(n9887), .A(n7384), .ZN(n7386) );
  AOI21_X1 U9216 ( .B1(n9872), .B2(n7387), .A(n7386), .ZN(n7388) );
  OAI21_X1 U9217 ( .B1(n7389), .B2(n8224), .A(n7388), .ZN(P2_U3193) );
  INV_X1 U9218 ( .A(n7359), .ZN(n7390) );
  AOI22_X1 U9219 ( .A1(n7392), .A2(n7391), .B1(n8440), .B2(n7390), .ZN(n7394)
         );
  XNOR2_X1 U9220 ( .A(n7394), .B(n7393), .ZN(n7400) );
  NOR2_X1 U9221 ( .A1(n8063), .A2(n8441), .ZN(n7395) );
  AOI211_X1 U9222 ( .C1(n8061), .C2(n8080), .A(n7396), .B(n7395), .ZN(n7397)
         );
  OAI21_X1 U9223 ( .B1(n8442), .B2(n8040), .A(n7397), .ZN(n7398) );
  AOI21_X1 U9224 ( .B1(n9971), .B2(n8042), .A(n7398), .ZN(n7399) );
  OAI21_X1 U9225 ( .B1(n7400), .B2(n8056), .A(n7399), .ZN(P2_U3176) );
  AOI211_X1 U9226 ( .C1(n7403), .C2(n9836), .A(n7402), .B(n7401), .ZN(n7409)
         );
  NOR2_X1 U9227 ( .A1(n9691), .A2(n5988), .ZN(n7404) );
  AOI21_X1 U9228 ( .B1(n8843), .B2(n7405), .A(n7404), .ZN(n7406) );
  OAI21_X1 U9229 ( .B1(n7409), .B2(n9838), .A(n7406), .ZN(P1_U3492) );
  AOI22_X1 U9230 ( .A1(n8843), .A2(n7407), .B1(n9843), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7408) );
  OAI21_X1 U9231 ( .B1(n7409), .B2(n9843), .A(n7408), .ZN(P1_U3535) );
  XNOR2_X1 U9232 ( .A(n8593), .B(n6674), .ZN(n7411) );
  INV_X1 U9233 ( .A(n7411), .ZN(n7410) );
  NAND2_X1 U9234 ( .A1(n7410), .A2(n8395), .ZN(n7440) );
  NAND2_X1 U9235 ( .A1(n7411), .A2(n8430), .ZN(n7438) );
  NAND2_X1 U9236 ( .A1(n7440), .A2(n7438), .ZN(n7416) );
  NAND2_X1 U9237 ( .A1(n7413), .A2(n8409), .ZN(n7414) );
  XOR2_X1 U9238 ( .A(n7416), .B(n7439), .Z(n7421) );
  NOR2_X1 U9239 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10200), .ZN(n8096) );
  NOR2_X1 U9240 ( .A1(n8063), .A2(n7877), .ZN(n7417) );
  AOI211_X1 U9241 ( .C1(n8061), .C2(n8409), .A(n8096), .B(n7417), .ZN(n7418)
         );
  OAI21_X1 U9242 ( .B1(n8406), .B2(n8040), .A(n7418), .ZN(n7419) );
  AOI21_X1 U9243 ( .B1(n8593), .B2(n8042), .A(n7419), .ZN(n7420) );
  OAI21_X1 U9244 ( .B1(n7421), .B2(n8056), .A(n7420), .ZN(P2_U3174) );
  INV_X1 U9245 ( .A(n7422), .ZN(n7436) );
  OAI222_X1 U9246 ( .A1(n7861), .A2(n7436), .B1(P2_U3151), .B2(n7424), .C1(
        n7423), .C2(n8612), .ZN(P2_U3271) );
  XOR2_X1 U9247 ( .A(n7553), .B(n7425), .Z(n7426) );
  OAI222_X1 U9248 ( .A1(n9909), .A2(n8429), .B1(n9910), .B2(n7427), .C1(n9907), 
        .C2(n7426), .ZN(n9963) );
  INV_X1 U9249 ( .A(n9963), .ZN(n7435) );
  OAI21_X1 U9250 ( .B1(n7428), .B2(n7640), .A(n7553), .ZN(n7430) );
  NAND2_X1 U9251 ( .A1(n7430), .A2(n7429), .ZN(n9965) );
  AOI22_X1 U9252 ( .A1(n8421), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8389), .B2(
        n7431), .ZN(n7432) );
  OAI21_X1 U9253 ( .B1(n9962), .B2(n8352), .A(n7432), .ZN(n7433) );
  AOI21_X1 U9254 ( .B1(n9965), .B2(n8419), .A(n7433), .ZN(n7434) );
  OAI21_X1 U9255 ( .B1(n7435), .B2(n8421), .A(n7434), .ZN(P2_U3223) );
  OAI222_X1 U9256 ( .A1(n7437), .A2(P1_U3086), .B1(n9707), .B2(n7436), .C1(
        n10079), .C2(n9709), .ZN(P1_U3331) );
  XNOR2_X1 U9257 ( .A(n8399), .B(n6674), .ZN(n7876) );
  XNOR2_X1 U9258 ( .A(n7876), .B(n8411), .ZN(n7879) );
  XOR2_X1 U9259 ( .A(n7879), .B(n7880), .Z(n7445) );
  AOI22_X1 U9260 ( .A1(n8030), .A2(n8396), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7442) );
  NAND2_X1 U9261 ( .A1(n8061), .A2(n8395), .ZN(n7441) );
  OAI211_X1 U9262 ( .C1(n8398), .C2(n8040), .A(n7442), .B(n7441), .ZN(n7443)
         );
  AOI21_X1 U9263 ( .B1(n8587), .B2(n8042), .A(n7443), .ZN(n7444) );
  OAI21_X1 U9264 ( .B1(n7445), .B2(n8056), .A(n7444), .ZN(P2_U3155) );
  INV_X1 U9265 ( .A(n7446), .ZN(n7450) );
  OAI222_X1 U9266 ( .A1(n7861), .A2(n7450), .B1(P2_U3151), .B2(n7448), .C1(
        n7447), .C2(n8612), .ZN(P2_U3270) );
  OAI222_X1 U9267 ( .A1(n7451), .A2(P1_U3086), .B1(n9707), .B2(n7450), .C1(
        n7449), .C2(n9709), .ZN(P1_U3330) );
  INV_X1 U9268 ( .A(n7452), .ZN(n7456) );
  OAI222_X1 U9269 ( .A1(n7861), .A2(n7456), .B1(P2_U3151), .B2(n7454), .C1(
        n7453), .C2(n8612), .ZN(P2_U3269) );
  OAI222_X1 U9270 ( .A1(n7457), .A2(P1_U3086), .B1(n9707), .B2(n7456), .C1(
        n7455), .C2(n9709), .ZN(P1_U3329) );
  INV_X1 U9271 ( .A(n7458), .ZN(n7763) );
  AOI21_X1 U9272 ( .B1(n8606), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7459), .ZN(
        n7460) );
  OAI21_X1 U9273 ( .B1(n7763), .B2(n8608), .A(n7460), .ZN(P2_U3268) );
  NOR2_X1 U9274 ( .A1(n7468), .A2(n7461), .ZN(n7463) );
  NAND2_X1 U9275 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7495), .ZN(n7464) );
  OAI21_X1 U9276 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7495), .A(n7464), .ZN(
        n7465) );
  AOI21_X1 U9277 ( .B1(n7466), .B2(n7465), .A(n7494), .ZN(n7488) );
  NOR2_X1 U9278 ( .A1(n7468), .A2(n7467), .ZN(n7470) );
  NAND2_X1 U9279 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7495), .ZN(n7471) );
  OAI21_X1 U9280 ( .B1(n7495), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7471), .ZN(
        n7472) );
  AOI21_X1 U9281 ( .B1(n7473), .B2(n7472), .A(n7489), .ZN(n7474) );
  NOR2_X1 U9282 ( .A1(n7474), .A2(n8221), .ZN(n7486) );
  INV_X1 U9283 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10163) );
  OAI22_X1 U9284 ( .A1(n8184), .A2(n7495), .B1(n9887), .B2(n10163), .ZN(n7484)
         );
  OAI21_X1 U9285 ( .B1(n7477), .B2(n7476), .A(n7475), .ZN(n7482) );
  MUX2_X1 U9286 ( .A(n8432), .B(n8510), .S(n8208), .Z(n7478) );
  NOR2_X1 U9287 ( .A1(n7478), .A2(n7479), .ZN(n7503) );
  AOI21_X1 U9288 ( .B1(n7479), .B2(n7478), .A(n7503), .ZN(n7480) );
  INV_X1 U9289 ( .A(n7480), .ZN(n7481) );
  NOR2_X1 U9290 ( .A1(n7481), .A2(n7482), .ZN(n7502) );
  AOI211_X1 U9291 ( .C1(n7482), .C2(n7481), .A(n9848), .B(n7502), .ZN(n7483)
         );
  NOR4_X1 U9292 ( .A1(n7486), .A2(n7485), .A3(n7484), .A4(n7483), .ZN(n7487)
         );
  OAI21_X1 U9293 ( .B1(n7488), .B2(n8224), .A(n7487), .ZN(P2_U3194) );
  NOR2_X1 U9294 ( .A1(n8097), .A2(n7490), .ZN(n7491) );
  NAND2_X1 U9295 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8111), .ZN(n7492) );
  OAI21_X1 U9296 ( .B1(n8111), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7492), .ZN(
        n7493) );
  AOI21_X1 U9297 ( .B1(n4490), .B2(n7493), .A(n8110), .ZN(n7515) );
  NOR2_X1 U9298 ( .A1(n8097), .A2(n7496), .ZN(n7497) );
  NAND2_X1 U9299 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8111), .ZN(n7498) );
  OAI21_X1 U9300 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8111), .A(n7498), .ZN(
        n7499) );
  NOR2_X1 U9301 ( .A1(n7500), .A2(n7499), .ZN(n8103) );
  AOI21_X1 U9302 ( .B1(n7500), .B2(n7499), .A(n8103), .ZN(n7501) );
  OR2_X1 U9303 ( .A1(n7501), .A2(n8224), .ZN(n7514) );
  MUX2_X1 U9304 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8208), .Z(n7505) );
  XNOR2_X1 U9305 ( .A(n7505), .B(n8097), .ZN(n8091) );
  NAND2_X1 U9306 ( .A1(n8090), .A2(n8091), .ZN(n8089) );
  OAI21_X1 U9307 ( .B1(n7505), .B2(n7504), .A(n8089), .ZN(n7508) );
  MUX2_X1 U9308 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8208), .Z(n8105) );
  XNOR2_X1 U9309 ( .A(n8105), .B(n7506), .ZN(n7507) );
  NAND2_X1 U9310 ( .A1(n7507), .A2(n7508), .ZN(n8106) );
  OAI21_X1 U9311 ( .B1(n7508), .B2(n7507), .A(n8106), .ZN(n7512) );
  INV_X1 U9312 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7509) );
  NOR2_X1 U9313 ( .A1(n9887), .A2(n7509), .ZN(n7511) );
  INV_X1 U9314 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10084) );
  OAI22_X1 U9315 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10084), .B1(n8184), .B2(
        n8111), .ZN(n7510) );
  AOI211_X1 U9316 ( .C1(n9872), .C2(n7512), .A(n7511), .B(n7510), .ZN(n7513)
         );
  OAI211_X1 U9317 ( .C1(n7515), .C2(n8221), .A(n7514), .B(n7513), .ZN(P2_U3196) );
  OAI222_X1 U9318 ( .A1(n9709), .A2(n7517), .B1(n9707), .B2(n7516), .C1(
        P1_U3086), .C2(n6153), .ZN(P1_U3336) );
  INV_X1 U9319 ( .A(n7518), .ZN(n9702) );
  OAI222_X1 U9320 ( .A1(n8608), .A2(n9702), .B1(n7519), .B2(P2_U3151), .C1(
        n10078), .C2(n8612), .ZN(P2_U3266) );
  INV_X1 U9321 ( .A(SI_29_), .ZN(n7523) );
  OR2_X1 U9322 ( .A1(n7521), .A2(n7520), .ZN(n7522) );
  INV_X1 U9323 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7862) );
  INV_X1 U9324 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8995) );
  MUX2_X1 U9325 ( .A(n7862), .B(n8995), .S(n5133), .Z(n7526) );
  INV_X1 U9326 ( .A(SI_30_), .ZN(n7525) );
  NAND2_X1 U9327 ( .A1(n7526), .A2(n7525), .ZN(n7529) );
  INV_X1 U9328 ( .A(n7526), .ZN(n7527) );
  NAND2_X1 U9329 ( .A1(n7527), .A2(SI_30_), .ZN(n7528) );
  NAND2_X1 U9330 ( .A1(n7529), .A2(n7528), .ZN(n7535) );
  MUX2_X1 U9331 ( .A(n6348), .B(n10195), .S(n5133), .Z(n7530) );
  XNOR2_X1 U9332 ( .A(n7530), .B(SI_31_), .ZN(n7531) );
  MUX2_X1 U9333 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n8999), .S(n7533), .Z(n7534) );
  NAND2_X1 U9334 ( .A1(n8515), .A2(n7569), .ZN(n7743) );
  INV_X1 U9335 ( .A(n7743), .ZN(n7576) );
  OR2_X1 U9336 ( .A1(n7538), .A2(n7862), .ZN(n7539) );
  INV_X1 U9337 ( .A(n7570), .ZN(n8071) );
  NAND2_X1 U9338 ( .A1(n8518), .A2(n8071), .ZN(n7578) );
  INV_X1 U9339 ( .A(n7730), .ZN(n7568) );
  INV_X1 U9340 ( .A(n7541), .ZN(n7726) );
  INV_X1 U9341 ( .A(n7843), .ZN(n7567) );
  INV_X1 U9342 ( .A(n7722), .ZN(n7542) );
  NAND2_X1 U9343 ( .A1(n7713), .A2(n7711), .ZN(n8278) );
  INV_X1 U9344 ( .A(n7543), .ZN(n8311) );
  INV_X1 U9345 ( .A(n8321), .ZN(n7562) );
  INV_X1 U9346 ( .A(n8359), .ZN(n8361) );
  INV_X1 U9347 ( .A(n8371), .ZN(n8373) );
  AND2_X1 U9348 ( .A1(n7681), .A2(n7682), .ZN(n8393) );
  INV_X1 U9349 ( .A(n8393), .ZN(n8402) );
  INV_X1 U9350 ( .A(n7677), .ZN(n7544) );
  OR2_X1 U9351 ( .A1(n7673), .A2(n7544), .ZN(n8418) );
  NAND4_X1 U9352 ( .A1(n7546), .A2(n7757), .A3(n9897), .A4(n5694), .ZN(n7552)
         );
  NAND4_X1 U9353 ( .A1(n7549), .A2(n7618), .A3(n7548), .A4(n7547), .ZN(n7551)
         );
  NOR4_X1 U9354 ( .A1(n7553), .A2(n7552), .A3(n7551), .A4(n7550), .ZN(n7554)
         );
  NAND4_X1 U9355 ( .A1(n8418), .A2(n7555), .A3(n5696), .A4(n7554), .ZN(n7556)
         );
  NOR3_X1 U9356 ( .A1(n8402), .A2(n7556), .A3(n8423), .ZN(n7560) );
  INV_X1 U9357 ( .A(n7557), .ZN(n7558) );
  OR2_X1 U9358 ( .A1(n7559), .A2(n7558), .ZN(n8385) );
  NAND4_X1 U9359 ( .A1(n8361), .A2(n8373), .A3(n7560), .A4(n8385), .ZN(n7561)
         );
  NOR4_X1 U9360 ( .A1(n7562), .A2(n8331), .A3(n8351), .A4(n7561), .ZN(n7563)
         );
  NAND4_X1 U9361 ( .A1(n8285), .A2(n8311), .A3(n7563), .A4(n8295), .ZN(n7564)
         );
  NOR4_X1 U9362 ( .A1(n8251), .A2(n8267), .A3(n8278), .A4(n7564), .ZN(n7566)
         );
  NAND4_X1 U9363 ( .A1(n7568), .A2(n7567), .A3(n7566), .A4(n8234), .ZN(n7573)
         );
  INV_X1 U9364 ( .A(n7569), .ZN(n8227) );
  NAND2_X1 U9365 ( .A1(n7579), .A2(n8227), .ZN(n7740) );
  INV_X1 U9366 ( .A(n7740), .ZN(n7572) );
  NAND2_X1 U9367 ( .A1(n7577), .A2(n7570), .ZN(n7737) );
  NAND2_X1 U9368 ( .A1(n7737), .A2(n7571), .ZN(n7731) );
  NOR4_X1 U9369 ( .A1(n7576), .A2(n7573), .A3(n7572), .A4(n7731), .ZN(n7583)
         );
  NOR2_X1 U9370 ( .A1(n7574), .A2(n7732), .ZN(n7575) );
  OAI21_X1 U9371 ( .B1(n7575), .B2(n7731), .A(n7740), .ZN(n7581) );
  AOI21_X1 U9372 ( .B1(n8515), .B2(n7577), .A(n7576), .ZN(n7580) );
  INV_X1 U9373 ( .A(n7578), .ZN(n7736) );
  AOI22_X1 U9374 ( .A1(n7581), .A2(n7580), .B1(n7579), .B2(n7736), .ZN(n7582)
         );
  MUX2_X1 U9375 ( .A(n7583), .B(n7582), .S(n7598), .Z(n7585) );
  XNOR2_X1 U9376 ( .A(n7585), .B(n7584), .ZN(n7749) );
  MUX2_X1 U9377 ( .A(n7586), .B(n7590), .S(n7739), .Z(n7587) );
  INV_X1 U9378 ( .A(n7587), .ZN(n7588) );
  NOR2_X1 U9379 ( .A1(n8299), .A2(n7588), .ZN(n7708) );
  INV_X1 U9380 ( .A(n7708), .ZN(n7593) );
  AND2_X1 U9381 ( .A1(n7590), .A2(n7589), .ZN(n7592) );
  INV_X1 U9382 ( .A(n7594), .ZN(n7699) );
  NAND2_X1 U9383 ( .A1(n7600), .A2(n7597), .ZN(n7599) );
  MUX2_X1 U9384 ( .A(n6629), .B(n7599), .S(n7598), .Z(n7603) );
  INV_X1 U9385 ( .A(n7600), .ZN(n7601) );
  NAND2_X1 U9386 ( .A1(n5692), .A2(n7739), .ZN(n7606) );
  NAND2_X1 U9387 ( .A1(n7603), .A2(n7602), .ZN(n7610) );
  INV_X1 U9388 ( .A(n5692), .ZN(n7604) );
  NAND2_X1 U9389 ( .A1(n7604), .A2(n7738), .ZN(n7605) );
  OAI211_X1 U9390 ( .C1(n7607), .C2(n7606), .A(n9897), .B(n7605), .ZN(n7608)
         );
  INV_X1 U9391 ( .A(n7608), .ZN(n7609) );
  NAND2_X1 U9392 ( .A1(n7610), .A2(n7609), .ZN(n7617) );
  NAND2_X1 U9393 ( .A1(n7611), .A2(n7626), .ZN(n7614) );
  NAND2_X1 U9394 ( .A1(n7620), .A2(n7612), .ZN(n7613) );
  MUX2_X1 U9395 ( .A(n7614), .B(n7613), .S(n7738), .Z(n7615) );
  INV_X1 U9396 ( .A(n7615), .ZN(n7616) );
  NAND2_X1 U9397 ( .A1(n7617), .A2(n7616), .ZN(n7619) );
  NAND2_X1 U9398 ( .A1(n7619), .A2(n7618), .ZN(n7630) );
  INV_X1 U9399 ( .A(n7620), .ZN(n7622) );
  OAI21_X1 U9400 ( .B1(n7630), .B2(n7622), .A(n7621), .ZN(n7624) );
  INV_X1 U9401 ( .A(n7631), .ZN(n7623) );
  AOI21_X1 U9402 ( .B1(n7624), .B2(n7628), .A(n7623), .ZN(n7636) );
  INV_X1 U9403 ( .A(n7625), .ZN(n7634) );
  INV_X1 U9404 ( .A(n7626), .ZN(n7629) );
  OAI211_X1 U9405 ( .C1(n7630), .C2(n7629), .A(n7628), .B(n7627), .ZN(n7632)
         );
  OAI211_X1 U9406 ( .C1(n7634), .C2(n7633), .A(n7632), .B(n7631), .ZN(n7635)
         );
  MUX2_X1 U9407 ( .A(n7636), .B(n7635), .S(n7738), .Z(n7660) );
  NAND2_X1 U9408 ( .A1(n7653), .A2(n7648), .ZN(n7639) );
  INV_X1 U9409 ( .A(n7637), .ZN(n7638) );
  MUX2_X1 U9410 ( .A(n7639), .B(n7638), .S(n7738), .Z(n7641) );
  NOR2_X1 U9411 ( .A1(n7641), .A2(n7640), .ZN(n7652) );
  INV_X1 U9412 ( .A(n7652), .ZN(n7643) );
  NOR2_X1 U9413 ( .A1(n7643), .A2(n7642), .ZN(n7659) );
  INV_X1 U9414 ( .A(n7644), .ZN(n7645) );
  NAND3_X1 U9415 ( .A1(n7645), .A2(n7653), .A3(n7648), .ZN(n7647) );
  NAND3_X1 U9416 ( .A1(n7647), .A2(n7646), .A3(n7662), .ZN(n7657) );
  INV_X1 U9417 ( .A(n7648), .ZN(n7649) );
  NAND2_X1 U9418 ( .A1(n7652), .A2(n7649), .ZN(n7655) );
  INV_X1 U9419 ( .A(n7650), .ZN(n7651) );
  NAND2_X1 U9420 ( .A1(n7652), .A2(n7651), .ZN(n7654) );
  NAND4_X1 U9421 ( .A1(n7655), .A2(n7654), .A3(n7653), .A4(n7661), .ZN(n7656)
         );
  MUX2_X1 U9422 ( .A(n7657), .B(n7656), .S(n7738), .Z(n7658) );
  AOI21_X1 U9423 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n7669) );
  NAND2_X1 U9424 ( .A1(n7666), .A2(n7661), .ZN(n7664) );
  NAND2_X1 U9425 ( .A1(n7665), .A2(n7662), .ZN(n7663) );
  MUX2_X1 U9426 ( .A(n7664), .B(n7663), .S(n7738), .Z(n7668) );
  MUX2_X1 U9427 ( .A(n7666), .B(n7665), .S(n7739), .Z(n7667) );
  OAI211_X1 U9428 ( .C1(n7669), .C2(n7668), .A(n5699), .B(n7667), .ZN(n7676)
         );
  OR2_X1 U9429 ( .A1(n7670), .A2(n8409), .ZN(n7672) );
  MUX2_X1 U9430 ( .A(n7672), .B(n7671), .S(n7738), .Z(n7675) );
  MUX2_X1 U9431 ( .A(n8395), .B(n8593), .S(n7739), .Z(n7678) );
  NOR2_X1 U9432 ( .A1(n7678), .A2(n7673), .ZN(n7674) );
  AOI21_X1 U9433 ( .B1(n7676), .B2(n7675), .A(n7674), .ZN(n7680) );
  AND2_X1 U9434 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  OAI21_X1 U9435 ( .B1(n7680), .B2(n7679), .A(n8393), .ZN(n7684) );
  MUX2_X1 U9436 ( .A(n7682), .B(n7681), .S(n7738), .Z(n7683) );
  NAND3_X1 U9437 ( .A1(n7684), .A2(n8385), .A3(n7683), .ZN(n7685) );
  NAND2_X1 U9438 ( .A1(n8361), .A2(n7686), .ZN(n7692) );
  INV_X1 U9439 ( .A(n7687), .ZN(n7688) );
  NOR2_X1 U9440 ( .A1(n7692), .A2(n7688), .ZN(n7694) );
  INV_X1 U9441 ( .A(n7689), .ZN(n7691) );
  OAI211_X1 U9442 ( .C1(n7692), .C2(n7691), .A(n7702), .B(n7690), .ZN(n7693)
         );
  NAND3_X1 U9443 ( .A1(n7705), .A2(n7707), .A3(n7701), .ZN(n7695) );
  NAND3_X1 U9444 ( .A1(n7695), .A2(n8321), .A3(n7703), .ZN(n7697) );
  NAND2_X1 U9445 ( .A1(n8309), .A2(n7738), .ZN(n7696) );
  NAND2_X1 U9446 ( .A1(n7701), .A2(n7700), .ZN(n7704) );
  OAI211_X1 U9447 ( .C1(n7705), .C2(n7704), .A(n7703), .B(n7702), .ZN(n7706)
         );
  INV_X1 U9448 ( .A(n7709), .ZN(n8276) );
  OAI211_X1 U9449 ( .C1(n7715), .C2(n8276), .A(n7713), .B(n7710), .ZN(n7712)
         );
  INV_X1 U9450 ( .A(n7713), .ZN(n7714) );
  AOI21_X1 U9451 ( .B1(n7715), .B2(n4461), .A(n7714), .ZN(n7716) );
  MUX2_X1 U9452 ( .A(n7718), .B(n7717), .S(n7739), .Z(n7719) );
  INV_X1 U9453 ( .A(n7721), .ZN(n7723) );
  MUX2_X1 U9454 ( .A(n7723), .B(n7722), .S(n7739), .Z(n7724) );
  AOI211_X1 U9455 ( .C1(n7725), .C2(n8253), .A(n7724), .B(n7843), .ZN(n7729)
         );
  MUX2_X1 U9456 ( .A(n7727), .B(n7726), .S(n7738), .Z(n7728) );
  MUX2_X1 U9457 ( .A(n8072), .B(n8520), .S(n7739), .Z(n7735) );
  MUX2_X1 U9458 ( .A(n8072), .B(n8520), .S(n7738), .Z(n7733) );
  AOI21_X1 U9459 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7741) );
  INV_X1 U9460 ( .A(n7744), .ZN(n7746) );
  NAND3_X1 U9461 ( .A1(n7751), .A2(n7750), .A3(n8208), .ZN(n7752) );
  OAI211_X1 U9462 ( .C1(n7753), .C2(n7755), .A(n7752), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7754) );
  OAI21_X1 U9463 ( .B1(n7756), .B2(n7755), .A(n7754), .ZN(P2_U3296) );
  INV_X1 U9464 ( .A(n7757), .ZN(n7759) );
  AOI22_X1 U9465 ( .A1(n8048), .A2(n7759), .B1(n7758), .B2(n8042), .ZN(n7762)
         );
  NAND2_X1 U9466 ( .A1(n7760), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7761) );
  OAI211_X1 U9467 ( .C1(n5197), .C2(n8063), .A(n7762), .B(n7761), .ZN(P2_U3172) );
  OAI222_X1 U9468 ( .A1(n9709), .A2(n7764), .B1(n9707), .B2(n7763), .C1(n9183), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U9469 ( .A1(n8843), .A2(n8735), .ZN(n7766) );
  NAND2_X1 U9470 ( .A1(n9160), .A2(n8741), .ZN(n7765) );
  NAND2_X1 U9471 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  XNOR2_X1 U9472 ( .A(n7767), .B(n8674), .ZN(n7794) );
  AOI22_X1 U9473 ( .A1(n8843), .A2(n8741), .B1(n8740), .B2(n9160), .ZN(n7792)
         );
  INV_X1 U9474 ( .A(n7768), .ZN(n7769) );
  AOI22_X1 U9475 ( .A1(n8731), .A2(n8645), .B1(n8741), .B2(n9163), .ZN(n7772)
         );
  XNOR2_X1 U9476 ( .A(n7772), .B(n8674), .ZN(n7773) );
  OAI22_X1 U9477 ( .A1(n5954), .A2(n8651), .B1(n5953), .B2(n8680), .ZN(n8726)
         );
  INV_X1 U9478 ( .A(n8726), .ZN(n7775) );
  NAND2_X1 U9479 ( .A1(n8862), .A2(n8735), .ZN(n7778) );
  NAND2_X1 U9480 ( .A1(n9162), .A2(n8741), .ZN(n7777) );
  NAND2_X1 U9481 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  XNOR2_X1 U9482 ( .A(n7779), .B(n8674), .ZN(n7782) );
  NAND2_X1 U9483 ( .A1(n8862), .A2(n8741), .ZN(n7781) );
  NAND2_X1 U9484 ( .A1(n8740), .A2(n9162), .ZN(n7780) );
  NAND2_X1 U9485 ( .A1(n7781), .A2(n7780), .ZN(n7783) );
  NAND2_X1 U9486 ( .A1(n7782), .A2(n7783), .ZN(n8857) );
  INV_X1 U9487 ( .A(n7782), .ZN(n7785) );
  INV_X1 U9488 ( .A(n7783), .ZN(n7784) );
  NAND2_X1 U9489 ( .A1(n7785), .A2(n7784), .ZN(n8856) );
  NAND2_X1 U9490 ( .A1(n8768), .A2(n8735), .ZN(n7787) );
  NAND2_X1 U9491 ( .A1(n9161), .A2(n8741), .ZN(n7786) );
  NAND2_X1 U9492 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  XNOR2_X1 U9493 ( .A(n7788), .B(n8674), .ZN(n7791) );
  AOI22_X1 U9494 ( .A1(n8768), .A2(n8741), .B1(n8740), .B2(n9161), .ZN(n7789)
         );
  XNOR2_X1 U9495 ( .A(n7791), .B(n7789), .ZN(n8762) );
  INV_X1 U9496 ( .A(n7789), .ZN(n7790) );
  XNOR2_X1 U9497 ( .A(n7794), .B(n7792), .ZN(n8838) );
  NAND2_X1 U9498 ( .A1(n8837), .A2(n8838), .ZN(n7793) );
  AOI22_X1 U9499 ( .A1(n9647), .A2(n8735), .B1(n8741), .B2(n9529), .ZN(n7795)
         );
  XNOR2_X1 U9500 ( .A(n7795), .B(n8674), .ZN(n7796) );
  AOI22_X1 U9501 ( .A1(n9647), .A2(n8741), .B1(n8740), .B2(n9529), .ZN(n8709)
         );
  NAND2_X1 U9502 ( .A1(n9637), .A2(n8735), .ZN(n7798) );
  NAND2_X1 U9503 ( .A1(n9527), .A2(n8741), .ZN(n7797) );
  NAND2_X1 U9504 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  XNOR2_X1 U9505 ( .A(n7799), .B(n8674), .ZN(n8788) );
  NAND2_X1 U9506 ( .A1(n9637), .A2(n8741), .ZN(n7801) );
  NAND2_X1 U9507 ( .A1(n8740), .A2(n9527), .ZN(n7800) );
  NAND2_X1 U9508 ( .A1(n7801), .A2(n7800), .ZN(n7809) );
  NAND2_X1 U9509 ( .A1(n9535), .A2(n8735), .ZN(n7803) );
  NAND2_X1 U9510 ( .A1(n9159), .A2(n8736), .ZN(n7802) );
  NAND2_X1 U9511 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  XNOR2_X1 U9512 ( .A(n7804), .B(n8678), .ZN(n8786) );
  NOR2_X1 U9513 ( .A1(n9550), .A2(n8680), .ZN(n7805) );
  AOI21_X1 U9514 ( .B1(n9535), .B2(n8741), .A(n7805), .ZN(n8784) );
  NAND2_X1 U9515 ( .A1(n8786), .A2(n8784), .ZN(n7808) );
  INV_X1 U9516 ( .A(n7808), .ZN(n7811) );
  INV_X1 U9517 ( .A(n7809), .ZN(n8787) );
  AOI21_X1 U9518 ( .B1(n7809), .B2(n7808), .A(n8788), .ZN(n7810) );
  AOI21_X1 U9519 ( .B1(n7811), .B2(n8787), .A(n7810), .ZN(n8809) );
  NAND2_X1 U9520 ( .A1(n9498), .A2(n8735), .ZN(n7813) );
  NAND2_X1 U9521 ( .A1(n9158), .A2(n8741), .ZN(n7812) );
  NAND2_X1 U9522 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  XNOR2_X1 U9523 ( .A(n7814), .B(n8674), .ZN(n7823) );
  INV_X1 U9524 ( .A(n7823), .ZN(n7815) );
  AOI22_X1 U9525 ( .A1(n9498), .A2(n8741), .B1(n8740), .B2(n9158), .ZN(n7822)
         );
  NAND2_X1 U9526 ( .A1(n7815), .A2(n7822), .ZN(n7821) );
  AND2_X1 U9527 ( .A1(n8809), .A2(n7821), .ZN(n8866) );
  NAND2_X1 U9528 ( .A1(n9625), .A2(n8735), .ZN(n7817) );
  NAND2_X1 U9529 ( .A1(n9492), .A2(n8741), .ZN(n7816) );
  NAND2_X1 U9530 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  XNOR2_X1 U9531 ( .A(n7818), .B(n8674), .ZN(n7826) );
  INV_X1 U9532 ( .A(n7826), .ZN(n7819) );
  AOI22_X1 U9533 ( .A1(n9625), .A2(n8741), .B1(n8740), .B2(n9492), .ZN(n7825)
         );
  NAND2_X1 U9534 ( .A1(n7819), .A2(n7825), .ZN(n7820) );
  AND2_X1 U9535 ( .A1(n8866), .A2(n7820), .ZN(n8626) );
  NAND2_X1 U9536 ( .A1(n8867), .A2(n8626), .ZN(n7829) );
  INV_X1 U9537 ( .A(n7820), .ZN(n7828) );
  INV_X1 U9538 ( .A(n7821), .ZN(n7824) );
  XNOR2_X1 U9539 ( .A(n7823), .B(n7822), .ZN(n8811) );
  OR2_X1 U9540 ( .A1(n7824), .A2(n8811), .ZN(n8868) );
  XNOR2_X1 U9541 ( .A(n7826), .B(n7825), .ZN(n8871) );
  AND2_X1 U9542 ( .A1(n8868), .A2(n8871), .ZN(n7827) );
  AND2_X1 U9543 ( .A1(n7829), .A2(n8628), .ZN(n7836) );
  NAND2_X1 U9544 ( .A1(n9470), .A2(n8735), .ZN(n7831) );
  NAND2_X1 U9545 ( .A1(n9453), .A2(n8741), .ZN(n7830) );
  NAND2_X1 U9546 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  XNOR2_X1 U9547 ( .A(n7832), .B(n8674), .ZN(n8631) );
  NAND2_X1 U9548 ( .A1(n9470), .A2(n8741), .ZN(n7834) );
  NAND2_X1 U9549 ( .A1(n9453), .A2(n8740), .ZN(n7833) );
  NAND2_X1 U9550 ( .A1(n7834), .A2(n7833), .ZN(n8630) );
  XNOR2_X1 U9551 ( .A(n8631), .B(n8630), .ZN(n7835) );
  XNOR2_X1 U9552 ( .A(n7836), .B(n7835), .ZN(n7841) );
  AOI22_X1 U9553 ( .A1(n8801), .A2(n9492), .B1(n8800), .B2(n9471), .ZN(n7837)
         );
  NAND2_X1 U9554 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9282) );
  OAI211_X1 U9555 ( .C1(n7838), .C2(n8890), .A(n7837), .B(n9282), .ZN(n7839)
         );
  AOI21_X1 U9556 ( .B1(n9470), .B2(n8897), .A(n7839), .ZN(n7840) );
  OAI21_X1 U9557 ( .B1(n7841), .B2(n8899), .A(n7840), .ZN(P1_U3219) );
  XOR2_X1 U9558 ( .A(n7843), .B(n7842), .Z(n8458) );
  OR2_X1 U9559 ( .A1(n9975), .A2(n9967), .ZN(n8602) );
  INV_X1 U9560 ( .A(n7875), .ZN(n8246) );
  INV_X1 U9561 ( .A(n8264), .ZN(n8073) );
  AOI21_X2 U9562 ( .B1(n7848), .B2(n8413), .A(n7847), .ZN(n8250) );
  OAI21_X1 U9563 ( .B1(n8246), .B2(n9961), .A(n8250), .ZN(n8455) );
  MUX2_X1 U9564 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8455), .S(n9973), .Z(n7849)
         );
  INV_X1 U9565 ( .A(n7849), .ZN(n7850) );
  OAI21_X1 U9566 ( .B1(n8458), .B2(n8602), .A(n7850), .ZN(P2_U3454) );
  INV_X1 U9567 ( .A(n8994), .ZN(n7860) );
  OAI222_X1 U9568 ( .A1(n9709), .A2(n8995), .B1(n9707), .B2(n7860), .C1(
        P1_U3086), .C2(n7851), .ZN(P1_U3325) );
  NAND2_X1 U9569 ( .A1(n7853), .A2(n8389), .ZN(n8228) );
  NAND2_X1 U9570 ( .A1(n8421), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7854) );
  OAI211_X1 U9571 ( .C1(n7855), .C2(n8352), .A(n8228), .B(n7854), .ZN(n7856)
         );
  AOI21_X1 U9572 ( .B1(n7857), .B2(n8419), .A(n7856), .ZN(n7858) );
  OAI21_X1 U9573 ( .B1(n7852), .B2(n8421), .A(n7858), .ZN(P2_U3204) );
  OAI222_X1 U9574 ( .A1(n8612), .A2(n7862), .B1(n7861), .B2(n7860), .C1(
        P2_U3151), .C2(n7859), .ZN(P2_U3265) );
  OAI21_X1 U9575 ( .B1(n7865), .B2(n7864), .A(n7863), .ZN(n7866) );
  NAND2_X1 U9576 ( .A1(n7866), .A2(n8048), .ZN(n7874) );
  AOI21_X1 U9577 ( .B1(n8042), .B2(n7868), .A(n7867), .ZN(n7873) );
  AOI22_X1 U9578 ( .A1(n8030), .A2(n8081), .B1(n8061), .B2(n8083), .ZN(n7872)
         );
  INV_X1 U9579 ( .A(n7869), .ZN(n7870) );
  NAND2_X1 U9580 ( .A1(n8066), .A2(n7870), .ZN(n7871) );
  NAND4_X1 U9581 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(
        P2_U3153) );
  INV_X1 U9582 ( .A(n8042), .ZN(n8069) );
  XNOR2_X1 U9583 ( .A(n7875), .B(n4414), .ZN(n7941) );
  XNOR2_X1 U9584 ( .A(n7941), .B(n8256), .ZN(n7912) );
  INV_X1 U9585 ( .A(n7912), .ZN(n7914) );
  XNOR2_X1 U9586 ( .A(n8532), .B(n4414), .ZN(n7906) );
  INV_X1 U9587 ( .A(n7906), .ZN(n7907) );
  INV_X1 U9588 ( .A(n7876), .ZN(n7878) );
  XNOR2_X1 U9589 ( .A(n8581), .B(n4414), .ZN(n7881) );
  XNOR2_X1 U9590 ( .A(n7881), .B(n8396), .ZN(n8057) );
  OR2_X2 U9591 ( .A1(n8055), .A2(n8057), .ZN(n8058) );
  NAND2_X1 U9592 ( .A1(n7881), .A2(n8396), .ZN(n7882) );
  XNOR2_X1 U9593 ( .A(n8576), .B(n4414), .ZN(n7968) );
  NAND2_X1 U9594 ( .A1(n7970), .A2(n7968), .ZN(n7884) );
  INV_X1 U9595 ( .A(n8064), .ZN(n8386) );
  XNOR2_X1 U9596 ( .A(n8570), .B(n6674), .ZN(n7885) );
  NAND2_X1 U9597 ( .A1(n7885), .A2(n8346), .ZN(n7987) );
  INV_X1 U9598 ( .A(n7885), .ZN(n7886) );
  INV_X1 U9599 ( .A(n8346), .ZN(n8375) );
  NAND2_X1 U9600 ( .A1(n7886), .A2(n8375), .ZN(n7988) );
  XNOR2_X1 U9601 ( .A(n8567), .B(n4414), .ZN(n7889) );
  XNOR2_X1 U9602 ( .A(n7889), .B(n8335), .ZN(n8037) );
  XNOR2_X1 U9603 ( .A(n8559), .B(n6674), .ZN(n7888) );
  INV_X1 U9604 ( .A(n7888), .ZN(n7887) );
  INV_X1 U9605 ( .A(n8347), .ZN(n8078) );
  OR2_X1 U9606 ( .A1(n8037), .A2(n4438), .ZN(n7891) );
  XNOR2_X1 U9607 ( .A(n7888), .B(n8347), .ZN(n7929) );
  INV_X1 U9608 ( .A(n7929), .ZN(n7890) );
  NAND2_X1 U9609 ( .A1(n7889), .A2(n8335), .ZN(n7928) );
  AND2_X1 U9610 ( .A1(n7890), .A2(n7928), .ZN(n7931) );
  XNOR2_X1 U9611 ( .A(n8323), .B(n4414), .ZN(n7892) );
  NAND2_X1 U9612 ( .A1(n7892), .A2(n8077), .ZN(n8017) );
  NAND2_X1 U9613 ( .A1(n8020), .A2(n8017), .ZN(n7894) );
  INV_X1 U9614 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U9615 ( .A1(n7893), .A2(n8334), .ZN(n8018) );
  NAND2_X1 U9616 ( .A1(n7894), .A2(n8018), .ZN(n7952) );
  XNOR2_X1 U9617 ( .A(n5530), .B(n4414), .ZN(n7895) );
  XNOR2_X1 U9618 ( .A(n7895), .B(n8320), .ZN(n7953) );
  INV_X1 U9619 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9620 ( .A1(n7896), .A2(n8320), .ZN(n7897) );
  XNOR2_X1 U9621 ( .A(n8026), .B(n4414), .ZN(n7898) );
  XNOR2_X1 U9622 ( .A(n7898), .B(n8076), .ZN(n8027) );
  XNOR2_X1 U9623 ( .A(n8290), .B(n4414), .ZN(n7900) );
  NOR2_X1 U9624 ( .A1(n7899), .A2(n7900), .ZN(n7920) );
  INV_X1 U9625 ( .A(n7900), .ZN(n7901) );
  XNOR2_X1 U9626 ( .A(n8537), .B(n4414), .ZN(n7903) );
  NAND2_X1 U9627 ( .A1(n7903), .A2(n8284), .ZN(n7959) );
  INV_X1 U9628 ( .A(n7903), .ZN(n7904) );
  INV_X1 U9629 ( .A(n8284), .ZN(n8074) );
  NAND2_X1 U9630 ( .A1(n7904), .A2(n8074), .ZN(n7905) );
  XNOR2_X1 U9631 ( .A(n7906), .B(n8255), .ZN(n7960) );
  XNOR2_X1 U9632 ( .A(n8054), .B(n4414), .ZN(n7908) );
  XNOR2_X1 U9633 ( .A(n7910), .B(n7908), .ZN(n8047) );
  NAND2_X1 U9634 ( .A1(n8047), .A2(n8264), .ZN(n8046) );
  INV_X1 U9635 ( .A(n7908), .ZN(n7909) );
  OR2_X2 U9636 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  INV_X1 U9637 ( .A(n7943), .ZN(n7913) );
  AOI22_X1 U9638 ( .A1(n8073), .A2(n8061), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7915) );
  OAI21_X1 U9639 ( .B1(n7916), .B2(n8063), .A(n7915), .ZN(n7917) );
  AOI21_X1 U9640 ( .B1(n8244), .B2(n8066), .A(n7917), .ZN(n7918) );
  OAI211_X1 U9641 ( .C1(n8246), .C2(n8069), .A(n7919), .B(n7918), .ZN(P2_U3154) );
  INV_X1 U9642 ( .A(n7999), .ZN(n7922) );
  OAI21_X1 U9643 ( .B1(n7920), .B2(n7998), .A(n8075), .ZN(n7921) );
  OAI21_X1 U9644 ( .B1(n7922), .B2(n7998), .A(n7921), .ZN(n7923) );
  NAND2_X1 U9645 ( .A1(n7923), .A2(n8048), .ZN(n7927) );
  AOI22_X1 U9646 ( .A1(n8074), .A2(n8030), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7924) );
  OAI21_X1 U9647 ( .B1(n8308), .B2(n8032), .A(n7924), .ZN(n7925) );
  AOI21_X1 U9648 ( .B1(n8288), .B2(n8066), .A(n7925), .ZN(n7926) );
  OAI211_X1 U9649 ( .C1(n8290), .C2(n8069), .A(n7927), .B(n7926), .ZN(P2_U3156) );
  OR2_X1 U9650 ( .A1(n8036), .A2(n8037), .ZN(n7932) );
  NAND2_X1 U9651 ( .A1(n7932), .A2(n7928), .ZN(n7930) );
  AOI21_X1 U9652 ( .B1(n7930), .B2(n7929), .A(n8056), .ZN(n7934) );
  NAND2_X1 U9653 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U9654 ( .A1(n7934), .A2(n7933), .ZN(n7939) );
  INV_X1 U9655 ( .A(n7935), .ZN(n8340) );
  INV_X1 U9656 ( .A(n8335), .ZN(n8363) );
  NAND2_X1 U9657 ( .A1(n8061), .A2(n8363), .ZN(n7936) );
  NAND2_X1 U9658 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8214) );
  OAI211_X1 U9659 ( .C1(n8334), .C2(n8063), .A(n7936), .B(n8214), .ZN(n7937)
         );
  AOI21_X1 U9660 ( .B1(n8340), .B2(n8066), .A(n7937), .ZN(n7938) );
  OAI211_X1 U9661 ( .C1(n7940), .C2(n8069), .A(n7939), .B(n7938), .ZN(P2_U3159) );
  XNOR2_X1 U9662 ( .A(n8234), .B(n4414), .ZN(n7944) );
  XNOR2_X1 U9663 ( .A(n7945), .B(n7944), .ZN(n7950) );
  AOI22_X1 U9664 ( .A1(n8256), .A2(n8061), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7947) );
  NAND2_X1 U9665 ( .A1(n8241), .A2(n8066), .ZN(n7946) );
  OAI211_X1 U9666 ( .C1(n8237), .C2(n8063), .A(n7947), .B(n7946), .ZN(n7948)
         );
  AOI21_X1 U9667 ( .B1(n8520), .B2(n8042), .A(n7948), .ZN(n7949) );
  OAI21_X1 U9668 ( .B1(n7950), .B2(n8056), .A(n7949), .ZN(P2_U3160) );
  OAI21_X1 U9669 ( .B1(n7953), .B2(n7952), .A(n7951), .ZN(n7954) );
  NAND2_X1 U9670 ( .A1(n7954), .A2(n8048), .ZN(n7958) );
  AOI22_X1 U9671 ( .A1(n8030), .A2(n8076), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7955) );
  OAI21_X1 U9672 ( .B1(n8334), .B2(n8032), .A(n7955), .ZN(n7956) );
  AOI21_X1 U9673 ( .B1(n8313), .B2(n8066), .A(n7956), .ZN(n7957) );
  OAI211_X1 U9674 ( .C1(n8552), .C2(n8069), .A(n7958), .B(n7957), .ZN(P2_U3163) );
  INV_X1 U9675 ( .A(n8532), .ZN(n7967) );
  AND3_X1 U9676 ( .A1(n7996), .A2(n7960), .A3(n7959), .ZN(n7961) );
  OAI21_X1 U9677 ( .B1(n7962), .B2(n7961), .A(n8048), .ZN(n7966) );
  AOI22_X1 U9678 ( .A1(n8073), .A2(n8030), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7963) );
  OAI21_X1 U9679 ( .B1(n8284), .B2(n8032), .A(n7963), .ZN(n7964) );
  AOI21_X1 U9680 ( .B1(n8265), .B2(n8066), .A(n7964), .ZN(n7965) );
  OAI211_X1 U9681 ( .C1(n7967), .C2(n8069), .A(n7966), .B(n7965), .ZN(P2_U3165) );
  XNOR2_X1 U9682 ( .A(n7968), .B(n8064), .ZN(n7969) );
  XNOR2_X1 U9683 ( .A(n7970), .B(n7969), .ZN(n7976) );
  NAND2_X1 U9684 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8136) );
  OAI21_X1 U9685 ( .B1(n8032), .B2(n7971), .A(n8136), .ZN(n7972) );
  AOI21_X1 U9686 ( .B1(n8030), .B2(n8375), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9687 ( .B1(n8378), .B2(n8040), .A(n7973), .ZN(n7974) );
  AOI21_X1 U9688 ( .B1(n8576), .B2(n8042), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9689 ( .B1(n7976), .B2(n8056), .A(n7975), .ZN(P2_U3166) );
  XNOR2_X1 U9690 ( .A(n7978), .B(n7977), .ZN(n7979) );
  NAND2_X1 U9691 ( .A1(n7979), .A2(n8048), .ZN(n7986) );
  AOI22_X1 U9692 ( .A1(n8042), .A2(n7980), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3151), .ZN(n7985) );
  AOI22_X1 U9693 ( .A1(n8030), .A2(n8083), .B1(n8061), .B2(n8085), .ZN(n7984)
         );
  INV_X1 U9694 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U9695 ( .A1(n8066), .A2(n7982), .ZN(n7983) );
  NAND4_X1 U9696 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(
        P2_U3167) );
  NAND2_X1 U9697 ( .A1(n7988), .A2(n7987), .ZN(n7990) );
  XOR2_X1 U9698 ( .A(n7990), .B(n7989), .Z(n7995) );
  AND2_X1 U9699 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8161) );
  NOR2_X1 U9700 ( .A1(n8063), .A2(n8335), .ZN(n7991) );
  AOI211_X1 U9701 ( .C1(n8061), .C2(n8386), .A(n8161), .B(n7991), .ZN(n7992)
         );
  OAI21_X1 U9702 ( .B1(n8366), .B2(n8040), .A(n7992), .ZN(n7993) );
  AOI21_X1 U9703 ( .B1(n8570), .B2(n8042), .A(n7993), .ZN(n7994) );
  OAI21_X1 U9704 ( .B1(n7995), .B2(n8056), .A(n7994), .ZN(P2_U3168) );
  INV_X1 U9705 ( .A(n7996), .ZN(n8001) );
  NOR3_X1 U9706 ( .A1(n7999), .A2(n7998), .A3(n7997), .ZN(n8000) );
  OAI21_X1 U9707 ( .B1(n8001), .B2(n8000), .A(n8048), .ZN(n8005) );
  AOI22_X1 U9708 ( .A1(n8255), .A2(n8030), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8002) );
  OAI21_X1 U9709 ( .B1(n8298), .B2(n8032), .A(n8002), .ZN(n8003) );
  AOI21_X1 U9710 ( .B1(n8275), .B2(n8066), .A(n8003), .ZN(n8004) );
  OAI211_X1 U9711 ( .C1(n8537), .C2(n8069), .A(n8005), .B(n8004), .ZN(P2_U3169) );
  OAI21_X1 U9712 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n8009) );
  NAND2_X1 U9713 ( .A1(n8009), .A2(n8048), .ZN(n8016) );
  AOI21_X1 U9714 ( .B1(n8042), .B2(n8011), .A(n8010), .ZN(n8015) );
  AOI22_X1 U9715 ( .A1(n8030), .A2(n8084), .B1(n8061), .B2(n5246), .ZN(n8014)
         );
  NAND2_X1 U9716 ( .A1(n8066), .A2(n8012), .ZN(n8013) );
  NAND4_X1 U9717 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(
        P2_U3170) );
  NAND2_X1 U9718 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  XNOR2_X1 U9719 ( .A(n8020), .B(n8019), .ZN(n8025) );
  AOI22_X1 U9720 ( .A1(n8061), .A2(n8078), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8022) );
  NAND2_X1 U9721 ( .A1(n8066), .A2(n8324), .ZN(n8021) );
  OAI211_X1 U9722 ( .C1(n8320), .C2(n8063), .A(n8022), .B(n8021), .ZN(n8023)
         );
  AOI21_X1 U9723 ( .B1(n8323), .B2(n8042), .A(n8023), .ZN(n8024) );
  OAI21_X1 U9724 ( .B1(n8025), .B2(n8056), .A(n8024), .ZN(P2_U3173) );
  INV_X1 U9725 ( .A(n8026), .ZN(n8548) );
  AOI21_X1 U9726 ( .B1(n8028), .B2(n8027), .A(n8056), .ZN(n8029) );
  NAND2_X1 U9727 ( .A1(n8029), .A2(n4488), .ZN(n8035) );
  AOI22_X1 U9728 ( .A1(n8075), .A2(n8030), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8031) );
  OAI21_X1 U9729 ( .B1(n8320), .B2(n8032), .A(n8031), .ZN(n8033) );
  AOI21_X1 U9730 ( .B1(n8301), .B2(n8066), .A(n8033), .ZN(n8034) );
  OAI211_X1 U9731 ( .C1(n8548), .C2(n8069), .A(n8035), .B(n8034), .ZN(P2_U3175) );
  XOR2_X1 U9732 ( .A(n8037), .B(n8036), .Z(n8045) );
  INV_X1 U9733 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8187) );
  OAI22_X1 U9734 ( .A1(n8063), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8187), .ZN(n8038) );
  AOI21_X1 U9735 ( .B1(n8061), .B2(n8375), .A(n8038), .ZN(n8039) );
  OAI21_X1 U9736 ( .B1(n8353), .B2(n8040), .A(n8039), .ZN(n8041) );
  AOI21_X1 U9737 ( .B1(n8043), .B2(n8042), .A(n8041), .ZN(n8044) );
  OAI21_X1 U9738 ( .B1(n8045), .B2(n8056), .A(n8044), .ZN(P2_U3178) );
  OAI21_X1 U9739 ( .B1(n8264), .B2(n8047), .A(n8046), .ZN(n8049) );
  NAND2_X1 U9740 ( .A1(n8049), .A2(n8048), .ZN(n8053) );
  AOI22_X1 U9741 ( .A1(n8255), .A2(n8061), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8050) );
  OAI21_X1 U9742 ( .B1(n8236), .B2(n8063), .A(n8050), .ZN(n8051) );
  AOI21_X1 U9743 ( .B1(n8259), .B2(n8066), .A(n8051), .ZN(n8052) );
  OAI211_X1 U9744 ( .C1(n8054), .C2(n8069), .A(n8053), .B(n8052), .ZN(P2_U3180) );
  INV_X1 U9745 ( .A(n8581), .ZN(n8070) );
  AOI21_X1 U9746 ( .B1(n8055), .B2(n8057), .A(n8056), .ZN(n8059) );
  NAND2_X1 U9747 ( .A1(n8059), .A2(n8058), .ZN(n8068) );
  INV_X1 U9748 ( .A(n8060), .ZN(n8388) );
  NAND2_X1 U9749 ( .A1(n8061), .A2(n8411), .ZN(n8062) );
  NAND2_X1 U9750 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8114) );
  OAI211_X1 U9751 ( .C1(n8064), .C2(n8063), .A(n8062), .B(n8114), .ZN(n8065)
         );
  AOI21_X1 U9752 ( .B1(n8388), .B2(n8066), .A(n8065), .ZN(n8067) );
  OAI211_X1 U9753 ( .C1(n8070), .C2(n8069), .A(n8068), .B(n8067), .ZN(P2_U3181) );
  MUX2_X1 U9754 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8071), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9755 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8072), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9756 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8256), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9757 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8073), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9758 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8255), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9759 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8074), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9760 ( .A(n8075), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8185), .Z(
        P2_U3514) );
  MUX2_X1 U9761 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8076), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9762 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8077), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9763 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8078), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9764 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8363), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9765 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8375), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9766 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8386), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9767 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8396), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9768 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8411), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9769 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8409), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9770 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8079), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9771 ( .A(n8080), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8185), .Z(
        P2_U3501) );
  MUX2_X1 U9772 ( .A(n8081), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8185), .Z(
        P2_U3499) );
  MUX2_X1 U9773 ( .A(n8082), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8185), .Z(
        P2_U3498) );
  MUX2_X1 U9774 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8083), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9775 ( .A(n8084), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8185), .Z(
        P2_U3496) );
  MUX2_X1 U9776 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8085), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9777 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n5246), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9778 ( .A(n5229), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8185), .Z(
        P2_U3493) );
  MUX2_X1 U9779 ( .A(n8086), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8185), .Z(
        P2_U3492) );
  AOI21_X1 U9780 ( .B1(n8503), .B2(n8088), .A(n8087), .ZN(n8102) );
  OAI21_X1 U9781 ( .B1(n8091), .B2(n8090), .A(n8089), .ZN(n8100) );
  INV_X1 U9782 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10155) );
  AOI21_X1 U9783 ( .B1(n8093), .B2(n5396), .A(n8092), .ZN(n8094) );
  NOR2_X1 U9784 ( .A1(n8221), .A2(n8094), .ZN(n8095) );
  AOI211_X1 U9785 ( .C1(n8097), .C2(n9881), .A(n8096), .B(n8095), .ZN(n8098)
         );
  OAI21_X1 U9786 ( .B1(n10155), .B2(n9887), .A(n8098), .ZN(n8099) );
  AOI21_X1 U9787 ( .B1(n9872), .B2(n8100), .A(n8099), .ZN(n8101) );
  OAI21_X1 U9788 ( .B1(n8102), .B2(n8224), .A(n8101), .ZN(P2_U3195) );
  AOI21_X1 U9789 ( .B1(n10199), .B2(n8104), .A(n8124), .ZN(n8122) );
  MUX2_X1 U9790 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8208), .Z(n8129) );
  XNOR2_X1 U9791 ( .A(n8129), .B(n8138), .ZN(n8109) );
  OR2_X1 U9792 ( .A1(n8105), .A2(n8111), .ZN(n8107) );
  NAND2_X1 U9793 ( .A1(n8107), .A2(n8106), .ZN(n8108) );
  NAND2_X1 U9794 ( .A1(n8109), .A2(n8108), .ZN(n8131) );
  OAI21_X1 U9795 ( .B1(n8109), .B2(n8108), .A(n8131), .ZN(n8120) );
  INV_X1 U9796 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8112) );
  AOI21_X1 U9797 ( .B1(n8113), .B2(n8112), .A(n8139), .ZN(n8116) );
  NAND2_X1 U9798 ( .A1(n9881), .A2(n8138), .ZN(n8115) );
  OAI211_X1 U9799 ( .C1(n8116), .C2(n8221), .A(n8115), .B(n8114), .ZN(n8119)
         );
  NOR2_X1 U9800 ( .A1(n9887), .A2(n8117), .ZN(n8118) );
  AOI211_X1 U9801 ( .C1(n9872), .C2(n8120), .A(n8119), .B(n8118), .ZN(n8121)
         );
  OAI21_X1 U9802 ( .B1(n8122), .B2(n8224), .A(n8121), .ZN(P2_U3197) );
  NAND2_X1 U9803 ( .A1(n8155), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8164) );
  INV_X1 U9804 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U9805 ( .A1(n8141), .A2(n8495), .ZN(n8125) );
  NAND2_X1 U9806 ( .A1(n8164), .A2(n8125), .ZN(n8127) );
  INV_X1 U9807 ( .A(n8165), .ZN(n8126) );
  AOI21_X1 U9808 ( .B1(n8128), .B2(n8127), .A(n8126), .ZN(n8150) );
  MUX2_X1 U9809 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8208), .Z(n8156) );
  XNOR2_X1 U9810 ( .A(n8156), .B(n8141), .ZN(n8134) );
  INV_X1 U9811 ( .A(n8129), .ZN(n8130) );
  NAND2_X1 U9812 ( .A1(n8138), .A2(n8130), .ZN(n8132) );
  NAND2_X1 U9813 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  NAND2_X1 U9814 ( .A1(n8134), .A2(n8133), .ZN(n8157) );
  OAI21_X1 U9815 ( .B1(n8134), .B2(n8133), .A(n8157), .ZN(n8148) );
  INV_X1 U9816 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U9817 ( .A1(n9881), .A2(n8141), .ZN(n8135) );
  OAI211_X1 U9818 ( .C1(n9887), .C2(n10269), .A(n8136), .B(n8135), .ZN(n8147)
         );
  NOR2_X1 U9819 ( .A1(n8138), .A2(n8137), .ZN(n8140) );
  NOR2_X1 U9820 ( .A1(n8140), .A2(n8139), .ZN(n8144) );
  NAND2_X1 U9821 ( .A1(n8155), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U9822 ( .A1(n8141), .A2(n8377), .ZN(n8142) );
  NAND2_X1 U9823 ( .A1(n8151), .A2(n8142), .ZN(n8143) );
  OR2_X1 U9824 ( .A1(n8144), .A2(n8143), .ZN(n8152) );
  NAND2_X1 U9825 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  AOI21_X1 U9826 ( .B1(n8152), .B2(n8145), .A(n8221), .ZN(n8146) );
  AOI211_X1 U9827 ( .C1(n9872), .C2(n8148), .A(n8147), .B(n8146), .ZN(n8149)
         );
  OAI21_X1 U9828 ( .B1(n8150), .B2(n8224), .A(n8149), .ZN(P2_U3198) );
  XNOR2_X1 U9829 ( .A(n8190), .B(n8191), .ZN(n8153) );
  NOR2_X1 U9830 ( .A1(n8365), .A2(n8153), .ZN(n8192) );
  AOI21_X1 U9831 ( .B1(n8153), .B2(n8365), .A(n8192), .ZN(n8172) );
  MUX2_X1 U9832 ( .A(n8365), .B(n8492), .S(n8208), .Z(n8180) );
  XNOR2_X1 U9833 ( .A(n8180), .B(n8154), .ZN(n8160) );
  OR2_X1 U9834 ( .A1(n8156), .A2(n8155), .ZN(n8158) );
  NAND2_X1 U9835 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U9836 ( .A1(n8160), .A2(n8159), .ZN(n8178) );
  OAI21_X1 U9837 ( .B1(n8160), .B2(n8159), .A(n8178), .ZN(n8170) );
  AOI21_X1 U9838 ( .B1(n9881), .B2(n8191), .A(n8161), .ZN(n8162) );
  OAI21_X1 U9839 ( .B1(n9887), .B2(n8163), .A(n8162), .ZN(n8169) );
  XNOR2_X1 U9840 ( .A(n8191), .B(n8173), .ZN(n8166) );
  NOR2_X1 U9841 ( .A1(n8167), .A2(n8224), .ZN(n8168) );
  AOI211_X1 U9842 ( .C1(n9872), .C2(n8170), .A(n8169), .B(n8168), .ZN(n8171)
         );
  OAI21_X1 U9843 ( .B1(n8172), .B2(n8221), .A(n8171), .ZN(P2_U3199) );
  NOR2_X1 U9844 ( .A1(n8191), .A2(n8173), .ZN(n8175) );
  NOR2_X1 U9845 ( .A1(n8175), .A2(n8174), .ZN(n8177) );
  NAND2_X1 U9846 ( .A1(n8194), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8200) );
  OAI21_X1 U9847 ( .B1(n8194), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8200), .ZN(
        n8176) );
  NOR2_X1 U9848 ( .A1(n8177), .A2(n8176), .ZN(n8202) );
  AOI21_X1 U9849 ( .B1(n8177), .B2(n8176), .A(n8202), .ZN(n8199) );
  INV_X1 U9850 ( .A(n8178), .ZN(n8179) );
  MUX2_X1 U9851 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8208), .Z(n8181) );
  INV_X1 U9852 ( .A(n8205), .ZN(n8183) );
  NAND2_X1 U9853 ( .A1(n8182), .A2(n8181), .ZN(n8206) );
  NAND2_X1 U9854 ( .A1(n8183), .A2(n8206), .ZN(n8186) );
  OAI21_X1 U9855 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(n8198) );
  NAND3_X1 U9856 ( .A1(n8186), .A2(n9872), .A3(n8194), .ZN(n8189) );
  OR2_X1 U9857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8187), .ZN(n8188) );
  OAI211_X1 U9858 ( .C1(n10292), .C2(n9887), .A(n8189), .B(n8188), .ZN(n8197)
         );
  NOR2_X1 U9859 ( .A1(n8191), .A2(n8190), .ZN(n8193) );
  NOR2_X1 U9860 ( .A1(n8193), .A2(n8192), .ZN(n8196) );
  NAND2_X1 U9861 ( .A1(n8194), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8216) );
  OAI21_X1 U9862 ( .B1(n8194), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8216), .ZN(
        n8195) );
  NOR2_X1 U9863 ( .A1(n8196), .A2(n8195), .ZN(n8218) );
  INV_X1 U9864 ( .A(n8200), .ZN(n8201) );
  NOR2_X1 U9865 ( .A1(n8202), .A2(n8201), .ZN(n8204) );
  XNOR2_X1 U9866 ( .A(n8212), .B(n8484), .ZN(n8209) );
  INV_X1 U9867 ( .A(n8209), .ZN(n8203) );
  XNOR2_X1 U9868 ( .A(n8204), .B(n8203), .ZN(n8225) );
  MUX2_X1 U9869 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8339), .S(n8212), .Z(n8220)
         );
  MUX2_X1 U9870 ( .A(n8220), .B(n8209), .S(n8208), .Z(n8210) );
  XNOR2_X1 U9871 ( .A(n8211), .B(n8210), .ZN(n8223) );
  INV_X1 U9872 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U9873 ( .A1(n9881), .A2(n8212), .ZN(n8213) );
  OAI211_X1 U9874 ( .C1(n9887), .C2(n8215), .A(n8214), .B(n8213), .ZN(n8222)
         );
  INV_X1 U9875 ( .A(n8216), .ZN(n8217) );
  NOR2_X1 U9876 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  OR2_X1 U9877 ( .A1(n8227), .A2(n8226), .ZN(n8513) );
  OAI21_X1 U9878 ( .B1(n8421), .B2(n8513), .A(n8228), .ZN(n8230) );
  AOI21_X1 U9879 ( .B1(n8421), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8230), .ZN(
        n8229) );
  OAI21_X1 U9880 ( .B1(n8515), .B2(n8352), .A(n8229), .ZN(P2_U3202) );
  AOI21_X1 U9881 ( .B1(n8421), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8230), .ZN(
        n8231) );
  OAI21_X1 U9882 ( .B1(n8518), .B2(n8352), .A(n8231), .ZN(P2_U3203) );
  INV_X1 U9883 ( .A(n8234), .ZN(n8232) );
  INV_X1 U9884 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U9885 ( .A(n8235), .B(n8234), .ZN(n8239) );
  OAI22_X1 U9886 ( .A1(n8237), .A2(n9909), .B1(n8236), .B2(n9910), .ZN(n8238)
         );
  MUX2_X1 U9887 ( .A(n8240), .B(n8519), .S(n9913), .Z(n8243) );
  AOI22_X1 U9888 ( .A1(n8520), .A2(n8445), .B1(n8389), .B2(n8241), .ZN(n8242)
         );
  OAI211_X1 U9889 ( .C1(n8523), .C2(n8448), .A(n8243), .B(n8242), .ZN(P2_U3205) );
  INV_X1 U9890 ( .A(n8458), .ZN(n8248) );
  AOI22_X1 U9891 ( .A1(n8244), .A2(n8389), .B1(n8421), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8245) );
  OAI21_X1 U9892 ( .B1(n8246), .B2(n8352), .A(n8245), .ZN(n8247) );
  AOI21_X1 U9893 ( .B1(n8248), .B2(n8419), .A(n8247), .ZN(n8249) );
  OAI21_X1 U9894 ( .B1(n8250), .B2(n8421), .A(n8249), .ZN(P2_U3206) );
  XNOR2_X1 U9895 ( .A(n8252), .B(n8251), .ZN(n8529) );
  XNOR2_X1 U9896 ( .A(n8254), .B(n8253), .ZN(n8257) );
  AOI222_X1 U9897 ( .A1(n8413), .A2(n8257), .B1(n8256), .B2(n8410), .C1(n8255), 
        .C2(n8408), .ZN(n8524) );
  MUX2_X1 U9898 ( .A(n8258), .B(n8524), .S(n9913), .Z(n8261) );
  AOI22_X1 U9899 ( .A1(n8526), .A2(n8445), .B1(n8389), .B2(n8259), .ZN(n8260)
         );
  OAI211_X1 U9900 ( .C1(n8529), .C2(n8448), .A(n8261), .B(n8260), .ZN(P2_U3207) );
  XOR2_X1 U9901 ( .A(n8267), .B(n8262), .Z(n8263) );
  OAI222_X1 U9902 ( .A1(n9909), .A2(n8264), .B1(n9910), .B2(n8284), .C1(n9907), 
        .C2(n8263), .ZN(n8462) );
  AOI21_X1 U9903 ( .B1(n8416), .B2(n8532), .A(n8462), .ZN(n8270) );
  AOI22_X1 U9904 ( .A1(n8265), .A2(n8389), .B1(n8421), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U9905 ( .A1(n8533), .A2(n8419), .ZN(n8268) );
  OAI211_X1 U9906 ( .C1(n8270), .C2(n8421), .A(n8269), .B(n8268), .ZN(P2_U3208) );
  NOR2_X1 U9907 ( .A1(n8537), .A2(n9899), .ZN(n8274) );
  XNOR2_X1 U9908 ( .A(n8271), .B(n8278), .ZN(n8272) );
  OAI222_X1 U9909 ( .A1(n9909), .A2(n8273), .B1(n9910), .B2(n8298), .C1(n8272), 
        .C2(n9907), .ZN(n8536) );
  AOI211_X1 U9910 ( .C1(n8389), .C2(n8275), .A(n8274), .B(n8536), .ZN(n8281)
         );
  INV_X1 U9911 ( .A(n8538), .ZN(n8279) );
  AOI22_X1 U9912 ( .A1(n8279), .A2(n8419), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8421), .ZN(n8280) );
  OAI21_X1 U9913 ( .B1(n8281), .B2(n8421), .A(n8280), .ZN(P2_U3209) );
  XOR2_X1 U9914 ( .A(n8285), .B(n8282), .Z(n8283) );
  OAI222_X1 U9915 ( .A1(n9909), .A2(n8284), .B1(n9910), .B2(n8308), .C1(n9907), 
        .C2(n8283), .ZN(n8468) );
  INV_X1 U9916 ( .A(n8468), .ZN(n8294) );
  INV_X1 U9917 ( .A(n8285), .ZN(n8286) );
  XNOR2_X1 U9918 ( .A(n8287), .B(n8286), .ZN(n8544) );
  INV_X1 U9919 ( .A(n8544), .ZN(n8292) );
  AOI22_X1 U9920 ( .A1(n8421), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8389), .B2(
        n8288), .ZN(n8289) );
  OAI21_X1 U9921 ( .B1(n8290), .B2(n8352), .A(n8289), .ZN(n8291) );
  AOI21_X1 U9922 ( .B1(n8292), .B2(n8419), .A(n8291), .ZN(n8293) );
  OAI21_X1 U9923 ( .B1(n8294), .B2(n8421), .A(n8293), .ZN(P2_U3210) );
  XNOR2_X1 U9924 ( .A(n8296), .B(n8295), .ZN(n8297) );
  OAI22_X1 U9925 ( .A1(n8297), .A2(n9907), .B1(n8320), .B2(n9910), .ZN(n8472)
         );
  NOR2_X1 U9926 ( .A1(n8298), .A2(n9909), .ZN(n8473) );
  OAI21_X1 U9927 ( .B1(n8472), .B2(n8473), .A(n9913), .ZN(n8305) );
  XNOR2_X1 U9928 ( .A(n8300), .B(n8299), .ZN(n8474) );
  AOI22_X1 U9929 ( .A1(n8421), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8389), .B2(
        n8301), .ZN(n8302) );
  OAI21_X1 U9930 ( .B1(n8548), .B2(n8352), .A(n8302), .ZN(n8303) );
  AOI21_X1 U9931 ( .B1(n8474), .B2(n8419), .A(n8303), .ZN(n8304) );
  NAND2_X1 U9932 ( .A1(n8305), .A2(n8304), .ZN(P2_U3211) );
  XNOR2_X1 U9933 ( .A(n8306), .B(n8311), .ZN(n8307) );
  OAI222_X1 U9934 ( .A1(n9909), .A2(n8308), .B1(n9910), .B2(n8334), .C1(n9907), 
        .C2(n8307), .ZN(n8477) );
  INV_X1 U9935 ( .A(n8477), .ZN(n8317) );
  NAND2_X1 U9936 ( .A1(n8310), .A2(n8309), .ZN(n8312) );
  XNOR2_X1 U9937 ( .A(n8312), .B(n8311), .ZN(n8478) );
  AOI22_X1 U9938 ( .A1(n8421), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8389), .B2(
        n8313), .ZN(n8314) );
  OAI21_X1 U9939 ( .B1(n8552), .B2(n8352), .A(n8314), .ZN(n8315) );
  AOI21_X1 U9940 ( .B1(n8478), .B2(n8419), .A(n8315), .ZN(n8316) );
  OAI21_X1 U9941 ( .B1(n8317), .B2(n8421), .A(n8316), .ZN(P2_U3212) );
  AOI21_X1 U9942 ( .B1(n8321), .B2(n8318), .A(n4445), .ZN(n8319) );
  OAI222_X1 U9943 ( .A1(n9909), .A2(n8320), .B1(n9910), .B2(n8347), .C1(n9907), 
        .C2(n8319), .ZN(n8480) );
  INV_X1 U9944 ( .A(n8480), .ZN(n8328) );
  XNOR2_X1 U9945 ( .A(n8322), .B(n8321), .ZN(n8481) );
  INV_X1 U9946 ( .A(n8323), .ZN(n8556) );
  AOI22_X1 U9947 ( .A1(n8421), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8389), .B2(
        n8324), .ZN(n8325) );
  OAI21_X1 U9948 ( .B1(n8556), .B2(n8352), .A(n8325), .ZN(n8326) );
  AOI21_X1 U9949 ( .B1(n8481), .B2(n8419), .A(n8326), .ZN(n8327) );
  OAI21_X1 U9950 ( .B1(n8328), .B2(n8421), .A(n8327), .ZN(P2_U3213) );
  XNOR2_X1 U9951 ( .A(n8329), .B(n8331), .ZN(n8560) );
  INV_X1 U9952 ( .A(n8560), .ZN(n8343) );
  INV_X1 U9953 ( .A(n8330), .ZN(n8333) );
  INV_X1 U9954 ( .A(n8331), .ZN(n8332) );
  AOI21_X1 U9955 ( .B1(n8333), .B2(n8332), .A(n9907), .ZN(n8338) );
  OAI22_X1 U9956 ( .A1(n8335), .A2(n9910), .B1(n8334), .B2(n9909), .ZN(n8336)
         );
  AOI21_X1 U9957 ( .B1(n8338), .B2(n8337), .A(n8336), .ZN(n8557) );
  MUX2_X1 U9958 ( .A(n8339), .B(n8557), .S(n9913), .Z(n8342) );
  AOI22_X1 U9959 ( .A1(n8559), .A2(n8445), .B1(n8389), .B2(n8340), .ZN(n8341)
         );
  OAI211_X1 U9960 ( .C1(n8343), .C2(n8448), .A(n8342), .B(n8341), .ZN(P2_U3214) );
  XNOR2_X1 U9961 ( .A(n8344), .B(n8351), .ZN(n8345) );
  OAI222_X1 U9962 ( .A1(n9909), .A2(n8347), .B1(n9910), .B2(n8346), .C1(n8345), 
        .C2(n9907), .ZN(n8487) );
  INV_X1 U9963 ( .A(n8487), .ZN(n8358) );
  INV_X1 U9964 ( .A(n8348), .ZN(n8349) );
  AOI21_X1 U9965 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8488) );
  NOR2_X1 U9966 ( .A1(n8567), .A2(n8352), .ZN(n8356) );
  OAI22_X1 U9967 ( .A1(n9913), .A2(n8354), .B1(n8353), .B2(n9898), .ZN(n8355)
         );
  AOI211_X1 U9968 ( .C1(n8488), .C2(n8419), .A(n8356), .B(n8355), .ZN(n8357)
         );
  OAI21_X1 U9969 ( .B1(n8358), .B2(n8421), .A(n8357), .ZN(P2_U3215) );
  XNOR2_X1 U9970 ( .A(n8360), .B(n8359), .ZN(n8571) );
  INV_X1 U9971 ( .A(n8571), .ZN(n8370) );
  XNOR2_X1 U9972 ( .A(n8362), .B(n8361), .ZN(n8364) );
  AOI222_X1 U9973 ( .A1(n8413), .A2(n8364), .B1(n8363), .B2(n8410), .C1(n8386), 
        .C2(n8408), .ZN(n8568) );
  MUX2_X1 U9974 ( .A(n8365), .B(n8568), .S(n9913), .Z(n8369) );
  INV_X1 U9975 ( .A(n8366), .ZN(n8367) );
  AOI22_X1 U9976 ( .A1(n8570), .A2(n8445), .B1(n8389), .B2(n8367), .ZN(n8368)
         );
  OAI211_X1 U9977 ( .C1(n8370), .C2(n8448), .A(n8369), .B(n8368), .ZN(P2_U3216) );
  XNOR2_X1 U9978 ( .A(n8372), .B(n8371), .ZN(n8577) );
  INV_X1 U9979 ( .A(n8577), .ZN(n8382) );
  XNOR2_X1 U9980 ( .A(n8374), .B(n8373), .ZN(n8376) );
  AOI222_X1 U9981 ( .A1(n8413), .A2(n8376), .B1(n8375), .B2(n8410), .C1(n8396), 
        .C2(n8408), .ZN(n8574) );
  MUX2_X1 U9982 ( .A(n8377), .B(n8574), .S(n9913), .Z(n8381) );
  INV_X1 U9983 ( .A(n8378), .ZN(n8379) );
  AOI22_X1 U9984 ( .A1(n8576), .A2(n8445), .B1(n8389), .B2(n8379), .ZN(n8380)
         );
  OAI211_X1 U9985 ( .C1(n8382), .C2(n8448), .A(n8381), .B(n8380), .ZN(P2_U3217) );
  XOR2_X1 U9986 ( .A(n8385), .B(n8383), .Z(n8582) );
  INV_X1 U9987 ( .A(n8582), .ZN(n8392) );
  XOR2_X1 U9988 ( .A(n8385), .B(n8384), .Z(n8387) );
  AOI222_X1 U9989 ( .A1(n8413), .A2(n8387), .B1(n8386), .B2(n8410), .C1(n8411), 
        .C2(n8408), .ZN(n8580) );
  MUX2_X1 U9990 ( .A(n8112), .B(n8580), .S(n9913), .Z(n8391) );
  AOI22_X1 U9991 ( .A1(n8581), .A2(n8445), .B1(n8389), .B2(n8388), .ZN(n8390)
         );
  OAI211_X1 U9992 ( .C1(n8392), .C2(n8448), .A(n8391), .B(n8390), .ZN(P2_U3218) );
  XNOR2_X1 U9993 ( .A(n8394), .B(n8393), .ZN(n8397) );
  AOI222_X1 U9994 ( .A1(n8413), .A2(n8397), .B1(n8396), .B2(n8410), .C1(n8395), 
        .C2(n8408), .ZN(n8585) );
  INV_X1 U9995 ( .A(n8585), .ZN(n8401) );
  OAI22_X1 U9996 ( .A1(n8399), .A2(n9899), .B1(n8398), .B2(n9898), .ZN(n8400)
         );
  OAI21_X1 U9997 ( .B1(n8401), .B2(n8400), .A(n9913), .ZN(n8405) );
  XNOR2_X1 U9998 ( .A(n8403), .B(n8402), .ZN(n8588) );
  AOI22_X1 U9999 ( .A1(n8588), .A2(n8419), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8421), .ZN(n8404) );
  NAND2_X1 U10000 ( .A1(n8405), .A2(n8404), .ZN(P2_U3219) );
  NOR2_X1 U10001 ( .A1(n9898), .A2(n8406), .ZN(n8415) );
  XOR2_X1 U10002 ( .A(n8407), .B(n8418), .Z(n8412) );
  AOI222_X1 U10003 ( .A1(n8413), .A2(n8412), .B1(n8411), .B2(n8410), .C1(n8409), .C2(n8408), .ZN(n8591) );
  INV_X1 U10004 ( .A(n8591), .ZN(n8414) );
  AOI211_X1 U10005 ( .C1(n8416), .C2(n8593), .A(n8415), .B(n8414), .ZN(n8422)
         );
  XOR2_X1 U10006 ( .A(n8418), .B(n8417), .Z(n8596) );
  AOI22_X1 U10007 ( .A1(n8596), .A2(n8419), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8421), .ZN(n8420) );
  OAI21_X1 U10008 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(P2_U3220) );
  NAND2_X1 U10009 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  NAND2_X1 U10010 ( .A1(n8426), .A2(n8425), .ZN(n8603) );
  XNOR2_X1 U10011 ( .A(n8427), .B(n5699), .ZN(n8428) );
  OAI222_X1 U10012 ( .A1(n9909), .A2(n8430), .B1(n9910), .B2(n8429), .C1(n9907), .C2(n8428), .ZN(n8508) );
  NAND2_X1 U10013 ( .A1(n8508), .A2(n9913), .ZN(n8435) );
  OAI22_X1 U10014 ( .A1(n9913), .A2(n8432), .B1(n8431), .B2(n9898), .ZN(n8433)
         );
  AOI21_X1 U10015 ( .B1(n8509), .B2(n8445), .A(n8433), .ZN(n8434) );
  OAI211_X1 U10016 ( .C1(n8603), .C2(n8448), .A(n8435), .B(n8434), .ZN(
        P2_U3221) );
  XNOR2_X1 U10017 ( .A(n8436), .B(n8438), .ZN(n9968) );
  XNOR2_X1 U10018 ( .A(n8437), .B(n8438), .ZN(n8439) );
  OAI222_X1 U10019 ( .A1(n9909), .A2(n8441), .B1(n9910), .B2(n8440), .C1(n8439), .C2(n9907), .ZN(n9969) );
  NAND2_X1 U10020 ( .A1(n9969), .A2(n9913), .ZN(n8447) );
  OAI22_X1 U10021 ( .A1(n9913), .A2(n8443), .B1(n8442), .B2(n9898), .ZN(n8444)
         );
  AOI21_X1 U10022 ( .B1(n9971), .B2(n8445), .A(n8444), .ZN(n8446) );
  OAI211_X1 U10023 ( .C1(n8448), .C2(n9968), .A(n8447), .B(n8446), .ZN(
        P2_U3222) );
  NOR2_X1 U10024 ( .A1(n8513), .A2(n9990), .ZN(n8450) );
  AOI21_X1 U10025 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9990), .A(n8450), .ZN(
        n8449) );
  OAI21_X1 U10026 ( .B1(n8515), .B2(n8491), .A(n8449), .ZN(P2_U3490) );
  AOI21_X1 U10027 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9990), .A(n8450), .ZN(
        n8451) );
  OAI21_X1 U10028 ( .B1(n8518), .B2(n8491), .A(n8451), .ZN(P2_U3489) );
  NAND2_X1 U10029 ( .A1(n9992), .A2(n9966), .ZN(n8512) );
  INV_X1 U10030 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8452) );
  MUX2_X1 U10031 ( .A(n8452), .B(n8519), .S(n9992), .Z(n8454) );
  INV_X1 U10032 ( .A(n8491), .ZN(n8504) );
  NAND2_X1 U10033 ( .A1(n8520), .A2(n8504), .ZN(n8453) );
  OAI211_X1 U10034 ( .C1(n8523), .C2(n8512), .A(n8454), .B(n8453), .ZN(
        P2_U3487) );
  MUX2_X1 U10035 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8455), .S(n9992), .Z(n8456) );
  INV_X1 U10036 ( .A(n8456), .ZN(n8457) );
  OAI21_X1 U10037 ( .B1(n8458), .B2(n8512), .A(n8457), .ZN(P2_U3486) );
  INV_X1 U10038 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8459) );
  MUX2_X1 U10039 ( .A(n8459), .B(n8524), .S(n9992), .Z(n8461) );
  NAND2_X1 U10040 ( .A1(n8526), .A2(n8504), .ZN(n8460) );
  OAI211_X1 U10041 ( .C1(n8512), .C2(n8529), .A(n8461), .B(n8460), .ZN(
        P2_U3485) );
  INV_X1 U10042 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8463) );
  INV_X1 U10043 ( .A(n8462), .ZN(n8530) );
  MUX2_X1 U10044 ( .A(n8463), .B(n8530), .S(n9992), .Z(n8465) );
  INV_X1 U10045 ( .A(n8512), .ZN(n8505) );
  AOI22_X1 U10046 ( .A1(n8533), .A2(n8505), .B1(n8504), .B2(n8532), .ZN(n8464)
         );
  NAND2_X1 U10047 ( .A1(n8465), .A2(n8464), .ZN(P2_U3484) );
  MUX2_X1 U10048 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8536), .S(n9992), .Z(n8467) );
  OAI22_X1 U10049 ( .A1(n8538), .A2(n8512), .B1(n8537), .B2(n8491), .ZN(n8466)
         );
  OR2_X1 U10050 ( .A1(n8467), .A2(n8466), .ZN(P2_U3483) );
  INV_X1 U10051 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8470) );
  AOI21_X1 U10052 ( .B1(n9972), .B2(n8469), .A(n8468), .ZN(n8541) );
  MUX2_X1 U10053 ( .A(n8470), .B(n8541), .S(n9992), .Z(n8471) );
  OAI21_X1 U10054 ( .B1(n8544), .B2(n8512), .A(n8471), .ZN(P2_U3482) );
  INV_X1 U10055 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8475) );
  AOI211_X1 U10056 ( .C1(n8474), .C2(n9966), .A(n8473), .B(n8472), .ZN(n8545)
         );
  MUX2_X1 U10057 ( .A(n8475), .B(n8545), .S(n9992), .Z(n8476) );
  OAI21_X1 U10058 ( .B1(n8548), .B2(n8491), .A(n8476), .ZN(P2_U3481) );
  AOI21_X1 U10059 ( .B1(n8478), .B2(n9966), .A(n8477), .ZN(n8549) );
  MUX2_X1 U10060 ( .A(n10226), .B(n8549), .S(n9992), .Z(n8479) );
  OAI21_X1 U10061 ( .B1(n8552), .B2(n8491), .A(n8479), .ZN(P2_U3480) );
  AOI21_X1 U10062 ( .B1(n8481), .B2(n9966), .A(n8480), .ZN(n8553) );
  MUX2_X1 U10063 ( .A(n8482), .B(n8553), .S(n9992), .Z(n8483) );
  OAI21_X1 U10064 ( .B1(n8556), .B2(n8491), .A(n8483), .ZN(P2_U3479) );
  MUX2_X1 U10065 ( .A(n8484), .B(n8557), .S(n9992), .Z(n8486) );
  AOI22_X1 U10066 ( .A1(n8560), .A2(n8505), .B1(n8504), .B2(n8559), .ZN(n8485)
         );
  NAND2_X1 U10067 ( .A1(n8486), .A2(n8485), .ZN(P2_U3478) );
  INV_X1 U10068 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8489) );
  AOI21_X1 U10069 ( .B1(n8488), .B2(n9966), .A(n8487), .ZN(n8563) );
  MUX2_X1 U10070 ( .A(n8489), .B(n8563), .S(n9992), .Z(n8490) );
  OAI21_X1 U10071 ( .B1(n8567), .B2(n8491), .A(n8490), .ZN(P2_U3477) );
  MUX2_X1 U10072 ( .A(n8492), .B(n8568), .S(n9992), .Z(n8494) );
  AOI22_X1 U10073 ( .A1(n8571), .A2(n8505), .B1(n8504), .B2(n8570), .ZN(n8493)
         );
  NAND2_X1 U10074 ( .A1(n8494), .A2(n8493), .ZN(P2_U3476) );
  MUX2_X1 U10075 ( .A(n8495), .B(n8574), .S(n9992), .Z(n8497) );
  AOI22_X1 U10076 ( .A1(n8577), .A2(n8505), .B1(n8504), .B2(n8576), .ZN(n8496)
         );
  NAND2_X1 U10077 ( .A1(n8497), .A2(n8496), .ZN(P2_U3475) );
  MUX2_X1 U10078 ( .A(n10199), .B(n8580), .S(n9992), .Z(n8499) );
  AOI22_X1 U10079 ( .A1(n8582), .A2(n8505), .B1(n8504), .B2(n8581), .ZN(n8498)
         );
  NAND2_X1 U10080 ( .A1(n8499), .A2(n8498), .ZN(P2_U3474) );
  MUX2_X1 U10081 ( .A(n8500), .B(n8585), .S(n9992), .Z(n8502) );
  AOI22_X1 U10082 ( .A1(n8588), .A2(n8505), .B1(n8504), .B2(n8587), .ZN(n8501)
         );
  NAND2_X1 U10083 ( .A1(n8502), .A2(n8501), .ZN(P2_U3473) );
  MUX2_X1 U10084 ( .A(n8503), .B(n8591), .S(n9992), .Z(n8507) );
  AOI22_X1 U10085 ( .A1(n8596), .A2(n8505), .B1(n8504), .B2(n8593), .ZN(n8506)
         );
  NAND2_X1 U10086 ( .A1(n8507), .A2(n8506), .ZN(P2_U3472) );
  AOI21_X1 U10087 ( .B1(n9972), .B2(n8509), .A(n8508), .ZN(n8599) );
  MUX2_X1 U10088 ( .A(n8510), .B(n8599), .S(n9992), .Z(n8511) );
  OAI21_X1 U10089 ( .B1(n8512), .B2(n8603), .A(n8511), .ZN(P2_U3471) );
  NOR2_X1 U10090 ( .A1(n8513), .A2(n9975), .ZN(n8516) );
  AOI21_X1 U10091 ( .B1(n9975), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8516), .ZN(
        n8514) );
  OAI21_X1 U10092 ( .B1(n8515), .B2(n8566), .A(n8514), .ZN(P2_U3458) );
  AOI21_X1 U10093 ( .B1(n9975), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8516), .ZN(
        n8517) );
  OAI21_X1 U10094 ( .B1(n8518), .B2(n8566), .A(n8517), .ZN(P2_U3457) );
  MUX2_X1 U10095 ( .A(n10129), .B(n8519), .S(n9973), .Z(n8522) );
  INV_X1 U10096 ( .A(n8566), .ZN(n8594) );
  NAND2_X1 U10097 ( .A1(n8520), .A2(n8594), .ZN(n8521) );
  OAI211_X1 U10098 ( .C1(n8523), .C2(n8602), .A(n8522), .B(n8521), .ZN(
        P2_U3455) );
  INV_X1 U10099 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8525) );
  MUX2_X1 U10100 ( .A(n8525), .B(n8524), .S(n9973), .Z(n8528) );
  NAND2_X1 U10101 ( .A1(n8526), .A2(n8594), .ZN(n8527) );
  OAI211_X1 U10102 ( .C1(n8529), .C2(n8602), .A(n8528), .B(n8527), .ZN(
        P2_U3453) );
  INV_X1 U10103 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8531) );
  MUX2_X1 U10104 ( .A(n8531), .B(n8530), .S(n9973), .Z(n8535) );
  INV_X1 U10105 ( .A(n8602), .ZN(n8595) );
  AOI22_X1 U10106 ( .A1(n8533), .A2(n8595), .B1(n8594), .B2(n8532), .ZN(n8534)
         );
  NAND2_X1 U10107 ( .A1(n8535), .A2(n8534), .ZN(P2_U3452) );
  MUX2_X1 U10108 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8536), .S(n9973), .Z(n8540) );
  OAI22_X1 U10109 ( .A1(n8538), .A2(n8602), .B1(n8537), .B2(n8566), .ZN(n8539)
         );
  OR2_X1 U10110 ( .A1(n8540), .A2(n8539), .ZN(P2_U3451) );
  INV_X1 U10111 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U10112 ( .A(n8542), .B(n8541), .S(n9973), .Z(n8543) );
  OAI21_X1 U10113 ( .B1(n8544), .B2(n8602), .A(n8543), .ZN(P2_U3450) );
  INV_X1 U10114 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8546) );
  MUX2_X1 U10115 ( .A(n8546), .B(n8545), .S(n9973), .Z(n8547) );
  OAI21_X1 U10116 ( .B1(n8548), .B2(n8566), .A(n8547), .ZN(P2_U3449) );
  MUX2_X1 U10117 ( .A(n8550), .B(n8549), .S(n9973), .Z(n8551) );
  OAI21_X1 U10118 ( .B1(n8552), .B2(n8566), .A(n8551), .ZN(P2_U3448) );
  MUX2_X1 U10119 ( .A(n8554), .B(n8553), .S(n9973), .Z(n8555) );
  OAI21_X1 U10120 ( .B1(n8556), .B2(n8566), .A(n8555), .ZN(P2_U3447) );
  INV_X1 U10121 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8558) );
  MUX2_X1 U10122 ( .A(n8558), .B(n8557), .S(n9973), .Z(n8562) );
  AOI22_X1 U10123 ( .A1(n8560), .A2(n8595), .B1(n8594), .B2(n8559), .ZN(n8561)
         );
  NAND2_X1 U10124 ( .A1(n8562), .A2(n8561), .ZN(P2_U3446) );
  MUX2_X1 U10125 ( .A(n8564), .B(n8563), .S(n9973), .Z(n8565) );
  OAI21_X1 U10126 ( .B1(n8567), .B2(n8566), .A(n8565), .ZN(P2_U3444) );
  INV_X1 U10127 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8569) );
  MUX2_X1 U10128 ( .A(n8569), .B(n8568), .S(n9973), .Z(n8573) );
  AOI22_X1 U10129 ( .A1(n8571), .A2(n8595), .B1(n8594), .B2(n8570), .ZN(n8572)
         );
  NAND2_X1 U10130 ( .A1(n8573), .A2(n8572), .ZN(P2_U3441) );
  MUX2_X1 U10131 ( .A(n8575), .B(n8574), .S(n9973), .Z(n8579) );
  AOI22_X1 U10132 ( .A1(n8577), .A2(n8595), .B1(n8594), .B2(n8576), .ZN(n8578)
         );
  NAND2_X1 U10133 ( .A1(n8579), .A2(n8578), .ZN(P2_U3438) );
  MUX2_X1 U10134 ( .A(n10096), .B(n8580), .S(n9973), .Z(n8584) );
  AOI22_X1 U10135 ( .A1(n8582), .A2(n8595), .B1(n8594), .B2(n8581), .ZN(n8583)
         );
  NAND2_X1 U10136 ( .A1(n8584), .A2(n8583), .ZN(P2_U3435) );
  INV_X1 U10137 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8586) );
  MUX2_X1 U10138 ( .A(n8586), .B(n8585), .S(n9973), .Z(n8590) );
  AOI22_X1 U10139 ( .A1(n8588), .A2(n8595), .B1(n8594), .B2(n8587), .ZN(n8589)
         );
  NAND2_X1 U10140 ( .A1(n8590), .A2(n8589), .ZN(P2_U3432) );
  INV_X1 U10141 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8592) );
  MUX2_X1 U10142 ( .A(n8592), .B(n8591), .S(n9973), .Z(n8598) );
  AOI22_X1 U10143 ( .A1(n8596), .A2(n8595), .B1(n8594), .B2(n8593), .ZN(n8597)
         );
  NAND2_X1 U10144 ( .A1(n8598), .A2(n8597), .ZN(P2_U3429) );
  INV_X1 U10145 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10146 ( .A(n8600), .B(n8599), .S(n9973), .Z(n8601) );
  OAI21_X1 U10147 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(P2_U3426) );
  INV_X1 U10148 ( .A(n8999), .ZN(n9700) );
  NOR4_X1 U10149 ( .A1(n8604), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5073), .ZN(n8605) );
  AOI21_X1 U10150 ( .B1(n8606), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8605), .ZN(
        n8607) );
  OAI21_X1 U10151 ( .B1(n9700), .B2(n8608), .A(n8607), .ZN(P2_U3264) );
  NAND2_X1 U10152 ( .A1(n9704), .A2(n8609), .ZN(n8610) );
  OAI211_X1 U10153 ( .C1(n8612), .C2(n8611), .A(n8610), .B(n9849), .ZN(
        P2_U3267) );
  MUX2_X1 U10154 ( .A(n8613), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10155 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8617) );
  NAND2_X1 U10156 ( .A1(n8617), .A2(n5036), .ZN(n8624) );
  INV_X1 U10157 ( .A(n8618), .ZN(n9808) );
  AOI22_X1 U10158 ( .A1(n8801), .A2(n9167), .B1(n8800), .B2(n9808), .ZN(n8623)
         );
  NOR2_X1 U10159 ( .A1(n8890), .A2(n8619), .ZN(n8620) );
  AOI211_X1 U10160 ( .C1(n9804), .C2(n8897), .A(n8621), .B(n8620), .ZN(n8622)
         );
  NAND3_X1 U10161 ( .A1(n8624), .A2(n8623), .A3(n8622), .ZN(P1_U3213) );
  NOR2_X1 U10162 ( .A1(n8631), .A2(n8630), .ZN(n8629) );
  INV_X1 U10163 ( .A(n8629), .ZN(n8625) );
  NAND2_X1 U10164 ( .A1(n8867), .A2(n8627), .ZN(n8633) );
  AOI22_X1 U10165 ( .A1(n9614), .A2(n8645), .B1(n8741), .B2(n9464), .ZN(n8634)
         );
  XNOR2_X1 U10166 ( .A(n8634), .B(n8674), .ZN(n8636) );
  AOI22_X1 U10167 ( .A1(n9614), .A2(n8741), .B1(n8740), .B2(n9464), .ZN(n8635)
         );
  NAND2_X1 U10168 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  OAI21_X1 U10169 ( .B1(n8636), .B2(n8635), .A(n8637), .ZN(n8831) );
  NAND2_X1 U10170 ( .A1(n9437), .A2(n8735), .ZN(n8639) );
  NAND2_X1 U10171 ( .A1(n9454), .A2(n8741), .ZN(n8638) );
  NAND2_X1 U10172 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  XNOR2_X1 U10173 ( .A(n8640), .B(n8674), .ZN(n8641) );
  AOI22_X1 U10174 ( .A1(n9437), .A2(n8741), .B1(n8740), .B2(n9454), .ZN(n8642)
         );
  XNOR2_X1 U10175 ( .A(n8641), .B(n8642), .ZN(n8756) );
  INV_X1 U10176 ( .A(n8641), .ZN(n8643) );
  NAND2_X1 U10177 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  AOI22_X1 U10178 ( .A1(n9605), .A2(n8645), .B1(n8741), .B2(n9433), .ZN(n8646)
         );
  XNOR2_X1 U10179 ( .A(n8646), .B(n8674), .ZN(n8647) );
  OAI22_X1 U10180 ( .A1(n9420), .A2(n8651), .B1(n8650), .B2(n8680), .ZN(n8848)
         );
  NAND2_X1 U10181 ( .A1(n9407), .A2(n8735), .ZN(n8653) );
  NAND2_X1 U10182 ( .A1(n9424), .A2(n8736), .ZN(n8652) );
  NAND2_X1 U10183 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  XNOR2_X1 U10184 ( .A(n8654), .B(n8678), .ZN(n8656) );
  AND2_X1 U10185 ( .A1(n9424), .A2(n8740), .ZN(n8655) );
  AOI21_X1 U10186 ( .B1(n9407), .B2(n8741), .A(n8655), .ZN(n8657) );
  NAND2_X1 U10187 ( .A1(n8656), .A2(n8657), .ZN(n8817) );
  INV_X1 U10188 ( .A(n8656), .ZN(n8659) );
  INV_X1 U10189 ( .A(n8657), .ZN(n8658) );
  NAND2_X1 U10190 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  NAND2_X1 U10191 ( .A1(n8717), .A2(n8817), .ZN(n8670) );
  NAND2_X1 U10192 ( .A1(n9595), .A2(n8735), .ZN(n8662) );
  NAND2_X1 U10193 ( .A1(n9403), .A2(n8736), .ZN(n8661) );
  NAND2_X1 U10194 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  XNOR2_X1 U10195 ( .A(n8663), .B(n8678), .ZN(n8665) );
  AND2_X1 U10196 ( .A1(n9403), .A2(n8740), .ZN(n8664) );
  AOI21_X1 U10197 ( .B1(n9595), .B2(n8741), .A(n8664), .ZN(n8666) );
  NAND2_X1 U10198 ( .A1(n8665), .A2(n8666), .ZN(n8671) );
  INV_X1 U10199 ( .A(n8665), .ZN(n8668) );
  INV_X1 U10200 ( .A(n8666), .ZN(n8667) );
  NAND2_X1 U10201 ( .A1(n8668), .A2(n8667), .ZN(n8669) );
  NAND2_X1 U10202 ( .A1(n9375), .A2(n8735), .ZN(n8673) );
  NAND2_X1 U10203 ( .A1(n9393), .A2(n8736), .ZN(n8672) );
  NAND2_X1 U10204 ( .A1(n8673), .A2(n8672), .ZN(n8675) );
  XNOR2_X1 U10205 ( .A(n8675), .B(n8674), .ZN(n8684) );
  AOI22_X1 U10206 ( .A1(n9375), .A2(n8741), .B1(n8740), .B2(n9393), .ZN(n8682)
         );
  XNOR2_X1 U10207 ( .A(n8684), .B(n8682), .ZN(n8773) );
  NAND2_X1 U10208 ( .A1(n9585), .A2(n8735), .ZN(n8677) );
  NAND2_X1 U10209 ( .A1(n9371), .A2(n8736), .ZN(n8676) );
  NAND2_X1 U10210 ( .A1(n8677), .A2(n8676), .ZN(n8679) );
  XNOR2_X1 U10211 ( .A(n8679), .B(n8678), .ZN(n8686) );
  NOR2_X1 U10212 ( .A1(n8776), .A2(n8680), .ZN(n8681) );
  AOI21_X1 U10213 ( .B1(n9585), .B2(n8741), .A(n8681), .ZN(n8687) );
  XNOR2_X1 U10214 ( .A(n8686), .B(n8687), .ZN(n8876) );
  INV_X1 U10215 ( .A(n8682), .ZN(n8683) );
  NOR2_X1 U10216 ( .A1(n8684), .A2(n8683), .ZN(n8877) );
  NOR2_X1 U10217 ( .A1(n8876), .A2(n8877), .ZN(n8685) );
  INV_X1 U10218 ( .A(n8686), .ZN(n8689) );
  INV_X1 U10219 ( .A(n8687), .ZN(n8688) );
  NAND2_X1 U10220 ( .A1(n8689), .A2(n8688), .ZN(n8698) );
  NAND2_X1 U10221 ( .A1(n9341), .A2(n8735), .ZN(n8691) );
  NAND2_X1 U10222 ( .A1(n9360), .A2(n8736), .ZN(n8690) );
  NAND2_X1 U10223 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  XNOR2_X1 U10224 ( .A(n8692), .B(n8674), .ZN(n8696) );
  NAND2_X1 U10225 ( .A1(n9341), .A2(n8736), .ZN(n8694) );
  NAND2_X1 U10226 ( .A1(n8740), .A2(n9360), .ZN(n8693) );
  NAND2_X1 U10227 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  AOI21_X1 U10228 ( .B1(n8696), .B2(n8695), .A(n8748), .ZN(n8697) );
  AOI21_X1 U10229 ( .B1(n8702), .B2(n8698), .A(n8697), .ZN(n8703) );
  INV_X1 U10230 ( .A(n8697), .ZN(n8700) );
  INV_X1 U10231 ( .A(n8698), .ZN(n8699) );
  NOR2_X1 U10232 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  OAI21_X1 U10233 ( .B1(n8703), .B2(n8744), .A(n5036), .ZN(n8708) );
  AOI22_X1 U10234 ( .A1(n8861), .A2(n9337), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8707) );
  INV_X1 U10235 ( .A(n8704), .ZN(n9343) );
  AOI22_X1 U10236 ( .A1(n8801), .A2(n9371), .B1(n8800), .B2(n9343), .ZN(n8706)
         );
  NAND2_X1 U10237 ( .A1(n9341), .A2(n8897), .ZN(n8705) );
  NAND4_X1 U10238 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(
        P1_U3214) );
  XNOR2_X1 U10239 ( .A(n4523), .B(n8709), .ZN(n8710) );
  XNOR2_X1 U10240 ( .A(n8711), .B(n8710), .ZN(n8712) );
  NAND2_X1 U10241 ( .A1(n8712), .A2(n5036), .ZN(n8716) );
  AND2_X1 U10242 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9785) );
  INV_X1 U10243 ( .A(n9559), .ZN(n8713) );
  OAI22_X1 U10244 ( .A1(n8894), .A2(n8713), .B1(n5993), .B2(n8891), .ZN(n8714)
         );
  AOI211_X1 U10245 ( .C1(n8861), .C2(n9159), .A(n9785), .B(n8714), .ZN(n8715)
         );
  OAI211_X1 U10246 ( .C1(n9561), .C2(n8782), .A(n8716), .B(n8715), .ZN(
        P1_U3215) );
  NAND3_X1 U10247 ( .A1(n8718), .A2(n8719), .A3(n4486), .ZN(n8720) );
  AOI21_X1 U10248 ( .B1(n8717), .B2(n8720), .A(n8899), .ZN(n8724) );
  AOI22_X1 U10249 ( .A1(n9403), .A2(n8861), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8722) );
  AOI22_X1 U10250 ( .A1(n8801), .A2(n9433), .B1(n9408), .B2(n8800), .ZN(n8721)
         );
  OAI211_X1 U10251 ( .C1(n9673), .C2(n8782), .A(n8722), .B(n8721), .ZN(n8723)
         );
  OR2_X1 U10252 ( .A1(n8724), .A2(n8723), .ZN(P1_U3216) );
  AOI21_X1 U10253 ( .B1(n8726), .B2(n8725), .A(n4485), .ZN(n8734) );
  NOR2_X1 U10254 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8727), .ZN(n9723) );
  OAI22_X1 U10255 ( .A1(n8894), .A2(n8729), .B1(n8728), .B2(n8891), .ZN(n8730)
         );
  AOI211_X1 U10256 ( .C1(n8861), .C2(n9162), .A(n9723), .B(n8730), .ZN(n8733)
         );
  NAND2_X1 U10257 ( .A1(n8731), .A2(n8897), .ZN(n8732) );
  OAI211_X1 U10258 ( .C1(n8734), .C2(n8899), .A(n8733), .B(n8732), .ZN(
        P1_U3217) );
  NAND2_X1 U10259 ( .A1(n9574), .A2(n8735), .ZN(n8738) );
  NAND2_X1 U10260 ( .A1(n9337), .A2(n8736), .ZN(n8737) );
  NAND2_X1 U10261 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  XNOR2_X1 U10262 ( .A(n8739), .B(n8674), .ZN(n8743) );
  AOI22_X1 U10263 ( .A1(n9574), .A2(n8741), .B1(n8740), .B2(n9337), .ZN(n8742)
         );
  XNOR2_X1 U10264 ( .A(n8743), .B(n8742), .ZN(n8749) );
  NAND3_X1 U10265 ( .A1(n8744), .A2(n5036), .A3(n8749), .ZN(n8752) );
  OAI22_X1 U10266 ( .A1(n8890), .A2(n9053), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8745), .ZN(n8747) );
  OAI22_X1 U10267 ( .A1(n8894), .A2(n9323), .B1(n8980), .B2(n8891), .ZN(n8746)
         );
  AOI211_X1 U10268 ( .C1(n9574), .C2(n8897), .A(n8747), .B(n8746), .ZN(n8751)
         );
  NAND3_X1 U10269 ( .A1(n8749), .A2(n5036), .A3(n8748), .ZN(n8750) );
  NAND4_X1 U10270 ( .A1(n8753), .A2(n8752), .A3(n8751), .A4(n8750), .ZN(
        P1_U3220) );
  OAI21_X1 U10271 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8760) );
  AOI22_X1 U10272 ( .A1(n9433), .A2(n8861), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8758) );
  AOI22_X1 U10273 ( .A1(n8801), .A2(n9464), .B1(n8800), .B2(n9438), .ZN(n8757)
         );
  OAI211_X1 U10274 ( .C1(n4583), .C2(n8782), .A(n8758), .B(n8757), .ZN(n8759)
         );
  AOI21_X1 U10275 ( .B1(n8760), .B2(n5036), .A(n8759), .ZN(n8761) );
  INV_X1 U10276 ( .A(n8761), .ZN(P1_U3223) );
  XOR2_X1 U10277 ( .A(n8763), .B(n8762), .Z(n8770) );
  NAND2_X1 U10278 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9757) );
  OAI21_X1 U10279 ( .B1(n8890), .B2(n5993), .A(n9757), .ZN(n8767) );
  OAI22_X1 U10280 ( .A1(n8894), .A2(n8765), .B1(n8891), .B2(n8764), .ZN(n8766)
         );
  AOI211_X1 U10281 ( .C1(n8768), .C2(n8897), .A(n8767), .B(n8766), .ZN(n8769)
         );
  OAI21_X1 U10282 ( .B1(n8770), .B2(n8899), .A(n8769), .ZN(P1_U3224) );
  OAI21_X1 U10283 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(n8774) );
  NAND2_X1 U10284 ( .A1(n8774), .A2(n5036), .ZN(n8781) );
  INV_X1 U10285 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8775) );
  OAI22_X1 U10286 ( .A1(n8890), .A2(n8776), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8775), .ZN(n8779) );
  NOR2_X1 U10287 ( .A1(n8777), .A2(n8891), .ZN(n8778) );
  AOI211_X1 U10288 ( .C1(n8800), .C2(n9376), .A(n8779), .B(n8778), .ZN(n8780)
         );
  OAI211_X1 U10289 ( .C1(n9669), .C2(n8782), .A(n8781), .B(n8780), .ZN(
        P1_U3225) );
  XNOR2_X1 U10290 ( .A(n8785), .B(n8786), .ZN(n8887) );
  INV_X1 U10291 ( .A(n8784), .ZN(n8886) );
  NOR2_X1 U10292 ( .A1(n8887), .A2(n8886), .ZN(n8885) );
  AOI21_X1 U10293 ( .B1(n8786), .B2(n8785), .A(n8885), .ZN(n8790) );
  XNOR2_X1 U10294 ( .A(n8788), .B(n8787), .ZN(n8789) );
  XNOR2_X1 U10295 ( .A(n8790), .B(n8789), .ZN(n8794) );
  AOI22_X1 U10296 ( .A1(n8801), .A2(n9159), .B1(n8800), .B2(n9515), .ZN(n8791)
         );
  NAND2_X1 U10297 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9257) );
  OAI211_X1 U10298 ( .C1(n9510), .C2(n8890), .A(n8791), .B(n9257), .ZN(n8792)
         );
  AOI21_X1 U10299 ( .B1(n9637), .B2(n8897), .A(n8792), .ZN(n8793) );
  OAI21_X1 U10300 ( .B1(n8794), .B2(n8899), .A(n8793), .ZN(P1_U3226) );
  OAI21_X1 U10301 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8798) );
  NAND2_X1 U10302 ( .A1(n8798), .A2(n5036), .ZN(n8808) );
  AOI22_X1 U10303 ( .A1(n8801), .A2(n9169), .B1(n8800), .B2(n8799), .ZN(n8807)
         );
  OAI21_X1 U10304 ( .B1(n8890), .B2(n8803), .A(n8802), .ZN(n8804) );
  AOI21_X1 U10305 ( .B1(n8805), .B2(n8897), .A(n8804), .ZN(n8806) );
  NAND3_X1 U10306 ( .A1(n8808), .A2(n8807), .A3(n8806), .ZN(P1_U3227) );
  NAND2_X1 U10307 ( .A1(n8867), .A2(n8809), .ZN(n8810) );
  XOR2_X1 U10308 ( .A(n8811), .B(n8810), .Z(n8816) );
  NAND2_X1 U10309 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9276) );
  OAI21_X1 U10310 ( .B1(n8812), .B2(n8890), .A(n9276), .ZN(n8814) );
  OAI22_X1 U10311 ( .A1(n8894), .A2(n9500), .B1(n8889), .B2(n8891), .ZN(n8813)
         );
  AOI211_X1 U10312 ( .C1(n9498), .C2(n8897), .A(n8814), .B(n8813), .ZN(n8815)
         );
  OAI21_X1 U10313 ( .B1(n8816), .B2(n8899), .A(n8815), .ZN(P1_U3228) );
  INV_X1 U10314 ( .A(n8817), .ZN(n8818) );
  NOR2_X1 U10315 ( .A1(n8819), .A2(n8818), .ZN(n8822) );
  INV_X1 U10316 ( .A(n8820), .ZN(n8821) );
  AOI21_X1 U10317 ( .B1(n8822), .B2(n8717), .A(n8821), .ZN(n8827) );
  OAI22_X1 U10318 ( .A1(n8850), .A2(n8891), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8823), .ZN(n8825) );
  OAI22_X1 U10319 ( .A1(n8880), .A2(n8890), .B1(n8894), .B2(n9386), .ZN(n8824)
         );
  AOI211_X1 U10320 ( .C1(n9595), .C2(n8897), .A(n8825), .B(n8824), .ZN(n8826)
         );
  OAI21_X1 U10321 ( .B1(n8827), .B2(n8899), .A(n8826), .ZN(P1_U3229) );
  INV_X1 U10322 ( .A(n8828), .ZN(n8829) );
  AOI21_X1 U10323 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8836) );
  INV_X1 U10324 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8832) );
  OAI22_X1 U10325 ( .A1(n8961), .A2(n8890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8832), .ZN(n8834) );
  OAI22_X1 U10326 ( .A1(n9447), .A2(n8894), .B1(n8891), .B2(n9487), .ZN(n8833)
         );
  AOI211_X1 U10327 ( .C1(n9614), .C2(n8897), .A(n8834), .B(n8833), .ZN(n8835)
         );
  OAI21_X1 U10328 ( .B1(n8836), .B2(n8899), .A(n8835), .ZN(P1_U3233) );
  XOR2_X1 U10329 ( .A(n8838), .B(n8837), .Z(n8845) );
  NAND2_X1 U10330 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9772) );
  OAI21_X1 U10331 ( .B1(n8890), .B2(n8892), .A(n9772), .ZN(n8842) );
  OAI22_X1 U10332 ( .A1(n8894), .A2(n8840), .B1(n8891), .B2(n8839), .ZN(n8841)
         );
  AOI211_X1 U10333 ( .C1(n8843), .C2(n8897), .A(n8842), .B(n8841), .ZN(n8844)
         );
  OAI21_X1 U10334 ( .B1(n8845), .B2(n8899), .A(n8844), .ZN(P1_U3234) );
  INV_X1 U10335 ( .A(n8718), .ZN(n8846) );
  AOI21_X1 U10336 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8854) );
  OAI22_X1 U10337 ( .A1(n8850), .A2(n8890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8849), .ZN(n8852) );
  OAI22_X1 U10338 ( .A1(n8961), .A2(n8891), .B1(n8894), .B2(n9417), .ZN(n8851)
         );
  AOI211_X1 U10339 ( .C1(n9605), .C2(n8897), .A(n8852), .B(n8851), .ZN(n8853)
         );
  OAI21_X1 U10340 ( .B1(n8854), .B2(n8899), .A(n8853), .ZN(P1_U3235) );
  NAND2_X1 U10341 ( .A1(n8857), .A2(n8856), .ZN(n8858) );
  XNOR2_X1 U10342 ( .A(n8855), .B(n8858), .ZN(n8865) );
  NOR2_X1 U10343 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5959), .ZN(n9744) );
  OAI22_X1 U10344 ( .A1(n8894), .A2(n8859), .B1(n5953), .B2(n8891), .ZN(n8860)
         );
  AOI211_X1 U10345 ( .C1(n8861), .C2(n9161), .A(n9744), .B(n8860), .ZN(n8864)
         );
  NAND2_X1 U10346 ( .A1(n8862), .A2(n8897), .ZN(n8863) );
  OAI211_X1 U10347 ( .C1(n8865), .C2(n8899), .A(n8864), .B(n8863), .ZN(
        P1_U3236) );
  NAND2_X1 U10348 ( .A1(n8867), .A2(n8866), .ZN(n8869) );
  AND2_X1 U10349 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  XOR2_X1 U10350 ( .A(n8871), .B(n8870), .Z(n8875) );
  NAND2_X1 U10351 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9800) );
  OAI21_X1 U10352 ( .B1(n9487), .B2(n8890), .A(n9800), .ZN(n8873) );
  OAI22_X1 U10353 ( .A1(n8894), .A2(n9480), .B1(n8891), .B2(n9510), .ZN(n8872)
         );
  AOI211_X1 U10354 ( .C1(n9625), .C2(n8897), .A(n8873), .B(n8872), .ZN(n8874)
         );
  OAI21_X1 U10355 ( .B1(n8875), .B2(n8899), .A(n8874), .ZN(P1_U3238) );
  OAI21_X1 U10356 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8879) );
  NAND3_X1 U10357 ( .A1(n8879), .A2(n5036), .A3(n8702), .ZN(n8884) );
  INV_X1 U10358 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10306) );
  OAI22_X1 U10359 ( .A1(n8890), .A2(n8980), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10306), .ZN(n8882) );
  OAI22_X1 U10360 ( .A1(n8880), .A2(n8891), .B1(n9353), .B2(n8894), .ZN(n8881)
         );
  AOI211_X1 U10361 ( .C1(n9585), .C2(n8897), .A(n8882), .B(n8881), .ZN(n8883)
         );
  NAND2_X1 U10362 ( .A1(n8884), .A2(n8883), .ZN(P1_U3240) );
  AOI21_X1 U10363 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8900) );
  INV_X1 U10364 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8888) );
  OAI22_X1 U10365 ( .A1(n8890), .A2(n8889), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8888), .ZN(n8896) );
  OAI22_X1 U10366 ( .A1(n8894), .A2(n8893), .B1(n8892), .B2(n8891), .ZN(n8895)
         );
  AOI211_X1 U10367 ( .C1(n9535), .C2(n8897), .A(n8896), .B(n8895), .ZN(n8898)
         );
  OAI21_X1 U10368 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(P1_U3241) );
  AOI21_X1 U10369 ( .B1(n9076), .B2(n9159), .A(n9049), .ZN(n8948) );
  AND2_X1 U10370 ( .A1(n8928), .A2(n8901), .ZN(n8924) );
  AND2_X1 U10371 ( .A1(n8902), .A2(n8904), .ZN(n8903) );
  NAND2_X1 U10372 ( .A1(n8911), .A2(n8904), .ZN(n9065) );
  INV_X1 U10373 ( .A(n8907), .ZN(n8913) );
  INV_X1 U10374 ( .A(n8911), .ZN(n8912) );
  OAI22_X1 U10375 ( .A1(n8916), .A2(n8915), .B1(n9025), .B2(n9049), .ZN(n8919)
         );
  AOI21_X1 U10376 ( .B1(n9049), .B2(n8917), .A(n8919), .ZN(n8922) );
  INV_X1 U10377 ( .A(n8918), .ZN(n8921) );
  INV_X1 U10378 ( .A(n8919), .ZN(n8920) );
  OAI22_X1 U10379 ( .A1(n8922), .A2(n8921), .B1(n8920), .B2(n9049), .ZN(n8923)
         );
  OAI21_X1 U10380 ( .B1(n8924), .B2(n9049), .A(n8923), .ZN(n8929) );
  NAND2_X1 U10381 ( .A1(n9535), .A2(n9550), .ZN(n8945) );
  AND2_X1 U10382 ( .A1(n8945), .A2(n8926), .ZN(n9073) );
  OAI211_X1 U10383 ( .C1(n8948), .C2(n9535), .A(n8927), .B(n8947), .ZN(n8944)
         );
  OAI21_X1 U10384 ( .B1(n8929), .B2(n4675), .A(n8928), .ZN(n8932) );
  NAND2_X1 U10385 ( .A1(n8931), .A2(n8930), .ZN(n9066) );
  AOI21_X1 U10386 ( .B1(n8932), .B2(n9054), .A(n9066), .ZN(n8935) );
  NAND2_X1 U10387 ( .A1(n8934), .A2(n8933), .ZN(n9071) );
  OAI21_X1 U10388 ( .B1(n8935), .B2(n9071), .A(n9070), .ZN(n8938) );
  AOI211_X1 U10389 ( .C1(n8938), .C2(n8937), .A(n8936), .B(n9544), .ZN(n8942)
         );
  INV_X1 U10390 ( .A(n8939), .ZN(n8941) );
  NAND2_X1 U10391 ( .A1(n8947), .A2(n8940), .ZN(n9078) );
  NOR3_X1 U10392 ( .A1(n8942), .A2(n8941), .A3(n9078), .ZN(n8943) );
  MUX2_X1 U10393 ( .A(n8944), .B(n8943), .S(n9049), .Z(n8951) );
  INV_X1 U10394 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U10395 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  AOI21_X1 U10396 ( .B1(n9076), .B2(n8949), .A(n8948), .ZN(n8950) );
  AND2_X1 U10397 ( .A1(n9084), .A2(n8952), .ZN(n9082) );
  INV_X1 U10398 ( .A(n8954), .ZN(n9097) );
  NAND2_X1 U10399 ( .A1(n8960), .A2(n8954), .ZN(n8955) );
  AOI21_X1 U10400 ( .B1(n9510), .B2(n9498), .A(n4875), .ZN(n9079) );
  NAND3_X1 U10401 ( .A1(n9083), .A2(n9049), .A3(n9084), .ZN(n8956) );
  AOI21_X1 U10402 ( .B1(n8957), .B2(n9079), .A(n8956), .ZN(n8959) );
  AOI21_X1 U10403 ( .B1(n8964), .B2(n9083), .A(n9049), .ZN(n8958) );
  NAND2_X1 U10404 ( .A1(n8965), .A2(n8960), .ZN(n9102) );
  OR2_X1 U10405 ( .A1(n9437), .A2(n8961), .ZN(n9101) );
  OAI21_X1 U10406 ( .B1(n8966), .B2(n9102), .A(n9101), .ZN(n8963) );
  NAND2_X1 U10407 ( .A1(n8971), .A2(n8962), .ZN(n9088) );
  AOI21_X1 U10408 ( .B1(n8963), .B2(n9423), .A(n9088), .ZN(n8970) );
  NAND2_X1 U10409 ( .A1(n9101), .A2(n8964), .ZN(n9094) );
  OAI21_X1 U10410 ( .B1(n8966), .B2(n9094), .A(n8965), .ZN(n8968) );
  NAND2_X1 U10411 ( .A1(n9390), .A2(n8967), .ZN(n9103) );
  AOI21_X1 U10412 ( .B1(n8968), .B2(n9423), .A(n9103), .ZN(n8969) );
  MUX2_X1 U10413 ( .A(n8970), .B(n8969), .S(n9049), .Z(n8975) );
  MUX2_X1 U10414 ( .A(n9390), .B(n8971), .S(n9049), .Z(n8972) );
  NAND2_X1 U10415 ( .A1(n9391), .A2(n8972), .ZN(n8974) );
  MUX2_X1 U10416 ( .A(n9089), .B(n9104), .S(n9049), .Z(n8973) );
  NAND2_X1 U10417 ( .A1(n9108), .A2(n8976), .ZN(n9092) );
  NOR2_X1 U10418 ( .A1(n9360), .A2(n9049), .ZN(n8978) );
  INV_X1 U10419 ( .A(n8978), .ZN(n8977) );
  OAI22_X1 U10420 ( .A1(n9664), .A2(n8977), .B1(n9049), .B2(n9337), .ZN(n8986)
         );
  AOI21_X1 U10421 ( .B1(n8979), .B2(n8978), .A(n9664), .ZN(n8984) );
  NOR2_X1 U10422 ( .A1(n8980), .A2(n9004), .ZN(n8981) );
  AOI21_X1 U10423 ( .B1(n8981), .B2(n9337), .A(n9341), .ZN(n8983) );
  AOI22_X1 U10424 ( .A1(n9664), .A2(n8981), .B1(n9049), .B2(n9337), .ZN(n8982)
         );
  OAI22_X1 U10425 ( .A1(n8984), .A2(n8983), .B1(n8982), .B2(n9574), .ZN(n8985)
         );
  AOI21_X1 U10426 ( .B1(n9574), .B2(n8986), .A(n8985), .ZN(n8989) );
  INV_X1 U10427 ( .A(n9099), .ZN(n9120) );
  OAI21_X1 U10428 ( .B1(n9120), .B2(n4661), .A(n9108), .ZN(n8988) );
  NAND2_X1 U10429 ( .A1(n9053), .A2(n9049), .ZN(n8991) );
  MUX2_X1 U10430 ( .A(n9049), .B(n9053), .S(n9314), .Z(n8990) );
  AOI22_X1 U10431 ( .A1(n8993), .A2(n8992), .B1(n8991), .B2(n8990), .ZN(n9006)
         );
  NAND2_X1 U10432 ( .A1(n8994), .A2(n8998), .ZN(n8997) );
  OR2_X1 U10433 ( .A1(n9000), .A2(n8995), .ZN(n8996) );
  NAND2_X1 U10434 ( .A1(n8999), .A2(n8998), .ZN(n9002) );
  OR2_X1 U10435 ( .A1(n9000), .A2(n10195), .ZN(n9001) );
  NAND2_X1 U10436 ( .A1(n9002), .A2(n9001), .ZN(n9009) );
  NAND2_X1 U10437 ( .A1(n9009), .A2(n9126), .ZN(n9132) );
  NAND2_X1 U10438 ( .A1(n9003), .A2(n9132), .ZN(n9008) );
  INV_X1 U10439 ( .A(n9157), .ZN(n9011) );
  NAND2_X1 U10440 ( .A1(n9305), .A2(n9157), .ZN(n9005) );
  OR2_X1 U10441 ( .A1(n9305), .A2(n9011), .ZN(n9010) );
  OAI22_X1 U10442 ( .A1(n9006), .A2(n9005), .B1(n9004), .B2(n9010), .ZN(n9007)
         );
  AOI21_X1 U10443 ( .B1(n9048), .B2(n6154), .A(n9056), .ZN(n9156) );
  OR2_X1 U10444 ( .A1(n9009), .A2(n9126), .ZN(n9146) );
  NAND2_X1 U10445 ( .A1(n9146), .A2(n9132), .ZN(n9047) );
  INV_X1 U10446 ( .A(n9010), .ZN(n9129) );
  AND2_X1 U10447 ( .A1(n9305), .A2(n9011), .ZN(n9052) );
  INV_X1 U10448 ( .A(n9052), .ZN(n9044) );
  INV_X1 U10449 ( .A(n9391), .ZN(n9041) );
  NOR2_X1 U10450 ( .A1(n9012), .A2(n6288), .ZN(n9021) );
  INV_X1 U10451 ( .A(n9013), .ZN(n9020) );
  NOR2_X1 U10452 ( .A1(n9015), .A2(n9014), .ZN(n9019) );
  NOR2_X1 U10453 ( .A1(n4514), .A2(n9016), .ZN(n9018) );
  NAND4_X1 U10454 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(n9018), .ZN(n9023)
         );
  NOR2_X1 U10455 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  NAND3_X1 U10456 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9027) );
  OR3_X1 U10457 ( .A1(n9029), .A2(n9028), .A3(n9027), .ZN(n9030) );
  OR3_X1 U10458 ( .A1(n9032), .A2(n9031), .A3(n9030), .ZN(n9033) );
  NOR2_X1 U10459 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  NAND4_X1 U10460 ( .A1(n9511), .A2(n4862), .A3(n9035), .A4(n9525), .ZN(n9036)
         );
  NOR2_X1 U10461 ( .A1(n9485), .A2(n9036), .ZN(n9037) );
  NAND3_X1 U10462 ( .A1(n9462), .A2(n9037), .A3(n9495), .ZN(n9038) );
  NOR2_X1 U10463 ( .A1(n9452), .A2(n9038), .ZN(n9039) );
  NAND4_X1 U10464 ( .A1(n9401), .A2(n9423), .A3(n9039), .A4(n9430), .ZN(n9040)
         );
  OR3_X1 U10465 ( .A1(n9366), .A2(n9041), .A3(n9040), .ZN(n9042) );
  NOR2_X1 U10466 ( .A1(n9348), .A2(n9042), .ZN(n9043) );
  NAND4_X1 U10467 ( .A1(n9044), .A2(n9329), .A3(n9339), .A4(n9043), .ZN(n9045)
         );
  OR4_X1 U10468 ( .A1(n9047), .A2(n9046), .A3(n9129), .A4(n9045), .ZN(n9136)
         );
  NAND4_X1 U10469 ( .A1(n9136), .A2(n9143), .A3(n9140), .A4(n9137), .ZN(n9155)
         );
  NOR3_X1 U10470 ( .A1(n9142), .A2(n6154), .A3(n9050), .ZN(n9051) );
  AOI21_X1 U10471 ( .B1(n9053), .B2(n9314), .A(n9052), .ZN(n9131) );
  AND2_X1 U10472 ( .A1(n9055), .A2(n9054), .ZN(n9068) );
  AOI21_X1 U10473 ( .B1(n9171), .B2(n5848), .A(n9056), .ZN(n9060) );
  NAND2_X1 U10474 ( .A1(n9057), .A2(n4415), .ZN(n9058) );
  NAND4_X1 U10475 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n9064)
         );
  OAI211_X1 U10476 ( .C1(n9065), .C2(n9064), .A(n9063), .B(n9062), .ZN(n9067)
         );
  AOI21_X1 U10477 ( .B1(n9068), .B2(n9067), .A(n9066), .ZN(n9072) );
  OAI211_X1 U10478 ( .C1(n9072), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9075)
         );
  INV_X1 U10479 ( .A(n9073), .ZN(n9074) );
  AOI21_X1 U10480 ( .B1(n4484), .B2(n9075), .A(n9074), .ZN(n9077) );
  OAI21_X1 U10481 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9081) );
  INV_X1 U10482 ( .A(n9079), .ZN(n9080) );
  AOI21_X1 U10483 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9087) );
  INV_X1 U10484 ( .A(n9083), .ZN(n9086) );
  INV_X1 U10485 ( .A(n9084), .ZN(n9085) );
  NOR3_X1 U10486 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(n9096) );
  INV_X1 U10487 ( .A(n9088), .ZN(n9091) );
  INV_X1 U10488 ( .A(n9390), .ZN(n9090) );
  OAI21_X1 U10489 ( .B1(n9091), .B2(n9090), .A(n9089), .ZN(n9093) );
  AOI21_X1 U10490 ( .B1(n9104), .B2(n9093), .A(n9092), .ZN(n9110) );
  INV_X1 U10491 ( .A(n9110), .ZN(n9095) );
  NOR2_X1 U10492 ( .A1(n9095), .A2(n9094), .ZN(n9121) );
  OAI21_X1 U10493 ( .B1(n9097), .B2(n9096), .A(n9121), .ZN(n9100) );
  INV_X1 U10494 ( .A(n9098), .ZN(n9125) );
  AOI21_X1 U10495 ( .B1(n9100), .B2(n9099), .A(n9125), .ZN(n9116) );
  INV_X1 U10496 ( .A(n9101), .ZN(n9107) );
  INV_X1 U10497 ( .A(n9102), .ZN(n9106) );
  INV_X1 U10498 ( .A(n9103), .ZN(n9105) );
  OAI211_X1 U10499 ( .C1(n9107), .C2(n9106), .A(n9105), .B(n9104), .ZN(n9109)
         );
  AOI22_X1 U10500 ( .A1(n9110), .A2(n9109), .B1(n4661), .B2(n9108), .ZN(n9113)
         );
  OAI211_X1 U10501 ( .C1(n9113), .C2(n9125), .A(n9112), .B(n9111), .ZN(n9122)
         );
  INV_X1 U10502 ( .A(n9114), .ZN(n9115) );
  AOI21_X1 U10503 ( .B1(n6178), .B2(n9330), .A(n9115), .ZN(n9127) );
  OAI21_X1 U10504 ( .B1(n9116), .B2(n9122), .A(n9127), .ZN(n9118) );
  INV_X1 U10505 ( .A(n9132), .ZN(n9117) );
  AOI211_X1 U10506 ( .C1(n9131), .C2(n9118), .A(n9129), .B(n9117), .ZN(n9144)
         );
  NAND4_X1 U10507 ( .A1(n9530), .A2(n9729), .A3(n9693), .A4(n9147), .ZN(n9119)
         );
  OAI211_X1 U10508 ( .C1(n6154), .C2(n9142), .A(n9119), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9145) );
  NAND3_X1 U10509 ( .A1(n9144), .A2(n9143), .A3(n9145), .ZN(n9152) );
  AOI21_X1 U10510 ( .B1(n9121), .B2(n9451), .A(n9120), .ZN(n9124) );
  INV_X1 U10511 ( .A(n9122), .ZN(n9123) );
  OAI21_X1 U10512 ( .B1(n9125), .B2(n9124), .A(n9123), .ZN(n9128) );
  AOI22_X1 U10513 ( .A1(n9128), .A2(n9127), .B1(n9126), .B2(n9305), .ZN(n9130)
         );
  AOI22_X1 U10514 ( .A1(n9131), .A2(n9130), .B1(n9129), .B2(n9299), .ZN(n9135)
         );
  INV_X1 U10515 ( .A(n9146), .ZN(n9134) );
  OAI211_X1 U10516 ( .C1(n9135), .C2(n9134), .A(n9133), .B(n9132), .ZN(n9138)
         );
  NAND4_X1 U10517 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9145), .ZN(n9151)
         );
  NAND3_X1 U10518 ( .A1(n9146), .A2(n9140), .A3(n9139), .ZN(n9141) );
  OAI211_X1 U10519 ( .C1(n9143), .C2(n9142), .A(n9141), .B(n9145), .ZN(n9150)
         );
  INV_X1 U10520 ( .A(n9144), .ZN(n9148) );
  NAND4_X1 U10521 ( .A1(n9148), .A2(n9147), .A3(n9146), .A4(n9145), .ZN(n9149)
         );
  NAND4_X1 U10522 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n9153)
         );
  OAI211_X1 U10523 ( .C1(n9156), .C2(n9155), .A(n9154), .B(n9153), .ZN(
        P1_U3242) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9157), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9330), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9337), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9360), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9371), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10529 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9393), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9403), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9424), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9433), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10533 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9454), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9464), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9453), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9492), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9158), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9527), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9159), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9529), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9160), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9161), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9162), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9163), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9164), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9165), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9167), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9168), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9169), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9170), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10552 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3556) );
  OAI211_X1 U10553 ( .C1(n9173), .C2(n9185), .A(n9755), .B(n9172), .ZN(n9181)
         );
  AOI22_X1 U10554 ( .A1(n9731), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9180) );
  OAI211_X1 U10555 ( .C1(n9176), .C2(n9175), .A(n9764), .B(n9174), .ZN(n9179)
         );
  NAND2_X1 U10556 ( .A1(n10329), .A2(n9177), .ZN(n9178) );
  NAND4_X1 U10557 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(
        P1_U3244) );
  AOI21_X1 U10558 ( .B1(n9729), .B2(n10051), .A(n9705), .ZN(n9728) );
  INV_X1 U10559 ( .A(n9182), .ZN(n9184) );
  MUX2_X1 U10560 ( .A(n9185), .B(n9184), .S(n9183), .Z(n9187) );
  NAND2_X1 U10561 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  OAI211_X1 U10562 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9728), .A(n9188), .B(
        P1_U3973), .ZN(n9227) );
  INV_X1 U10563 ( .A(n9189), .ZN(n9193) );
  INV_X1 U10564 ( .A(n9731), .ZN(n10333) );
  INV_X1 U10565 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9191) );
  OAI22_X1 U10566 ( .A1(n10333), .A2(n9191), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9190), .ZN(n9192) );
  AOI21_X1 U10567 ( .B1(n9193), .B2(n10329), .A(n9192), .ZN(n9202) );
  OAI211_X1 U10568 ( .C1(n9196), .C2(n9195), .A(n9755), .B(n9194), .ZN(n9201)
         );
  OAI211_X1 U10569 ( .C1(n9199), .C2(n9198), .A(n9764), .B(n9197), .ZN(n9200)
         );
  NAND4_X1 U10570 ( .A1(n9227), .A2(n9202), .A3(n9201), .A4(n9200), .ZN(
        P1_U3245) );
  OAI211_X1 U10571 ( .C1(n9205), .C2(n9204), .A(n9755), .B(n9203), .ZN(n9214)
         );
  AOI21_X1 U10572 ( .B1(n9731), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9206), .ZN(
        n9213) );
  OAI211_X1 U10573 ( .C1(n9209), .C2(n9208), .A(n9764), .B(n9207), .ZN(n9212)
         );
  NAND2_X1 U10574 ( .A1(n10329), .A2(n9210), .ZN(n9211) );
  NAND4_X1 U10575 ( .A1(n9214), .A2(n9213), .A3(n9212), .A4(n9211), .ZN(
        P1_U3246) );
  NOR2_X1 U10576 ( .A1(n9769), .A2(n9215), .ZN(n9216) );
  AOI211_X1 U10577 ( .C1(n9731), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9217), .B(
        n9216), .ZN(n9226) );
  OAI211_X1 U10578 ( .C1(n9220), .C2(n9219), .A(n9755), .B(n9218), .ZN(n9225)
         );
  OAI211_X1 U10579 ( .C1(n9223), .C2(n9222), .A(n9764), .B(n9221), .ZN(n9224)
         );
  NAND4_X1 U10580 ( .A1(n9227), .A2(n9226), .A3(n9225), .A4(n9224), .ZN(
        P1_U3247) );
  XNOR2_X1 U10581 ( .A(n9784), .B(n9228), .ZN(n9776) );
  OR2_X1 U10582 ( .A1(n9248), .A2(n9229), .ZN(n9231) );
  INV_X1 U10583 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U10584 ( .A1(n9248), .A2(n9229), .ZN(n9230) );
  NAND2_X1 U10585 ( .A1(n9231), .A2(n9230), .ZN(n9765) );
  OR2_X1 U10586 ( .A1(n9754), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9237) );
  OR2_X1 U10587 ( .A1(n9245), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U10588 ( .A1(n9233), .A2(n9232), .ZN(n9711) );
  INV_X1 U10589 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9234) );
  MUX2_X1 U10590 ( .A(n9234), .B(P1_REG1_REG_10__SCAN_IN), .S(n9717), .Z(n9710) );
  NOR2_X1 U10591 ( .A1(n9711), .A2(n9710), .ZN(n9720) );
  AOI21_X1 U10592 ( .B1(n9717), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9720), .ZN(
        n9740) );
  MUX2_X1 U10593 ( .A(n9235), .B(P1_REG1_REG_11__SCAN_IN), .S(n9743), .Z(n9739) );
  NOR2_X1 U10594 ( .A1(n9740), .A2(n9739), .ZN(n9738) );
  AOI21_X1 U10595 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9743), .A(n9738), .ZN(
        n9752) );
  MUX2_X1 U10596 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9236), .S(n9754), .Z(n9751) );
  NAND2_X1 U10597 ( .A1(n9752), .A2(n9751), .ZN(n9750) );
  AND2_X1 U10598 ( .A1(n9237), .A2(n9750), .ZN(n9766) );
  NAND2_X1 U10599 ( .A1(n9765), .A2(n9766), .ZN(n9763) );
  NAND2_X1 U10600 ( .A1(n9248), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U10601 ( .A1(n9763), .A2(n9238), .ZN(n9775) );
  AND2_X1 U10602 ( .A1(n9776), .A2(n9775), .ZN(n9778) );
  AOI21_X1 U10603 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9784), .A(n9778), .ZN(
        n9239) );
  NOR2_X1 U10604 ( .A1(n9239), .A2(n9250), .ZN(n9240) );
  XNOR2_X1 U10605 ( .A(n9250), .B(n9239), .ZN(n10322) );
  NOR2_X1 U10606 ( .A1(n10321), .A2(n10322), .ZN(n10320) );
  NOR2_X1 U10607 ( .A1(n9240), .A2(n10320), .ZN(n9269) );
  XNOR2_X1 U10608 ( .A(n9258), .B(n9241), .ZN(n9271) );
  XNOR2_X1 U10609 ( .A(n9269), .B(n9271), .ZN(n9262) );
  XNOR2_X1 U10610 ( .A(n9248), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9761) );
  NOR2_X1 U10611 ( .A1(n9754), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9242) );
  AOI21_X1 U10612 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9754), .A(n9242), .ZN(
        n9749) );
  XNOR2_X1 U10613 ( .A(n9717), .B(n9243), .ZN(n9714) );
  OAI21_X1 U10614 ( .B1(n9245), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9244), .ZN(
        n9246) );
  INV_X1 U10615 ( .A(n9246), .ZN(n9713) );
  NAND2_X1 U10616 ( .A1(n9743), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9247) );
  OAI21_X1 U10617 ( .B1(n9743), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9247), .ZN(
        n9736) );
  NAND2_X1 U10618 ( .A1(n9749), .A2(n9748), .ZN(n9747) );
  OAI21_X1 U10619 ( .B1(n9754), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9747), .ZN(
        n9762) );
  NAND2_X1 U10620 ( .A1(n9784), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9249) );
  OAI21_X1 U10621 ( .B1(n9784), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9249), .ZN(
        n9780) );
  NOR2_X1 U10622 ( .A1(n9251), .A2(n9250), .ZN(n9252) );
  XOR2_X1 U10623 ( .A(n10328), .B(n9251), .Z(n10325) );
  NOR2_X1 U10624 ( .A1(n6016), .A2(n10325), .ZN(n10324) );
  NOR2_X1 U10625 ( .A1(n9252), .A2(n10324), .ZN(n9255) );
  XNOR2_X1 U10626 ( .A(n9258), .B(n9253), .ZN(n9254) );
  AOI21_X1 U10627 ( .B1(n9255), .B2(n9254), .A(n10323), .ZN(n9260) );
  NAND2_X1 U10628 ( .A1(n9731), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9256) );
  OAI211_X1 U10629 ( .C1(n9769), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9259)
         );
  AOI21_X1 U10630 ( .B1(n9260), .B2(n9264), .A(n9259), .ZN(n9261) );
  OAI21_X1 U10631 ( .B1(n9262), .B2(n10319), .A(n9261), .ZN(P1_U3259) );
  NAND2_X1 U10632 ( .A1(n9270), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9263) );
  NOR2_X1 U10633 ( .A1(n9288), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9265) );
  AOI21_X1 U10634 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9288), .A(n9265), .ZN(
        n9266) );
  NAND2_X1 U10635 ( .A1(n9266), .A2(n9267), .ZN(n9287) );
  OAI21_X1 U10636 ( .B1(n9267), .B2(n9266), .A(n9287), .ZN(n9268) );
  INV_X1 U10637 ( .A(n9268), .ZN(n9281) );
  INV_X1 U10638 ( .A(n9269), .ZN(n9272) );
  OAI22_X1 U10639 ( .A1(n9272), .A2(n9271), .B1(n9270), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n9274) );
  AOI22_X1 U10640 ( .A1(n9288), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9632), .B2(
        n9277), .ZN(n9273) );
  NAND2_X1 U10641 ( .A1(n9273), .A2(n9274), .ZN(n9283) );
  OAI21_X1 U10642 ( .B1(n9274), .B2(n9273), .A(n9283), .ZN(n9279) );
  NAND2_X1 U10643 ( .A1(n9731), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9275) );
  OAI211_X1 U10644 ( .C1(n9769), .C2(n9277), .A(n9276), .B(n9275), .ZN(n9278)
         );
  AOI21_X1 U10645 ( .B1(n9279), .B2(n9764), .A(n9278), .ZN(n9280) );
  OAI21_X1 U10646 ( .B1(n9281), .B2(n10323), .A(n9280), .ZN(P1_U3260) );
  INV_X1 U10647 ( .A(n9282), .ZN(n9296) );
  NAND2_X1 U10648 ( .A1(n9799), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9285) );
  OAI21_X1 U10649 ( .B1(n9799), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9285), .ZN(
        n9791) );
  OR2_X1 U10650 ( .A1(n9288), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U10651 ( .A1(n9284), .A2(n9283), .ZN(n9792) );
  OR2_X1 U10652 ( .A1(n9791), .A2(n9792), .ZN(n9789) );
  NAND2_X1 U10653 ( .A1(n9789), .A2(n9285), .ZN(n9286) );
  XNOR2_X1 U10654 ( .A(n9286), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9294) );
  INV_X1 U10655 ( .A(n9294), .ZN(n9293) );
  NAND2_X1 U10656 ( .A1(n9799), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9289) );
  OAI21_X1 U10657 ( .B1(n9799), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9289), .ZN(
        n9795) );
  OAI21_X1 U10658 ( .B1(n9288), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9287), .ZN(
        n9796) );
  OR2_X1 U10659 ( .A1(n9795), .A2(n9796), .ZN(n9793) );
  NAND2_X1 U10660 ( .A1(n9793), .A2(n9289), .ZN(n9290) );
  XNOR2_X1 U10661 ( .A(n9290), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U10662 ( .A1(n9291), .A2(n9295), .ZN(n9292) );
  NOR2_X1 U10663 ( .A1(n9304), .A2(n9305), .ZN(n9303) );
  XNOR2_X1 U10664 ( .A(n9303), .B(n9656), .ZN(n9297) );
  NOR2_X1 U10665 ( .A1(n9297), .A2(n9557), .ZN(n9566) );
  NAND2_X1 U10666 ( .A1(n9566), .A2(n9805), .ZN(n9302) );
  AND3_X1 U10667 ( .A1(n9528), .A2(n9299), .A3(n9298), .ZN(n9569) );
  INV_X1 U10668 ( .A(n9569), .ZN(n9300) );
  NOR2_X1 U10669 ( .A1(n9521), .A2(n9300), .ZN(n9306) );
  AOI21_X1 U10670 ( .B1(n9521), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9306), .ZN(
        n9301) );
  OAI211_X1 U10671 ( .C1(n9656), .C2(n9811), .A(n9302), .B(n9301), .ZN(
        P1_U3263) );
  INV_X1 U10672 ( .A(n9305), .ZN(n9660) );
  AOI211_X1 U10673 ( .C1(n9305), .C2(n9304), .A(n9557), .B(n9303), .ZN(n9570)
         );
  NAND2_X1 U10674 ( .A1(n9570), .A2(n9805), .ZN(n9308) );
  AOI21_X1 U10675 ( .B1(n9521), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9306), .ZN(
        n9307) );
  OAI211_X1 U10676 ( .C1(n9660), .C2(n9811), .A(n9308), .B(n9307), .ZN(
        P1_U3264) );
  NAND2_X1 U10677 ( .A1(n9521), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9310) );
  OAI21_X1 U10678 ( .B1(n9499), .B2(n9311), .A(n9310), .ZN(n9312) );
  AOI21_X1 U10679 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9315) );
  OAI21_X1 U10680 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9318) );
  AOI21_X1 U10681 ( .B1(n9319), .B2(n9513), .A(n9318), .ZN(n9320) );
  OAI21_X1 U10682 ( .B1(n9321), .B2(n9521), .A(n9320), .ZN(P1_U3356) );
  INV_X1 U10683 ( .A(n9574), .ZN(n9326) );
  INV_X1 U10684 ( .A(n9323), .ZN(n9324) );
  AOI22_X1 U10685 ( .A1(n9521), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9324), .B2(
        n9807), .ZN(n9325) );
  OAI21_X1 U10686 ( .B1(n9326), .B2(n9811), .A(n9325), .ZN(n9333) );
  OAI21_X1 U10687 ( .B1(n9329), .B2(n9328), .A(n9327), .ZN(n9331) );
  AOI211_X1 U10688 ( .C1(n9573), .C2(n9805), .A(n9333), .B(n9332), .ZN(n9334)
         );
  OAI21_X1 U10689 ( .B1(n9577), .B2(n9541), .A(n9334), .ZN(P1_U3265) );
  OAI21_X1 U10690 ( .B1(n9339), .B2(n9336), .A(n9335), .ZN(n9338) );
  AOI222_X1 U10691 ( .A1(n9523), .A2(n9338), .B1(n9371), .B2(n9530), .C1(n9337), .C2(n9528), .ZN(n9578) );
  NAND2_X1 U10692 ( .A1(n9581), .A2(n9513), .ZN(n9347) );
  AOI21_X1 U10693 ( .B1(n9350), .B2(n9341), .A(n9557), .ZN(n9342) );
  AOI22_X1 U10694 ( .A1(n9521), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9343), .B2(
        n9807), .ZN(n9344) );
  OAI21_X1 U10695 ( .B1(n9664), .B2(n9811), .A(n9344), .ZN(n9345) );
  AOI21_X1 U10696 ( .B1(n9580), .B2(n9805), .A(n9345), .ZN(n9346) );
  OAI211_X1 U10697 ( .C1(n9521), .C2(n9578), .A(n9347), .B(n9346), .ZN(
        P1_U3266) );
  XNOR2_X1 U10698 ( .A(n9349), .B(n9348), .ZN(n9588) );
  INV_X1 U10699 ( .A(n9374), .ZN(n9352) );
  INV_X1 U10700 ( .A(n9350), .ZN(n9351) );
  AOI211_X1 U10701 ( .C1(n9585), .C2(n9352), .A(n9557), .B(n9351), .ZN(n9584)
         );
  INV_X1 U10702 ( .A(n9353), .ZN(n9354) );
  AOI22_X1 U10703 ( .A1(n9521), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9354), .B2(
        n9807), .ZN(n9355) );
  OAI21_X1 U10704 ( .B1(n9356), .B2(n9811), .A(n9355), .ZN(n9363) );
  OAI21_X1 U10705 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9361) );
  AOI222_X1 U10706 ( .A1(n9523), .A2(n9361), .B1(n9393), .B2(n9530), .C1(n9360), .C2(n9528), .ZN(n9587) );
  NOR2_X1 U10707 ( .A1(n9587), .A2(n9521), .ZN(n9362) );
  AOI211_X1 U10708 ( .C1(n9584), .C2(n9805), .A(n9363), .B(n9362), .ZN(n9364)
         );
  OAI21_X1 U10709 ( .B1(n9588), .B2(n9541), .A(n9364), .ZN(P1_U3267) );
  XOR2_X1 U10710 ( .A(n9366), .B(n9365), .Z(n9591) );
  INV_X1 U10711 ( .A(n9591), .ZN(n9381) );
  NAND2_X1 U10712 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NAND2_X1 U10713 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U10714 ( .A1(n9370), .A2(n9523), .ZN(n9373) );
  AOI22_X1 U10715 ( .A1(n9403), .A2(n9530), .B1(n9528), .B2(n9371), .ZN(n9372)
         );
  NAND2_X1 U10716 ( .A1(n9373), .A2(n9372), .ZN(n9589) );
  AOI211_X1 U10717 ( .C1(n9375), .C2(n9384), .A(n9557), .B(n9374), .ZN(n9590)
         );
  NAND2_X1 U10718 ( .A1(n9590), .A2(n9805), .ZN(n9378) );
  AOI22_X1 U10719 ( .A1(n9376), .A2(n9807), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9521), .ZN(n9377) );
  OAI211_X1 U10720 ( .C1(n9669), .C2(n9811), .A(n9378), .B(n9377), .ZN(n9379)
         );
  AOI21_X1 U10721 ( .B1(n9502), .B2(n9589), .A(n9379), .ZN(n9380) );
  OAI21_X1 U10722 ( .B1(n9381), .B2(n9541), .A(n9380), .ZN(P1_U3268) );
  XNOR2_X1 U10723 ( .A(n9382), .B(n9391), .ZN(n9598) );
  INV_X1 U10724 ( .A(n9384), .ZN(n9385) );
  AOI211_X1 U10725 ( .C1(n9595), .C2(n9406), .A(n9557), .B(n9385), .ZN(n9594)
         );
  INV_X1 U10726 ( .A(n9595), .ZN(n9389) );
  INV_X1 U10727 ( .A(n9386), .ZN(n9387) );
  AOI22_X1 U10728 ( .A1(n9387), .A2(n9807), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9521), .ZN(n9388) );
  OAI21_X1 U10729 ( .B1(n9389), .B2(n9811), .A(n9388), .ZN(n9396) );
  NAND2_X1 U10730 ( .A1(n9399), .A2(n9390), .ZN(n9392) );
  XNOR2_X1 U10731 ( .A(n9392), .B(n9391), .ZN(n9394) );
  AOI222_X1 U10732 ( .A1(n9523), .A2(n9394), .B1(n9393), .B2(n9528), .C1(n9424), .C2(n9530), .ZN(n9597) );
  NOR2_X1 U10733 ( .A1(n9597), .A2(n9521), .ZN(n9395) );
  AOI211_X1 U10734 ( .C1(n9594), .C2(n9805), .A(n9396), .B(n9395), .ZN(n9397)
         );
  OAI21_X1 U10735 ( .B1(n9598), .B2(n9541), .A(n9397), .ZN(P1_U3269) );
  XNOR2_X1 U10736 ( .A(n9398), .B(n9401), .ZN(n9601) );
  INV_X1 U10737 ( .A(n9601), .ZN(n9413) );
  OAI21_X1 U10738 ( .B1(n9401), .B2(n9400), .A(n9399), .ZN(n9402) );
  NAND2_X1 U10739 ( .A1(n9402), .A2(n9523), .ZN(n9405) );
  AOI22_X1 U10740 ( .A1(n9403), .A2(n9528), .B1(n9530), .B2(n9433), .ZN(n9404)
         );
  NAND2_X1 U10741 ( .A1(n9405), .A2(n9404), .ZN(n9599) );
  AOI211_X1 U10742 ( .C1(n9407), .C2(n9415), .A(n9557), .B(n9383), .ZN(n9600)
         );
  NAND2_X1 U10743 ( .A1(n9600), .A2(n9805), .ZN(n9410) );
  AOI22_X1 U10744 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n9521), .B1(n9408), .B2(
        n9807), .ZN(n9409) );
  OAI211_X1 U10745 ( .C1(n9673), .C2(n9811), .A(n9410), .B(n9409), .ZN(n9411)
         );
  AOI21_X1 U10746 ( .B1(n9502), .B2(n9599), .A(n9411), .ZN(n9412) );
  OAI21_X1 U10747 ( .B1(n9413), .B2(n9541), .A(n9412), .ZN(P1_U3270) );
  XNOR2_X1 U10748 ( .A(n9414), .B(n9423), .ZN(n9608) );
  INV_X1 U10749 ( .A(n9415), .ZN(n9416) );
  AOI211_X1 U10750 ( .C1(n9605), .C2(n4585), .A(n9557), .B(n9416), .ZN(n9604)
         );
  INV_X1 U10751 ( .A(n9417), .ZN(n9418) );
  AOI22_X1 U10752 ( .A1(n9521), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9418), .B2(
        n9807), .ZN(n9419) );
  OAI21_X1 U10753 ( .B1(n9420), .B2(n9811), .A(n9419), .ZN(n9427) );
  OAI21_X1 U10754 ( .B1(n9423), .B2(n9422), .A(n9421), .ZN(n9425) );
  AOI222_X1 U10755 ( .A1(n9523), .A2(n9425), .B1(n9424), .B2(n9528), .C1(n9454), .C2(n9530), .ZN(n9607) );
  NOR2_X1 U10756 ( .A1(n9607), .A2(n9521), .ZN(n9426) );
  AOI211_X1 U10757 ( .C1(n9604), .C2(n9805), .A(n9427), .B(n9426), .ZN(n9428)
         );
  OAI21_X1 U10758 ( .B1(n9608), .B2(n9541), .A(n9428), .ZN(P1_U3271) );
  XOR2_X1 U10759 ( .A(n9430), .B(n4437), .Z(n9611) );
  INV_X1 U10760 ( .A(n9611), .ZN(n9443) );
  OAI21_X1 U10761 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  NAND2_X1 U10762 ( .A1(n9432), .A2(n9523), .ZN(n9435) );
  AOI22_X1 U10763 ( .A1(n9433), .A2(n9528), .B1(n9530), .B2(n9464), .ZN(n9434)
         );
  NAND2_X1 U10764 ( .A1(n9435), .A2(n9434), .ZN(n9609) );
  AOI211_X1 U10765 ( .C1(n9437), .C2(n9445), .A(n9557), .B(n9436), .ZN(n9610)
         );
  NAND2_X1 U10766 ( .A1(n9610), .A2(n9805), .ZN(n9440) );
  AOI22_X1 U10767 ( .A1(n9521), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9438), .B2(
        n9807), .ZN(n9439) );
  OAI211_X1 U10768 ( .C1(n4583), .C2(n9811), .A(n9440), .B(n9439), .ZN(n9441)
         );
  AOI21_X1 U10769 ( .B1(n9502), .B2(n9609), .A(n9441), .ZN(n9442) );
  OAI21_X1 U10770 ( .B1(n9443), .B2(n9541), .A(n9442), .ZN(P1_U3272) );
  XNOR2_X1 U10771 ( .A(n9444), .B(n9452), .ZN(n9617) );
  INV_X1 U10772 ( .A(n9445), .ZN(n9446) );
  AOI211_X1 U10773 ( .C1(n9614), .C2(n9468), .A(n9557), .B(n9446), .ZN(n9613)
         );
  INV_X1 U10774 ( .A(n9447), .ZN(n9448) );
  AOI22_X1 U10775 ( .A1(n9521), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9448), .B2(
        n9807), .ZN(n9449) );
  OAI21_X1 U10776 ( .B1(n9450), .B2(n9811), .A(n9449), .ZN(n9457) );
  XOR2_X1 U10777 ( .A(n9452), .B(n9451), .Z(n9455) );
  AOI222_X1 U10778 ( .A1(n9523), .A2(n9455), .B1(n9454), .B2(n9528), .C1(n9453), .C2(n9530), .ZN(n9616) );
  NOR2_X1 U10779 ( .A1(n9616), .A2(n9521), .ZN(n9456) );
  AOI211_X1 U10780 ( .C1(n9613), .C2(n9805), .A(n9457), .B(n9456), .ZN(n9458)
         );
  OAI21_X1 U10781 ( .B1(n9617), .B2(n9541), .A(n9458), .ZN(P1_U3273) );
  XNOR2_X1 U10782 ( .A(n9459), .B(n9462), .ZN(n9620) );
  INV_X1 U10783 ( .A(n9620), .ZN(n9476) );
  OAI21_X1 U10784 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9463) );
  NAND2_X1 U10785 ( .A1(n9463), .A2(n9523), .ZN(n9466) );
  AOI22_X1 U10786 ( .A1(n9464), .A2(n9528), .B1(n9530), .B2(n9492), .ZN(n9465)
         );
  NAND2_X1 U10787 ( .A1(n9466), .A2(n9465), .ZN(n9618) );
  INV_X1 U10788 ( .A(n9467), .ZN(n9478) );
  INV_X1 U10789 ( .A(n9468), .ZN(n9469) );
  AOI211_X1 U10790 ( .C1(n9470), .C2(n9478), .A(n9557), .B(n9469), .ZN(n9619)
         );
  NAND2_X1 U10791 ( .A1(n9619), .A2(n9805), .ZN(n9473) );
  AOI22_X1 U10792 ( .A1(n9521), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9471), .B2(
        n9807), .ZN(n9472) );
  OAI211_X1 U10793 ( .C1(n6177), .C2(n9811), .A(n9473), .B(n9472), .ZN(n9474)
         );
  AOI21_X1 U10794 ( .B1(n9502), .B2(n9618), .A(n9474), .ZN(n9475) );
  OAI21_X1 U10795 ( .B1(n9476), .B2(n9541), .A(n9475), .ZN(P1_U3274) );
  XNOR2_X1 U10796 ( .A(n9477), .B(n9485), .ZN(n9628) );
  AOI211_X1 U10797 ( .C1(n9625), .C2(n9496), .A(n9557), .B(n9467), .ZN(n9624)
         );
  NOR2_X1 U10798 ( .A1(n9479), .A2(n9811), .ZN(n9483) );
  INV_X1 U10799 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9481) );
  OAI22_X1 U10800 ( .A1(n9502), .A2(n9481), .B1(n9480), .B2(n9499), .ZN(n9482)
         );
  AOI211_X1 U10801 ( .C1(n9624), .C2(n9805), .A(n9483), .B(n9482), .ZN(n9489)
         );
  AOI21_X1 U10802 ( .B1(n9485), .B2(n9484), .A(n4487), .ZN(n9486) );
  OAI222_X1 U10803 ( .A1(n9549), .A2(n9487), .B1(n9551), .B2(n9510), .C1(n9546), .C2(n9486), .ZN(n9623) );
  NAND2_X1 U10804 ( .A1(n9623), .A2(n9502), .ZN(n9488) );
  OAI211_X1 U10805 ( .C1(n9628), .C2(n9541), .A(n9489), .B(n9488), .ZN(
        P1_U3275) );
  XNOR2_X1 U10806 ( .A(n9490), .B(n4876), .ZN(n9491) );
  NAND2_X1 U10807 ( .A1(n9491), .A2(n9523), .ZN(n9494) );
  AOI22_X1 U10808 ( .A1(n9492), .A2(n9528), .B1(n9530), .B2(n9527), .ZN(n9493)
         );
  NAND2_X1 U10809 ( .A1(n9494), .A2(n9493), .ZN(n9629) );
  INV_X1 U10810 ( .A(n9629), .ZN(n9507) );
  XOR2_X1 U10811 ( .A(n9495), .B(n4483), .Z(n9631) );
  NAND2_X1 U10812 ( .A1(n9631), .A2(n9513), .ZN(n9506) );
  INV_X1 U10813 ( .A(n9496), .ZN(n9497) );
  AOI211_X1 U10814 ( .C1(n9498), .C2(n4575), .A(n9557), .B(n9497), .ZN(n9630)
         );
  NOR2_X1 U10815 ( .A1(n9685), .A2(n9811), .ZN(n9504) );
  OAI22_X1 U10816 ( .A1(n9502), .A2(n9501), .B1(n9500), .B2(n9499), .ZN(n9503)
         );
  AOI211_X1 U10817 ( .C1(n9630), .C2(n9805), .A(n9504), .B(n9503), .ZN(n9505)
         );
  OAI211_X1 U10818 ( .C1(n9521), .C2(n9507), .A(n9506), .B(n9505), .ZN(
        P1_U3276) );
  XNOR2_X1 U10819 ( .A(n9508), .B(n9511), .ZN(n9509) );
  OAI222_X1 U10820 ( .A1(n9549), .A2(n9510), .B1(n9551), .B2(n9550), .C1(n9546), .C2(n9509), .ZN(n9635) );
  INV_X1 U10821 ( .A(n9635), .ZN(n9520) );
  NAND2_X1 U10822 ( .A1(n9512), .A2(n9511), .ZN(n9634) );
  NAND3_X1 U10823 ( .A1(n4851), .A2(n9513), .A3(n9634), .ZN(n9519) );
  AOI211_X1 U10824 ( .C1(n9637), .C2(n9533), .A(n9557), .B(n9514), .ZN(n9636)
         );
  AOI22_X1 U10825 ( .A1(n9521), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9515), .B2(
        n9807), .ZN(n9516) );
  OAI21_X1 U10826 ( .B1(n4573), .B2(n9811), .A(n9516), .ZN(n9517) );
  AOI21_X1 U10827 ( .B1(n9636), .B2(n9805), .A(n9517), .ZN(n9518) );
  OAI211_X1 U10828 ( .C1(n9521), .C2(n9520), .A(n9519), .B(n9518), .ZN(
        P1_U3277) );
  XNOR2_X1 U10829 ( .A(n9522), .B(n9525), .ZN(n9643) );
  INV_X1 U10830 ( .A(n9643), .ZN(n9542) );
  OAI211_X1 U10831 ( .C1(n9526), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9532)
         );
  AOI22_X1 U10832 ( .A1(n9530), .A2(n9529), .B1(n9528), .B2(n9527), .ZN(n9531)
         );
  NAND2_X1 U10833 ( .A1(n9532), .A2(n9531), .ZN(n9641) );
  INV_X1 U10834 ( .A(n9533), .ZN(n9534) );
  AOI211_X1 U10835 ( .C1(n9535), .C2(n9555), .A(n9557), .B(n9534), .ZN(n9642)
         );
  NAND2_X1 U10836 ( .A1(n9642), .A2(n9805), .ZN(n9538) );
  AOI22_X1 U10837 ( .A1(n9521), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9536), .B2(
        n9807), .ZN(n9537) );
  OAI211_X1 U10838 ( .C1(n9690), .C2(n9811), .A(n9538), .B(n9537), .ZN(n9539)
         );
  AOI21_X1 U10839 ( .B1(n9502), .B2(n9641), .A(n9539), .ZN(n9540) );
  OAI21_X1 U10840 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(P1_U3278) );
  XNOR2_X1 U10841 ( .A(n9543), .B(n9544), .ZN(n9562) );
  NAND2_X1 U10842 ( .A1(n9545), .A2(n9544), .ZN(n9547) );
  AOI21_X1 U10843 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9553) );
  OAI22_X1 U10844 ( .A1(n5993), .A2(n9551), .B1(n9550), .B2(n9549), .ZN(n9552)
         );
  AOI211_X1 U10845 ( .C1(n9562), .C2(n9554), .A(n9553), .B(n9552), .ZN(n9650)
         );
  INV_X1 U10846 ( .A(n9555), .ZN(n9556) );
  AOI211_X1 U10847 ( .C1(n9647), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9646)
         );
  AOI22_X1 U10848 ( .A1(n9521), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9559), .B2(
        n9807), .ZN(n9560) );
  OAI21_X1 U10849 ( .B1(n9561), .B2(n9811), .A(n9560), .ZN(n9564) );
  INV_X1 U10850 ( .A(n9562), .ZN(n9652) );
  NOR2_X1 U10851 ( .A1(n9652), .A2(n9803), .ZN(n9563) );
  AOI211_X1 U10852 ( .C1(n9646), .C2(n9805), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OAI21_X1 U10853 ( .B1(n9521), .B2(n9650), .A(n9565), .ZN(P1_U3279) );
  INV_X1 U10854 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9567) );
  NOR2_X1 U10855 ( .A1(n9566), .A2(n9569), .ZN(n9653) );
  MUX2_X1 U10856 ( .A(n9567), .B(n9653), .S(n9845), .Z(n9568) );
  OAI21_X1 U10857 ( .B1(n9656), .B2(n9645), .A(n9568), .ZN(P1_U3553) );
  INV_X1 U10858 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9571) );
  NOR2_X1 U10859 ( .A1(n9570), .A2(n9569), .ZN(n9657) );
  MUX2_X1 U10860 ( .A(n9571), .B(n9657), .S(n9845), .Z(n9572) );
  OAI21_X1 U10861 ( .B1(n9660), .B2(n9645), .A(n9572), .ZN(P1_U3552) );
  AOI21_X1 U10862 ( .B1(n9648), .B2(n9574), .A(n9573), .ZN(n9575) );
  OAI211_X1 U10863 ( .C1(n9577), .C2(n9627), .A(n9576), .B(n9575), .ZN(n9661)
         );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9661), .S(n9845), .Z(
        P1_U3550) );
  INV_X1 U10865 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9582) );
  INV_X1 U10866 ( .A(n9578), .ZN(n9579) );
  MUX2_X1 U10867 ( .A(n9582), .B(n9662), .S(n9845), .Z(n9583) );
  OAI21_X1 U10868 ( .B1(n9664), .B2(n9645), .A(n9583), .ZN(P1_U3549) );
  AOI21_X1 U10869 ( .B1(n9648), .B2(n9585), .A(n9584), .ZN(n9586) );
  OAI211_X1 U10870 ( .C1(n9588), .C2(n9627), .A(n9587), .B(n9586), .ZN(n9665)
         );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9665), .S(n9845), .Z(
        P1_U3548) );
  MUX2_X1 U10872 ( .A(n9592), .B(n9666), .S(n9845), .Z(n9593) );
  OAI21_X1 U10873 ( .B1(n9669), .B2(n9645), .A(n9593), .ZN(P1_U3547) );
  AOI21_X1 U10874 ( .B1(n9648), .B2(n9595), .A(n9594), .ZN(n9596) );
  OAI211_X1 U10875 ( .C1(n9598), .C2(n9627), .A(n9597), .B(n9596), .ZN(n9670)
         );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9670), .S(n9845), .Z(
        P1_U3546) );
  INV_X1 U10877 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9602) );
  AOI211_X1 U10878 ( .C1(n9601), .C2(n9836), .A(n9600), .B(n9599), .ZN(n9671)
         );
  MUX2_X1 U10879 ( .A(n9602), .B(n9671), .S(n9845), .Z(n9603) );
  OAI21_X1 U10880 ( .B1(n9673), .B2(n9645), .A(n9603), .ZN(P1_U3545) );
  AOI21_X1 U10881 ( .B1(n9648), .B2(n9605), .A(n9604), .ZN(n9606) );
  OAI211_X1 U10882 ( .C1(n9608), .C2(n9627), .A(n9607), .B(n9606), .ZN(n9674)
         );
  MUX2_X1 U10883 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9674), .S(n9845), .Z(
        P1_U3544) );
  AOI211_X1 U10884 ( .C1(n9611), .C2(n9836), .A(n9610), .B(n9609), .ZN(n9675)
         );
  MUX2_X1 U10885 ( .A(n10123), .B(n9675), .S(n9845), .Z(n9612) );
  OAI21_X1 U10886 ( .B1(n4583), .B2(n9645), .A(n9612), .ZN(P1_U3543) );
  AOI21_X1 U10887 ( .B1(n9648), .B2(n9614), .A(n9613), .ZN(n9615) );
  OAI211_X1 U10888 ( .C1(n9617), .C2(n9627), .A(n9616), .B(n9615), .ZN(n9678)
         );
  MUX2_X1 U10889 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9678), .S(n9845), .Z(
        P1_U3542) );
  INV_X1 U10890 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9621) );
  AOI211_X1 U10891 ( .C1(n9620), .C2(n9836), .A(n9619), .B(n9618), .ZN(n9679)
         );
  MUX2_X1 U10892 ( .A(n9621), .B(n9679), .S(n9845), .Z(n9622) );
  OAI21_X1 U10893 ( .B1(n6177), .B2(n9645), .A(n9622), .ZN(P1_U3541) );
  AOI211_X1 U10894 ( .C1(n9648), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9626)
         );
  OAI21_X1 U10895 ( .B1(n9628), .B2(n9627), .A(n9626), .ZN(n9681) );
  MUX2_X1 U10896 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9681), .S(n9845), .Z(
        P1_U3540) );
  AOI211_X1 U10897 ( .C1(n9631), .C2(n9836), .A(n9630), .B(n9629), .ZN(n9682)
         );
  MUX2_X1 U10898 ( .A(n9632), .B(n9682), .S(n9845), .Z(n9633) );
  OAI21_X1 U10899 ( .B1(n9685), .B2(n9645), .A(n9633), .ZN(P1_U3539) );
  NAND2_X1 U10900 ( .A1(n9634), .A2(n9836), .ZN(n9639) );
  AOI211_X1 U10901 ( .C1(n9648), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9638)
         );
  OAI21_X1 U10902 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9686) );
  MUX2_X1 U10903 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9686), .S(n9845), .Z(
        P1_U3538) );
  AOI211_X1 U10904 ( .C1(n9643), .C2(n9836), .A(n9642), .B(n9641), .ZN(n9687)
         );
  MUX2_X1 U10905 ( .A(n10321), .B(n9687), .S(n9845), .Z(n9644) );
  OAI21_X1 U10906 ( .B1(n9690), .B2(n9645), .A(n9644), .ZN(P1_U3537) );
  AOI21_X1 U10907 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  OAI211_X1 U10908 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9692)
         );
  MUX2_X1 U10909 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9692), .S(n9845), .Z(
        P1_U3536) );
  MUX2_X1 U10910 ( .A(n9654), .B(n9653), .S(n9691), .Z(n9655) );
  OAI21_X1 U10911 ( .B1(n9656), .B2(n9689), .A(n9655), .ZN(P1_U3521) );
  MUX2_X1 U10912 ( .A(n9658), .B(n9657), .S(n9839), .Z(n9659) );
  OAI21_X1 U10913 ( .B1(n9660), .B2(n9689), .A(n9659), .ZN(P1_U3520) );
  MUX2_X1 U10914 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9661), .S(n9839), .Z(
        P1_U3518) );
  MUX2_X1 U10915 ( .A(n10098), .B(n9662), .S(n9839), .Z(n9663) );
  OAI21_X1 U10916 ( .B1(n9664), .B2(n9689), .A(n9663), .ZN(P1_U3517) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9665), .S(n9839), .Z(
        P1_U3516) );
  INV_X1 U10918 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9667) );
  MUX2_X1 U10919 ( .A(n9667), .B(n9666), .S(n9839), .Z(n9668) );
  OAI21_X1 U10920 ( .B1(n9669), .B2(n9689), .A(n9668), .ZN(P1_U3515) );
  MUX2_X1 U10921 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9670), .S(n9839), .Z(
        P1_U3514) );
  MUX2_X1 U10922 ( .A(n10165), .B(n9671), .S(n9691), .Z(n9672) );
  OAI21_X1 U10923 ( .B1(n9673), .B2(n9689), .A(n9672), .ZN(P1_U3513) );
  MUX2_X1 U10924 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9674), .S(n9691), .Z(
        P1_U3512) );
  INV_X1 U10925 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9676) );
  MUX2_X1 U10926 ( .A(n9676), .B(n9675), .S(n9691), .Z(n9677) );
  OAI21_X1 U10927 ( .B1(n4583), .B2(n9689), .A(n9677), .ZN(P1_U3511) );
  MUX2_X1 U10928 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9678), .S(n9691), .Z(
        P1_U3510) );
  MUX2_X1 U10929 ( .A(n10236), .B(n9679), .S(n9691), .Z(n9680) );
  OAI21_X1 U10930 ( .B1(n6177), .B2(n9689), .A(n9680), .ZN(P1_U3509) );
  MUX2_X1 U10931 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9681), .S(n9691), .Z(
        P1_U3507) );
  INV_X1 U10932 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9683) );
  MUX2_X1 U10933 ( .A(n9683), .B(n9682), .S(n9691), .Z(n9684) );
  OAI21_X1 U10934 ( .B1(n9685), .B2(n9689), .A(n9684), .ZN(P1_U3504) );
  MUX2_X1 U10935 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9686), .S(n9691), .Z(
        P1_U3501) );
  MUX2_X1 U10936 ( .A(n10223), .B(n9687), .S(n9691), .Z(n9688) );
  OAI21_X1 U10937 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(P1_U3498) );
  MUX2_X1 U10938 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9692), .S(n9691), .Z(
        P1_U3495) );
  MUX2_X1 U10939 ( .A(P1_D_REG_0__SCAN_IN), .B(n9694), .S(n9693), .Z(P1_U3439)
         );
  INV_X1 U10940 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10296) );
  NAND4_X1 U10941 ( .A1(n10296), .A2(n9695), .A3(P1_IR_REG_31__SCAN_IN), .A4(
        P1_STATE_REG_SCAN_IN), .ZN(n9696) );
  OAI22_X1 U10942 ( .A1(n9697), .A2(n9696), .B1(n10195), .B2(n9709), .ZN(n9698) );
  INV_X1 U10943 ( .A(n9698), .ZN(n9699) );
  OAI21_X1 U10944 ( .B1(n9700), .B2(n9707), .A(n9699), .ZN(P1_U3324) );
  OAI222_X1 U10945 ( .A1(n9709), .A2(n9703), .B1(n9707), .B2(n9702), .C1(n9701), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U10946 ( .A(n9704), .ZN(n9706) );
  OAI222_X1 U10947 ( .A1(n9709), .A2(n9708), .B1(n9707), .B2(n9706), .C1(n9705), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U10948 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U10949 ( .A1(n9711), .A2(n9710), .ZN(n9712) );
  NAND2_X1 U10950 ( .A1(n9764), .A2(n9712), .ZN(n9721) );
  NOR2_X1 U10951 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  OR3_X1 U10952 ( .A1(n10323), .A2(n9716), .A3(n9715), .ZN(n9719) );
  NAND2_X1 U10953 ( .A1(n10329), .A2(n9717), .ZN(n9718) );
  OAI211_X1 U10954 ( .C1(n9721), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9722)
         );
  INV_X1 U10955 ( .A(n9722), .ZN(n9725) );
  INV_X1 U10956 ( .A(n9723), .ZN(n9724) );
  OAI211_X1 U10957 ( .C1(n10333), .C2(n9726), .A(n9725), .B(n9724), .ZN(
        P1_U3253) );
  XNOR2_X1 U10958 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U10959 ( .B1(n9729), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9728), .ZN(
        n9730) );
  XNOR2_X1 U10960 ( .A(n9730), .B(n5016), .ZN(n9733) );
  AOI22_X1 U10961 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9731), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9732) );
  OAI21_X1 U10962 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(P1_U3243) );
  AOI211_X1 U10963 ( .C1(n9737), .C2(n9736), .A(n9735), .B(n10323), .ZN(n9742)
         );
  AOI211_X1 U10964 ( .C1(n9740), .C2(n9739), .A(n10319), .B(n9738), .ZN(n9741)
         );
  AOI211_X1 U10965 ( .C1(n10329), .C2(n9743), .A(n9742), .B(n9741), .ZN(n9746)
         );
  INV_X1 U10966 ( .A(n9744), .ZN(n9745) );
  OAI211_X1 U10967 ( .C1(n10333), .C2(n10175), .A(n9746), .B(n9745), .ZN(
        P1_U3254) );
  INV_X1 U10968 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9759) );
  OAI21_X1 U10969 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9756) );
  OAI21_X1 U10970 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9753) );
  AOI222_X1 U10971 ( .A1(n9756), .A2(n9755), .B1(n9754), .B2(n10329), .C1(
        n9753), .C2(n9764), .ZN(n9758) );
  OAI211_X1 U10972 ( .C1(n10333), .C2(n9759), .A(n9758), .B(n9757), .ZN(
        P1_U3255) );
  INV_X1 U10973 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9774) );
  AOI211_X1 U10974 ( .C1(n9762), .C2(n9761), .A(n9760), .B(n10323), .ZN(n9771)
         );
  OAI211_X1 U10975 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9767)
         );
  OAI21_X1 U10976 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  NOR2_X1 U10977 ( .A1(n9771), .A2(n9770), .ZN(n9773) );
  OAI211_X1 U10978 ( .C1(n10333), .C2(n9774), .A(n9773), .B(n9772), .ZN(
        P1_U3256) );
  INV_X1 U10979 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9788) );
  NOR2_X1 U10980 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  NOR3_X1 U10981 ( .A1(n10319), .A2(n9778), .A3(n9777), .ZN(n9783) );
  AOI211_X1 U10982 ( .C1(n9781), .C2(n9780), .A(n9779), .B(n10323), .ZN(n9782)
         );
  AOI211_X1 U10983 ( .C1(n10329), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9787)
         );
  INV_X1 U10984 ( .A(n9785), .ZN(n9786) );
  OAI211_X1 U10985 ( .C1(n10333), .C2(n9788), .A(n9787), .B(n9786), .ZN(
        P1_U3257) );
  INV_X1 U10986 ( .A(n9789), .ZN(n9790) );
  AOI211_X1 U10987 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n10319), .ZN(n9798)
         );
  INV_X1 U10988 ( .A(n9793), .ZN(n9794) );
  AOI211_X1 U10989 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n10323), .ZN(n9797)
         );
  AOI211_X1 U10990 ( .C1(n10329), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9801)
         );
  OAI211_X1 U10991 ( .C1(n10333), .C2(n9802), .A(n9801), .B(n9800), .ZN(
        P1_U3261) );
  INV_X1 U10992 ( .A(n9803), .ZN(n9814) );
  INV_X1 U10993 ( .A(n9804), .ZN(n9812) );
  NAND2_X1 U10994 ( .A1(n9806), .A2(n9805), .ZN(n9810) );
  AOI22_X1 U10995 ( .A1(n9521), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9808), .B2(
        n9807), .ZN(n9809) );
  OAI211_X1 U10996 ( .C1(n9812), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9813)
         );
  AOI21_X1 U10997 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9816) );
  OAI21_X1 U10998 ( .B1(n9521), .B2(n9817), .A(n9816), .ZN(P1_U3286) );
  AND2_X1 U10999 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9818), .ZN(P1_U3294) );
  AND2_X1 U11000 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9818), .ZN(P1_U3295) );
  NOR2_X1 U11001 ( .A1(n9819), .A2(n10161), .ZN(P1_U3296) );
  AND2_X1 U11002 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9818), .ZN(P1_U3297) );
  NOR2_X1 U11003 ( .A1(n9819), .A2(n10206), .ZN(P1_U3298) );
  INV_X1 U11004 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11005 ( .A1(n9819), .A2(n10141), .ZN(P1_U3299) );
  AND2_X1 U11006 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9818), .ZN(P1_U3300) );
  INV_X1 U11007 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U11008 ( .A1(n9819), .A2(n10093), .ZN(P1_U3301) );
  INV_X1 U11009 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U11010 ( .A1(n9819), .A2(n10210), .ZN(P1_U3302) );
  AND2_X1 U11011 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9818), .ZN(P1_U3303) );
  INV_X1 U11012 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10243) );
  NOR2_X1 U11013 ( .A1(n9819), .A2(n10243), .ZN(P1_U3304) );
  AND2_X1 U11014 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9818), .ZN(P1_U3305) );
  AND2_X1 U11015 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9818), .ZN(P1_U3306) );
  INV_X1 U11016 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U11017 ( .A1(n9819), .A2(n10225), .ZN(P1_U3307) );
  AND2_X1 U11018 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9818), .ZN(P1_U3308) );
  AND2_X1 U11019 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9818), .ZN(P1_U3309) );
  AND2_X1 U11020 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9818), .ZN(P1_U3310) );
  INV_X1 U11021 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U11022 ( .A1(n9819), .A2(n10081), .ZN(P1_U3311) );
  INV_X1 U11023 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10241) );
  NOR2_X1 U11024 ( .A1(n9819), .A2(n10241), .ZN(P1_U3312) );
  AND2_X1 U11025 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9818), .ZN(P1_U3313) );
  INV_X1 U11026 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10197) );
  NOR2_X1 U11027 ( .A1(n9819), .A2(n10197), .ZN(P1_U3314) );
  INV_X1 U11028 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10176) );
  NOR2_X1 U11029 ( .A1(n9819), .A2(n10176), .ZN(P1_U3315) );
  AND2_X1 U11030 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9818), .ZN(P1_U3316) );
  AND2_X1 U11031 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9818), .ZN(P1_U3317) );
  INV_X1 U11032 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U11033 ( .A1(n9819), .A2(n10240), .ZN(P1_U3318) );
  AND2_X1 U11034 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9818), .ZN(P1_U3319) );
  AND2_X1 U11035 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9818), .ZN(P1_U3320) );
  INV_X1 U11036 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U11037 ( .A1(n9819), .A2(n10119), .ZN(P1_U3321) );
  INV_X1 U11038 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U11039 ( .A1(n9819), .A2(n10253), .ZN(P1_U3322) );
  INV_X1 U11040 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U11041 ( .A1(n9819), .A2(n10150), .ZN(P1_U3323) );
  OAI21_X1 U11042 ( .B1(n9821), .B2(n9833), .A(n9820), .ZN(n9823) );
  AOI211_X1 U11043 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9841)
         );
  AOI22_X1 U11044 ( .A1(n9839), .A2(n9841), .B1(n5914), .B2(n9838), .ZN(
        P1_U3477) );
  OAI21_X1 U11045 ( .B1(n9827), .B2(n9833), .A(n9826), .ZN(n9829) );
  AOI211_X1 U11046 ( .C1(n9836), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9842)
         );
  INV_X1 U11047 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U11048 ( .A1(n9839), .A2(n9842), .B1(n9831), .B2(n9838), .ZN(
        P1_U3480) );
  OAI21_X1 U11049 ( .B1(n5954), .B2(n9833), .A(n9832), .ZN(n9835) );
  AOI211_X1 U11050 ( .C1(n9837), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9844)
         );
  AOI22_X1 U11051 ( .A1(n9839), .A2(n9844), .B1(n5948), .B2(n9838), .ZN(
        P1_U3483) );
  AOI22_X1 U11052 ( .A1(n9845), .A2(n9841), .B1(n9840), .B2(n9843), .ZN(
        P1_U3530) );
  AOI22_X1 U11053 ( .A1(n9845), .A2(n9842), .B1(n5926), .B2(n9843), .ZN(
        P1_U3531) );
  AOI22_X1 U11054 ( .A1(n9845), .A2(n9844), .B1(n9234), .B2(n9843), .ZN(
        P1_U3532) );
  AOI22_X1 U11055 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n9881), .B1(n9846), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n9855) );
  INV_X1 U11056 ( .A(n9847), .ZN(n9850) );
  OAI21_X1 U11057 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9853) );
  XNOR2_X1 U11058 ( .A(n9851), .B(P2_IR_REG_0__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U11059 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  OAI211_X1 U11060 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5198), .A(n9855), .B(
        n9854), .ZN(P2_U3182) );
  XNOR2_X1 U11061 ( .A(n9857), .B(n9856), .ZN(n9859) );
  AOI22_X1 U11062 ( .A1(n9883), .A2(n9859), .B1(n9881), .B2(n9858), .ZN(n9864)
         );
  OAI211_X1 U11063 ( .C1(n9862), .C2(n9861), .A(n9860), .B(n9872), .ZN(n9863)
         );
  OAI211_X1 U11064 ( .C1(n10091), .C2(n9887), .A(n9864), .B(n9863), .ZN(n9865)
         );
  INV_X1 U11065 ( .A(n9865), .ZN(n9871) );
  INV_X1 U11066 ( .A(n9866), .ZN(n9869) );
  AND2_X1 U11067 ( .A1(n9867), .A2(n10182), .ZN(n9868) );
  OAI21_X1 U11068 ( .B1(n9869), .B2(n9868), .A(n9893), .ZN(n9870) );
  OAI211_X1 U11069 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6983), .A(n9871), .B(
        n9870), .ZN(P2_U3183) );
  INV_X1 U11070 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9886) );
  OAI21_X1 U11071 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(n9875) );
  OR2_X1 U11072 ( .A1(n9876), .A2(n9875), .ZN(n9885) );
  OAI21_X1 U11073 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9882) );
  AOI22_X1 U11074 ( .A1(n9883), .A2(n9882), .B1(n9881), .B2(n9880), .ZN(n9884)
         );
  OAI211_X1 U11075 ( .C1(n9887), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9888)
         );
  INV_X1 U11076 ( .A(n9888), .ZN(n9895) );
  OAI21_X1 U11077 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9892) );
  NAND2_X1 U11078 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  OAI211_X1 U11079 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5209), .A(n9895), .B(
        n9894), .ZN(P2_U3184) );
  OAI22_X1 U11080 ( .A1(n9923), .A2(n9899), .B1(n5209), .B2(n9898), .ZN(n9911)
         );
  INV_X1 U11081 ( .A(n9900), .ZN(n9905) );
  NOR3_X1 U11082 ( .A1(n9903), .A2(n9902), .A3(n9901), .ZN(n9904) );
  NOR2_X1 U11083 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  OAI222_X1 U11084 ( .A1(n9910), .A2(n5197), .B1(n9909), .B2(n9908), .C1(n9907), .C2(n9906), .ZN(n9924) );
  AOI211_X1 U11085 ( .C1(n9912), .C2(n9926), .A(n9911), .B(n9924), .ZN(n9914)
         );
  AOI22_X1 U11086 ( .A1(n8421), .A2(n9915), .B1(n9914), .B2(n9913), .ZN(
        P2_U3231) );
  INV_X1 U11087 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U11088 ( .A1(n9975), .A2(n9917), .B1(n9916), .B2(n9973), .ZN(
        P2_U3390) );
  INV_X1 U11089 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U11090 ( .A1(n9918), .A2(n9961), .ZN(n9920) );
  AOI211_X1 U11091 ( .C1(n9958), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9976)
         );
  AOI22_X1 U11092 ( .A1(n9975), .A2(n9922), .B1(n9976), .B2(n9973), .ZN(
        P2_U3393) );
  NOR2_X1 U11093 ( .A1(n9923), .A2(n9961), .ZN(n9925) );
  AOI211_X1 U11094 ( .C1(n9966), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9978)
         );
  AOI22_X1 U11095 ( .A1(n9975), .A2(n5207), .B1(n9978), .B2(n9973), .ZN(
        P2_U3396) );
  INV_X1 U11096 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U11097 ( .A1(n9927), .A2(n9961), .ZN(n9929) );
  AOI211_X1 U11098 ( .C1(n9966), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9979)
         );
  AOI22_X1 U11099 ( .A1(n9975), .A2(n9931), .B1(n9979), .B2(n9973), .ZN(
        P2_U3399) );
  INV_X1 U11100 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9937) );
  INV_X1 U11101 ( .A(n9932), .ZN(n9936) );
  OAI21_X1 U11102 ( .B1(n9934), .B2(n9961), .A(n9933), .ZN(n9935) );
  AOI21_X1 U11103 ( .B1(n9936), .B2(n9966), .A(n9935), .ZN(n9980) );
  AOI22_X1 U11104 ( .A1(n9975), .A2(n9937), .B1(n9980), .B2(n9973), .ZN(
        P2_U3402) );
  INV_X1 U11105 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U11106 ( .A1(n9938), .A2(n9961), .ZN(n9940) );
  AOI211_X1 U11107 ( .C1(n9958), .C2(n9941), .A(n9940), .B(n9939), .ZN(n9981)
         );
  AOI22_X1 U11108 ( .A1(n9975), .A2(n10281), .B1(n9981), .B2(n9973), .ZN(
        P2_U3405) );
  OAI22_X1 U11109 ( .A1(n9943), .A2(n9967), .B1(n9942), .B2(n9961), .ZN(n9944)
         );
  NOR2_X1 U11110 ( .A1(n9945), .A2(n9944), .ZN(n9983) );
  AOI22_X1 U11111 ( .A1(n9975), .A2(n5280), .B1(n9983), .B2(n9973), .ZN(
        P2_U3408) );
  OAI22_X1 U11112 ( .A1(n9948), .A2(n9947), .B1(n9946), .B2(n9961), .ZN(n9949)
         );
  NOR2_X1 U11113 ( .A1(n9950), .A2(n9949), .ZN(n9985) );
  AOI22_X1 U11114 ( .A1(n9975), .A2(n5300), .B1(n9985), .B2(n9973), .ZN(
        P2_U3411) );
  OAI22_X1 U11115 ( .A1(n9952), .A2(n9967), .B1(n9951), .B2(n9961), .ZN(n9953)
         );
  NOR2_X1 U11116 ( .A1(n9954), .A2(n9953), .ZN(n9987) );
  AOI22_X1 U11117 ( .A1(n9975), .A2(n5316), .B1(n9987), .B2(n9973), .ZN(
        P2_U3414) );
  INV_X1 U11118 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U11119 ( .A1(n9955), .A2(n9961), .ZN(n9957) );
  AOI211_X1 U11120 ( .C1(n9959), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9988)
         );
  AOI22_X1 U11121 ( .A1(n9975), .A2(n9960), .B1(n9988), .B2(n9973), .ZN(
        P2_U3417) );
  INV_X1 U11122 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10290) );
  NOR2_X1 U11123 ( .A1(n9962), .A2(n9961), .ZN(n9964) );
  AOI211_X1 U11124 ( .C1(n9966), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9989)
         );
  AOI22_X1 U11125 ( .A1(n9975), .A2(n10290), .B1(n9989), .B2(n9973), .ZN(
        P2_U3420) );
  INV_X1 U11126 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U11127 ( .A1(n9968), .A2(n9967), .ZN(n9970) );
  AOI211_X1 U11128 ( .C1(n9972), .C2(n9971), .A(n9970), .B(n9969), .ZN(n9991)
         );
  AOI22_X1 U11129 ( .A1(n9975), .A2(n9974), .B1(n9991), .B2(n9973), .ZN(
        P2_U3423) );
  AOI22_X1 U11130 ( .A1(n9992), .A2(n9976), .B1(n10182), .B2(n9990), .ZN(
        P2_U3460) );
  AOI22_X1 U11131 ( .A1(n9992), .A2(n9978), .B1(n9977), .B2(n9990), .ZN(
        P2_U3461) );
  AOI22_X1 U11132 ( .A1(n9992), .A2(n9979), .B1(n6224), .B2(n9990), .ZN(
        P2_U3462) );
  AOI22_X1 U11133 ( .A1(n9992), .A2(n9980), .B1(n6248), .B2(n9990), .ZN(
        P2_U3463) );
  AOI22_X1 U11134 ( .A1(n9992), .A2(n9981), .B1(n5263), .B2(n9990), .ZN(
        P2_U3464) );
  AOI22_X1 U11135 ( .A1(n9992), .A2(n9983), .B1(n9982), .B2(n9990), .ZN(
        P2_U3465) );
  AOI22_X1 U11136 ( .A1(n9992), .A2(n9985), .B1(n9984), .B2(n9990), .ZN(
        P2_U3466) );
  AOI22_X1 U11137 ( .A1(n9992), .A2(n9987), .B1(n9986), .B2(n9990), .ZN(
        P2_U3467) );
  AOI22_X1 U11138 ( .A1(n9992), .A2(n9988), .B1(n5342), .B2(n9990), .ZN(
        P2_U3468) );
  AOI22_X1 U11139 ( .A1(n9992), .A2(n9989), .B1(n5361), .B2(n9990), .ZN(
        P2_U3469) );
  AOI22_X1 U11140 ( .A1(n9992), .A2(n9991), .B1(n5381), .B2(n9990), .ZN(
        P2_U3470) );
  OAI222_X1 U11141 ( .A1(n10091), .A2(n9996), .B1(n10091), .B2(n9995), .C1(
        n9994), .C2(n9993), .ZN(ADD_1068_U5) );
  XOR2_X1 U11142 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11143 ( .A(n9999), .ZN(n9998) );
  OAI222_X1 U11144 ( .A1(n10292), .A2(n10000), .B1(n10292), .B2(n9999), .C1(
        n9998), .C2(n9997), .ZN(ADD_1068_U55) );
  OAI21_X1 U11145 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(ADD_1068_U56) );
  OAI21_X1 U11146 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(ADD_1068_U57) );
  OAI21_X1 U11147 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(ADD_1068_U58) );
  OAI21_X1 U11148 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(ADD_1068_U59) );
  OAI21_X1 U11149 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(ADD_1068_U60) );
  OAI21_X1 U11150 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(ADD_1068_U61) );
  OAI21_X1 U11151 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1068_U62) );
  OAI21_X1 U11152 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1068_U63) );
  NOR2_X1 U11153 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .ZN(
        n10026) );
  NOR4_X1 U11154 ( .A1(SI_11_), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(
        P2_REG1_REG_21__SCAN_IN), .A4(P2_ADDR_REG_13__SCAN_IN), .ZN(n10025) );
  NAND4_X1 U11155 ( .A1(n10026), .A2(n10025), .A3(n10284), .A4(n10125), .ZN(
        n10034) );
  NAND4_X1 U11156 ( .A1(n10120), .A2(n10223), .A3(n5961), .A4(n5884), .ZN(
        n10033) );
  NAND4_X1 U11157 ( .A1(n10161), .A2(n10099), .A3(n10098), .A4(n10123), .ZN(
        n10032) );
  NOR4_X1 U11158 ( .A1(P1_D_REG_27__SCAN_IN), .A2(SI_13_), .A3(
        P1_REG3_REG_21__SCAN_IN), .A4(P1_REG3_REG_10__SCAN_IN), .ZN(n10030) );
  NOR4_X1 U11159 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_31__SCAN_IN), .A4(n6016), .ZN(n10029) );
  NOR4_X1 U11160 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(P2_REG1_REG_11__SCAN_IN), .A4(P2_REG1_REG_0__SCAN_IN), .ZN(n10028)
         );
  NOR4_X1 U11161 ( .A1(SI_16_), .A2(P2_REG3_REG_10__SCAN_IN), .A3(
        P2_IR_REG_4__SCAN_IN), .A4(P2_REG0_REG_5__SCAN_IN), .ZN(n10027) );
  NAND4_X1 U11162 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n10031) );
  NOR4_X1 U11163 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10074) );
  NAND4_X1 U11164 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(P2_IR_REG_17__SCAN_IN), .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n10038)
         );
  NAND4_X1 U11165 ( .A1(P1_D_REG_13__SCAN_IN), .A2(SI_23_), .A3(
        P2_DATAO_REG_10__SCAN_IN), .A4(P2_REG2_REG_10__SCAN_IN), .ZN(n10037)
         );
  NAND4_X1 U11166 ( .A1(SI_24_), .A2(P1_REG3_REG_26__SCAN_IN), .A3(
        P1_REG3_REG_11__SCAN_IN), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n10036) );
  NAND4_X1 U11167 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), 
        .A3(P2_REG2_REG_19__SCAN_IN), .A4(P2_REG0_REG_10__SCAN_IN), .ZN(n10035) );
  NOR4_X1 U11168 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10073) );
  NAND4_X1 U11169 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .A3(P2_IR_REG_19__SCAN_IN), .A4(P2_IR_REG_22__SCAN_IN), .ZN(n10042) );
  NAND4_X1 U11170 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(P2_DATAO_REG_31__SCAN_IN), .ZN(n10041) );
  NAND4_X1 U11171 ( .A1(SI_20_), .A2(P2_DATAO_REG_16__SCAN_IN), .A3(
        P1_REG0_REG_19__SCAN_IN), .A4(P1_ADDR_REG_17__SCAN_IN), .ZN(n10040) );
  NAND4_X1 U11172 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(P1_DATAO_REG_0__SCAN_IN), .A3(P1_REG0_REG_12__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n10039) );
  NOR4_X1 U11173 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10072) );
  INV_X1 U11174 ( .A(n10043), .ZN(n10059) );
  NOR4_X1 U11175 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .A3(P1_ADDR_REG_6__SCAN_IN), .A4(n10122), .ZN(n10044) );
  NAND4_X1 U11176 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10045), .A3(n10044), 
        .A4(n10105), .ZN(n10058) );
  NOR3_X1 U11177 ( .A1(n10046), .A2(n6180), .A3(n6007), .ZN(n10048) );
  NAND3_X1 U11178 ( .A1(n10048), .A2(P1_IR_REG_11__SCAN_IN), .A3(n10047), .ZN(
        n10049) );
  NOR3_X1 U11179 ( .A1(n10049), .A2(P1_REG1_REG_13__SCAN_IN), .A3(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n10056) );
  INV_X1 U11180 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10050) );
  NOR4_X1 U11181 ( .A1(n10050), .A2(n10285), .A3(P1_IR_REG_6__SCAN_IN), .A4(
        P1_IR_REG_23__SCAN_IN), .ZN(n10055) );
  NOR4_X1 U11182 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(
        P1_REG2_REG_7__SCAN_IN), .ZN(n10054) );
  NAND3_X1 U11183 ( .A1(n10056), .A2(n10055), .A3(n10054), .ZN(n10057) );
  OR4_X1 U11184 ( .A1(n10059), .A2(n10058), .A3(n10307), .A4(n10057), .ZN(
        n10070) );
  NAND4_X1 U11185 ( .A1(SI_27_), .A2(P2_IR_REG_14__SCAN_IN), .A3(
        P2_IR_REG_5__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n10069) );
  NAND4_X1 U11186 ( .A1(P1_D_REG_0__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P1_DATAO_REG_29__SCAN_IN), .A4(P2_REG2_REG_11__SCAN_IN), .ZN(
        n10068) );
  NOR4_X1 U11187 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P2_REG0_REG_15__SCAN_IN), .A4(n10079), .ZN(n10066) );
  NOR4_X1 U11188 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_IR_REG_30__SCAN_IN), .A3(
        P2_REG1_REG_14__SCAN_IN), .A4(SI_30_), .ZN(n10065) );
  NAND4_X1 U11189 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(SI_2_), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_IR_REG_27__SCAN_IN), .ZN(n10063) );
  NAND4_X1 U11190 ( .A1(P1_D_REG_4__SCAN_IN), .A2(SI_8_), .A3(
        P2_REG3_REG_28__SCAN_IN), .A4(P2_REG0_REG_28__SCAN_IN), .ZN(n10062) );
  NAND4_X1 U11191 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_DATAO_REG_7__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(P1_ADDR_REG_11__SCAN_IN), .ZN(n10061)
         );
  NAND4_X1 U11192 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .A3(P2_REG1_REG_5__SCAN_IN), .A4(P2_ADDR_REG_12__SCAN_IN), .ZN(n10060)
         );
  NOR4_X1 U11193 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10064) );
  NAND3_X1 U11194 ( .A1(n10066), .A2(n10065), .A3(n10064), .ZN(n10067) );
  NOR4_X1 U11195 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        n10071) );
  NAND4_X1 U11196 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10337) );
  AOI22_X1 U11197 ( .A1(n5902), .A2(keyinput101), .B1(keyinput18), .B2(n10076), 
        .ZN(n10075) );
  OAI221_X1 U11198 ( .B1(n5902), .B2(keyinput101), .C1(n10076), .C2(keyinput18), .A(n10075), .ZN(n10088) );
  AOI22_X1 U11199 ( .A1(n10079), .A2(keyinput17), .B1(keyinput1), .B2(n10078), 
        .ZN(n10077) );
  OAI221_X1 U11200 ( .B1(n10079), .B2(keyinput17), .C1(n10078), .C2(keyinput1), 
        .A(n10077), .ZN(n10087) );
  AOI22_X1 U11201 ( .A1(n10081), .A2(keyinput100), .B1(keyinput40), .B2(n8443), 
        .ZN(n10080) );
  OAI221_X1 U11202 ( .B1(n10081), .B2(keyinput100), .C1(n8443), .C2(keyinput40), .A(n10080), .ZN(n10086) );
  AOI22_X1 U11203 ( .A1(n10084), .A2(keyinput119), .B1(n10083), .B2(keyinput60), .ZN(n10082) );
  OAI221_X1 U11204 ( .B1(n10084), .B2(keyinput119), .C1(n10083), .C2(
        keyinput60), .A(n10082), .ZN(n10085) );
  NOR4_X1 U11205 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10137) );
  AOI22_X1 U11206 ( .A1(n10091), .A2(keyinput111), .B1(n10090), .B2(
        keyinput104), .ZN(n10089) );
  OAI221_X1 U11207 ( .B1(n10091), .B2(keyinput111), .C1(n10090), .C2(
        keyinput104), .A(n10089), .ZN(n10103) );
  AOI22_X1 U11208 ( .A1(n10094), .A2(keyinput28), .B1(n10093), .B2(keyinput31), 
        .ZN(n10092) );
  OAI221_X1 U11209 ( .B1(n10094), .B2(keyinput28), .C1(n10093), .C2(keyinput31), .A(n10092), .ZN(n10102) );
  AOI22_X1 U11210 ( .A1(n10096), .A2(keyinput41), .B1(n5102), .B2(keyinput105), 
        .ZN(n10095) );
  OAI221_X1 U11211 ( .B1(n10096), .B2(keyinput41), .C1(n5102), .C2(keyinput105), .A(n10095), .ZN(n10101) );
  AOI22_X1 U11212 ( .A1(n10099), .A2(keyinput35), .B1(keyinput14), .B2(n10098), 
        .ZN(n10097) );
  OAI221_X1 U11213 ( .B1(n10099), .B2(keyinput35), .C1(n10098), .C2(keyinput14), .A(n10097), .ZN(n10100) );
  NOR4_X1 U11214 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10136) );
  AOI22_X1 U11215 ( .A1(n10106), .A2(keyinput51), .B1(keyinput94), .B2(n10105), 
        .ZN(n10104) );
  OAI221_X1 U11216 ( .B1(n10106), .B2(keyinput51), .C1(n10105), .C2(keyinput94), .A(n10104), .ZN(n10117) );
  AOI22_X1 U11217 ( .A1(n5272), .A2(keyinput36), .B1(keyinput110), .B2(n10108), 
        .ZN(n10107) );
  OAI221_X1 U11218 ( .B1(n5272), .B2(keyinput36), .C1(n10108), .C2(keyinput110), .A(n10107), .ZN(n10116) );
  AOI22_X1 U11219 ( .A1(n5422), .A2(keyinput45), .B1(keyinput63), .B2(n10110), 
        .ZN(n10109) );
  OAI221_X1 U11220 ( .B1(n5422), .B2(keyinput45), .C1(n10110), .C2(keyinput63), 
        .A(n10109), .ZN(n10115) );
  INV_X1 U11221 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11222 ( .A1(n10113), .A2(keyinput19), .B1(keyinput33), .B2(n10112), 
        .ZN(n10111) );
  OAI221_X1 U11223 ( .B1(n10113), .B2(keyinput19), .C1(n10112), .C2(keyinput33), .A(n10111), .ZN(n10114) );
  NOR4_X1 U11224 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10135) );
  AOI22_X1 U11225 ( .A1(n10120), .A2(keyinput108), .B1(n10119), .B2(keyinput23), .ZN(n10118) );
  OAI221_X1 U11226 ( .B1(n10120), .B2(keyinput108), .C1(n10119), .C2(
        keyinput23), .A(n10118), .ZN(n10133) );
  AOI22_X1 U11227 ( .A1(n10123), .A2(keyinput72), .B1(keyinput15), .B2(n10122), 
        .ZN(n10121) );
  OAI221_X1 U11228 ( .B1(n10123), .B2(keyinput72), .C1(n10122), .C2(keyinput15), .A(n10121), .ZN(n10132) );
  INV_X1 U11229 ( .A(SI_16_), .ZN(n10126) );
  AOI22_X1 U11230 ( .A1(n10126), .A2(keyinput126), .B1(keyinput69), .B2(n10125), .ZN(n10124) );
  OAI221_X1 U11231 ( .B1(n10126), .B2(keyinput126), .C1(n10125), .C2(
        keyinput69), .A(n10124), .ZN(n10131) );
  AOI22_X1 U11232 ( .A1(n10129), .A2(keyinput70), .B1(n10128), .B2(keyinput49), 
        .ZN(n10127) );
  OAI221_X1 U11233 ( .B1(n10129), .B2(keyinput70), .C1(n10128), .C2(keyinput49), .A(n10127), .ZN(n10130) );
  NOR4_X1 U11234 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  NAND4_X1 U11235 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10318) );
  AOI22_X1 U11236 ( .A1(n5894), .A2(keyinput50), .B1(keyinput39), .B2(n10139), 
        .ZN(n10138) );
  OAI221_X1 U11237 ( .B1(n5894), .B2(keyinput50), .C1(n10139), .C2(keyinput39), 
        .A(n10138), .ZN(n10148) );
  AOI22_X1 U11238 ( .A1(n6007), .A2(keyinput118), .B1(keyinput25), .B2(n10141), 
        .ZN(n10140) );
  OAI221_X1 U11239 ( .B1(n6007), .B2(keyinput118), .C1(n10141), .C2(keyinput25), .A(n10140), .ZN(n10147) );
  XOR2_X1 U11240 ( .A(n6236), .B(keyinput79), .Z(n10145) );
  XNOR2_X1 U11241 ( .A(SI_30_), .B(keyinput8), .ZN(n10144) );
  XNOR2_X1 U11242 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput74), .ZN(n10143) );
  XNOR2_X1 U11243 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput16), .ZN(n10142) );
  NAND4_X1 U11244 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10146) );
  NOR3_X1 U11245 ( .A1(n10148), .A2(n10147), .A3(n10146), .ZN(n10191) );
  AOI22_X1 U11246 ( .A1(n10150), .A2(keyinput57), .B1(keyinput71), .B2(n5198), 
        .ZN(n10149) );
  OAI221_X1 U11247 ( .B1(n10150), .B2(keyinput57), .C1(n5198), .C2(keyinput71), 
        .A(n10149), .ZN(n10159) );
  AOI22_X1 U11248 ( .A1(n9481), .A2(keyinput67), .B1(keyinput62), .B2(n10052), 
        .ZN(n10151) );
  OAI221_X1 U11249 ( .B1(n9481), .B2(keyinput67), .C1(n10052), .C2(keyinput62), 
        .A(n10151), .ZN(n10158) );
  XNOR2_X1 U11250 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput123), .ZN(n10154) );
  XNOR2_X1 U11251 ( .A(SI_2_), .B(keyinput13), .ZN(n10153) );
  XNOR2_X1 U11252 ( .A(P2_REG1_REG_14__SCAN_IN), .B(keyinput77), .ZN(n10152)
         );
  NAND3_X1 U11253 ( .A1(n10154), .A2(n10153), .A3(n10152), .ZN(n10157) );
  XNOR2_X1 U11254 ( .A(n10155), .B(keyinput58), .ZN(n10156) );
  NOR4_X1 U11255 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10190) );
  AOI22_X1 U11256 ( .A1(n10161), .A2(keyinput120), .B1(keyinput102), .B2(
        n10051), .ZN(n10160) );
  OAI221_X1 U11257 ( .B1(n10161), .B2(keyinput120), .C1(n10051), .C2(
        keyinput102), .A(n10160), .ZN(n10172) );
  AOI22_X1 U11258 ( .A1(n10163), .A2(keyinput75), .B1(n5263), .B2(keyinput7), 
        .ZN(n10162) );
  OAI221_X1 U11259 ( .B1(n10163), .B2(keyinput75), .C1(n5263), .C2(keyinput7), 
        .A(n10162), .ZN(n10171) );
  AOI22_X1 U11260 ( .A1(n10166), .A2(keyinput29), .B1(n10165), .B2(keyinput59), 
        .ZN(n10164) );
  OAI221_X1 U11261 ( .B1(n10166), .B2(keyinput29), .C1(n10165), .C2(keyinput59), .A(n10164), .ZN(n10170) );
  XNOR2_X1 U11262 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput81), .ZN(n10168) );
  XNOR2_X1 U11263 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput93), .ZN(n10167)
         );
  NAND2_X1 U11264 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NOR4_X1 U11265 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10189) );
  INV_X1 U11266 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11267 ( .A1(n10175), .A2(keyinput0), .B1(n10174), .B2(keyinput5), 
        .ZN(n10173) );
  OAI221_X1 U11268 ( .B1(n10175), .B2(keyinput0), .C1(n10174), .C2(keyinput5), 
        .A(n10173), .ZN(n10180) );
  XNOR2_X1 U11269 ( .A(n10176), .B(keyinput86), .ZN(n10179) );
  XNOR2_X1 U11270 ( .A(n10177), .B(keyinput98), .ZN(n10178) );
  OR3_X1 U11271 ( .A1(n10180), .A2(n10179), .A3(n10178), .ZN(n10187) );
  AOI22_X1 U11272 ( .A1(n10182), .A2(keyinput106), .B1(n5914), .B2(keyinput52), 
        .ZN(n10181) );
  OAI221_X1 U11273 ( .B1(n10182), .B2(keyinput106), .C1(n5914), .C2(keyinput52), .A(n10181), .ZN(n10186) );
  AOI22_X1 U11274 ( .A1(n5381), .A2(keyinput122), .B1(n10184), .B2(keyinput95), 
        .ZN(n10183) );
  OAI221_X1 U11275 ( .B1(n5381), .B2(keyinput122), .C1(n10184), .C2(keyinput95), .A(n10183), .ZN(n10185) );
  NOR3_X1 U11276 ( .A1(n10187), .A2(n10186), .A3(n10185), .ZN(n10188) );
  NAND4_X1 U11277 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10317) );
  INV_X1 U11278 ( .A(P2_B_REG_SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11279 ( .A1(n5300), .A2(keyinput112), .B1(n10193), .B2(keyinput22), 
        .ZN(n10192) );
  OAI221_X1 U11280 ( .B1(n5300), .B2(keyinput112), .C1(n10193), .C2(keyinput22), .A(n10192), .ZN(n10204) );
  AOI22_X1 U11281 ( .A1(n6183), .A2(keyinput80), .B1(keyinput11), .B2(n10195), 
        .ZN(n10194) );
  OAI221_X1 U11282 ( .B1(n6183), .B2(keyinput80), .C1(n10195), .C2(keyinput11), 
        .A(n10194), .ZN(n10203) );
  AOI22_X1 U11283 ( .A1(n6016), .A2(keyinput121), .B1(n10197), .B2(keyinput66), 
        .ZN(n10196) );
  OAI221_X1 U11284 ( .B1(n6016), .B2(keyinput121), .C1(n10197), .C2(keyinput66), .A(n10196), .ZN(n10202) );
  AOI22_X1 U11285 ( .A1(n10200), .A2(keyinput68), .B1(keyinput88), .B2(n10199), 
        .ZN(n10198) );
  OAI221_X1 U11286 ( .B1(n10200), .B2(keyinput68), .C1(n10199), .C2(keyinput88), .A(n10198), .ZN(n10201) );
  NOR4_X1 U11287 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        n10251) );
  AOI22_X1 U11288 ( .A1(n10207), .A2(keyinput82), .B1(n10206), .B2(keyinput26), 
        .ZN(n10205) );
  OAI221_X1 U11289 ( .B1(n10207), .B2(keyinput82), .C1(n10206), .C2(keyinput26), .A(n10205), .ZN(n10218) );
  INV_X1 U11290 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U11291 ( .A1(n10210), .A2(keyinput99), .B1(keyinput9), .B2(n10209), 
        .ZN(n10208) );
  OAI221_X1 U11292 ( .B1(n10210), .B2(keyinput99), .C1(n10209), .C2(keyinput9), 
        .A(n10208), .ZN(n10217) );
  AOI22_X1 U11293 ( .A1(n10212), .A2(keyinput46), .B1(n10047), .B2(keyinput84), 
        .ZN(n10211) );
  OAI221_X1 U11294 ( .B1(n10212), .B2(keyinput46), .C1(n10047), .C2(keyinput84), .A(n10211), .ZN(n10216) );
  XNOR2_X1 U11295 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput30), .ZN(n10214) );
  XNOR2_X1 U11296 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput42), .ZN(n10213)
         );
  NAND2_X1 U11297 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  NOR4_X1 U11298 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10250) );
  AOI22_X1 U11299 ( .A1(n10220), .A2(keyinput91), .B1(keyinput47), .B2(n5961), 
        .ZN(n10219) );
  OAI221_X1 U11300 ( .B1(n10220), .B2(keyinput91), .C1(n5961), .C2(keyinput47), 
        .A(n10219), .ZN(n10233) );
  AOI22_X1 U11301 ( .A1(n10223), .A2(keyinput78), .B1(n10222), .B2(keyinput3), 
        .ZN(n10221) );
  OAI221_X1 U11302 ( .B1(n10223), .B2(keyinput78), .C1(n10222), .C2(keyinput3), 
        .A(n10221), .ZN(n10232) );
  AOI22_X1 U11303 ( .A1(n10226), .A2(keyinput90), .B1(n10225), .B2(keyinput87), 
        .ZN(n10224) );
  OAI221_X1 U11304 ( .B1(n10226), .B2(keyinput90), .C1(n10225), .C2(keyinput87), .A(n10224), .ZN(n10231) );
  INV_X1 U11305 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U11306 ( .A1(n10229), .A2(keyinput37), .B1(n10228), .B2(keyinput53), 
        .ZN(n10227) );
  OAI221_X1 U11307 ( .B1(n10229), .B2(keyinput37), .C1(n10228), .C2(keyinput53), .A(n10227), .ZN(n10230) );
  NOR4_X1 U11308 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10249) );
  AOI22_X1 U11309 ( .A1(n10236), .A2(keyinput61), .B1(n10235), .B2(keyinput24), 
        .ZN(n10234) );
  OAI221_X1 U11310 ( .B1(n10236), .B2(keyinput61), .C1(n10235), .C2(keyinput24), .A(n10234), .ZN(n10247) );
  AOI22_X1 U11311 ( .A1(n5673), .A2(keyinput92), .B1(keyinput73), .B2(n10238), 
        .ZN(n10237) );
  OAI221_X1 U11312 ( .B1(n5673), .B2(keyinput92), .C1(n10238), .C2(keyinput73), 
        .A(n10237), .ZN(n10246) );
  AOI22_X1 U11313 ( .A1(n10241), .A2(keyinput27), .B1(n10240), .B2(keyinput4), 
        .ZN(n10239) );
  OAI221_X1 U11314 ( .B1(n10241), .B2(keyinput27), .C1(n10240), .C2(keyinput4), 
        .A(n10239), .ZN(n10245) );
  AOI22_X1 U11315 ( .A1(n10243), .A2(keyinput10), .B1(keyinput96), .B2(n5884), 
        .ZN(n10242) );
  OAI221_X1 U11316 ( .B1(n10243), .B2(keyinput10), .C1(n5884), .C2(keyinput96), 
        .A(n10242), .ZN(n10244) );
  NOR4_X1 U11317 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  NAND4_X1 U11318 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10316) );
  AOI22_X1 U11319 ( .A1(n10254), .A2(keyinput89), .B1(n10253), .B2(keyinput115), .ZN(n10252) );
  OAI221_X1 U11320 ( .B1(n10254), .B2(keyinput89), .C1(n10253), .C2(
        keyinput115), .A(n10252), .ZN(n10264) );
  AOI22_X1 U11321 ( .A1(n6180), .A2(keyinput12), .B1(keyinput48), .B2(n5078), 
        .ZN(n10255) );
  OAI221_X1 U11322 ( .B1(n6180), .B2(keyinput12), .C1(n5078), .C2(keyinput48), 
        .A(n10255), .ZN(n10263) );
  AOI22_X1 U11323 ( .A1(n10258), .A2(keyinput114), .B1(keyinput55), .B2(n10257), .ZN(n10256) );
  OAI221_X1 U11324 ( .B1(n10258), .B2(keyinput114), .C1(n10257), .C2(
        keyinput55), .A(n10256), .ZN(n10262) );
  XOR2_X1 U11325 ( .A(n5364), .B(keyinput127), .Z(n10260) );
  XNOR2_X1 U11326 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput56), .ZN(n10259) );
  NAND2_X1 U11327 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  NOR4_X1 U11328 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10314) );
  AOI22_X1 U11329 ( .A1(n10267), .A2(keyinput124), .B1(keyinput76), .B2(n10266), .ZN(n10265) );
  OAI221_X1 U11330 ( .B1(n10267), .B2(keyinput124), .C1(n10266), .C2(
        keyinput76), .A(n10265), .ZN(n10279) );
  INV_X1 U11331 ( .A(SI_11_), .ZN(n10270) );
  AOI22_X1 U11332 ( .A1(n10270), .A2(keyinput97), .B1(keyinput20), .B2(n10269), 
        .ZN(n10268) );
  OAI221_X1 U11333 ( .B1(n10270), .B2(keyinput97), .C1(n10269), .C2(keyinput20), .A(n10268), .ZN(n10278) );
  INV_X1 U11334 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U11335 ( .A1(n10273), .A2(keyinput64), .B1(n10272), .B2(keyinput43), 
        .ZN(n10271) );
  OAI221_X1 U11336 ( .B1(n10273), .B2(keyinput64), .C1(n10272), .C2(keyinput43), .A(n10271), .ZN(n10277) );
  XNOR2_X1 U11337 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput34), .ZN(n10275) );
  XNOR2_X1 U11338 ( .A(keyinput65), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10274)
         );
  NAND2_X1 U11339 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NOR4_X1 U11340 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10313) );
  AOI22_X1 U11341 ( .A1(n8339), .A2(keyinput113), .B1(keyinput2), .B2(n10281), 
        .ZN(n10280) );
  OAI221_X1 U11342 ( .B1(n8339), .B2(keyinput113), .C1(n10281), .C2(keyinput2), 
        .A(n10280), .ZN(n10288) );
  AOI22_X1 U11343 ( .A1(n10284), .A2(keyinput21), .B1(n10283), .B2(keyinput125), .ZN(n10282) );
  OAI221_X1 U11344 ( .B1(n10284), .B2(keyinput21), .C1(n10283), .C2(
        keyinput125), .A(n10282), .ZN(n10287) );
  XNOR2_X1 U11345 ( .A(n10285), .B(keyinput32), .ZN(n10286) );
  OR3_X1 U11346 ( .A1(n10288), .A2(n10287), .A3(n10286), .ZN(n10295) );
  INV_X1 U11347 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U11348 ( .A1(n10291), .A2(keyinput54), .B1(keyinput103), .B2(n10290), .ZN(n10289) );
  OAI221_X1 U11349 ( .B1(n10291), .B2(keyinput54), .C1(n10290), .C2(
        keyinput103), .A(n10289), .ZN(n10294) );
  XNOR2_X1 U11350 ( .A(n10292), .B(keyinput44), .ZN(n10293) );
  NOR3_X1 U11351 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(n10312) );
  XOR2_X1 U11352 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput116), .Z(n10299) );
  XNOR2_X1 U11353 ( .A(n10296), .B(keyinput38), .ZN(n10298) );
  XNOR2_X1 U11354 ( .A(keyinput83), .B(n5959), .ZN(n10297) );
  NOR3_X1 U11355 ( .A1(n10299), .A2(n10298), .A3(n10297), .ZN(n10303) );
  XOR2_X1 U11356 ( .A(n10300), .B(keyinput6), .Z(n10302) );
  XNOR2_X1 U11357 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput85), .ZN(n10301) );
  NAND3_X1 U11358 ( .A1(n10303), .A2(n10302), .A3(n10301), .ZN(n10310) );
  AOI22_X1 U11359 ( .A1(n10306), .A2(keyinput107), .B1(keyinput109), .B2(
        n10305), .ZN(n10304) );
  OAI221_X1 U11360 ( .B1(n10306), .B2(keyinput107), .C1(n10305), .C2(
        keyinput109), .A(n10304), .ZN(n10309) );
  XNOR2_X1 U11361 ( .A(n10307), .B(keyinput117), .ZN(n10308) );
  NOR3_X1 U11362 ( .A1(n10310), .A2(n10309), .A3(n10308), .ZN(n10311) );
  NAND4_X1 U11363 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10315) );
  NOR4_X1 U11364 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10335) );
  AOI211_X1 U11365 ( .C1(n10322), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10327) );
  AOI211_X1 U11366 ( .C1(n10325), .C2(n6016), .A(n10324), .B(n10323), .ZN(
        n10326) );
  AOI211_X1 U11367 ( .C1(n10329), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10331) );
  NAND2_X1 U11368 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10330)
         );
  OAI211_X1 U11369 ( .C1(n10333), .C2(n10332), .A(n10331), .B(n10330), .ZN(
        n10334) );
  XOR2_X1 U11370 ( .A(n10335), .B(n10334), .Z(n10336) );
  XNOR2_X1 U11371 ( .A(n10337), .B(n10336), .ZN(P1_U3258) );
  OAI21_X1 U11372 ( .B1(n10340), .B2(n10339), .A(n10338), .ZN(ADD_1068_U50) );
  OAI21_X1 U11373 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(ADD_1068_U51) );
  OAI21_X1 U11374 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(ADD_1068_U47) );
  OAI21_X1 U11375 ( .B1(n10349), .B2(n10348), .A(n10347), .ZN(ADD_1068_U49) );
  OAI21_X1 U11376 ( .B1(n10352), .B2(n10351), .A(n10350), .ZN(ADD_1068_U48) );
  AOI21_X1 U11377 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(ADD_1068_U54) );
  AOI21_X1 U11378 ( .B1(n10358), .B2(n10357), .A(n10356), .ZN(ADD_1068_U53) );
  OAI21_X1 U11379 ( .B1(n10361), .B2(n10360), .A(n10359), .ZN(ADD_1068_U52) );
  OR2_X1 U6597 ( .A1(n5362), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5378) );
  CLKBUF_X1 U4922 ( .A(n8645), .Z(n8735) );
  CLKBUF_X1 U4979 ( .A(n5857), .Z(n9000) );
  CLKBUF_X1 U4982 ( .A(n5837), .Z(n5979) );
  CLKBUF_X1 U5179 ( .A(n6926), .Z(n4418) );
endmodule

