

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273;

  INV_X2 U4881 ( .A(n9692), .ZN(n4381) );
  OR2_X1 U4882 ( .A1(n9220), .A2(n9146), .ZN(n4562) );
  INV_X4 U4883 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4884 ( .A(n4379), .ZN(n4380) );
  BUF_X2 U4885 ( .A(n4382), .Z(n4403) );
  INV_X1 U4886 ( .A(n5080), .ZN(n5114) );
  INV_X2 U4887 ( .A(n5686), .ZN(n5581) );
  OAI21_X1 U4888 ( .B1(n4830), .B2(n4829), .A(n4827), .ZN(n5218) );
  CLKBUF_X1 U4889 ( .A(n8727), .Z(n4410) );
  AND4_X1 U4890 ( .A1(n5919), .A2(n5757), .A3(n5756), .A4(n5945), .ZN(n4414)
         );
  INV_X1 U4891 ( .A(n5992), .ZN(n4382) );
  INV_X1 U4893 ( .A(n5874), .ZN(n5992) );
  OAI211_X1 U4894 ( .C1(n4399), .C2(n6843), .A(n5862), .B(n5861), .ZN(n7298)
         );
  INV_X1 U4896 ( .A(n6529), .ZN(n6979) );
  AND3_X1 U4898 ( .A1(n5850), .A2(n5849), .A3(n5848), .ZN(n7294) );
  AND3_X1 U4899 ( .A1(n5825), .A2(n5824), .A3(n5823), .ZN(n7224) );
  AND2_X1 U4900 ( .A1(n8969), .A2(n5637), .ZN(n8971) );
  INV_X1 U4901 ( .A(n7994), .ZN(n6388) );
  INV_X2 U4902 ( .A(n6362), .ZN(n7169) );
  NOR2_X1 U4903 ( .A1(n7110), .A2(n7988), .ZN(n9678) );
  INV_X1 U4904 ( .A(n8094), .ZN(n9736) );
  INV_X1 U4905 ( .A(n7160), .ZN(n9709) );
  OAI21_X1 U4906 ( .B1(n5264), .B2(n4863), .A(n4861), .ZN(n5311) );
  INV_X1 U4907 ( .A(n8727), .ZN(n4625) );
  OAI211_X1 U4908 ( .C1(n5294), .C2(n6714), .A(n5135), .B(n5134), .ZN(n7160)
         );
  NAND2_X1 U4909 ( .A1(n5442), .A2(n5441), .ZN(n7905) );
  INV_X1 U4910 ( .A(n9376), .ZN(n5726) );
  INV_X1 U4911 ( .A(n7995), .ZN(n5690) );
  NAND4_X1 U4912 ( .A1(n5006), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(n7117)
         );
  AOI21_X1 U4913 ( .B1(n7467), .B2(n7466), .A(n4433), .ZN(n7469) );
  NAND2_X1 U4914 ( .A1(n5097), .A2(n5096), .ZN(n7122) );
  AOI211_X1 U4916 ( .C1(n8407), .C2(n8406), .A(n8478), .B(n8405), .ZN(n8411)
         );
  INV_X1 U4918 ( .A(n4391), .ZN(n7935) );
  XNOR2_X1 U4919 ( .A(n5073), .B(n5071), .ZN(n5728) );
  AND2_X1 U4920 ( .A1(n4930), .A2(n4931), .ZN(n4376) );
  INV_X2 U4921 ( .A(n5093), .ZN(n6628) );
  INV_X1 U4922 ( .A(n6538), .ZN(n4379) );
  AND3_X2 U4924 ( .A1(n5020), .A2(n5023), .A3(n4924), .ZN(n5368) );
  INV_X1 U4925 ( .A(n6628), .ZN(n4377) );
  NAND2_X2 U4926 ( .A1(n4883), .A2(n4882), .ZN(n5093) );
  INV_X1 U4927 ( .A(n4377), .ZN(n4397) );
  XNOR2_X1 U4928 ( .A(n5065), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5747) );
  OAI222_X1 U4929 ( .A1(n9479), .A2(n7936), .B1(P1_U3084), .B2(n5038), .C1(
        n8002), .C2(n7945), .ZN(P1_U3324) );
  INV_X1 U4930 ( .A(n5038), .ZN(n5036) );
  INV_X1 U4931 ( .A(n5724), .ZN(n5049) );
  AND2_X1 U4932 ( .A1(n9214), .A2(n9202), .ZN(n9196) );
  NAND2_X1 U4933 ( .A1(n7729), .A2(n4922), .ZN(n9511) );
  NAND2_X2 U4934 ( .A1(n7068), .A2(n6208), .ZN(n7021) );
  AOI22_X1 U4935 ( .A1(n9055), .A2(n5098), .B1(n7122), .B2(n6359), .ZN(n5100)
         );
  BUF_X2 U4936 ( .A(n6415), .Z(n4401) );
  AND2_X1 U4937 ( .A1(n4394), .A2(n4377), .ZN(n5874) );
  INV_X2 U4938 ( .A(n6135), .ZN(n6147) );
  NAND2_X2 U4939 ( .A1(n5049), .A2(n5728), .ZN(n5080) );
  NAND2_X1 U4940 ( .A1(n4392), .A2(n5786), .ZN(n4987) );
  INV_X1 U4941 ( .A(n5784), .ZN(n5786) );
  NOR2_X2 U4942 ( .A1(n6191), .A2(n6401), .ZN(n6399) );
  NAND2_X2 U4943 ( .A1(n5747), .A2(n9603), .ZN(n5294) );
  XNOR2_X1 U4944 ( .A(n5200), .B(SI_5_), .ZN(n5198) );
  XNOR2_X1 U4945 ( .A(n6336), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U4946 ( .A1(n5033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5066) );
  NOR2_X1 U4947 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5919) );
  AND2_X1 U4948 ( .A1(n4619), .A2(n4618), .ZN(n9383) );
  AND2_X1 U4949 ( .A1(n8600), .A2(n8599), .ZN(n8602) );
  OR2_X1 U4950 ( .A1(n8926), .A2(n5593), .ZN(n8929) );
  OR2_X1 U4951 ( .A1(n9379), .A2(n9753), .ZN(n4619) );
  AOI21_X1 U4952 ( .B1(n9222), .B2(n9161), .A(n9160), .ZN(n9209) );
  INV_X1 U4953 ( .A(n9387), .ZN(n4734) );
  AOI211_X1 U4954 ( .C1(n4625), .C2(n8764), .A(n9808), .B(n8763), .ZN(n8765)
         );
  INV_X1 U4955 ( .A(n8176), .ZN(n4517) );
  NAND2_X1 U4956 ( .A1(n7993), .A2(n7992), .ZN(n9558) );
  AND2_X1 U4957 ( .A1(n4756), .A2(n6054), .ZN(n4755) );
  AOI21_X1 U4958 ( .B1(n4932), .B2(n4940), .A(n4453), .ZN(n4931) );
  NAND2_X1 U4959 ( .A1(n7646), .A2(n6479), .ZN(n7650) );
  OR2_X1 U4960 ( .A1(n9528), .A2(n4740), .ZN(n4736) );
  NAND2_X1 U4961 ( .A1(n5605), .A2(n5604), .ZN(n9412) );
  NAND2_X1 U4962 ( .A1(n6044), .A2(n6043), .ZN(n8827) );
  XNOR2_X1 U4963 ( .A(n5603), .B(n5602), .ZN(n7721) );
  NAND2_X1 U4964 ( .A1(n6032), .A2(n6031), .ZN(n8832) );
  NAND2_X1 U4965 ( .A1(n5553), .A2(n5552), .ZN(n9422) );
  OR2_X1 U4966 ( .A1(n4796), .A2(n7909), .ZN(n9349) );
  AOI21_X1 U4967 ( .B1(n4723), .B2(n4413), .A(n8139), .ZN(n4722) );
  NAND2_X1 U4968 ( .A1(n5233), .A2(n5232), .ZN(n7439) );
  NAND2_X1 U4969 ( .A1(n8137), .A2(n8069), .ZN(n8135) );
  NAND2_X1 U4970 ( .A1(n9747), .A2(n7364), .ZN(n7394) );
  NAND2_X1 U4971 ( .A1(n5973), .A2(n5972), .ZN(n8861) );
  OR2_X1 U4972 ( .A1(n7270), .A2(n8018), .ZN(n9747) );
  XNOR2_X1 U4973 ( .A(n5454), .B(n5453), .ZN(n7081) );
  OAI21_X1 U4974 ( .B1(n9660), .B2(n9671), .A(n7165), .ZN(n7168) );
  AND2_X1 U4975 ( .A1(n8097), .A2(n8100), .ZN(n8101) );
  XNOR2_X1 U4976 ( .A(n5199), .B(n5198), .ZN(n6638) );
  XNOR2_X1 U4977 ( .A(n5218), .B(n5217), .ZN(n6641) );
  XNOR2_X1 U4978 ( .A(n6415), .B(n9851), .ZN(n6410) );
  NAND4_X2 U4979 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n9053)
         );
  AND3_X2 U4980 ( .A1(n5814), .A2(n5813), .A3(n5812), .ZN(n9851) );
  AND3_X1 U4981 ( .A1(n5795), .A2(n5796), .A3(n5797), .ZN(n4805) );
  INV_X2 U4982 ( .A(n6061), .ZN(n6153) );
  INV_X1 U4983 ( .A(n6421), .ZN(n6415) );
  OAI211_X1 U4984 ( .C1(n5294), .C2(n9587), .A(n5109), .B(n5108), .ZN(n7988)
         );
  NAND2_X1 U4985 ( .A1(n6402), .A2(n7027), .ZN(n6421) );
  INV_X1 U4986 ( .A(n5828), .ZN(n6061) );
  AOI21_X1 U4987 ( .B1(n5198), .B2(n4828), .A(n4459), .ZN(n4827) );
  BUF_X4 U4988 ( .A(n5995), .Z(n6093) );
  NAND2_X1 U4989 ( .A1(n4880), .A2(n5157), .ZN(n5175) );
  OR2_X1 U4990 ( .A1(n5173), .A2(n6630), .ZN(n5109) );
  INV_X2 U4991 ( .A(n4987), .ZN(n6079) );
  INV_X2 U4992 ( .A(n4404), .ZN(n4405) );
  AND2_X1 U4993 ( .A1(n4393), .A2(n4397), .ZN(n5995) );
  INV_X1 U4994 ( .A(n4400), .ZN(n5821) );
  NAND2_X1 U4995 ( .A1(n6191), .A2(n4625), .ZN(n7032) );
  AND2_X2 U4996 ( .A1(n5036), .A2(n9477), .ZN(n7994) );
  NAND2_X1 U4997 ( .A1(n5786), .A2(n7935), .ZN(n4986) );
  INV_X2 U4998 ( .A(n5827), .ZN(n6135) );
  NAND2_X1 U4999 ( .A1(n5792), .A2(n5791), .ZN(n7840) );
  AND2_X1 U5000 ( .A1(n5784), .A2(n5785), .ZN(n5827) );
  MUX2_X1 U5001 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9480), .S(n5294), .Z(n7150) );
  XNOR2_X1 U5002 ( .A(n5782), .B(n5781), .ZN(n5784) );
  MUX2_X1 U5003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5789), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5792) );
  OR2_X1 U5004 ( .A1(n5054), .A2(n4595), .ZN(n5052) );
  OR2_X1 U5005 ( .A1(n8889), .A2(n10207), .ZN(n5782) );
  XNOR2_X1 U5006 ( .A(n5035), .B(n5034), .ZN(n9477) );
  CLKBUF_X1 U5007 ( .A(n6346), .Z(n4389) );
  XNOR2_X1 U5008 ( .A(n5066), .B(n5067), .ZN(n9603) );
  NOR2_X1 U5009 ( .A1(n4426), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U5010 ( .A1(n5066), .A2(n5027), .ZN(n5065) );
  NAND2_X1 U5011 ( .A1(n4678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6336) );
  NAND2_X2 U5012 ( .A1(n4377), .A2(P1_U3084), .ZN(n7945) );
  AND2_X2 U5013 ( .A1(n5970), .A2(n5763), .ZN(n5765) );
  NAND2_X1 U5014 ( .A1(n5060), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U5015 ( .A1(n4799), .A2(n5058), .ZN(n4883) );
  INV_X1 U5016 ( .A(n5171), .ZN(n5020) );
  AND2_X1 U5017 ( .A1(n4419), .A2(n4682), .ZN(n4681) );
  NOR2_X1 U5018 ( .A1(n4615), .A2(n4614), .ZN(n5050) );
  AND2_X1 U5019 ( .A1(n4926), .A2(n4925), .ZN(n4924) );
  NOR2_X1 U5020 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4616) );
  INV_X1 U5021 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5295) );
  INV_X1 U5022 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5071) );
  INV_X1 U5023 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5486) );
  NOR2_X1 U5024 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4617) );
  NOR2_X2 U5025 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5834) );
  INV_X1 U5026 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5762) );
  INV_X1 U5027 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5857) );
  INV_X1 U5028 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5051) );
  INV_X1 U5029 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5438) );
  INV_X1 U5030 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5945) );
  INV_X1 U5031 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5240) );
  INV_X1 U5032 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5102) );
  INV_X1 U5033 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U5034 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5018) );
  INV_X1 U5035 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5019) );
  INV_X4 U5036 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  XNOR2_X1 U5037 ( .A(n5100), .B(n6362), .ZN(n6928) );
  OAI21_X2 U5038 ( .B1(n9011), .B2(n9013), .A(n9012), .ZN(n8896) );
  NOR3_X2 U5039 ( .A1(n9353), .A2(n4602), .A3(n9427), .ZN(n4601) );
  NAND2_X1 U5040 ( .A1(n7057), .A2(n6423), .ZN(n4383) );
  NAND2_X1 U5041 ( .A1(n7279), .A2(n4387), .ZN(n4384) );
  AND2_X1 U5042 ( .A1(n4384), .A2(n4385), .ZN(n6465) );
  OR2_X1 U5043 ( .A1(n4386), .A2(n4993), .ZN(n4385) );
  INV_X1 U5044 ( .A(n6460), .ZN(n4386) );
  AND2_X1 U5045 ( .A1(n6450), .A2(n6460), .ZN(n4387) );
  AOI22_X1 U5047 ( .A1(n8414), .A2(n8413), .B1(n6528), .B2(n6527), .ZN(n4390)
         );
  XNOR2_X1 U5048 ( .A(n4777), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4391) );
  XNOR2_X1 U5049 ( .A(n4777), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U5050 ( .A1(n7057), .A2(n6423), .ZN(n7082) );
  NAND4_X1 U5051 ( .A1(n5800), .A2(n5802), .A3(n5801), .A4(n5803), .ZN(n6403)
         );
  AOI22_X1 U5052 ( .A1(n8414), .A2(n8413), .B1(n6528), .B2(n6527), .ZN(n8393)
         );
  XNOR2_X1 U5053 ( .A(n4777), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U5054 ( .A1(n7275), .A2(n6443), .ZN(n6448) );
  OAI222_X1 U5055 ( .A1(n7935), .A2(P2_U3152), .B1(n8894), .B2(n7936), .C1(
        n7934), .C2(n8311), .ZN(P2_U3329) );
  AND2_X1 U5056 ( .A1(n5784), .A2(n7935), .ZN(n5815) );
  INV_X4 U5057 ( .A(n5080), .ZN(n6365) );
  NAND2_X1 U5058 ( .A1(n6353), .A2(n7840), .ZN(n4393) );
  NAND2_X1 U5059 ( .A1(n6353), .A2(n7840), .ZN(n4394) );
  INV_X1 U5060 ( .A(n4986), .ZN(n4395) );
  INV_X2 U5061 ( .A(n4986), .ZN(n5828) );
  INV_X1 U5062 ( .A(n4377), .ZN(n4396) );
  INV_X1 U5063 ( .A(n4987), .ZN(n4398) );
  NAND2_X1 U5064 ( .A1(n6353), .A2(n7840), .ZN(n4399) );
  NAND2_X1 U5065 ( .A1(n6353), .A2(n7840), .ZN(n4400) );
  NAND2_X2 U5066 ( .A1(n6477), .A2(n8430), .ZN(n7646) );
  AND2_X4 U5067 ( .A1(n6365), .A2(n5719), .ZN(n5098) );
  NAND2_X2 U5068 ( .A1(n5057), .A2(n5707), .ZN(n5719) );
  NAND2_X1 U5069 ( .A1(n7094), .A2(n6434), .ZN(n7095) );
  NAND2_X1 U5070 ( .A1(n4992), .A2(n7082), .ZN(n7094) );
  NAND2_X2 U5071 ( .A1(n6485), .A2(n6486), .ZN(n8266) );
  NAND2_X2 U5072 ( .A1(n7650), .A2(n6483), .ZN(n6485) );
  AND3_X2 U5073 ( .A1(n5840), .A2(n5839), .A3(n5838), .ZN(n7230) );
  AOI21_X2 U5074 ( .B1(n8335), .B2(n8338), .A(n8333), .ZN(n6525) );
  NAND2_X1 U5075 ( .A1(n7054), .A2(n6414), .ZN(n6420) );
  NAND2_X1 U5076 ( .A1(n5995), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U5077 ( .A1(n5769), .A2(n5768), .ZN(n7526) );
  NAND2_X1 U5078 ( .A1(n5768), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5766) );
  AND2_X1 U5079 ( .A1(n4414), .A2(n4804), .ZN(n5970) );
  NAND2_X1 U5080 ( .A1(n8313), .A2(n8312), .ZN(n7275) );
  NAND2_X1 U5081 ( .A1(n6972), .A2(n4991), .ZN(n7054) );
  NAND2_X1 U5082 ( .A1(n6406), .A2(n6405), .ZN(n6972) );
  NAND2_X1 U5083 ( .A1(n4830), .A2(n5178), .ZN(n5199) );
  NAND2_X1 U5084 ( .A1(n6420), .A2(n7055), .ZN(n7057) );
  AND2_X4 U5085 ( .A1(n5080), .A2(n5719), .ZN(n6359) );
  NAND2_X1 U5086 ( .A1(n7279), .A2(n6450), .ZN(n7317) );
  NAND2_X1 U5087 ( .A1(n6448), .A2(n7276), .ZN(n7279) );
  NAND3_X2 U5088 ( .A1(n8268), .A2(n8267), .A3(n6489), .ZN(n7883) );
  INV_X1 U5089 ( .A(n5173), .ZN(n4404) );
  INV_X2 U5090 ( .A(n6501), .ZN(n8466) );
  NAND2_X2 U5091 ( .A1(n7883), .A2(n6494), .ZN(n8407) );
  AND2_X1 U5092 ( .A1(n5784), .A2(n7935), .ZN(n4407) );
  AND2_X1 U5093 ( .A1(n5784), .A2(n7935), .ZN(n4408) );
  INV_X1 U5094 ( .A(n5974), .ZN(n4409) );
  XNOR2_X1 U5095 ( .A(n5772), .B(n5771), .ZN(n8727) );
  XNOR2_X2 U5096 ( .A(n5766), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6401) );
  INV_X1 U5097 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4925) );
  AOI21_X1 U5098 ( .B1(n4861), .B2(n4863), .A(n4860), .ZN(n4857) );
  INV_X1 U5099 ( .A(n4999), .ZN(n4860) );
  OR2_X1 U5100 ( .A1(n8799), .A2(n8328), .ZN(n6313) );
  NAND2_X1 U5101 ( .A1(n4944), .A2(n4942), .ZN(n4941) );
  INV_X1 U5102 ( .A(n9029), .ZN(n4942) );
  INV_X1 U5103 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5021) );
  AND2_X1 U5104 ( .A1(n6191), .A2(n6401), .ZN(n6765) );
  NOR2_X1 U5105 ( .A1(n4816), .A2(n8804), .ZN(n4814) );
  OR2_X1 U5106 ( .A1(n8794), .A2(n8799), .ZN(n4816) );
  AOI211_X1 U5107 ( .C1(n8106), .C2(n8105), .A(n8104), .B(n8103), .ZN(n8118)
         );
  NAND2_X1 U5108 ( .A1(n6290), .A2(n6324), .ZN(n4664) );
  AND2_X1 U5109 ( .A1(n6294), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5110 ( .A1(n6288), .A2(n6285), .ZN(n4662) );
  AOI21_X1 U5111 ( .B1(n8165), .B2(n8164), .A(n8163), .ZN(n8177) );
  NAND2_X1 U5112 ( .A1(n4520), .A2(n4519), .ZN(n8165) );
  INV_X1 U5113 ( .A(n6151), .ZN(n6152) );
  OAI21_X1 U5114 ( .B1(n8556), .B2(n6156), .A(n6317), .ZN(n6151) );
  AND2_X1 U5115 ( .A1(n6550), .A2(n9810), .ZN(n7025) );
  INV_X1 U5116 ( .A(n5614), .ZN(n5619) );
  AOI21_X1 U5117 ( .B1(n4866), .B2(n5265), .A(n4865), .ZN(n4864) );
  INV_X1 U5118 ( .A(n5005), .ZN(n4865) );
  OAI22_X1 U5119 ( .A1(n4988), .A2(n4987), .B1(n4986), .B2(n7046), .ZN(n4985)
         );
  OAI21_X1 U5120 ( .B1(n8602), .B2(n6105), .A(n6308), .ZN(n8570) );
  OR2_X1 U5121 ( .A1(n8804), .A2(n8604), .ZN(n6308) );
  NAND2_X1 U5122 ( .A1(n8719), .A2(n6022), .ZN(n6023) );
  NOR2_X1 U5123 ( .A1(n8772), .A2(n4742), .ZN(n4741) );
  INV_X1 U5124 ( .A(n6260), .ZN(n4742) );
  OR2_X1 U5125 ( .A1(n8295), .A2(n8471), .ZN(n6266) );
  OR2_X1 U5126 ( .A1(n8818), .A2(n8635), .ZN(n8620) );
  OAI21_X1 U5127 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n6542), .A(n9834), .ZN(n7289)
         );
  INV_X1 U5128 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5787) );
  AND2_X1 U5129 ( .A1(n4681), .A2(n4680), .ZN(n4679) );
  INV_X1 U5130 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4680) );
  NOR2_X1 U5131 ( .A1(n9158), .A2(n4708), .ZN(n4707) );
  INV_X1 U5132 ( .A(n9140), .ZN(n4589) );
  OR2_X1 U5133 ( .A1(n9412), .A2(n9261), .ZN(n9143) );
  NAND2_X1 U5134 ( .A1(n4790), .A2(n4792), .ZN(n4789) );
  NAND2_X1 U5135 ( .A1(n4790), .A2(n4588), .ZN(n4587) );
  NOR2_X1 U5136 ( .A1(n4590), .A2(n9141), .ZN(n4588) );
  AOI21_X1 U5137 ( .B1(n9307), .B2(n4427), .A(n9142), .ZN(n4793) );
  OR2_X1 U5138 ( .A1(n9434), .A2(n9437), .ZN(n4604) );
  NAND2_X1 U5139 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  NOR2_X1 U5140 ( .A1(n4415), .A2(n4577), .ZN(n4572) );
  NOR2_X1 U5141 ( .A1(n8135), .A2(n4439), .ZN(n7909) );
  NAND2_X1 U5142 ( .A1(n7475), .A2(n8044), .ZN(n4699) );
  INV_X1 U5143 ( .A(n7114), .ZN(n6943) );
  XNOR2_X1 U5144 ( .A(n6163), .B(n6161), .ZN(n6160) );
  AND2_X1 U5145 ( .A1(n6088), .A2(n5680), .ZN(n6086) );
  AOI21_X1 U5146 ( .B1(n5674), .B2(n5673), .A(n4839), .ZN(n4838) );
  INV_X1 U5147 ( .A(n5676), .ZN(n4839) );
  NOR2_X1 U5148 ( .A1(n5651), .A2(n5650), .ZN(n5674) );
  AND2_X1 U5149 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  NOR2_X1 U5150 ( .A1(n5647), .A2(n5646), .ZN(n5675) );
  OR2_X1 U5151 ( .A1(n5645), .A2(n5651), .ZN(n5646) );
  AND2_X1 U5152 ( .A1(n5551), .A2(n5537), .ZN(n5549) );
  INV_X1 U5153 ( .A(SI_19_), .ZN(n5509) );
  OAI21_X1 U5154 ( .B1(n5485), .B2(n5484), .A(n5483), .ZN(n5505) );
  NAND2_X1 U5155 ( .A1(n4778), .A2(n4779), .ZN(n5382) );
  INV_X1 U5156 ( .A(n4780), .ZN(n4779) );
  OAI21_X1 U5157 ( .B1(n4785), .B2(n4781), .A(n5361), .ZN(n4780) );
  OAI211_X1 U5158 ( .C1(n4883), .C2(P1_DATAO_REG_8__SCAN_IN), .A(n4801), .B(
        n4800), .ZN(n5254) );
  OR2_X1 U5159 ( .A1(n4882), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U5160 ( .A1(n6015), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5161 ( .A1(n6325), .A2(n6324), .ZN(n4689) );
  AND2_X1 U5162 ( .A1(n6085), .A2(n6084), .ZN(n8400) );
  OR2_X1 U5163 ( .A1(n8804), .A2(n8572), .ZN(n8293) );
  NAND2_X1 U5164 ( .A1(n4770), .A2(n4768), .ZN(n8719) );
  NOR2_X1 U5165 ( .A1(n4771), .A2(n4769), .ZN(n4768) );
  INV_X1 U5166 ( .A(n6273), .ZN(n4769) );
  NAND2_X1 U5167 ( .A1(n8741), .A2(n6272), .ZN(n4770) );
  AND2_X1 U5168 ( .A1(n6765), .A2(n6571), .ZN(n9787) );
  INV_X1 U5169 ( .A(n9535), .ZN(n9785) );
  NAND2_X1 U5170 ( .A1(n7032), .A2(n7031), .ZN(n9790) );
  NAND2_X1 U5171 ( .A1(n6112), .A2(n6111), .ZN(n8799) );
  NAND2_X1 U5172 ( .A1(n5765), .A2(n4681), .ZN(n5768) );
  NAND2_X1 U5173 ( .A1(n4947), .A2(n4939), .ZN(n4938) );
  INV_X1 U5174 ( .A(n4950), .ZN(n4939) );
  AND2_X1 U5175 ( .A1(n4943), .A2(n4941), .ZN(n4940) );
  INV_X1 U5176 ( .A(n4947), .ZN(n4943) );
  NAND2_X1 U5177 ( .A1(n5186), .A2(n5188), .ZN(n4913) );
  NOR2_X1 U5178 ( .A1(n9507), .A2(n4923), .ZN(n4922) );
  INV_X1 U5179 ( .A(n5333), .ZN(n4923) );
  NAND2_X1 U5180 ( .A1(n8004), .A2(n8003), .ZN(n9380) );
  NAND2_X1 U5181 ( .A1(n6586), .A2(n6585), .ZN(n9388) );
  AND2_X1 U5182 ( .A1(n9163), .A2(n9164), .ZN(n9187) );
  NAND2_X1 U5183 ( .A1(n9227), .A2(n4559), .ZN(n4558) );
  AOI21_X1 U5184 ( .B1(n4707), .B2(n4705), .A(n4704), .ZN(n4703) );
  INV_X1 U5185 ( .A(n4710), .ZN(n4705) );
  INV_X1 U5186 ( .A(n9245), .ZN(n9273) );
  INV_X1 U5187 ( .A(n4405), .ZN(n5513) );
  NAND2_X1 U5188 ( .A1(n4607), .A2(n7742), .ZN(n4606) );
  NOR2_X1 U5189 ( .A1(n4608), .A2(n7905), .ZN(n4607) );
  INV_X1 U5190 ( .A(n4724), .ZN(n4723) );
  OAI21_X1 U5191 ( .B1(n7666), .B2(n4413), .A(n8068), .ZN(n4724) );
  INV_X1 U5192 ( .A(n5128), .ZN(n8035) );
  NAND2_X1 U5193 ( .A1(n5294), .A2(n4377), .ZN(n5173) );
  AND2_X1 U5194 ( .A1(n5050), .A2(n4454), .ZN(n5026) );
  NAND2_X1 U5195 ( .A1(n4696), .A2(n4695), .ZN(n4694) );
  INV_X1 U5196 ( .A(n6216), .ZN(n4696) );
  NAND2_X1 U5197 ( .A1(n4499), .A2(n4496), .ZN(n4495) );
  INV_X1 U5198 ( .A(n8131), .ZN(n4493) );
  NAND2_X1 U5199 ( .A1(n8129), .A2(n4490), .ZN(n4489) );
  INV_X1 U5200 ( .A(n8128), .ZN(n4491) );
  INV_X1 U5201 ( .A(n8136), .ZN(n4488) );
  INV_X1 U5202 ( .A(n8135), .ZN(n4487) );
  OAI22_X1 U5203 ( .A1(n7704), .A2(n4667), .B1(n6324), .B2(n6249), .ZN(n4666)
         );
  NOR2_X1 U5204 ( .A1(n4764), .A2(n6316), .ZN(n4667) );
  NOR2_X1 U5205 ( .A1(n7704), .A2(n4669), .ZN(n4668) );
  INV_X1 U5206 ( .A(n6248), .ZN(n4669) );
  NAND2_X1 U5207 ( .A1(n4672), .A2(n6316), .ZN(n4671) );
  INV_X1 U5208 ( .A(n6255), .ZN(n4672) );
  NOR2_X1 U5209 ( .A1(n8145), .A2(n8144), .ZN(n8152) );
  AND2_X1 U5210 ( .A1(n9155), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U5211 ( .A1(n4437), .A2(n9154), .ZN(n4531) );
  AOI21_X1 U5212 ( .B1(n4530), .B2(n8156), .A(n9156), .ZN(n4529) );
  AOI21_X1 U5213 ( .B1(n4529), .B2(n4525), .A(n8188), .ZN(n4524) );
  INV_X1 U5214 ( .A(n4530), .ZN(n4525) );
  NOR2_X1 U5215 ( .A1(n4528), .A2(n4535), .ZN(n4527) );
  NOR2_X1 U5216 ( .A1(n8236), .A2(n4708), .ZN(n4528) );
  NOR2_X1 U5217 ( .A1(n4676), .A2(n8753), .ZN(n4675) );
  INV_X1 U5218 ( .A(n6271), .ZN(n4676) );
  INV_X1 U5219 ( .A(n6274), .ZN(n6281) );
  NAND2_X1 U5220 ( .A1(n4463), .A2(n8180), .ZN(n4516) );
  NAND2_X1 U5221 ( .A1(n4847), .A2(n4843), .ZN(n4842) );
  INV_X1 U5222 ( .A(n6142), .ZN(n4843) );
  INV_X1 U5223 ( .A(n4664), .ZN(n4657) );
  INV_X1 U5224 ( .A(n4661), .ZN(n4660) );
  AOI21_X1 U5225 ( .B1(n4661), .B2(n4659), .A(n6293), .ZN(n4658) );
  NAND2_X1 U5226 ( .A1(n8659), .A2(n4664), .ZN(n4656) );
  INV_X1 U5227 ( .A(n6288), .ZN(n4659) );
  INV_X1 U5228 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5759) );
  INV_X1 U5229 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5760) );
  INV_X1 U5230 ( .A(n4516), .ZN(n4514) );
  NOR2_X1 U5231 ( .A1(n4518), .A2(n4517), .ZN(n4511) );
  AOI21_X1 U5232 ( .B1(n4518), .B2(n4510), .A(n4507), .ZN(n4506) );
  AND2_X1 U5233 ( .A1(n5644), .A2(SI_24_), .ZN(n5651) );
  INV_X1 U5234 ( .A(n4853), .ZN(n4852) );
  OAI21_X1 U5235 ( .B1(n4855), .B2(n4854), .A(n5549), .ZN(n4853) );
  INV_X1 U5236 ( .A(n5531), .ZN(n4854) );
  NAND2_X1 U5237 ( .A1(n8300), .A2(n6152), .ZN(n6159) );
  OR2_X1 U5238 ( .A1(n8822), .A2(n8398), .ZN(n6296) );
  NAND2_X1 U5239 ( .A1(n6042), .A2(n4757), .ZN(n4756) );
  INV_X1 U5240 ( .A(n4760), .ZN(n4757) );
  NOR2_X1 U5241 ( .A1(n8827), .A2(n4823), .ZN(n4822) );
  INV_X1 U5242 ( .A(n4824), .ZN(n4823) );
  NOR2_X1 U5243 ( .A1(n8695), .A2(n4761), .ZN(n4760) );
  NOR2_X1 U5244 ( .A1(n8295), .A2(n8861), .ZN(n4812) );
  AND2_X1 U5245 ( .A1(n4766), .A2(n6248), .ZN(n4765) );
  NAND2_X1 U5246 ( .A1(n6245), .A2(n7545), .ZN(n4766) );
  NAND2_X1 U5247 ( .A1(n5893), .A2(n6234), .ZN(n7531) );
  NAND2_X1 U5248 ( .A1(n7401), .A2(n7299), .ZN(n4537) );
  INV_X1 U5249 ( .A(n7399), .ZN(n7401) );
  NAND2_X1 U5250 ( .A1(n7294), .A2(n7230), .ZN(n4820) );
  AOI21_X1 U5251 ( .B1(n4904), .B2(n7783), .A(n4452), .ZN(n4903) );
  NOR2_X1 U5252 ( .A1(n7025), .A2(n7024), .ZN(n7290) );
  INV_X1 U5253 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5780) );
  INV_X1 U5254 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4825) );
  INV_X1 U5255 ( .A(n6350), .ZN(n5779) );
  INV_X1 U5256 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5778) );
  NOR2_X1 U5257 ( .A1(n5429), .A2(n4951), .ZN(n4945) );
  NOR2_X1 U5258 ( .A1(n7498), .A2(n4478), .ZN(n7695) );
  NOR2_X1 U5259 ( .A1(n9208), .A2(n4555), .ZN(n4554) );
  INV_X1 U5260 ( .A(n4561), .ZN(n4555) );
  OR2_X1 U5261 ( .A1(n9427), .A2(n9299), .ZN(n9140) );
  OR2_X1 U5262 ( .A1(n9437), .A2(n9335), .ZN(n8146) );
  INV_X1 U5263 ( .A(n7739), .ZN(n4574) );
  AND2_X1 U5264 ( .A1(n8146), .A2(n9330), .ZN(n8028) );
  OR2_X1 U5265 ( .A1(n7982), .A2(n9044), .ZN(n7739) );
  INV_X1 U5266 ( .A(n7663), .ZN(n4578) );
  OR2_X1 U5267 ( .A1(n7982), .A2(n7662), .ZN(n4608) );
  OAI21_X1 U5268 ( .B1(n7166), .B2(n4582), .A(n8016), .ZN(n4581) );
  INV_X1 U5269 ( .A(n8101), .ZN(n7166) );
  NAND2_X1 U5270 ( .A1(n4603), .A2(n9123), .ZN(n4602) );
  INV_X1 U5271 ( .A(n4604), .ZN(n4603) );
  NOR2_X1 U5272 ( .A1(n9353), .A2(n9437), .ZN(n9337) );
  AOI21_X1 U5273 ( .B1(n6667), .B2(n6648), .A(n6646), .ZN(n7107) );
  AND2_X1 U5274 ( .A1(n5729), .A2(n6647), .ZN(n7108) );
  INV_X1 U5275 ( .A(n6124), .ZN(n4847) );
  AOI21_X1 U5276 ( .B1(n4838), .B2(n5672), .A(n4836), .ZN(n4835) );
  INV_X1 U5277 ( .A(n6086), .ZN(n4836) );
  INV_X1 U5278 ( .A(n4838), .ZN(n4837) );
  INV_X1 U5279 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5721) );
  AOI21_X1 U5280 ( .B1(n4875), .B2(n4873), .A(n4872), .ZN(n4871) );
  NOR2_X1 U5281 ( .A1(n5434), .A2(n4878), .ZN(n4877) );
  INV_X1 U5282 ( .A(n5404), .ZN(n4878) );
  AND2_X1 U5283 ( .A1(n5455), .A2(n5437), .ZN(n5453) );
  AOI21_X1 U5284 ( .B1(n4877), .B2(n5405), .A(n4876), .ZN(n4875) );
  INV_X1 U5285 ( .A(n5433), .ZN(n4876) );
  NAND2_X1 U5286 ( .A1(n5384), .A2(n5383), .ZN(n5406) );
  NOR2_X1 U5287 ( .A1(n5338), .A2(n4786), .ZN(n4785) );
  INV_X1 U5288 ( .A(n5312), .ZN(n4786) );
  NAND2_X1 U5289 ( .A1(n4857), .A2(n4858), .ZN(n4787) );
  AND2_X1 U5290 ( .A1(n4859), .A2(n5289), .ZN(n4861) );
  INV_X1 U5291 ( .A(n5265), .ZN(n4862) );
  NAND2_X1 U5292 ( .A1(n5020), .A2(n4926), .ZN(n4929) );
  INV_X1 U5293 ( .A(n5178), .ZN(n4828) );
  NAND2_X1 U5294 ( .A1(n5093), .A2(n4451), .ZN(n4500) );
  NOR2_X1 U5295 ( .A1(n4971), .A2(n4970), .ZN(n4969) );
  INV_X1 U5296 ( .A(n6531), .ZN(n4970) );
  NOR2_X1 U5297 ( .A1(n4977), .A2(n4972), .ZN(n4971) );
  INV_X1 U5298 ( .A(n4973), .ZN(n4972) );
  XNOR2_X1 U5299 ( .A(n4401), .B(n7224), .ZN(n7084) );
  XNOR2_X1 U5300 ( .A(n7230), .B(n6538), .ZN(n6426) );
  AND2_X1 U5301 ( .A1(n6459), .A2(n6454), .ZN(n4993) );
  NOR2_X1 U5302 ( .A1(n8479), .A2(n4974), .ZN(n4973) );
  INV_X1 U5303 ( .A(n4976), .ZN(n4974) );
  NAND2_X1 U5304 ( .A1(n4690), .A2(n4688), .ZN(n4687) );
  INV_X1 U5305 ( .A(n6311), .ZN(n4688) );
  NAND2_X1 U5306 ( .A1(n4685), .A2(n4689), .ZN(n4683) );
  AOI21_X1 U5307 ( .B1(n4460), .B2(n4690), .A(n6323), .ZN(n4686) );
  AND2_X1 U5308 ( .A1(n6122), .A2(n6121), .ZN(n8328) );
  OR2_X1 U5309 ( .A1(n6580), .A2(n6132), .ZN(n6122) );
  OR3_X1 U5310 ( .A1(n7726), .A2(n7816), .A3(n7813), .ZN(n6762) );
  AND4_X1 U5311 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n7400)
         );
  NAND2_X1 U5312 ( .A1(n5827), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4990) );
  INV_X1 U5313 ( .A(n4985), .ZN(n4984) );
  NAND2_X1 U5314 ( .A1(n4408), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U5315 ( .A1(n4645), .A2(n4644), .ZN(n4643) );
  OR2_X1 U5316 ( .A1(n6846), .A2(n6845), .ZN(n4636) );
  AND2_X1 U5317 ( .A1(n4636), .A2(n4635), .ZN(n6835) );
  NAND2_X1 U5318 ( .A1(n6784), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4635) );
  OR2_X1 U5319 ( .A1(n6835), .A2(n6834), .ZN(n4634) );
  NOR2_X1 U5320 ( .A1(n8810), .A2(n8620), .ZN(n8610) );
  AOI21_X1 U5321 ( .B1(n8595), .B2(n4887), .A(n4475), .ZN(n4886) );
  INV_X1 U5322 ( .A(n8292), .ZN(n4887) );
  OAI21_X1 U5323 ( .B1(n8668), .B2(n4891), .A(n4420), .ZN(n8618) );
  OR2_X1 U5324 ( .A1(n8822), .A2(n8663), .ZN(n8291) );
  NAND2_X1 U5325 ( .A1(n4893), .A2(n4896), .ZN(n4892) );
  AOI21_X1 U5326 ( .B1(n4897), .B2(n8677), .A(n4447), .ZN(n4895) );
  INV_X1 U5327 ( .A(n4897), .ZN(n4896) );
  INV_X1 U5328 ( .A(n8668), .ZN(n8290) );
  AND2_X1 U5329 ( .A1(n8659), .A2(n4440), .ZN(n4897) );
  AND2_X1 U5330 ( .A1(n6053), .A2(n6288), .ZN(n8677) );
  INV_X1 U5331 ( .A(n6023), .ZN(n4759) );
  NAND2_X1 U5332 ( .A1(n6023), .A2(n4760), .ZN(n8696) );
  NOR2_X1 U5333 ( .A1(n8718), .A2(n8842), .ZN(n8705) );
  AND4_X1 U5334 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n9534)
         );
  INV_X1 U5335 ( .A(n4741), .ZN(n4740) );
  AOI21_X1 U5336 ( .B1(n4741), .B2(n4739), .A(n4738), .ZN(n4737) );
  INV_X1 U5337 ( .A(n6261), .ZN(n4739) );
  INV_X1 U5338 ( .A(n6264), .ZN(n4738) );
  NAND2_X1 U5339 ( .A1(n9528), .A2(n6261), .ZN(n4743) );
  AND2_X1 U5340 ( .A1(n6257), .A2(n6256), .ZN(n8278) );
  AND4_X1 U5341 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n8280)
         );
  NAND2_X1 U5342 ( .A1(n4906), .A2(n7704), .ZN(n7786) );
  NAND2_X1 U5343 ( .A1(n4901), .A2(n4900), .ZN(n7554) );
  AND2_X1 U5344 ( .A1(n6253), .A2(n6251), .ZN(n7702) );
  NAND2_X1 U5345 ( .A1(n7531), .A2(n7532), .ZN(n7618) );
  NOR2_X1 U5346 ( .A1(n7955), .A2(n9881), .ZN(n7957) );
  AND2_X1 U5347 ( .A1(n6227), .A2(n6228), .ZN(n7399) );
  NAND2_X1 U5348 ( .A1(n7071), .A2(n4745), .ZN(n4748) );
  NOR2_X1 U5349 ( .A1(n6199), .A2(n4749), .ZN(n4745) );
  NAND2_X1 U5350 ( .A1(n6194), .A2(n6218), .ZN(n9803) );
  OR2_X1 U5351 ( .A1(n6572), .A2(n6571), .ZN(n9535) );
  INV_X1 U5352 ( .A(n9787), .ZN(n9533) );
  NAND2_X1 U5353 ( .A1(n6131), .A2(n6130), .ZN(n8794) );
  NAND2_X1 U5354 ( .A1(n6006), .A2(n6005), .ZN(n8849) );
  NAND2_X1 U5355 ( .A1(n5997), .A2(n5996), .ZN(n8852) );
  AND2_X1 U5356 ( .A1(n8764), .A2(n8760), .ZN(n8858) );
  NOR2_X1 U5357 ( .A1(n9519), .A2(n8861), .ZN(n8759) );
  AND2_X1 U5358 ( .A1(n6399), .A2(n7526), .ZN(n9883) );
  NOR2_X1 U5359 ( .A1(n6541), .A2(n7816), .ZN(n9810) );
  AND2_X1 U5360 ( .A1(n5780), .A2(n5787), .ZN(n4997) );
  INV_X1 U5361 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5763) );
  AND2_X1 U5362 ( .A1(n5954), .A2(n5947), .ZN(n7848) );
  AND2_X1 U5363 ( .A1(n5810), .A2(n5834), .ZN(n5835) );
  NAND2_X1 U5364 ( .A1(n5502), .A2(n8999), .ZN(n4909) );
  AND2_X1 U5365 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  INV_X1 U5366 ( .A(n4959), .ZN(n4958) );
  AOI21_X1 U5367 ( .B1(n4959), .B2(n4957), .A(n4956), .ZN(n4955) );
  AOI21_X1 U5368 ( .B1(n7601), .B2(n5287), .A(n4960), .ZN(n4959) );
  AND2_X1 U5369 ( .A1(n8970), .A2(n8940), .ZN(n4914) );
  NAND2_X1 U5370 ( .A1(n5726), .A2(n5049), .ZN(n8198) );
  OR2_X1 U5371 ( .A1(n5730), .A2(n8259), .ZN(n5744) );
  NOR2_X1 U5372 ( .A1(n5432), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U5373 ( .A1(n4462), .A2(n4954), .ZN(n4944) );
  NAND2_X1 U5374 ( .A1(n5381), .A2(n5380), .ZN(n4952) );
  NAND2_X1 U5375 ( .A1(n7894), .A2(n4945), .ZN(n4934) );
  AND2_X1 U5376 ( .A1(n4948), .A2(n4953), .ZN(n4947) );
  NAND2_X1 U5377 ( .A1(n5427), .A2(n4949), .ZN(n4948) );
  AND2_X1 U5378 ( .A1(n5381), .A2(n5380), .ZN(n4949) );
  AND2_X1 U5379 ( .A1(n5728), .A2(n9305), .ZN(n8255) );
  NAND2_X1 U5380 ( .A1(n5726), .A2(n9305), .ZN(n6946) );
  AND2_X1 U5381 ( .A1(n9613), .A2(n9612), .ZN(n9615) );
  XNOR2_X1 U5382 ( .A(n7695), .B(n7694), .ZN(n7500) );
  NOR2_X1 U5383 ( .A1(n7500), .A2(n7673), .ZN(n7696) );
  XNOR2_X1 U5384 ( .A(n9168), .B(n9167), .ZN(n9169) );
  OAI21_X1 U5385 ( .B1(n9188), .B2(n9165), .A(n9164), .ZN(n9168) );
  INV_X1 U5386 ( .A(n9041), .ZN(n9191) );
  INV_X1 U5387 ( .A(n4558), .ZN(n4557) );
  AOI21_X1 U5388 ( .B1(n9297), .B2(n4703), .A(n4701), .ZN(n4700) );
  NAND2_X1 U5389 ( .A1(n4702), .A2(n9260), .ZN(n4701) );
  NAND2_X1 U5390 ( .A1(n4703), .A2(n4706), .ZN(n4702) );
  AND2_X1 U5391 ( .A1(n8241), .A2(n9242), .ZN(n9260) );
  NOR2_X1 U5392 ( .A1(n9156), .A2(n8156), .ZN(n4710) );
  INV_X1 U5393 ( .A(n4793), .ZN(n4792) );
  INV_X1 U5394 ( .A(n4427), .ZN(n4791) );
  OR2_X1 U5395 ( .A1(n9158), .A2(n4704), .ZN(n9267) );
  OAI21_X1 U5396 ( .B1(n9313), .B2(n9141), .A(n9140), .ZN(n9308) );
  NAND2_X1 U5397 ( .A1(n4714), .A2(n4712), .ZN(n9298) );
  NAND2_X1 U5398 ( .A1(n4713), .A2(n4715), .ZN(n4712) );
  NAND2_X1 U5399 ( .A1(n4716), .A2(n9153), .ZN(n4713) );
  AND2_X1 U5400 ( .A1(n4718), .A2(n9151), .ZN(n4716) );
  NAND2_X1 U5401 ( .A1(n9150), .A2(n4431), .ZN(n4717) );
  NAND2_X1 U5402 ( .A1(n4717), .A2(n4718), .ZN(n9331) );
  NAND2_X1 U5403 ( .A1(n4795), .A2(n7907), .ZN(n7914) );
  NAND2_X1 U5404 ( .A1(n9349), .A2(n4429), .ZN(n4795) );
  OR2_X1 U5405 ( .A1(n9348), .A2(n7910), .ZN(n7913) );
  INV_X1 U5406 ( .A(n8062), .ZN(n4725) );
  OR2_X1 U5407 ( .A1(n8133), .A2(n8134), .ZN(n8131) );
  NAND2_X1 U5408 ( .A1(n7668), .A2(n7666), .ZN(n7746) );
  NOR2_X1 U5409 ( .A1(n8113), .A2(n4698), .ZN(n4697) );
  INV_X1 U5410 ( .A(n8057), .ZN(n4698) );
  AND2_X1 U5411 ( .A1(n8056), .A2(n8043), .ZN(n8023) );
  NAND2_X1 U5412 ( .A1(n5346), .A2(n5345), .ZN(n7563) );
  NAND2_X1 U5413 ( .A1(n5316), .A2(n5315), .ZN(n7476) );
  OAI211_X1 U5414 ( .C1(n5294), .C2(n6748), .A(n5223), .B(n5222), .ZN(n8094)
         );
  OAI21_X1 U5415 ( .B1(n4567), .B2(n4566), .A(n4563), .ZN(n7241) );
  AND2_X1 U5416 ( .A1(n4564), .A2(n7162), .ZN(n4563) );
  NAND2_X1 U5417 ( .A1(n6939), .A2(n6938), .ZN(n8216) );
  INV_X1 U5418 ( .A(n9685), .ZN(n9363) );
  OR2_X1 U5419 ( .A1(n9603), .A2(n4965), .ZN(n4963) );
  NAND2_X1 U5420 ( .A1(n4377), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4965) );
  XNOR2_X1 U5421 ( .A(n9055), .B(n7122), .ZN(n6942) );
  OR2_X1 U5422 ( .A1(n8198), .A2(n9606), .ZN(n9683) );
  OR2_X1 U5423 ( .A1(n8198), .A2(n4378), .ZN(n9685) );
  INV_X1 U5424 ( .A(n9683), .ZN(n9664) );
  NOR2_X1 U5425 ( .A1(n9382), .A2(n9381), .ZN(n4618) );
  NAND2_X1 U5426 ( .A1(n5657), .A2(n5656), .ZN(n9400) );
  NOR2_X1 U5427 ( .A1(n5704), .A2(n7720), .ZN(n5057) );
  XNOR2_X1 U5428 ( .A(n6168), .B(n6167), .ZN(n8888) );
  XNOR2_X1 U5429 ( .A(n6160), .B(n6144), .ZN(n8310) );
  NAND2_X1 U5430 ( .A1(n6107), .A2(n6106), .ZN(n6109) );
  XNOR2_X1 U5431 ( .A(n5056), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U5432 ( .A1(n5055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U5433 ( .A1(n5054), .A2(n5051), .ZN(n5055) );
  NAND2_X1 U5434 ( .A1(n4834), .A2(n4838), .ZN(n6087) );
  NAND2_X1 U5435 ( .A1(n5675), .A2(n5673), .ZN(n4834) );
  XNOR2_X1 U5436 ( .A(n5621), .B(n5649), .ZN(n7719) );
  NAND2_X1 U5437 ( .A1(n4851), .A2(n5531), .ZN(n5550) );
  NOR2_X1 U5438 ( .A1(n5043), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U5439 ( .A1(n5256), .A2(n5265), .ZN(n4866) );
  NAND2_X1 U5440 ( .A1(n4879), .A2(n5221), .ZN(n5248) );
  NAND2_X1 U5441 ( .A1(n5175), .A2(n5174), .ZN(n4830) );
  AND4_X1 U5442 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n7709)
         );
  AND3_X1 U5443 ( .A1(n6020), .A2(n6019), .A3(n6018), .ZN(n8373) );
  NAND2_X1 U5444 ( .A1(n6068), .A2(n6067), .ZN(n8818) );
  NAND2_X1 U5445 ( .A1(n4383), .A2(n6427), .ZN(n7140) );
  NAND2_X1 U5446 ( .A1(n5934), .A2(n5933), .ZN(n8866) );
  AND2_X1 U5447 ( .A1(n6041), .A2(n6040), .ZN(n8372) );
  AND4_X1 U5448 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(n8471)
         );
  NAND2_X1 U5449 ( .A1(n5957), .A2(n5956), .ZN(n8294) );
  NAND2_X1 U5450 ( .A1(n5009), .A2(n4650), .ZN(n4647) );
  NOR2_X1 U5451 ( .A1(n6342), .A2(n4651), .ZN(n4650) );
  INV_X1 U5452 ( .A(n8372), .ZN(n8698) );
  INV_X1 U5453 ( .A(n8373), .ZN(n8697) );
  AND2_X1 U5454 ( .A1(n6779), .A2(n6778), .ZN(n9773) );
  NAND2_X1 U5455 ( .A1(n6805), .A2(n6804), .ZN(n9776) );
  AND2_X1 U5456 ( .A1(n4817), .A2(n4815), .ZN(n8795) );
  NAND2_X1 U5457 ( .A1(n8564), .A2(n8794), .ZN(n4817) );
  AOI21_X1 U5458 ( .B1(n8306), .B2(n9790), .A(n8305), .ZN(n8797) );
  NAND2_X1 U5459 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  AND2_X1 U5460 ( .A1(n4775), .A2(n4774), .ZN(n8802) );
  AOI21_X1 U5461 ( .B1(n8571), .B2(n9785), .A(n4473), .ZN(n4774) );
  NAND2_X1 U5462 ( .A1(n4776), .A2(n9790), .ZN(n4775) );
  AND2_X1 U5463 ( .A1(n7968), .A2(n9883), .ZN(n9521) );
  NAND2_X1 U5464 ( .A1(n9791), .A2(n9537), .ZN(n8748) );
  NAND3_X1 U5465 ( .A1(n4547), .A2(n4545), .A3(n4544), .ZN(n8798) );
  NAND2_X1 U5466 ( .A1(n4423), .A2(n4471), .ZN(n4544) );
  OR2_X1 U5467 ( .A1(n8562), .A2(n4692), .ZN(n4547) );
  NAND2_X1 U5468 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  NAND2_X1 U5469 ( .A1(n7729), .A2(n5333), .ZN(n9508) );
  AND2_X1 U5470 ( .A1(n5179), .A2(n4501), .ZN(n9722) );
  AND2_X1 U5471 ( .A1(n5180), .A2(n4436), .ZN(n4501) );
  NAND2_X1 U5472 ( .A1(n5574), .A2(n5573), .ZN(n9417) );
  NAND2_X1 U5473 ( .A1(n4908), .A2(n4907), .ZN(n7985) );
  NAND2_X1 U5474 ( .A1(n5014), .A2(n6928), .ZN(n4907) );
  INV_X1 U5475 ( .A(n6926), .ZN(n5099) );
  NAND2_X1 U5476 ( .A1(n5664), .A2(n5663), .ZN(n9262) );
  OR2_X1 U5477 ( .A1(n9238), .A2(n5581), .ZN(n5664) );
  NAND2_X1 U5478 ( .A1(n5633), .A2(n5632), .ZN(n9245) );
  OR2_X1 U5479 ( .A1(n9254), .A2(n5581), .ZN(n5633) );
  NAND2_X1 U5480 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
  NAND2_X1 U5481 ( .A1(n4731), .A2(n9389), .ZN(n9458) );
  NOR2_X1 U5482 ( .A1(n9386), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5483 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  OR2_X1 U5484 ( .A1(n5033), .A2(n5032), .ZN(n9472) );
  INV_X1 U5485 ( .A(n8119), .ZN(n4498) );
  NAND2_X1 U5486 ( .A1(n8122), .A2(n8121), .ZN(n4497) );
  AOI21_X1 U5487 ( .B1(n6213), .B2(n6316), .A(n4693), .ZN(n6215) );
  NOR2_X1 U5488 ( .A1(n4694), .A2(n6212), .ZN(n4693) );
  AOI21_X1 U5489 ( .B1(n4494), .B2(n4441), .A(n4486), .ZN(n8141) );
  NAND2_X1 U5490 ( .A1(n4488), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U5491 ( .A1(n4495), .A2(n8132), .ZN(n4494) );
  AND2_X1 U5492 ( .A1(n8278), .A2(n4671), .ZN(n4670) );
  AOI21_X1 U5493 ( .B1(n6252), .B2(n4668), .A(n4666), .ZN(n4665) );
  INV_X1 U5494 ( .A(n4524), .ZN(n4523) );
  NAND2_X1 U5495 ( .A1(n4532), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U5496 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  NAND2_X1 U5497 ( .A1(n4534), .A2(n4533), .ZN(n4532) );
  INV_X1 U5498 ( .A(n4527), .ZN(n4522) );
  AOI21_X1 U5499 ( .B1(n4524), .B2(n4526), .A(n4455), .ZN(n4519) );
  INV_X1 U5500 ( .A(n4529), .ZN(n4526) );
  NAND2_X1 U5501 ( .A1(n4674), .A2(n4673), .ZN(n6274) );
  INV_X1 U5502 ( .A(n6270), .ZN(n4673) );
  NAND2_X1 U5503 ( .A1(n4677), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5504 ( .A1(n8180), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U5505 ( .A1(n4517), .A2(n4509), .ZN(n4504) );
  NAND2_X1 U5506 ( .A1(n8180), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5507 ( .A1(n4517), .A2(n4509), .ZN(n4508) );
  INV_X1 U5508 ( .A(n8170), .ZN(n4518) );
  NAND2_X1 U5509 ( .A1(n7549), .A2(n4899), .ZN(n7548) );
  INV_X1 U5510 ( .A(n7705), .ZN(n4905) );
  NAND2_X1 U5511 ( .A1(n4512), .A2(n4516), .ZN(n8191) );
  OAI21_X1 U5512 ( .B1(n8177), .B2(n4505), .A(n4502), .ZN(n4512) );
  AOI21_X1 U5513 ( .B1(n4518), .B2(n4510), .A(n4503), .ZN(n4502) );
  NOR2_X1 U5514 ( .A1(n4518), .A2(n4517), .ZN(n4505) );
  AND2_X1 U5515 ( .A1(n9260), .A2(n9269), .ZN(n8164) );
  NAND2_X1 U5516 ( .A1(n7170), .A2(n8212), .ZN(n9682) );
  AOI21_X1 U5517 ( .B1(n6109), .B2(n4844), .A(n4841), .ZN(n4840) );
  NOR2_X1 U5518 ( .A1(n4846), .A2(n6142), .ZN(n4844) );
  OAI21_X1 U5519 ( .B1(n4846), .B2(n4842), .A(n6141), .ZN(n4841) );
  INV_X1 U5520 ( .A(SI_21_), .ZN(n10076) );
  NOR2_X1 U5521 ( .A1(n4874), .A2(n4869), .ZN(n4868) );
  INV_X1 U5522 ( .A(n5383), .ZN(n4869) );
  INV_X1 U5523 ( .A(n4875), .ZN(n4874) );
  INV_X1 U5524 ( .A(n4877), .ZN(n4873) );
  INV_X1 U5525 ( .A(n5453), .ZN(n4872) );
  INV_X1 U5526 ( .A(n5337), .ZN(n4783) );
  XNOR2_X1 U5527 ( .A(n4805), .B(n6421), .ZN(n6408) );
  NAND2_X1 U5528 ( .A1(n7019), .A2(n6529), .ZN(n6407) );
  OR2_X1 U5529 ( .A1(n8395), .A2(n8394), .ZN(n4977) );
  OR2_X1 U5530 ( .A1(n6292), .A2(n4657), .ZN(n4654) );
  AND2_X1 U5531 ( .A1(n4663), .A2(n4469), .ZN(n4655) );
  OR2_X1 U5532 ( .A1(n6300), .A2(n6327), .ZN(n4663) );
  NOR2_X1 U5533 ( .A1(n4692), .A2(n4691), .ZN(n4690) );
  INV_X1 U5534 ( .A(n6315), .ZN(n4691) );
  AND2_X1 U5535 ( .A1(n6328), .A2(n6321), .ZN(n6322) );
  AOI21_X1 U5536 ( .B1(n8623), .B2(n6298), .A(n6301), .ZN(n8600) );
  NOR2_X1 U5537 ( .A1(n8832), .A2(n8837), .ZN(n4824) );
  NAND2_X1 U5538 ( .A1(n4812), .A2(n8739), .ZN(n4811) );
  NAND2_X1 U5539 ( .A1(n7019), .A2(n4805), .ZN(n6203) );
  NAND2_X1 U5540 ( .A1(n5798), .A2(n9844), .ZN(n6176) );
  INV_X1 U5541 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5542 ( .A1(n6337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U5543 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  INV_X1 U5544 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6338) );
  INV_X1 U5545 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5546 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5757) );
  NOR2_X1 U5547 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5756) );
  INV_X1 U5548 ( .A(n5761), .ZN(n4983) );
  AND3_X1 U5549 ( .A1(n5810), .A2(n5762), .A3(n5834), .ZN(n5858) );
  NAND2_X1 U5550 ( .A1(n7117), .A2(n5098), .ZN(n5069) );
  AOI21_X1 U5551 ( .B1(n6359), .B2(n7150), .A(n5003), .ZN(n5068) );
  INV_X1 U5552 ( .A(n7629), .ZN(n4960) );
  INV_X1 U5553 ( .A(n7628), .ZN(n4956) );
  INV_X1 U5554 ( .A(n5287), .ZN(n4957) );
  NOR2_X1 U5555 ( .A1(n5476), .A2(n4937), .ZN(n4932) );
  NOR2_X1 U5556 ( .A1(n8182), .A2(n8181), .ZN(n8195) );
  AND2_X1 U5557 ( .A1(n4515), .A2(n4513), .ZN(n8187) );
  NAND2_X1 U5558 ( .A1(n4514), .A2(n4430), .ZN(n4513) );
  INV_X1 U5559 ( .A(SI_15_), .ZN(n10088) );
  INV_X1 U5560 ( .A(SI_13_), .ZN(n10219) );
  INV_X1 U5561 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5024) );
  INV_X1 U5562 ( .A(SI_16_), .ZN(n10216) );
  NAND2_X1 U5563 ( .A1(n4613), .A2(n9241), .ZN(n4612) );
  NOR2_X1 U5564 ( .A1(n9406), .A2(n9412), .ZN(n4613) );
  NOR2_X1 U5565 ( .A1(n5391), .A2(n7496), .ZN(n5415) );
  NAND2_X1 U5566 ( .A1(n9722), .A2(n9051), .ZN(n8013) );
  INV_X1 U5567 ( .A(n4569), .ZN(n4565) );
  NAND2_X1 U5568 ( .A1(n9686), .A2(n6937), .ZN(n4569) );
  INV_X1 U5569 ( .A(n6670), .ZN(n6667) );
  OR2_X1 U5570 ( .A1(n5619), .A2(n5618), .ZN(n5648) );
  OR2_X1 U5571 ( .A1(n5615), .A2(n5619), .ZN(n5645) );
  NAND2_X1 U5572 ( .A1(n4850), .A2(n4848), .ZN(n5563) );
  AOI21_X1 U5573 ( .B1(n4852), .B2(n4854), .A(n4849), .ZN(n4848) );
  INV_X1 U5574 ( .A(n5551), .ZN(n4849) );
  NOR2_X1 U5575 ( .A1(n5532), .A2(n4856), .ZN(n4855) );
  INV_X1 U5576 ( .A(n5507), .ZN(n4856) );
  OAI21_X1 U5577 ( .B1(n6628), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5158), .ZN(
        n5176) );
  NOR2_X2 U5578 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5101) );
  INV_X1 U5579 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5059) );
  INV_X1 U5580 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4802) );
  AND2_X1 U5581 ( .A1(n5851), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5867) );
  INV_X1 U5582 ( .A(n5999), .ZN(n5998) );
  OR2_X1 U5583 ( .A1(n5986), .A2(n8516), .ZN(n5999) );
  NAND2_X1 U5584 ( .A1(n8466), .A2(n4980), .ZN(n4979) );
  NOR2_X1 U5585 ( .A1(n8356), .A2(n4981), .ZN(n4980) );
  INV_X1 U5586 ( .A(n6505), .ZN(n4981) );
  NAND2_X1 U5587 ( .A1(n6033), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U5588 ( .A1(n8395), .A2(n8394), .ZN(n4976) );
  NAND2_X2 U5589 ( .A1(n6488), .A2(n6487), .ZN(n8267) );
  INV_X1 U5590 ( .A(n6485), .ZN(n6488) );
  AND3_X1 U5591 ( .A1(n6150), .A2(n6149), .A3(n6148), .ZN(n6681) );
  AND4_X1 U5592 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n8444)
         );
  AND2_X1 U5593 ( .A1(n4643), .A2(n4642), .ZN(n6811) );
  INV_X1 U5594 ( .A(n6812), .ZN(n4642) );
  NOR2_X1 U5595 ( .A1(n6811), .A2(n4641), .ZN(n6824) );
  AND2_X1 U5596 ( .A1(n6787), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4641) );
  AND2_X1 U5597 ( .A1(n4634), .A2(n4633), .ZN(n6895) );
  NAND2_X1 U5598 ( .A1(n6775), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U5599 ( .A1(n6893), .A2(n4638), .ZN(n6781) );
  AND2_X1 U5600 ( .A1(n6898), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5601 ( .A1(n6781), .A2(n6780), .ZN(n6955) );
  NOR2_X1 U5602 ( .A1(n6955), .A2(n4637), .ZN(n6958) );
  AND2_X1 U5603 ( .A1(n6961), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5604 ( .A1(n6958), .A2(n6957), .ZN(n7125) );
  NOR2_X1 U5605 ( .A1(n7354), .A2(n4640), .ZN(n7358) );
  AND2_X1 U5606 ( .A1(n7355), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4640) );
  NOR2_X1 U5607 ( .A1(n7358), .A2(n7357), .ZN(n7417) );
  NOR2_X1 U5608 ( .A1(n7417), .A2(n4639), .ZN(n7420) );
  AND2_X1 U5609 ( .A1(n7418), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4639) );
  NAND2_X1 U5610 ( .A1(n7420), .A2(n7419), .ZN(n7515) );
  INV_X1 U5611 ( .A(n8509), .ZN(n4623) );
  INV_X1 U5612 ( .A(n4815), .ZN(n8555) );
  AOI21_X1 U5613 ( .B1(n8570), .B2(n6310), .A(n6123), .ZN(n8301) );
  NAND2_X1 U5614 ( .A1(n8589), .A2(n9787), .ZN(n8304) );
  NOR2_X1 U5615 ( .A1(n8799), .A2(n8804), .ZN(n4813) );
  NAND2_X1 U5616 ( .A1(n6313), .A2(n6314), .ZN(n8569) );
  AOI21_X1 U5617 ( .B1(n4886), .B2(n8599), .A(n6306), .ZN(n4885) );
  AND2_X1 U5618 ( .A1(n6104), .A2(n6103), .ZN(n8604) );
  OR2_X1 U5619 ( .A1(n8581), .A2(n6132), .ZN(n6104) );
  NAND2_X1 U5620 ( .A1(n8705), .A2(n4443), .ZN(n8635) );
  INV_X1 U5621 ( .A(n6042), .ZN(n4758) );
  AND2_X1 U5622 ( .A1(n8705), .A2(n4822), .ZN(n8654) );
  NAND2_X1 U5623 ( .A1(n8705), .A2(n4824), .ZN(n8670) );
  NAND2_X1 U5624 ( .A1(n8705), .A2(n8694), .ZN(n8688) );
  INV_X1 U5625 ( .A(n4812), .ZN(n4810) );
  AOI21_X1 U5626 ( .B1(n4542), .B2(n8282), .A(n4474), .ZN(n4541) );
  OR2_X1 U5627 ( .A1(n9518), .A2(n8294), .ZN(n9519) );
  NAND2_X1 U5628 ( .A1(n5949), .A2(n5948), .ZN(n8277) );
  NAND2_X1 U5629 ( .A1(n7790), .A2(n9548), .ZN(n9518) );
  NOR2_X1 U5630 ( .A1(n7791), .A2(n8866), .ZN(n7790) );
  AOI21_X1 U5631 ( .B1(n4765), .B2(n4767), .A(n4764), .ZN(n4763) );
  INV_X1 U5632 ( .A(n6245), .ZN(n4767) );
  AND4_X1 U5633 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n9532)
         );
  NAND2_X1 U5634 ( .A1(n4807), .A2(n4806), .ZN(n7791) );
  AND4_X1 U5635 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5889), .ZN(n7533)
         );
  AND2_X1 U5636 ( .A1(n7947), .A2(n7402), .ZN(n7403) );
  AND2_X1 U5637 ( .A1(n7957), .A2(n7414), .ZN(n7540) );
  NAND2_X1 U5638 ( .A1(n4537), .A2(n4434), .ZN(n4536) );
  NAND2_X1 U5639 ( .A1(n7946), .A2(n7948), .ZN(n7947) );
  AND2_X1 U5640 ( .A1(n5867), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5879) );
  NOR2_X1 U5641 ( .A1(n4820), .A2(n8317), .ZN(n4818) );
  NAND2_X1 U5642 ( .A1(n7334), .A2(n9877), .ZN(n7336) );
  NAND2_X1 U5643 ( .A1(n4750), .A2(n6200), .ZN(n7340) );
  NAND2_X1 U5644 ( .A1(n4748), .A2(n4746), .ZN(n4750) );
  NOR2_X1 U5645 ( .A1(n6219), .A2(n4747), .ZN(n4746) );
  INV_X1 U5646 ( .A(n6218), .ZN(n4747) );
  NOR2_X1 U5647 ( .A1(n4820), .A2(n9795), .ZN(n7334) );
  AND3_X1 U5648 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5851) );
  NOR2_X1 U5649 ( .A1(n9795), .A2(n9799), .ZN(n9797) );
  NAND2_X1 U5650 ( .A1(n9883), .A2(n4625), .ZN(n7288) );
  NAND3_X1 U5651 ( .A1(n7039), .A2(n7020), .A3(n7021), .ZN(n7067) );
  OR2_X1 U5652 ( .A1(n7026), .A2(n7289), .ZN(n7029) );
  NAND2_X1 U5653 ( .A1(n9837), .A2(n5804), .ZN(n7044) );
  NOR2_X1 U5654 ( .A1(n4423), .A2(n4471), .ZN(n4546) );
  INV_X1 U5655 ( .A(n9883), .ZN(n9900) );
  INV_X1 U5656 ( .A(n4997), .ZN(n4994) );
  NAND2_X1 U5657 ( .A1(n6339), .A2(n6338), .ZN(n6343) );
  OR2_X1 U5658 ( .A1(n5863), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5875) );
  OR2_X1 U5659 ( .A1(n5810), .A2(n10207), .ZN(n5811) );
  INV_X1 U5660 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U5661 ( .A1(n5624), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U5662 ( .A1(n4962), .A2(n4961), .ZN(n7598) );
  INV_X1 U5663 ( .A(n7601), .ZN(n4961) );
  INV_X1 U5664 ( .A(n7600), .ZN(n4962) );
  AND2_X1 U5665 ( .A1(n5083), .A2(n5082), .ZN(n6915) );
  NAND2_X1 U5666 ( .A1(n7117), .A2(n6590), .ZN(n5083) );
  AOI22_X1 U5667 ( .A1(n5098), .A2(n7150), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5081), .ZN(n5082) );
  NAND2_X1 U5668 ( .A1(n6915), .A2(n5084), .ZN(n6916) );
  NAND2_X1 U5669 ( .A1(n5516), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U5670 ( .A1(n8998), .A2(n9000), .ZN(n4910) );
  INV_X1 U5671 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5372) );
  OR2_X1 U5672 ( .A1(n5373), .A2(n5372), .ZN(n5391) );
  INV_X1 U5673 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10149) );
  OR2_X1 U5674 ( .A1(n5492), .A2(n10149), .ZN(n5518) );
  NAND2_X1 U5675 ( .A1(n5462), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5492) );
  INV_X1 U5676 ( .A(n5464), .ZN(n5462) );
  NAND2_X1 U5677 ( .A1(n4918), .A2(n4916), .ZN(n5703) );
  AND2_X1 U5678 ( .A1(n4917), .A2(n8940), .ZN(n4916) );
  NAND2_X1 U5679 ( .A1(n9371), .A2(n9127), .ZN(n8253) );
  NAND2_X1 U5680 ( .A1(n8000), .A2(n7999), .ZN(n8248) );
  INV_X1 U5681 ( .A(n9558), .ZN(n8000) );
  AND2_X1 U5682 ( .A1(n9065), .A2(n6716), .ZN(n9613) );
  NAND2_X1 U5683 ( .A1(n6731), .A2(n4450), .ZN(n6723) );
  NOR2_X1 U5684 ( .A1(n6723), .A2(n6722), .ZN(n6741) );
  NOR2_X1 U5685 ( .A1(n9646), .A2(n4593), .ZN(n6876) );
  AND2_X1 U5686 ( .A1(n9655), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4593) );
  NAND2_X1 U5687 ( .A1(n6876), .A2(n6875), .ZN(n6990) );
  NAND2_X1 U5688 ( .A1(n6990), .A2(n4592), .ZN(n6994) );
  OR2_X1 U5689 ( .A1(n6991), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U5690 ( .A1(n6994), .A2(n6993), .ZN(n7185) );
  NOR2_X1 U5691 ( .A1(n7696), .A2(n7697), .ZN(n7817) );
  NOR2_X1 U5692 ( .A1(n9097), .A2(n4600), .ZN(n9101) );
  AND2_X1 U5693 ( .A1(n9098), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4600) );
  NOR2_X1 U5694 ( .A1(n9101), .A2(n9100), .ZN(n9107) );
  XNOR2_X1 U5695 ( .A(n4598), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9117) );
  OR2_X1 U5696 ( .A1(n9107), .A2(n4599), .ZN(n4598) );
  AND2_X1 U5697 ( .A1(n9111), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U5698 ( .A1(n9397), .A2(n9246), .ZN(n4561) );
  OR2_X1 U5699 ( .A1(n9400), .A2(n9226), .ZN(n9221) );
  AND2_X1 U5700 ( .A1(n8005), .A2(n8173), .ZN(n9223) );
  NOR2_X1 U5701 ( .A1(n9283), .A2(n9412), .ZN(n9274) );
  NOR2_X1 U5702 ( .A1(n9283), .A2(n4611), .ZN(n9252) );
  INV_X1 U5703 ( .A(n4613), .ZN(n4611) );
  INV_X1 U5704 ( .A(n4586), .ZN(n4584) );
  NOR2_X1 U5705 ( .A1(n9313), .A2(n4587), .ZN(n4585) );
  OAI21_X1 U5706 ( .B1(n4411), .B2(n4418), .A(n5000), .ZN(n4586) );
  NOR2_X1 U5707 ( .A1(n9353), .A2(n4604), .ZN(n9338) );
  NOR3_X1 U5708 ( .A1(n9353), .A2(n9427), .A3(n4604), .ZN(n9314) );
  NAND2_X1 U5709 ( .A1(n4571), .A2(n4570), .ZN(n9136) );
  OR2_X1 U5710 ( .A1(n4573), .A2(n4415), .ZN(n4570) );
  NOR2_X1 U5711 ( .A1(n4448), .A2(n4574), .ZN(n4573) );
  OR2_X1 U5712 ( .A1(n8006), .A2(n8042), .ZN(n9351) );
  NOR2_X1 U5713 ( .A1(n4797), .A2(n4439), .ZN(n4796) );
  INV_X1 U5714 ( .A(n7908), .ZN(n4797) );
  NAND2_X1 U5715 ( .A1(n7664), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5716 ( .A1(n5371), .A2(n5370), .ZN(n7662) );
  NOR2_X1 U5717 ( .A1(n7572), .A2(n7662), .ZN(n7672) );
  INV_X1 U5718 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5347) );
  OR2_X1 U5719 ( .A1(n5348), .A2(n5347), .ZN(n5373) );
  NAND2_X1 U5720 ( .A1(n5318), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U5721 ( .A1(n7452), .A2(n8109), .ZN(n7453) );
  OR2_X1 U5722 ( .A1(n5234), .A2(n10214), .ZN(n5274) );
  INV_X1 U5723 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U5724 ( .A1(n7260), .A2(n4711), .ZN(n7382) );
  AND2_X1 U5725 ( .A1(n8018), .A2(n8096), .ZN(n4711) );
  INV_X1 U5726 ( .A(n4581), .ZN(n4580) );
  NAND2_X1 U5727 ( .A1(n8096), .A2(n8219), .ZN(n8016) );
  NAND2_X1 U5728 ( .A1(n4583), .A2(n7166), .ZN(n7206) );
  INV_X1 U5729 ( .A(n7168), .ZN(n4583) );
  AND2_X1 U5730 ( .A1(n7207), .A2(n8013), .ZN(n9671) );
  NAND2_X1 U5731 ( .A1(n7112), .A2(n6945), .ZN(n7159) );
  NOR2_X1 U5732 ( .A1(n7111), .A2(n7117), .ZN(n7118) );
  NAND2_X1 U5733 ( .A1(n9388), .A2(n9727), .ZN(n4733) );
  NAND2_X1 U5734 ( .A1(n5461), .A2(n5460), .ZN(n9442) );
  INV_X1 U5735 ( .A(n9753), .ZN(n9728) );
  INV_X1 U5736 ( .A(n9742), .ZN(n9727) );
  INV_X1 U5737 ( .A(n9755), .ZN(n9740) );
  OR2_X1 U5738 ( .A1(n6936), .A2(n6935), .ZN(n9753) );
  AND2_X1 U5739 ( .A1(n6664), .A2(n7108), .ZN(n6694) );
  INV_X1 U5740 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U5741 ( .A(n6143), .B(n6129), .ZN(n8001) );
  OAI21_X1 U5742 ( .B1(n6109), .B2(n4847), .A(n4845), .ZN(n6143) );
  NAND2_X1 U5743 ( .A1(n4833), .A2(n4831), .ZN(n6107) );
  AOI21_X1 U5744 ( .B1(n4835), .B2(n4837), .A(n4832), .ZN(n4831) );
  INV_X1 U5745 ( .A(n6088), .ZN(n4832) );
  AND2_X1 U5746 ( .A1(n6108), .A2(n6092), .ZN(n6106) );
  XNOR2_X1 U5747 ( .A(n5012), .B(n5672), .ZN(n7812) );
  NAND2_X1 U5748 ( .A1(n5047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5048) );
  OAI21_X2 U5749 ( .B1(n5076), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U5750 ( .A1(n5508), .A2(n5507), .ZN(n5533) );
  INV_X1 U5751 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U5752 ( .A1(n4870), .A2(n4875), .ZN(n5454) );
  NAND2_X1 U5753 ( .A1(n5406), .A2(n4877), .ZN(n4870) );
  XNOR2_X1 U5754 ( .A(n4798), .B(n5434), .ZN(n7062) );
  OAI21_X1 U5755 ( .B1(n5406), .B2(n5405), .A(n5404), .ZN(n4798) );
  INV_X1 U5756 ( .A(n5023), .ZN(n4928) );
  NAND2_X1 U5757 ( .A1(n4784), .A2(n5337), .ZN(n5363) );
  NAND2_X1 U5758 ( .A1(n4787), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5759 ( .A1(n4787), .A2(n5312), .ZN(n5339) );
  OAI21_X1 U5760 ( .B1(n5264), .B2(n4866), .A(n5265), .ZN(n5288) );
  AND2_X1 U5761 ( .A1(n5244), .A2(n5243), .ZN(n5296) );
  NAND2_X1 U5762 ( .A1(n4596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5151) );
  INV_X1 U5763 ( .A(n5101), .ZN(n4596) );
  NAND2_X1 U5764 ( .A1(n4968), .A2(n4966), .ZN(n8326) );
  AOI21_X1 U5765 ( .B1(n4969), .B2(n4972), .A(n4967), .ZN(n4966) );
  INV_X1 U5766 ( .A(n8322), .ZN(n4967) );
  NAND2_X1 U5767 ( .A1(n7317), .A2(n6454), .ZN(n8346) );
  INV_X1 U5768 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U5769 ( .A1(n8466), .A2(n6505), .ZN(n8360) );
  INV_X1 U5770 ( .A(n4805), .ZN(n9844) );
  AND2_X1 U5771 ( .A1(n6065), .A2(n6064), .ZN(n8398) );
  AND2_X1 U5772 ( .A1(n6052), .A2(n6051), .ZN(n8681) );
  NAND2_X1 U5773 ( .A1(n6056), .A2(n6055), .ZN(n8822) );
  AND4_X1 U5774 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n7318)
         );
  AND4_X1 U5775 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8425)
         );
  NAND2_X1 U5776 ( .A1(n4979), .A2(n8359), .ZN(n8422) );
  NAND2_X1 U5777 ( .A1(n6014), .A2(n6013), .ZN(n8842) );
  INV_X1 U5778 ( .A(n6522), .ZN(n6519) );
  OR2_X1 U5779 ( .A1(n8478), .A2(n6979), .ZN(n8464) );
  AND2_X1 U5780 ( .A1(n6972), .A2(n6409), .ZN(n8458) );
  INV_X1 U5781 ( .A(n8482), .ZN(n8472) );
  AND2_X1 U5782 ( .A1(n6078), .A2(n6097), .ZN(n8611) );
  AND2_X1 U5783 ( .A1(n6579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8481) );
  AND2_X1 U5784 ( .A1(n8315), .A2(n9787), .ZN(n8482) );
  NAND2_X1 U5785 ( .A1(n6569), .A2(n6559), .ZN(n8478) );
  INV_X1 U5786 ( .A(n8464), .ZN(n8412) );
  INV_X1 U5787 ( .A(n8478), .ZN(n8456) );
  NAND2_X1 U5788 ( .A1(n6557), .A2(n9793), .ZN(n8455) );
  NAND2_X1 U5789 ( .A1(n8268), .A2(n8267), .ZN(n8275) );
  OAI21_X1 U5790 ( .B1(n6312), .B2(n4684), .A(n4683), .ZN(n6330) );
  NAND2_X1 U5791 ( .A1(n4457), .A2(n4689), .ZN(n4684) );
  NAND2_X1 U5792 ( .A1(n6356), .A2(n6761), .ZN(n4649) );
  INV_X1 U5793 ( .A(n8328), .ZN(n8589) );
  INV_X1 U5794 ( .A(n8604), .ZN(n8572) );
  INV_X1 U5795 ( .A(n8400), .ZN(n8624) );
  OR2_X1 U5796 ( .A1(n6762), .A2(n9833), .ZN(n8491) );
  INV_X1 U5797 ( .A(n8425), .ZN(n8743) );
  CLKBUF_X1 U5798 ( .A(n7019), .Z(n8506) );
  INV_X1 U5799 ( .A(n4636), .ZN(n6844) );
  INV_X1 U5800 ( .A(n4634), .ZN(n6833) );
  NOR2_X1 U5801 ( .A1(n7858), .A2(n7859), .ZN(n8507) );
  NAND2_X1 U5802 ( .A1(n4622), .A2(n4620), .ZN(n8510) );
  NAND2_X1 U5803 ( .A1(n8513), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5804 ( .A1(n8507), .A2(n4623), .ZN(n4622) );
  INV_X1 U5805 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U5806 ( .A1(n8510), .A2(n8511), .ZN(n8528) );
  NAND2_X1 U5807 ( .A1(n8545), .A2(n4627), .ZN(n4626) );
  INV_X1 U5808 ( .A(n4628), .ZN(n4627) );
  OAI21_X1 U5809 ( .B1(n8547), .B2(n9776), .A(n9777), .ZN(n4628) );
  OAI21_X1 U5810 ( .B1(n8546), .B2(n9778), .A(n4632), .ZN(n4631) );
  NAND2_X1 U5811 ( .A1(n8547), .A2(n9774), .ZN(n4632) );
  NAND2_X1 U5812 ( .A1(n6170), .A2(n6169), .ZN(n8787) );
  AND2_X1 U5813 ( .A1(n6146), .A2(n6145), .ZN(n8556) );
  NAND2_X1 U5814 ( .A1(n8617), .A2(n8292), .ZN(n8596) );
  NAND2_X1 U5815 ( .A1(n6074), .A2(n6073), .ZN(n8810) );
  NAND2_X1 U5816 ( .A1(n4894), .A2(n4895), .ZN(n8634) );
  OR2_X1 U5817 ( .A1(n8290), .A2(n4896), .ZN(n4894) );
  NAND2_X1 U5818 ( .A1(n4898), .A2(n4897), .ZN(n8652) );
  AND2_X1 U5819 ( .A1(n4898), .A2(n4440), .ZN(n8653) );
  NAND2_X1 U5820 ( .A1(n8290), .A2(n8669), .ZN(n4898) );
  NOR2_X1 U5821 ( .A1(n4759), .A2(n4761), .ZN(n4998) );
  NAND2_X1 U5822 ( .A1(n4770), .A2(n6273), .ZN(n8721) );
  NAND2_X1 U5823 ( .A1(n4543), .A2(n4542), .ZN(n8750) );
  NAND2_X1 U5824 ( .A1(n4736), .A2(n4737), .ZN(n8754) );
  NAND2_X1 U5825 ( .A1(n4743), .A2(n6260), .ZN(n8769) );
  NAND2_X1 U5826 ( .A1(n7786), .A2(n7705), .ZN(n8279) );
  NAND2_X1 U5827 ( .A1(n7618), .A2(n6245), .ZN(n7555) );
  NAND2_X1 U5828 ( .A1(n4538), .A2(n7299), .ZN(n7398) );
  NAND2_X1 U5829 ( .A1(n4539), .A2(n4416), .ZN(n4538) );
  INV_X1 U5830 ( .A(n7332), .ZN(n4539) );
  NAND2_X1 U5831 ( .A1(n4748), .A2(n6218), .ZN(n7232) );
  NAND2_X1 U5832 ( .A1(n7071), .A2(n6198), .ZN(n9784) );
  NOR2_X1 U5833 ( .A1(n9844), .A2(n9837), .ZN(n9841) );
  NOR2_X1 U5834 ( .A1(n7041), .A2(n4805), .ZN(n9842) );
  OAI22_X1 U5835 ( .A1(n8748), .A2(n9847), .B1(n8781), .B2(n4805), .ZN(n7043)
         );
  INV_X1 U5836 ( .A(n9793), .ZN(n8778) );
  NAND2_X1 U5837 ( .A1(n9922), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4551) );
  AND2_X1 U5838 ( .A1(n8796), .A2(n8797), .ZN(n4890) );
  NAND2_X1 U5839 ( .A1(n4997), .A2(n4996), .ZN(n4995) );
  NOR2_X1 U5840 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4996) );
  NAND2_X1 U5841 ( .A1(n6349), .A2(n4826), .ZN(n7816) );
  INV_X1 U5842 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10031) );
  XNOR2_X1 U5843 ( .A(n6345), .B(n6344), .ZN(n7726) );
  INV_X1 U5844 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U5845 ( .A1(n6343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6345) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9970) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U5848 ( .A1(n5765), .A2(n5764), .ZN(n5770) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7158) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7154) );
  INV_X1 U5851 ( .A(n7848), .ZN(n7845) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6925) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6868) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10188) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6662) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6654) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10204) );
  OR2_X1 U5858 ( .A1(n5719), .A2(n6611), .ZN(n6683) );
  NAND2_X1 U5859 ( .A1(n4946), .A2(n5380), .ZN(n7975) );
  OR2_X1 U5860 ( .A1(n7894), .A2(n5381), .ZN(n4946) );
  OR2_X1 U5861 ( .A1(n5128), .A2(n6631), .ZN(n5134) );
  AND2_X1 U5862 ( .A1(n6367), .A2(n6366), .ZN(n6593) );
  INV_X1 U5863 ( .A(n9500), .ZN(n9003) );
  OR2_X1 U5864 ( .A1(n7894), .A2(n4940), .ZN(n4933) );
  NAND2_X1 U5865 ( .A1(n4912), .A2(n5189), .ZN(n6618) );
  INV_X1 U5866 ( .A(n4913), .ZN(n4912) );
  OR2_X1 U5867 ( .A1(n5749), .A2(n4378), .ZN(n9503) );
  INV_X1 U5868 ( .A(n7476), .ZN(n9576) );
  NAND2_X1 U5869 ( .A1(n5329), .A2(n5328), .ZN(n7729) );
  INV_X1 U5870 ( .A(n9503), .ZN(n9005) );
  NAND2_X1 U5871 ( .A1(n8940), .A2(n4921), .ZN(n4920) );
  NOR2_X1 U5872 ( .A1(n5744), .A2(n5727), .ZN(n9016) );
  INV_X1 U5873 ( .A(n9020), .ZN(n9038) );
  NAND2_X1 U5874 ( .A1(n4935), .A2(n4947), .ZN(n9028) );
  NAND2_X1 U5875 ( .A1(n7894), .A2(n4950), .ZN(n4935) );
  INV_X1 U5876 ( .A(n9016), .ZN(n9509) );
  OR2_X1 U5877 ( .A1(n6946), .A2(n5080), .ZN(n8260) );
  OR2_X1 U5878 ( .A1(n9215), .A2(n5581), .ZN(n5743) );
  NAND2_X1 U5879 ( .A1(n7995), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5880 ( .A1(n9592), .A2(n6713), .ZN(n9066) );
  NOR2_X1 U5881 ( .A1(n6741), .A2(n4591), .ZN(n6744) );
  NOR2_X1 U5882 ( .A1(n6747), .A2(n6718), .ZN(n4591) );
  NAND2_X1 U5883 ( .A1(n6744), .A2(n6743), .ZN(n6871) );
  AOI21_X1 U5884 ( .B1(n8888), .B2(n8035), .A(n8034), .ZN(n9129) );
  INV_X1 U5885 ( .A(n9380), .ZN(n9180) );
  NAND2_X1 U5886 ( .A1(n9174), .A2(n9173), .ZN(n9382) );
  NAND2_X1 U5887 ( .A1(n9169), .A2(n9189), .ZN(n9174) );
  NAND2_X1 U5888 ( .A1(n4553), .A2(n4552), .ZN(n9148) );
  NAND2_X1 U5889 ( .A1(n4432), .A2(n4417), .ZN(n4552) );
  NAND2_X1 U5890 ( .A1(n9195), .A2(n9194), .ZN(n9386) );
  NOR2_X1 U5891 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  NOR2_X1 U5892 ( .A1(n4556), .A2(n4432), .ZN(n9185) );
  NAND2_X1 U5893 ( .A1(n4560), .A2(n4558), .ZN(n9186) );
  INV_X1 U5894 ( .A(n4556), .ZN(n4560) );
  OAI21_X1 U5895 ( .B1(n9297), .B2(n4706), .A(n4703), .ZN(n9259) );
  NAND2_X1 U5896 ( .A1(n4709), .A2(n9155), .ZN(n9270) );
  NAND2_X1 U5897 ( .A1(n9297), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U5898 ( .A1(n4788), .A2(n4790), .ZN(n9268) );
  OR2_X1 U5899 ( .A1(n9308), .A2(n4792), .ZN(n4788) );
  NAND2_X1 U5900 ( .A1(n9297), .A2(n9154), .ZN(n9291) );
  AND2_X1 U5901 ( .A1(n4794), .A2(n4427), .ZN(n9282) );
  AND2_X1 U5902 ( .A1(n4717), .A2(n4716), .ZN(n9321) );
  NAND2_X1 U5903 ( .A1(n9150), .A2(n9149), .ZN(n9332) );
  NAND2_X1 U5904 ( .A1(n5491), .A2(n5490), .ZN(n9437) );
  OAI21_X1 U5905 ( .B1(n7668), .B2(n4413), .A(n4723), .ZN(n7916) );
  NAND2_X1 U5906 ( .A1(n7746), .A2(n8062), .ZN(n7805) );
  AND2_X1 U5907 ( .A1(n7260), .A2(n8096), .ZN(n7368) );
  NAND2_X1 U5908 ( .A1(n9692), .A2(n5008), .ZN(n9694) );
  INV_X1 U5909 ( .A(n9722), .ZN(n9668) );
  AND2_X1 U5910 ( .A1(n8260), .A2(n7169), .ZN(n9675) );
  OR2_X1 U5911 ( .A1(n7676), .A2(n9753), .ZN(n9176) );
  INV_X1 U5912 ( .A(n5092), .ZN(n5097) );
  OR2_X1 U5913 ( .A1(n7109), .A2(n8259), .ZN(n9693) );
  INV_X1 U5914 ( .A(n9694), .ZN(n9309) );
  AND2_X2 U5915 ( .A1(n6694), .A2(n7106), .ZN(n9759) );
  AND2_X1 U5916 ( .A1(n7811), .A2(n5704), .ZN(n6646) );
  AND2_X1 U5917 ( .A1(n7811), .A2(n7720), .ZN(n6668) );
  AND2_X1 U5918 ( .A1(n5719), .A2(n5723), .ZN(n6647) );
  INV_X1 U5919 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U5920 ( .A1(n9472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5035) );
  NOR2_X1 U5921 ( .A1(n5065), .A2(n5028), .ZN(n5030) );
  AND2_X1 U5922 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5028) );
  XNOR2_X1 U5923 ( .A(n6125), .B(n6124), .ZN(n7879) );
  NAND2_X1 U5924 ( .A1(n6109), .A2(n6108), .ZN(n6125) );
  XNOR2_X1 U5925 ( .A(n6107), .B(n6106), .ZN(n7839) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7944) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9958) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10022) );
  AND2_X1 U5929 ( .A1(n4397), .A2(P1_U3084), .ZN(n7878) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7642) );
  CLKBUF_X1 U5931 ( .A(n5724), .Z(n5725) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7506) );
  INV_X1 U5933 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7435) );
  INV_X1 U5934 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5077) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10235) );
  INV_X1 U5936 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10112) );
  INV_X1 U5937 ( .A(n7688), .ZN(n7694) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6870) );
  INV_X1 U5939 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6679) );
  INV_X1 U5940 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6650) );
  INV_X1 U5941 ( .A(n4866), .ZN(n5004) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U5943 ( .A1(n5125), .A2(n4597), .ZN(n9587) );
  NAND2_X1 U5944 ( .A1(n4596), .A2(n4594), .ZN(n4597) );
  NOR2_X1 U5945 ( .A1(n5102), .A2(n4595), .ZN(n4594) );
  NOR2_X1 U5946 ( .A1(n7773), .A2(n10263), .ZN(n9952) );
  AOI21_X1 U5947 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9950), .ZN(n9949) );
  NOR2_X1 U5948 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  AOI21_X1 U5949 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9947), .ZN(n9946) );
  OAI21_X1 U5950 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9944), .ZN(n9942) );
  NOR2_X1 U5951 ( .A1(n9940), .A2(n9939), .ZN(n9938) );
  NAND2_X1 U5952 ( .A1(n4629), .A2(n4624), .ZN(P2_U3264) );
  AOI21_X1 U5953 ( .B1(n4631), .B2(n4410), .A(n4630), .ZN(n4629) );
  NAND2_X1 U5954 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5955 ( .A(n8549), .ZN(n4630) );
  AOI211_X1 U5956 ( .C1(n8795), .C2(n9521), .A(n8308), .B(n8307), .ZN(n8309)
         );
  OAI21_X1 U5957 ( .B1(n8802), .B2(n9808), .A(n4773), .ZN(n4772) );
  AOI21_X1 U5958 ( .B1(n8800), .B2(n9521), .A(n8573), .ZN(n4773) );
  OAI21_X1 U5959 ( .B1(n8798), .B2(n4550), .A(n4548), .ZN(P2_U3549) );
  NAND2_X1 U5960 ( .A1(n9924), .A2(n9904), .ZN(n4550) );
  INV_X1 U5961 ( .A(n4549), .ZN(n4548) );
  OAI21_X1 U5962 ( .B1(n4890), .B2(n9922), .A(n4551), .ZN(n4549) );
  NAND2_X1 U5963 ( .A1(n4889), .A2(n4888), .ZN(P2_U3517) );
  NAND2_X1 U5964 ( .A1(n9906), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5965 ( .A1(n8873), .A2(n9908), .ZN(n4889) );
  OAI21_X1 U5966 ( .B1(n8798), .B2(n9871), .A(n4890), .ZN(n8873) );
  NAND2_X1 U5967 ( .A1(n4730), .A2(n4479), .ZN(P1_U3519) );
  NAND2_X1 U5968 ( .A1(n9458), .A2(n9759), .ZN(n4730) );
  INV_X1 U5969 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5970 ( .A1(n4789), .A2(n9143), .ZN(n4411) );
  AND2_X1 U5971 ( .A1(n6298), .A2(n6297), .ZN(n4412) );
  INV_X1 U5972 ( .A(n6327), .ZN(n6316) );
  AND2_X2 U5973 ( .A1(n6946), .A2(n5080), .ZN(n6362) );
  OR2_X1 U5974 ( .A1(n4725), .A2(n8133), .ZN(n4413) );
  INV_X1 U5975 ( .A(n9152), .ZN(n4715) );
  INV_X1 U5976 ( .A(n5380), .ZN(n4951) );
  INV_X1 U5977 ( .A(n8505), .ZN(n4752) );
  NOR2_X1 U5978 ( .A1(n7914), .A2(n8028), .ZN(n4415) );
  OR2_X1 U5979 ( .A1(n8503), .A2(n7298), .ZN(n4416) );
  INV_X1 U5980 ( .A(n8282), .ZN(n8772) );
  INV_X1 U5981 ( .A(n9329), .ZN(n4720) );
  NAND2_X1 U5982 ( .A1(n9388), .A2(n9210), .ZN(n4417) );
  AND2_X1 U5983 ( .A1(n4790), .A2(n4589), .ZN(n4418) );
  AND2_X1 U5984 ( .A1(n5764), .A2(n5771), .ZN(n4419) );
  NAND2_X1 U5985 ( .A1(n4919), .A2(n4442), .ZN(n6379) );
  NAND2_X1 U5986 ( .A1(n6250), .A2(n7554), .ZN(n7615) );
  INV_X1 U5987 ( .A(n7615), .ZN(n4899) );
  AND4_X1 U5988 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8381)
         );
  INV_X1 U5989 ( .A(n8381), .ZN(n4900) );
  INV_X1 U5990 ( .A(n8677), .ZN(n8669) );
  AND2_X1 U5991 ( .A1(n6265), .A2(n6264), .ZN(n8282) );
  AOI21_X1 U5992 ( .B1(n4793), .B2(n4791), .A(n4461), .ZN(n4790) );
  AND2_X1 U5993 ( .A1(n4892), .A2(n8291), .ZN(n4420) );
  NOR2_X1 U5994 ( .A1(n4744), .A2(n5015), .ZN(n4542) );
  NOR2_X1 U5995 ( .A1(n8421), .A2(n4978), .ZN(n4421) );
  AND2_X1 U5996 ( .A1(n5778), .A2(n4825), .ZN(n4422) );
  AND2_X1 U5997 ( .A1(n6318), .A2(n6317), .ZN(n4423) );
  OR2_X1 U5998 ( .A1(n7572), .A2(n4608), .ZN(n4424) );
  OR2_X1 U5999 ( .A1(n9519), .A2(n4810), .ZN(n4425) );
  INV_X1 U6000 ( .A(n9155), .ZN(n4708) );
  INV_X1 U6001 ( .A(n9246), .ZN(n9213) );
  NAND2_X1 U6002 ( .A1(n5694), .A2(n5693), .ZN(n9246) );
  XNOR2_X1 U6003 ( .A(n5075), .B(n10177), .ZN(n9376) );
  NAND2_X1 U6004 ( .A1(n5924), .A2(n5923), .ZN(n8388) );
  INV_X1 U6005 ( .A(n8388), .ZN(n4806) );
  AND2_X1 U6006 ( .A1(n5779), .A2(n4422), .ZN(n6348) );
  INV_X1 U6007 ( .A(n6348), .ZN(n4826) );
  INV_X1 U6008 ( .A(n6356), .ZN(n4651) );
  OR2_X1 U6009 ( .A1(n5720), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6010 ( .A1(n9422), .A2(n9323), .ZN(n4427) );
  NAND2_X1 U6011 ( .A1(n5294), .A2(n4397), .ZN(n5128) );
  AND2_X1 U6012 ( .A1(n8696), .A2(n6042), .ZN(n4428) );
  INV_X1 U6013 ( .A(n9146), .ZN(n4509) );
  NAND2_X1 U6014 ( .A1(n5539), .A2(n5538), .ZN(n9427) );
  NAND2_X1 U6015 ( .A1(n5414), .A2(n5413), .ZN(n9453) );
  AND2_X1 U6016 ( .A1(n6255), .A2(n6249), .ZN(n7783) );
  INV_X1 U6017 ( .A(n7783), .ZN(n7704) );
  NAND2_X1 U6018 ( .A1(n9442), .A2(n9042), .ZN(n4429) );
  NAND4_X1 U6019 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n9054)
         );
  INV_X1 U6020 ( .A(n9054), .ZN(n9686) );
  AND2_X1 U6021 ( .A1(n8184), .A2(n9380), .ZN(n4430) );
  AND2_X1 U6022 ( .A1(n4720), .A2(n9149), .ZN(n4431) );
  OR2_X1 U6023 ( .A1(n9187), .A2(n4557), .ZN(n4432) );
  NOR2_X1 U6024 ( .A1(n7476), .A2(n9046), .ZN(n4433) );
  XNOR2_X1 U6025 ( .A(n5030), .B(n5029), .ZN(n5038) );
  NAND2_X1 U6026 ( .A1(n7400), .A2(n7964), .ZN(n4434) );
  NOR2_X1 U6027 ( .A1(n6322), .A2(n6324), .ZN(n4435) );
  NAND2_X1 U6028 ( .A1(n8289), .A2(n8288), .ZN(n8668) );
  INV_X1 U6029 ( .A(n4929), .ZN(n5215) );
  INV_X1 U6030 ( .A(n9157), .ZN(n4704) );
  OR2_X1 U6031 ( .A1(n5294), .A2(n6737), .ZN(n4436) );
  OR2_X1 U6032 ( .A1(n8158), .A2(n9152), .ZN(n4437) );
  NAND2_X1 U6033 ( .A1(n4975), .A2(n4976), .ZN(n8476) );
  NAND2_X1 U6034 ( .A1(n5390), .A2(n5389), .ZN(n7982) );
  OR3_X1 U6035 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4438) );
  OAI21_X1 U6036 ( .B1(n8617), .B2(n8599), .A(n4886), .ZN(n8575) );
  AND2_X1 U6037 ( .A1(n7905), .A2(n9364), .ZN(n4439) );
  OR2_X1 U6038 ( .A1(n8832), .A2(n8698), .ZN(n4440) );
  AND3_X1 U6039 ( .A1(n4493), .A2(n4492), .A3(n4489), .ZN(n4441) );
  AND2_X1 U6040 ( .A1(n9162), .A2(n8178), .ZN(n9208) );
  INV_X1 U6041 ( .A(n9208), .ZN(n4510) );
  NOR3_X1 U6042 ( .A1(n9283), .A2(n9397), .A3(n4612), .ZN(n4609) );
  NAND2_X1 U6043 ( .A1(n8596), .A2(n8595), .ZN(n8594) );
  NAND2_X1 U6044 ( .A1(n5020), .A2(n5019), .ZN(n5196) );
  OR2_X1 U6045 ( .A1(n9788), .A2(n7224), .ZN(n6198) );
  INV_X1 U6046 ( .A(n6198), .ZN(n4749) );
  NAND2_X1 U6047 ( .A1(n5623), .A2(n5622), .ZN(n9406) );
  NAND2_X1 U6048 ( .A1(n6025), .A2(n6024), .ZN(n8837) );
  AND2_X1 U6049 ( .A1(n5702), .A2(n4920), .ZN(n4442) );
  INV_X1 U6050 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U6051 ( .A1(n4915), .A2(n5642), .ZN(n8939) );
  AND2_X1 U6052 ( .A1(n4822), .A2(n8641), .ZN(n4443) );
  NOR2_X1 U6053 ( .A1(n5594), .A2(n5595), .ZN(n4444) );
  AND2_X1 U6054 ( .A1(n6296), .A2(n6297), .ZN(n8642) );
  INV_X1 U6055 ( .A(n8642), .ZN(n8633) );
  AND3_X1 U6056 ( .A1(n6254), .A2(n6253), .A3(n6316), .ZN(n4445) );
  AND2_X1 U6057 ( .A1(n4656), .A2(n4658), .ZN(n4446) );
  AND2_X1 U6058 ( .A1(n8827), .A2(n8492), .ZN(n4447) );
  AND2_X1 U6059 ( .A1(n6279), .A2(n8710), .ZN(n8284) );
  INV_X1 U6060 ( .A(n8284), .ZN(n4771) );
  OR2_X1 U6061 ( .A1(n7913), .A2(n8028), .ZN(n4448) );
  OR2_X1 U6062 ( .A1(n4708), .A2(n8158), .ZN(n4449) );
  INV_X1 U6063 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5771) );
  INV_X1 U6064 ( .A(n5429), .ZN(n4954) );
  OR2_X1 U6065 ( .A1(n6717), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4450) );
  AND2_X1 U6066 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4451) );
  NOR2_X1 U6067 ( .A1(n8277), .A2(n8496), .ZN(n4452) );
  NOR2_X1 U6068 ( .A1(n5475), .A2(n8960), .ZN(n4453) );
  INV_X1 U6069 ( .A(n4937), .ZN(n4936) );
  OAI21_X1 U6070 ( .B1(n4941), .B2(n4945), .A(n4938), .ZN(n4937) );
  AND4_X1 U6071 ( .A1(n10082), .A2(n5025), .A3(n5721), .A4(n5051), .ZN(n4454)
         );
  AND2_X1 U6072 ( .A1(n4527), .A2(n4449), .ZN(n4455) );
  INV_X1 U6073 ( .A(n4577), .ZN(n4576) );
  OR2_X1 U6074 ( .A1(n7740), .A2(n4578), .ZN(n4577) );
  NAND2_X1 U6075 ( .A1(n4434), .A2(n4416), .ZN(n4456) );
  NOR2_X1 U6076 ( .A1(n4435), .A2(n4687), .ZN(n4457) );
  NAND2_X1 U6077 ( .A1(n5765), .A2(n4419), .ZN(n4458) );
  AND2_X1 U6078 ( .A1(n5201), .A2(SI_5_), .ZN(n4459) );
  INV_X1 U6079 ( .A(n4891), .ZN(n4893) );
  NAND2_X1 U6080 ( .A1(n4895), .A2(n8633), .ZN(n4891) );
  INV_X1 U6081 ( .A(n5000), .ZN(n4590) );
  OR2_X1 U6082 ( .A1(n9279), .A2(n9294), .ZN(n5000) );
  NAND2_X1 U6083 ( .A1(n6310), .A2(n6309), .ZN(n4460) );
  NOR2_X1 U6084 ( .A1(n9285), .A2(n9272), .ZN(n4461) );
  OAI21_X1 U6085 ( .B1(n4435), .B2(n4686), .A(n6326), .ZN(n4685) );
  NAND2_X1 U6086 ( .A1(n4952), .A2(n5431), .ZN(n4462) );
  NAND2_X1 U6087 ( .A1(n9187), .A2(n8179), .ZN(n4463) );
  OR2_X1 U6088 ( .A1(n7905), .A2(n7798), .ZN(n8137) );
  AND2_X1 U6089 ( .A1(n4737), .A2(n4744), .ZN(n4464) );
  NAND2_X1 U6090 ( .A1(n5515), .A2(n5514), .ZN(n9434) );
  OR2_X1 U6091 ( .A1(n9417), .A2(n9272), .ZN(n9155) );
  AND2_X1 U6092 ( .A1(n4554), .A2(n4417), .ZN(n4465) );
  INV_X1 U6093 ( .A(n7205), .ZN(n4582) );
  NOR2_X1 U6094 ( .A1(n8278), .A2(n4905), .ZN(n4904) );
  AND2_X1 U6095 ( .A1(n4430), .A2(n4506), .ZN(n4466) );
  AND2_X1 U6096 ( .A1(n8107), .A2(n7381), .ZN(n8018) );
  INV_X1 U6097 ( .A(n4782), .ZN(n4781) );
  NOR2_X1 U6098 ( .A1(n5362), .A2(n4783), .ZN(n4782) );
  AND2_X1 U6099 ( .A1(n4431), .A2(n4715), .ZN(n4467) );
  AND2_X1 U6100 ( .A1(n4412), .A2(n4446), .ZN(n4468) );
  NAND2_X1 U6101 ( .A1(n4412), .A2(n6299), .ZN(n4469) );
  INV_X1 U6102 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5042) );
  OR2_X1 U6103 ( .A1(n9122), .A2(n9121), .ZN(P1_U3260) );
  INV_X1 U6104 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U6105 ( .A1(n6176), .A2(n6203), .ZN(n7018) );
  AND2_X1 U6106 ( .A1(n7530), .A2(n7529), .ZN(n7547) );
  INV_X1 U6107 ( .A(n6251), .ZN(n4764) );
  INV_X1 U6108 ( .A(n6135), .ZN(n6117) );
  NOR2_X1 U6109 ( .A1(n8799), .A2(n8589), .ZN(n4471) );
  INV_X1 U6110 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U6111 ( .B1(n6108), .B2(n4847), .A(n6128), .ZN(n4846) );
  NAND2_X1 U6112 ( .A1(n4933), .A2(n4936), .ZN(n8947) );
  INV_X1 U6113 ( .A(n8753), .ZN(n4744) );
  NAND2_X1 U6114 ( .A1(n7598), .A2(n5287), .ZN(n7627) );
  NAND2_X1 U6115 ( .A1(n4699), .A2(n8057), .ZN(n7566) );
  AND2_X1 U6116 ( .A1(n4909), .A2(n4910), .ZN(n8917) );
  NAND2_X1 U6117 ( .A1(n7664), .A2(n7663), .ZN(n7741) );
  INV_X1 U6118 ( .A(n9330), .ZN(n4719) );
  INV_X1 U6119 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U6120 ( .A1(n4575), .A2(n7739), .ZN(n7912) );
  INV_X1 U6121 ( .A(n5642), .ZN(n4921) );
  INV_X1 U6122 ( .A(n4707), .ZN(n4706) );
  NOR3_X1 U6123 ( .A1(n9519), .A2(n8849), .A3(n4811), .ZN(n4808) );
  OR2_X1 U6124 ( .A1(n8842), .A2(n8373), .ZN(n6284) );
  INV_X1 U6125 ( .A(n6284), .ZN(n4761) );
  INV_X1 U6126 ( .A(n4605), .ZN(n7800) );
  NOR3_X1 U6127 ( .A1(n7572), .A2(n9453), .A3(n4608), .ZN(n4605) );
  NOR2_X1 U6128 ( .A1(n8852), .A2(n8493), .ZN(n4472) );
  NOR2_X1 U6129 ( .A1(n7572), .A2(n4606), .ZN(n7928) );
  INV_X1 U6130 ( .A(n8804), .ZN(n8584) );
  NAND2_X1 U6131 ( .A1(n6095), .A2(n6094), .ZN(n8804) );
  INV_X1 U6132 ( .A(n8295), .ZN(n8860) );
  NAND2_X1 U6133 ( .A1(n5985), .A2(n5984), .ZN(n8295) );
  INV_X1 U6134 ( .A(n4543), .ZN(n8771) );
  NAND2_X1 U6135 ( .A1(n8773), .A2(n8772), .ZN(n4543) );
  AND2_X1 U6136 ( .A1(n8572), .A2(n9787), .ZN(n4473) );
  NOR2_X1 U6137 ( .A1(n8295), .A2(n8742), .ZN(n4474) );
  INV_X1 U6138 ( .A(n4809), .ZN(n8736) );
  NOR2_X1 U6139 ( .A1(n9519), .A2(n4811), .ZN(n4809) );
  INV_X1 U6140 ( .A(n4610), .ZN(n9236) );
  NOR2_X1 U6141 ( .A1(n9283), .A2(n4612), .ZN(n4610) );
  INV_X1 U6142 ( .A(n9397), .ZN(n9232) );
  NAND2_X1 U6143 ( .A1(n5682), .A2(n5681), .ZN(n9397) );
  NOR2_X1 U6144 ( .A1(n8810), .A2(n8624), .ZN(n4475) );
  AND2_X1 U6145 ( .A1(n4934), .A2(n4944), .ZN(n4476) );
  NAND2_X1 U6146 ( .A1(n9523), .A2(n8281), .ZN(n8770) );
  OR2_X1 U6147 ( .A1(n9308), .A2(n9307), .ZN(n4794) );
  INV_X1 U6148 ( .A(n4423), .ZN(n4692) );
  OR2_X1 U6149 ( .A1(n4929), .A2(n4928), .ZN(n4477) );
  XNOR2_X1 U6150 ( .A(n5053), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5717) );
  NOR2_X1 U6151 ( .A1(n7621), .A2(n8449), .ZN(n4807) );
  INV_X2 U6152 ( .A(n9906), .ZN(n9908) );
  AND2_X1 U6153 ( .A1(n7499), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U6154 ( .A1(n4913), .A2(n5189), .ZN(n9011) );
  NAND2_X1 U6155 ( .A1(n7206), .A2(n7205), .ZN(n7266) );
  INV_X1 U6156 ( .A(n8359), .ZN(n4978) );
  NAND2_X1 U6157 ( .A1(n6358), .A2(n6357), .ZN(n9392) );
  INV_X1 U6158 ( .A(n9392), .ZN(n4559) );
  XNOR2_X1 U6159 ( .A(n5052), .B(n5051), .ZN(n5704) );
  OAI21_X1 U6160 ( .B1(n7332), .B2(n4456), .A(n4536), .ZN(n7946) );
  AOI21_X1 U6161 ( .B1(n7394), .B2(n7366), .A(n7365), .ZN(n7367) );
  NAND2_X1 U6162 ( .A1(n5186), .A2(n5189), .ZN(n6615) );
  INV_X1 U6163 ( .A(n7294), .ZN(n4821) );
  NOR2_X1 U6164 ( .A1(n7985), .A2(n7986), .ZN(n7009) );
  INV_X1 U6165 ( .A(n9795), .ZN(n4819) );
  NAND2_X1 U6166 ( .A1(n5912), .A2(n5911), .ZN(n8449) );
  INV_X1 U6167 ( .A(n8449), .ZN(n4901) );
  AND2_X1 U6168 ( .A1(n8212), .A2(n8214), .ZN(n8010) );
  INV_X1 U6169 ( .A(n8010), .ZN(n4568) );
  OAI21_X1 U6170 ( .B1(n7009), .B2(n7011), .A(n7010), .ZN(n7008) );
  OR2_X1 U6171 ( .A1(n9759), .A2(n4729), .ZN(n4479) );
  XNOR2_X1 U6172 ( .A(n6407), .B(n6408), .ZN(n6973) );
  AND2_X1 U6173 ( .A1(n8774), .A2(n9890), .ZN(n9871) );
  AND2_X1 U6174 ( .A1(n7039), .A2(n7020), .ZN(n4480) );
  INV_X1 U6175 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4988) );
  INV_X1 U6176 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5781) );
  INV_X1 U6177 ( .A(n9851), .ZN(n4751) );
  INV_X1 U6178 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5070) );
  INV_X1 U6179 ( .A(n9305), .ZN(n9670) );
  XNOR2_X1 U6180 ( .A(n5078), .B(n5077), .ZN(n9305) );
  NOR2_X1 U6181 ( .A1(n6346), .A2(n4995), .ZN(n8889) );
  NAND2_X1 U6182 ( .A1(n9483), .A2(n9482), .ZN(n4645) );
  AND2_X1 U6183 ( .A1(n5971), .A2(n5982), .ZN(n8508) );
  INV_X1 U6184 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4803) );
  INV_X1 U6185 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n4754) );
  INV_X2 U6186 ( .A(n9791), .ZN(n9808) );
  NAND2_X1 U6187 ( .A1(n7029), .A2(n9793), .ZN(n9791) );
  MUX2_X1 U6188 ( .A(n8190), .B(n8189), .S(n8188), .Z(n8197) );
  INV_X1 U6189 ( .A(n8188), .ZN(n4535) );
  OR2_X1 U6190 ( .A1(n8120), .A2(n8188), .ZN(n4499) );
  NAND2_X1 U6191 ( .A1(n8130), .A2(n8188), .ZN(n4492) );
  NOR2_X1 U6192 ( .A1(n4491), .A2(n8188), .ZN(n4490) );
  AOI21_X1 U6193 ( .B1(n4498), .B2(n8188), .A(n4497), .ZN(n4496) );
  INV_X1 U6194 ( .A(n5765), .ZN(n5993) );
  NAND2_X1 U6195 ( .A1(n8757), .A2(n6266), .ZN(n8741) );
  NAND2_X1 U6196 ( .A1(n4647), .A2(n4649), .ZN(n4646) );
  NAND4_X2 U6197 ( .A1(n5806), .A2(n5808), .A3(n5807), .A4(n4753), .ZN(n8505)
         );
  AND2_X2 U6198 ( .A1(n4975), .A2(n4973), .ZN(n8477) );
  NOR2_X1 U6199 ( .A1(n4481), .A2(n8205), .ZN(n8265) );
  NAND2_X1 U6200 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  AOI21_X1 U6201 ( .B1(n8202), .B2(n9305), .A(n5728), .ZN(n4482) );
  NAND2_X1 U6202 ( .A1(n4484), .A2(n9670), .ZN(n4483) );
  NAND2_X1 U6203 ( .A1(n4485), .A2(n8201), .ZN(n4484) );
  NAND2_X1 U6204 ( .A1(n8204), .A2(n5001), .ZN(n4485) );
  XNOR2_X1 U6205 ( .A(n5105), .B(n5095), .ZN(n5104) );
  NAND2_X1 U6206 ( .A1(n4500), .A2(n5094), .ZN(n5105) );
  OAI21_X1 U6207 ( .B1(n8177), .B2(n4511), .A(n4466), .ZN(n4515) );
  NAND2_X1 U6208 ( .A1(n8153), .A2(n8188), .ZN(n4533) );
  NAND2_X1 U6209 ( .A1(n8154), .A2(n4535), .ZN(n4534) );
  NOR2_X4 U6210 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5810) );
  NAND2_X1 U6211 ( .A1(n7067), .A2(n7066), .ZN(n7223) );
  NAND2_X1 U6212 ( .A1(n7223), .A2(n7222), .ZN(n7227) );
  AND2_X2 U6213 ( .A1(n6348), .A2(n5780), .ZN(n5790) );
  NAND2_X1 U6214 ( .A1(n8770), .A2(n4542), .ZN(n4540) );
  NAND2_X1 U6215 ( .A1(n4540), .A2(n4541), .ZN(n8735) );
  NOR2_X1 U6216 ( .A1(n8771), .A2(n5015), .ZN(n8749) );
  NAND2_X1 U6217 ( .A1(n8562), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U6218 ( .A1(n4562), .A2(n4465), .ZN(n4553) );
  AND2_X1 U6219 ( .A1(n4562), .A2(n4554), .ZN(n4556) );
  NAND2_X1 U6220 ( .A1(n4562), .A2(n4561), .ZN(n9206) );
  NAND2_X1 U6221 ( .A1(n4567), .A2(n4569), .ZN(n9681) );
  NAND2_X1 U6222 ( .A1(n7171), .A2(n4565), .ZN(n4564) );
  INV_X1 U6223 ( .A(n7171), .ZN(n4566) );
  NAND3_X1 U6224 ( .A1(n7112), .A2(n4568), .A3(n6945), .ZN(n4567) );
  NAND2_X1 U6225 ( .A1(n7664), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U6226 ( .A1(n7168), .A2(n7205), .ZN(n4579) );
  NAND2_X1 U6227 ( .A1(n4580), .A2(n4579), .ZN(n7268) );
  NOR2_X1 U6228 ( .A1(n4585), .A2(n4584), .ZN(n9251) );
  NAND3_X1 U6229 ( .A1(n5101), .A2(n5102), .A3(n5018), .ZN(n5171) );
  INV_X1 U6230 ( .A(n4601), .ZN(n9302) );
  INV_X1 U6231 ( .A(n4609), .ZN(n9228) );
  NAND4_X1 U6232 ( .A1(n5070), .A2(n10177), .A3(n5438), .A4(n5042), .ZN(n4614)
         );
  NAND4_X1 U6233 ( .A1(n4617), .A2(n4616), .A3(n5071), .A4(n5486), .ZN(n4615)
         );
  INV_X1 U6234 ( .A(n4643), .ZN(n6813) );
  NAND2_X1 U6235 ( .A1(n6789), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U6236 ( .A1(n4648), .A2(n4646), .ZN(P2_U3244) );
  NAND2_X1 U6237 ( .A1(n6334), .A2(n6341), .ZN(n4648) );
  NAND2_X1 U6238 ( .A1(n4652), .A2(n4655), .ZN(n6305) );
  NAND3_X1 U6239 ( .A1(n4653), .A2(n4468), .A3(n4654), .ZN(n4652) );
  OR2_X1 U6240 ( .A1(n6278), .A2(n4660), .ZN(n4653) );
  OAI21_X1 U6241 ( .B1(n4665), .B2(n4445), .A(n4670), .ZN(n6259) );
  NOR2_X2 U6242 ( .A1(n4735), .A2(n5761), .ZN(n4804) );
  NAND3_X1 U6243 ( .A1(n6263), .A2(n6262), .A3(n8282), .ZN(n4677) );
  NAND2_X1 U6244 ( .A1(n5765), .A2(n4679), .ZN(n4678) );
  INV_X1 U6245 ( .A(n7222), .ZN(n4695) );
  MUX2_X1 U6246 ( .A(n6196), .B(n6197), .S(n6327), .Z(n6216) );
  NAND2_X1 U6247 ( .A1(n4699), .A2(n4697), .ZN(n7567) );
  INV_X1 U6248 ( .A(n4700), .ZN(n9258) );
  NAND2_X1 U6249 ( .A1(n7382), .A2(n8108), .ZN(n7452) );
  NAND2_X1 U6250 ( .A1(n9150), .A2(n4467), .ZN(n4714) );
  NAND2_X1 U6251 ( .A1(n7668), .A2(n4723), .ZN(n4721) );
  NAND2_X1 U6252 ( .A1(n4721), .A2(n4722), .ZN(n7917) );
  OAI21_X1 U6253 ( .B1(n4727), .B2(n4726), .A(n8009), .ZN(n7213) );
  AND2_X1 U6254 ( .A1(n7246), .A2(n8012), .ZN(n4726) );
  OAI21_X1 U6255 ( .B1(n7246), .B2(n7173), .A(n8012), .ZN(n7208) );
  NAND2_X1 U6256 ( .A1(n8223), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U6257 ( .A1(n7173), .A2(n8012), .ZN(n4728) );
  NAND2_X1 U6258 ( .A1(n7568), .A2(n8023), .ZN(n7668) );
  NAND2_X1 U6259 ( .A1(n7172), .A2(n8217), .ZN(n7246) );
  NAND2_X1 U6260 ( .A1(n9207), .A2(n9162), .ZN(n9188) );
  NAND2_X1 U6261 ( .A1(n7917), .A2(n8069), .ZN(n9362) );
  NAND2_X1 U6262 ( .A1(n9258), .A2(n9159), .ZN(n9222) );
  OAI21_X1 U6263 ( .B1(n7174), .B2(n9659), .A(n8013), .ZN(n8102) );
  NOR2_X1 U6264 ( .A1(n8197), .A2(n8196), .ZN(n8204) );
  NAND2_X1 U6265 ( .A1(n4803), .A2(n4802), .ZN(n4799) );
  INV_X1 U6266 ( .A(n5198), .ZN(n4829) );
  NAND2_X1 U6267 ( .A1(n7211), .A2(n7210), .ZN(n7260) );
  NAND2_X1 U6268 ( .A1(n7567), .A2(n8121), .ZN(n7568) );
  INV_X1 U6269 ( .A(n7213), .ZN(n7211) );
  NAND3_X1 U6270 ( .A1(n4804), .A2(n5777), .A3(n4414), .ZN(n6350) );
  NAND4_X1 U6271 ( .A1(n5759), .A2(n5760), .A3(n5857), .A4(n5758), .ZN(n5761)
         );
  NAND4_X1 U6272 ( .A1(n5810), .A2(n5834), .A3(n4982), .A4(n5762), .ZN(n4735)
         );
  NAND2_X1 U6273 ( .A1(n4736), .A2(n4464), .ZN(n8757) );
  NAND2_X1 U6274 ( .A1(n5826), .A2(n4695), .ZN(n7071) );
  NAND2_X1 U6275 ( .A1(n4752), .A2(n4751), .ZN(n7068) );
  OR2_X1 U6276 ( .A1(n4987), .A2(n4754), .ZN(n4753) );
  OAI21_X2 U6277 ( .B1(n6023), .B2(n4758), .A(n4755), .ZN(n8661) );
  NAND2_X1 U6278 ( .A1(n7531), .A2(n4765), .ZN(n4762) );
  NAND2_X1 U6279 ( .A1(n4762), .A2(n4763), .ZN(n7782) );
  INV_X1 U6280 ( .A(n4772), .ZN(n8574) );
  XNOR2_X1 U6281 ( .A(n8570), .B(n8569), .ZN(n4776) );
  NAND2_X2 U6282 ( .A1(n5783), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4777) );
  NAND3_X1 U6283 ( .A1(n4857), .A2(n4858), .A3(n4782), .ZN(n4778) );
  INV_X1 U6284 ( .A(n4794), .ZN(n9426) );
  NAND3_X1 U6285 ( .A1(n4883), .A2(n4882), .A3(n6650), .ZN(n4800) );
  INV_X1 U6286 ( .A(n4808), .ZN(n8718) );
  NAND2_X1 U6287 ( .A1(n8610), .A2(n4814), .ZN(n4815) );
  NAND2_X1 U6288 ( .A1(n8610), .A2(n4813), .ZN(n8564) );
  NAND2_X1 U6289 ( .A1(n8610), .A2(n8584), .ZN(n8578) );
  NAND3_X1 U6290 ( .A1(n4819), .A2(n9877), .A3(n4818), .ZN(n7955) );
  NAND2_X1 U6291 ( .A1(n5779), .A2(n5778), .ZN(n6346) );
  NAND2_X1 U6292 ( .A1(n4826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5789) );
  MUX2_X1 U6293 ( .A(n6630), .B(n6624), .S(n5093), .Z(n5131) );
  MUX2_X1 U6294 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5093), .Z(n5103) );
  MUX2_X1 U6295 ( .A(n6632), .B(n6626), .S(n5093), .Z(n5155) );
  NAND2_X1 U6296 ( .A1(n5675), .A2(n4835), .ZN(n4833) );
  INV_X1 U6297 ( .A(n4840), .ZN(n6163) );
  NAND2_X1 U6298 ( .A1(n5508), .A2(n4852), .ZN(n4850) );
  NAND2_X1 U6299 ( .A1(n5508), .A2(n4855), .ZN(n4851) );
  INV_X1 U6300 ( .A(n4864), .ZN(n4863) );
  NAND2_X1 U6301 ( .A1(n5264), .A2(n4861), .ZN(n4858) );
  NAND2_X1 U6302 ( .A1(n4864), .A2(n4862), .ZN(n4859) );
  NAND2_X1 U6303 ( .A1(n5384), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U6304 ( .A1(n4867), .A2(n4871), .ZN(n5456) );
  NAND2_X1 U6305 ( .A1(n5218), .A2(n5217), .ZN(n4879) );
  NAND2_X1 U6306 ( .A1(n5154), .A2(n5153), .ZN(n4880) );
  NAND2_X1 U6307 ( .A1(n4881), .A2(n5133), .ZN(n5154) );
  NAND2_X1 U6308 ( .A1(n5130), .A2(n5129), .ZN(n4881) );
  NAND3_X1 U6309 ( .A1(n4883), .A2(n4882), .A3(n5063), .ZN(n5094) );
  NAND2_X1 U6310 ( .A1(n8617), .A2(n4886), .ZN(n4884) );
  NAND2_X1 U6311 ( .A1(n4884), .A2(n4885), .ZN(n8576) );
  NAND2_X2 U6312 ( .A1(n5252), .A2(n5251), .ZN(n5264) );
  INV_X1 U6313 ( .A(n7784), .ZN(n4906) );
  NAND2_X1 U6314 ( .A1(n4902), .A2(n4903), .ZN(n9525) );
  NAND2_X1 U6315 ( .A1(n7784), .A2(n4904), .ZN(n4902) );
  OAI21_X1 U6316 ( .B1(n5014), .B2(n6928), .A(n5099), .ZN(n4908) );
  AND2_X1 U6317 ( .A1(n5085), .A2(n6916), .ZN(n5014) );
  NAND3_X1 U6318 ( .A1(n4910), .A2(n4909), .A3(n5529), .ZN(n4911) );
  NAND2_X2 U6319 ( .A1(n4911), .A2(n5530), .ZN(n8926) );
  NAND2_X1 U6320 ( .A1(n8971), .A2(n4914), .ZN(n4919) );
  NAND2_X1 U6321 ( .A1(n8971), .A2(n8970), .ZN(n4915) );
  OR2_X1 U6322 ( .A1(n8970), .A2(n4921), .ZN(n4917) );
  OR2_X1 U6323 ( .A1(n8971), .A2(n4921), .ZN(n4918) );
  AND2_X2 U6324 ( .A1(n5019), .A2(n4927), .ZN(n4926) );
  NAND2_X1 U6325 ( .A1(n7894), .A2(n4932), .ZN(n4930) );
  AND2_X1 U6326 ( .A1(n5431), .A2(n5430), .ZN(n4953) );
  OAI21_X1 U6327 ( .B1(n7600), .B2(n4958), .A(n4955), .ZN(n7728) );
  OAI211_X1 U6328 ( .C1(n4965), .C2(n4378), .A(n4964), .B(n4963), .ZN(n5092)
         );
  NAND3_X1 U6329 ( .A1(n4378), .A2(n9057), .A3(n9603), .ZN(n4964) );
  NAND2_X1 U6330 ( .A1(n4390), .A2(n4969), .ZN(n4968) );
  NAND2_X1 U6331 ( .A1(n8393), .A2(n4977), .ZN(n4975) );
  NAND2_X1 U6332 ( .A1(n4979), .A2(n4421), .ZN(n6514) );
  NAND3_X1 U6333 ( .A1(n4414), .A2(n5858), .A3(n4983), .ZN(n5968) );
  NAND3_X1 U6334 ( .A1(n4990), .A2(n4989), .A3(n4984), .ZN(n7019) );
  AND2_X1 U6335 ( .A1(n8457), .A2(n6409), .ZN(n4991) );
  AND2_X1 U6336 ( .A1(n6432), .A2(n6427), .ZN(n4992) );
  NAND2_X2 U6337 ( .A1(n8266), .A2(n6484), .ZN(n8268) );
  NAND2_X1 U6338 ( .A1(n7317), .A2(n4993), .ZN(n8347) );
  OR3_X2 U6339 ( .A1(n6346), .A2(n4994), .A3(P2_IR_REG_26__SCAN_IN), .ZN(n5783) );
  NOR2_X2 U6340 ( .A1(n9662), .A2(n9726), .ZN(n7215) );
  OR2_X2 U6341 ( .A1(n9661), .A2(n9668), .ZN(n9662) );
  NAND2_X1 U6342 ( .A1(n5456), .A2(n5455), .ZN(n5485) );
  OAI21_X1 U6343 ( .B1(n8325), .B2(n8478), .A(n8324), .ZN(n8327) );
  AOI21_X1 U6344 ( .B1(n8191), .B2(n8186), .A(n8195), .ZN(n8183) );
  NAND2_X1 U6345 ( .A1(n7928), .A2(n9360), .ZN(n9353) );
  NAND2_X1 U6346 ( .A1(n6379), .A2(n9016), .ZN(n5755) );
  OAI21_X1 U6347 ( .B1(n6607), .B2(n6380), .A(n9016), .ZN(n6397) );
  NAND2_X1 U6348 ( .A1(n5703), .A2(n5671), .ZN(n5699) );
  NAND2_X1 U6349 ( .A1(n5185), .A2(n5184), .ZN(n5189) );
  INV_X1 U6350 ( .A(n9477), .ZN(n5037) );
  NAND2_X1 U6351 ( .A1(n5368), .A2(n5046), .ZN(n5076) );
  INV_X1 U6352 ( .A(n6401), .ZN(n7581) );
  INV_X1 U6353 ( .A(n8695), .ZN(n6030) );
  AND2_X1 U6354 ( .A1(n8125), .A2(n8121), .ZN(n8022) );
  AND2_X1 U6355 ( .A1(n5312), .A2(n5293), .ZN(n4999) );
  AND2_X1 U6356 ( .A1(n8200), .A2(n8199), .ZN(n5001) );
  AND2_X1 U6357 ( .A1(n6524), .A2(n6523), .ZN(n5002) );
  AND2_X1 U6358 ( .A1(n5081), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5003) );
  AND2_X1 U6359 ( .A1(n5289), .A2(n5269), .ZN(n5005) );
  INV_X1 U6360 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6335) );
  INV_X1 U6361 ( .A(n9882), .ZN(n9899) );
  NAND2_X1 U6362 ( .A1(n5686), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5006) );
  INV_X1 U6363 ( .A(n6761), .ZN(n6341) );
  AND2_X1 U6364 ( .A1(n5383), .A2(n5367), .ZN(n5007) );
  NOR2_X1 U6365 ( .A1(n6936), .A2(n5728), .ZN(n5008) );
  INV_X1 U6366 ( .A(n7139), .ZN(n6432) );
  NAND2_X1 U6367 ( .A1(n6331), .A2(n6333), .ZN(n5009) );
  AND2_X4 U6368 ( .A1(n9477), .A2(n5038), .ZN(n5010) );
  OR2_X1 U6369 ( .A1(n7199), .A2(n7198), .ZN(P1_U3289) );
  NOR2_X1 U6370 ( .A1(n5675), .A2(n5674), .ZN(n5012) );
  AND2_X1 U6371 ( .A1(n5699), .A2(n5701), .ZN(n5013) );
  NAND2_X1 U6372 ( .A1(n9791), .A2(n9526), .ZN(n8781) );
  AND2_X1 U6373 ( .A1(n8861), .A2(n8494), .ZN(n5015) );
  INV_X1 U6374 ( .A(n7885), .ZN(n6489) );
  OR2_X1 U6375 ( .A1(n8406), .A2(n8462), .ZN(n5016) );
  AND2_X1 U6376 ( .A1(n7399), .A2(n6224), .ZN(n5017) );
  INV_X1 U6377 ( .A(n9672), .ZN(n9189) );
  OR2_X1 U6378 ( .A1(n6223), .A2(n6324), .ZN(n6224) );
  OAI21_X1 U6379 ( .B1(n6226), .B2(n6225), .A(n5017), .ZN(n6230) );
  INV_X1 U6380 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5758) );
  AND4_X1 U6381 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5777)
         );
  NAND2_X1 U6382 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  NAND2_X1 U6383 ( .A1(n4376), .A2(n5501), .ZN(n5502) );
  INV_X1 U6384 ( .A(n10250), .ZN(n7999) );
  INV_X1 U6385 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10082) );
  INV_X1 U6386 ( .A(n8042), .ZN(n7918) );
  INV_X1 U6387 ( .A(n8016), .ZN(n7210) );
  AND4_X1 U6388 ( .A1(n5022), .A2(n5021), .A3(n5240), .A4(n5295), .ZN(n5023)
         );
  INV_X1 U6389 ( .A(n8345), .ZN(n6459) );
  INV_X1 U6390 ( .A(n6034), .ZN(n6033) );
  INV_X1 U6391 ( .A(n6016), .ZN(n6015) );
  OAI21_X1 U6392 ( .B1(n7707), .B2(n7706), .A(n6257), .ZN(n9528) );
  INV_X1 U6393 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10208) );
  INV_X1 U6394 ( .A(n8897), .ZN(n5229) );
  NAND2_X1 U6395 ( .A1(n5330), .A2(n5332), .ZN(n5333) );
  OR2_X1 U6396 ( .A1(n8918), .A2(n8919), .ZN(n5529) );
  INV_X1 U6397 ( .A(n5518), .ZN(n5516) );
  INV_X1 U6398 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7496) );
  AND2_X1 U6399 ( .A1(n9380), .A2(n9727), .ZN(n9381) );
  INV_X1 U6400 ( .A(n5672), .ZN(n5673) );
  INV_X1 U6401 ( .A(SI_20_), .ZN(n5534) );
  INV_X1 U6402 ( .A(SI_10_), .ZN(n10120) );
  AND2_X1 U6403 ( .A1(n6537), .A2(n6536), .ZN(n8322) );
  INV_X1 U6404 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5925) );
  INV_X1 U6405 ( .A(n6974), .ZN(n6405) );
  OR2_X1 U6406 ( .A1(n6077), .A2(n6076), .ZN(n6097) );
  OR2_X1 U6407 ( .A1(n6057), .A2(n10225), .ZN(n6077) );
  NAND2_X1 U6408 ( .A1(n5998), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6007) );
  INV_X1 U6409 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8516) );
  INV_X1 U6410 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5935) );
  INV_X1 U6411 ( .A(n6403), .ZN(n5804) );
  OAI22_X1 U6412 ( .A1(n7703), .A2(n7702), .B1(n8388), .B2(n8498), .ZN(n7784)
         );
  OR3_X1 U6413 ( .A1(n5921), .A2(P2_IR_REG_11__SCAN_IN), .A3(n5920), .ZN(n5932) );
  INV_X1 U6414 ( .A(n5098), .ZN(n5187) );
  NAND2_X1 U6415 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  OR2_X1 U6416 ( .A1(n5684), .A2(n5683), .ZN(n5736) );
  INV_X1 U6417 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8983) );
  AND2_X1 U6418 ( .A1(n5300), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5318) );
  INV_X1 U6419 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7829) );
  AND2_X1 U6420 ( .A1(n9406), .A2(n9245), .ZN(n9144) );
  NAND2_X1 U6421 ( .A1(n5576), .A2(n5575), .ZN(n5606) );
  NAND2_X1 U6422 ( .A1(n5415), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5443) );
  NOR2_X1 U6423 ( .A1(n5274), .A2(n5273), .ZN(n5300) );
  OR2_X1 U6424 ( .A1(n8198), .A2(n8255), .ZN(n5729) );
  AND2_X1 U6425 ( .A1(n5045), .A2(n5044), .ZN(n5046) );
  NAND2_X1 U6426 ( .A1(n6628), .A2(n6636), .ZN(n5158) );
  OR2_X1 U6427 ( .A1(n6007), .A2(n8364), .ZN(n6016) );
  OR2_X1 U6428 ( .A1(n5926), .A2(n5925), .ZN(n5936) );
  INV_X1 U6429 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10225) );
  OR2_X1 U6430 ( .A1(n6026), .A2(n8371), .ZN(n6034) );
  NOR2_X1 U6431 ( .A1(n5936), .A2(n5935), .ZN(n5959) );
  INV_X1 U6432 ( .A(n8294), .ZN(n9542) );
  INV_X1 U6433 ( .A(n9790), .ZN(n9531) );
  AND2_X1 U6434 ( .A1(n7813), .A2(n6540), .ZN(n6541) );
  INV_X1 U6435 ( .A(n6590), .ZN(n5613) );
  NAND2_X1 U6436 ( .A1(n8896), .A2(n5231), .ZN(n5233) );
  AND2_X1 U6437 ( .A1(n5736), .A2(n5685), .ZN(n9229) );
  OR2_X1 U6438 ( .A1(n5540), .A2(n8983), .ZN(n5579) );
  INV_X1 U6439 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6707) );
  INV_X1 U6440 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10214) );
  OR2_X1 U6441 ( .A1(n6705), .A2(n7880), .ZN(n6719) );
  INV_X1 U6442 ( .A(n9147), .ZN(n9227) );
  INV_X1 U6443 ( .A(n8022), .ZN(n7468) );
  OR2_X1 U6444 ( .A1(n6936), .A2(n9374), .ZN(n7109) );
  AND3_X1 U6445 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n9127) );
  AND2_X1 U6446 ( .A1(n8155), .A2(n9154), .ZN(n9307) );
  INV_X1 U6447 ( .A(n8018), .ZN(n7269) );
  AND2_X1 U6448 ( .A1(n6941), .A2(n6940), .ZN(n9672) );
  NAND2_X1 U6449 ( .A1(n9376), .A2(n5725), .ZN(n6936) );
  INV_X1 U6450 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5029) );
  XNOR2_X1 U6451 ( .A(n5048), .B(n5070), .ZN(n5724) );
  NOR2_X1 U6452 ( .A1(n6570), .A2(n6576), .ZN(n8315) );
  AND2_X1 U6453 ( .A1(n6574), .A2(n7023), .ZN(n6569) );
  AND2_X1 U6454 ( .A1(n8315), .A2(n9785), .ZN(n8480) );
  AND2_X1 U6455 ( .A1(n6138), .A2(n6137), .ZN(n6573) );
  INV_X1 U6456 ( .A(n6079), .ZN(n6132) );
  AND4_X1 U6457 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n8432)
         );
  INV_X1 U6458 ( .A(n9776), .ZN(n9774) );
  NAND2_X1 U6459 ( .A1(n8704), .A2(n8712), .ZN(n8703) );
  AND2_X1 U6460 ( .A1(n6273), .A2(n6272), .ZN(n8740) );
  INV_X1 U6461 ( .A(n9809), .ZN(n7023) );
  AND2_X1 U6462 ( .A1(n9791), .A2(n7077), .ZN(n8767) );
  INV_X1 U6463 ( .A(n8781), .ZN(n8598) );
  NAND2_X1 U6464 ( .A1(n9831), .A2(n6552), .ZN(n7291) );
  INV_X1 U6465 ( .A(n9871), .ZN(n9904) );
  INV_X1 U6466 ( .A(n7291), .ZN(n7309) );
  OR2_X1 U6467 ( .A1(n6578), .A2(P2_U3152), .ZN(n9809) );
  INV_X1 U6468 ( .A(n5294), .ZN(n6613) );
  OAI21_X1 U6469 ( .B1(n4559), .B2(n9020), .A(n6394), .ZN(n6395) );
  OR2_X1 U6470 ( .A1(n6936), .A2(n8255), .ZN(n9742) );
  AND2_X1 U6471 ( .A1(n5748), .A2(n4378), .ZN(n9500) );
  INV_X1 U6472 ( .A(n6647), .ZN(n8259) );
  OR2_X1 U6473 ( .A1(n9198), .A2(n5581), .ZN(n6391) );
  NAND2_X1 U6474 ( .A1(n5686), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5111) );
  AND2_X1 U6475 ( .A1(n9109), .A2(n6706), .ZN(n9654) );
  INV_X1 U6476 ( .A(n9647), .ZN(n9593) );
  INV_X1 U6477 ( .A(n9629), .ZN(n9656) );
  AND2_X1 U6478 ( .A1(n9221), .A2(n8171), .ZN(n9243) );
  INV_X1 U6479 ( .A(n7676), .ZN(n9340) );
  AOI21_X1 U6480 ( .B1(n6667), .B2(n5718), .A(n6668), .ZN(n6693) );
  AND2_X1 U6481 ( .A1(n7925), .A2(n7924), .ZN(n9440) );
  NAND2_X1 U6482 ( .A1(n9690), .A2(n9377), .ZN(n9755) );
  AND2_X1 U6483 ( .A1(n6672), .A2(n6671), .ZN(n7106) );
  NAND2_X1 U6484 ( .A1(n5706), .A2(n5707), .ZN(n6670) );
  NOR2_X1 U6485 ( .A1(n10257), .A2(n7762), .ZN(n7763) );
  OAI21_X1 U6486 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9929), .ZN(n10260) );
  AND2_X1 U6487 ( .A1(n6660), .A2(n6659), .ZN(n9775) );
  AND2_X1 U6488 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  INV_X1 U6489 ( .A(n8481), .ZN(n8470) );
  INV_X1 U6490 ( .A(n8480), .ZN(n8424) );
  INV_X1 U6491 ( .A(n8455), .ZN(n8485) );
  INV_X1 U6492 ( .A(n6573), .ZN(n8571) );
  INV_X1 U6493 ( .A(n8398), .ZN(n8663) );
  NAND2_X1 U6494 ( .A1(n6805), .A2(n6353), .ZN(n9777) );
  INV_X1 U6495 ( .A(n9773), .ZN(n9778) );
  NAND2_X1 U6496 ( .A1(n7023), .A2(n6556), .ZN(n9793) );
  INV_X1 U6497 ( .A(n8767), .ZN(n8783) );
  OR2_X1 U6498 ( .A1(n7310), .A2(n7291), .ZN(n9922) );
  INV_X2 U6499 ( .A(n9922), .ZN(n9924) );
  OR2_X1 U6500 ( .A1(n7310), .A2(n7309), .ZN(n9906) );
  NOR2_X1 U6501 ( .A1(n9810), .A2(n9809), .ZN(n9820) );
  CLKBUF_X1 U6502 ( .A(n9820), .Z(n9835) );
  INV_X1 U6503 ( .A(n6191), .ZN(n7643) );
  INV_X1 U6504 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7065) );
  INV_X1 U6505 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10011) );
  CLKBUF_X1 U6506 ( .A(n8894), .Z(n7582) );
  AND2_X1 U6507 ( .A1(n5734), .A2(n5733), .ZN(n9517) );
  OR2_X1 U6508 ( .A1(n6920), .A2(n9742), .ZN(n9020) );
  INV_X1 U6509 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U6510 ( .A1(n6391), .A2(n6390), .ZN(n9210) );
  NAND2_X1 U6511 ( .A1(n6721), .A2(n6720), .ZN(n9647) );
  OR2_X1 U6512 ( .A1(P1_U3083), .A2(n6684), .ZN(n9629) );
  NAND2_X1 U6513 ( .A1(n9692), .A2(n9675), .ZN(n9370) );
  INV_X1 U6514 ( .A(n9772), .ZN(n9770) );
  AND2_X2 U6515 ( .A1(n6694), .A2(n6693), .ZN(n9772) );
  INV_X1 U6516 ( .A(n9759), .ZN(n9757) );
  INV_X1 U6517 ( .A(n9700), .ZN(n9699) );
  NAND2_X1 U6518 ( .A1(n6647), .A2(n6670), .ZN(n9700) );
  INV_X1 U6519 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7810) );
  INV_X1 U6520 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7063) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U6522 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  OAI21_X1 U6523 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9941), .ZN(n9939) );
  INV_X2 U6524 ( .A(n8491), .ZN(P2_U3966) );
  NOR2_X1 U6525 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5022) );
  INV_X1 U6526 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6527 ( .A1(n5368), .A2(n5026), .ZN(n5033) );
  NAND2_X1 U6528 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5027) );
  INV_X1 U6529 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5031) );
  NAND3_X1 U6530 ( .A1(n5031), .A2(n5067), .A3(n5029), .ZN(n5032) );
  AND2_X2 U6531 ( .A1(n5036), .A2(n5037), .ZN(n5686) );
  NAND2_X1 U6532 ( .A1(n7994), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5041) );
  AND2_X4 U6533 ( .A1(n5037), .A2(n5038), .ZN(n7995) );
  NAND2_X1 U6534 ( .A1(n7995), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6535 ( .A1(n5010), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U6536 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5410) );
  AND2_X1 U6537 ( .A1(n5438), .A2(n5410), .ZN(n5045) );
  NAND2_X1 U6538 ( .A1(n5486), .A2(n5042), .ZN(n5043) );
  NAND2_X1 U6539 ( .A1(n5073), .A2(n5071), .ZN(n5047) );
  NAND2_X1 U6540 ( .A1(n5368), .A2(n5050), .ZN(n5720) );
  NAND2_X1 U6541 ( .A1(n4426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6542 ( .A1(n5059), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5060) );
  INV_X1 U6543 ( .A(SI_0_), .ZN(n5062) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U6545 ( .B1(n4377), .B2(n5062), .A(n5061), .ZN(n5064) );
  AND2_X1 U6546 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5063) );
  AND2_X1 U6547 ( .A1(n5064), .A2(n5094), .ZN(n9480) );
  INV_X1 U6548 ( .A(n5719), .ZN(n5081) );
  NAND2_X1 U6549 ( .A1(n5069), .A2(n5068), .ZN(n5084) );
  INV_X1 U6550 ( .A(n5084), .ZN(n6919) );
  AND2_X1 U6551 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NAND2_X1 U6552 ( .A1(n5073), .A2(n5072), .ZN(n5074) );
  NAND2_X1 U6553 ( .A1(n5074), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6554 ( .A1(n5076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6555 ( .A1(n6919), .A2(n7169), .ZN(n5085) );
  NAND2_X1 U6556 ( .A1(n9376), .A2(n8255), .ZN(n5079) );
  AND3_X4 U6557 ( .A1(n5080), .A2(n5719), .A3(n5079), .ZN(n6590) );
  NAND2_X1 U6558 ( .A1(n5010), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6559 ( .A1(n7994), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6560 ( .A1(n5686), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5086) );
  NAND4_X2 U6561 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n9055)
         );
  INV_X1 U6562 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6634) );
  INV_X1 U6563 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6564 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5090) );
  XNOR2_X1 U6565 ( .A(n5091), .B(n5090), .ZN(n6710) );
  INV_X1 U6566 ( .A(SI_1_), .ZN(n5095) );
  XNOR2_X1 U6567 ( .A(n5104), .B(n5103), .ZN(n6633) );
  OR2_X1 U6568 ( .A1(n5128), .A2(n6633), .ZN(n5096) );
  AOI22_X1 U6569 ( .A1(n9055), .A2(n6590), .B1(n7122), .B2(n5098), .ZN(n6926)
         );
  NAND2_X1 U6570 ( .A1(n5151), .A2(n5102), .ZN(n5125) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U6572 ( .A1(n5104), .A2(n5103), .ZN(n5107) );
  NAND2_X1 U6573 ( .A1(n5105), .A2(SI_1_), .ZN(n5106) );
  NAND2_X1 U6574 ( .A1(n5107), .A2(n5106), .ZN(n5130) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6624) );
  XNOR2_X1 U6576 ( .A(n5131), .B(SI_2_), .ZN(n5129) );
  XNOR2_X1 U6577 ( .A(n5130), .B(n5129), .ZN(n6629) );
  OR2_X1 U6578 ( .A1(n5128), .A2(n6629), .ZN(n5108) );
  NAND2_X1 U6579 ( .A1(n7988), .A2(n6359), .ZN(n5116) );
  NAND2_X1 U6580 ( .A1(n5010), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6581 ( .A1(n7995), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6582 ( .A1(n7994), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6583 ( .A1(n9054), .A2(n5114), .ZN(n5115) );
  NAND2_X1 U6584 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  XNOR2_X1 U6585 ( .A(n5117), .B(n6362), .ZN(n5119) );
  AOI22_X1 U6586 ( .A1(n9054), .A2(n6590), .B1(n7988), .B2(n5098), .ZN(n5118)
         );
  NAND2_X1 U6587 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  OAI21_X1 U6588 ( .B1(n5119), .B2(n5118), .A(n5120), .ZN(n7986) );
  INV_X1 U6589 ( .A(n5120), .ZN(n7011) );
  OR2_X1 U6590 ( .A1(n5581), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6591 ( .A1(n5010), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6592 ( .A1(n7995), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6593 ( .A1(n7994), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6594 ( .A1(n9053), .A2(n5114), .ZN(n5137) );
  NAND2_X1 U6595 ( .A1(n5125), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5127) );
  INV_X1 U6596 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6597 ( .A(n5127), .B(n5126), .ZN(n6714) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6632) );
  OR2_X1 U6599 ( .A1(n4405), .A2(n6632), .ZN(n5135) );
  INV_X1 U6600 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6601 ( .A1(n5132), .A2(SI_2_), .ZN(n5133) );
  INV_X1 U6602 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6626) );
  XNOR2_X1 U6603 ( .A(n5155), .B(SI_3_), .ZN(n5153) );
  XNOR2_X1 U6604 ( .A(n5154), .B(n5153), .ZN(n6631) );
  NAND2_X1 U6605 ( .A1(n7160), .A2(n6359), .ZN(n5136) );
  NAND2_X1 U6606 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  XNOR2_X1 U6607 ( .A(n5138), .B(n6362), .ZN(n5139) );
  AOI22_X1 U6608 ( .A1(n9053), .A2(n6590), .B1(n7160), .B2(n5098), .ZN(n5140)
         );
  NAND2_X1 U6609 ( .A1(n5139), .A2(n5140), .ZN(n5144) );
  INV_X1 U6610 ( .A(n5139), .ZN(n5142) );
  INV_X1 U6611 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6612 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  AND2_X1 U6613 ( .A1(n5144), .A2(n5143), .ZN(n7010) );
  NAND2_X1 U6614 ( .A1(n7008), .A2(n5144), .ZN(n7001) );
  NAND2_X1 U6615 ( .A1(n5010), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6616 ( .A1(n7995), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5148) );
  INV_X1 U6617 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6701) );
  OR2_X1 U6618 ( .A1(n6388), .A2(n6701), .ZN(n5147) );
  AND2_X2 U6619 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5165) );
  NOR2_X1 U6620 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5145) );
  NOR2_X1 U6621 ( .A1(n5165), .A2(n5145), .ZN(n7254) );
  NAND2_X1 U6622 ( .A1(n5686), .A2(n7254), .ZN(n5146) );
  NAND4_X1 U6623 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n9052)
         );
  OAI21_X1 U6624 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6625 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  XNOR2_X1 U6626 ( .A(n5152), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9620) );
  INV_X1 U6627 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6636) );
  OR2_X1 U6628 ( .A1(n4405), .A2(n6636), .ZN(n5160) );
  INV_X1 U6629 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6630 ( .A1(n5156), .A2(SI_3_), .ZN(n5157) );
  INV_X1 U6631 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6627) );
  XNOR2_X1 U6632 ( .A(n5176), .B(SI_4_), .ZN(n5174) );
  XNOR2_X1 U6633 ( .A(n5175), .B(n5174), .ZN(n6635) );
  OR2_X1 U6634 ( .A1(n5128), .A2(n6635), .ZN(n5159) );
  OAI211_X1 U6635 ( .C1(n9620), .C2(n5294), .A(n5160), .B(n5159), .ZN(n7255)
         );
  AOI22_X1 U6636 ( .A1(n9052), .A2(n6590), .B1(n7255), .B2(n5098), .ZN(n5162)
         );
  AOI22_X1 U6637 ( .A1(n9052), .A2(n5114), .B1(n7255), .B2(n6359), .ZN(n5161)
         );
  XNOR2_X1 U6638 ( .A(n5161), .B(n7169), .ZN(n5163) );
  XOR2_X1 U6639 ( .A(n5162), .B(n5163), .Z(n7002) );
  NAND2_X1 U6640 ( .A1(n7001), .A2(n7002), .ZN(n7000) );
  NAND2_X1 U6641 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  NAND2_X1 U6642 ( .A1(n7000), .A2(n5164), .ZN(n5185) );
  INV_X1 U6643 ( .A(n5185), .ZN(n5183) );
  NAND2_X1 U6644 ( .A1(n5010), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6645 ( .A1(n5165), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5190) );
  OAI21_X1 U6646 ( .B1(n5165), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5190), .ZN(
        n9666) );
  OR2_X1 U6647 ( .A1(n5581), .A2(n9666), .ZN(n5169) );
  INV_X1 U6648 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5166) );
  OR2_X1 U6649 ( .A1(n5690), .A2(n5166), .ZN(n5168) );
  NAND2_X1 U6650 ( .A1(n7994), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5167) );
  NAND4_X1 U6651 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n9051)
         );
  NAND2_X1 U6652 ( .A1(n5171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6653 ( .A(n5172), .B(n5019), .ZN(n6737) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6639) );
  OR2_X1 U6655 ( .A1(n4405), .A2(n6639), .ZN(n5180) );
  INV_X1 U6656 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6657 ( .A1(n5177), .A2(SI_4_), .ZN(n5178) );
  INV_X1 U6658 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U6659 ( .A(n6637), .B(n6639), .S(n6628), .Z(n5200) );
  OR2_X1 U6660 ( .A1(n5128), .A2(n6638), .ZN(n5179) );
  AOI22_X1 U6661 ( .A1(n9051), .A2(n5114), .B1(n9668), .B2(n6359), .ZN(n5181)
         );
  XNOR2_X1 U6662 ( .A(n5181), .B(n7169), .ZN(n5184) );
  INV_X1 U6663 ( .A(n5184), .ZN(n5182) );
  NAND2_X1 U6664 ( .A1(n5183), .A2(n5182), .ZN(n5186) );
  INV_X1 U6665 ( .A(n9051), .ZN(n9021) );
  OAI22_X1 U6666 ( .A1(n9021), .A2(n5613), .B1(n9722), .B2(n5187), .ZN(n6616)
         );
  INV_X1 U6667 ( .A(n6616), .ZN(n5188) );
  OR2_X1 U6668 ( .A1(n6388), .A2(n10012), .ZN(n5195) );
  INV_X1 U6669 ( .A(n5010), .ZN(n5687) );
  NAND2_X1 U6670 ( .A1(n5010), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5194) );
  AND2_X1 U6671 ( .A1(n5190), .A2(n6707), .ZN(n5191) );
  NOR2_X1 U6672 ( .A1(n5190), .A2(n6707), .ZN(n5209) );
  OR2_X1 U6673 ( .A1(n5191), .A2(n5209), .ZN(n9023) );
  OR2_X1 U6674 ( .A1(n5581), .A2(n9023), .ZN(n5193) );
  NAND2_X1 U6675 ( .A1(n7995), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5192) );
  NAND4_X1 U6676 ( .A1(n5195), .A2(n5194), .A3(n5193), .A4(n5192), .ZN(n9665)
         );
  NAND2_X1 U6677 ( .A1(n9665), .A2(n5114), .ZN(n5205) );
  NAND2_X1 U6678 ( .A1(n5196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6679 ( .A(n5197), .B(n4927), .ZN(n6747) );
  INV_X1 U6680 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6640) );
  OR2_X1 U6681 ( .A1(n4405), .A2(n6640), .ZN(n5203) );
  INV_X1 U6682 ( .A(n5200), .ZN(n5201) );
  INV_X1 U6683 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6642) );
  MUX2_X1 U6684 ( .A(n6642), .B(n6640), .S(n4396), .Z(n5219) );
  XNOR2_X1 U6685 ( .A(n5219), .B(SI_6_), .ZN(n5217) );
  OR2_X1 U6686 ( .A1(n5128), .A2(n6641), .ZN(n5202) );
  OAI211_X1 U6687 ( .C1(n5294), .C2(n6747), .A(n5203), .B(n5202), .ZN(n9726)
         );
  NAND2_X1 U6688 ( .A1(n9726), .A2(n6359), .ZN(n5204) );
  NAND2_X1 U6689 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  XNOR2_X1 U6690 ( .A(n5206), .B(n6362), .ZN(n5208) );
  AOI22_X1 U6691 ( .A1(n9665), .A2(n6590), .B1(n9726), .B2(n5098), .ZN(n5207)
         );
  AND2_X1 U6692 ( .A1(n5208), .A2(n5207), .ZN(n9013) );
  OR2_X1 U6693 ( .A1(n5208), .A2(n5207), .ZN(n9012) );
  NAND2_X1 U6694 ( .A1(n5010), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6695 ( .A1(n5209), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5234) );
  OR2_X1 U6696 ( .A1(n5209), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6697 ( .A1(n5234), .A2(n5210), .ZN(n8904) );
  OR2_X1 U6698 ( .A1(n5581), .A2(n8904), .ZN(n5213) );
  INV_X1 U6699 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6745) );
  OR2_X1 U6700 ( .A1(n6388), .A2(n6745), .ZN(n5212) );
  NAND2_X1 U6701 ( .A1(n7995), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5211) );
  NAND4_X1 U6702 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n9050)
         );
  NAND2_X1 U6703 ( .A1(n9050), .A2(n5114), .ZN(n5225) );
  OR2_X1 U6704 ( .A1(n5215), .A2(n4595), .ZN(n5216) );
  XNOR2_X1 U6705 ( .A(n5216), .B(n5240), .ZN(n6748) );
  OR2_X1 U6706 ( .A1(n4405), .A2(n10226), .ZN(n5223) );
  INV_X1 U6707 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6708 ( .A1(n5220), .A2(SI_6_), .ZN(n5221) );
  MUX2_X1 U6709 ( .A(n10204), .B(n10226), .S(n4396), .Z(n5249) );
  XNOR2_X1 U6710 ( .A(n5249), .B(SI_7_), .ZN(n5247) );
  XNOR2_X1 U6711 ( .A(n5248), .B(n5247), .ZN(n6644) );
  OR2_X1 U6712 ( .A1(n5128), .A2(n6644), .ZN(n5222) );
  NAND2_X1 U6713 ( .A1(n8094), .A2(n6359), .ZN(n5224) );
  NAND2_X1 U6714 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  XNOR2_X1 U6715 ( .A(n5226), .B(n7169), .ZN(n8898) );
  INV_X1 U6716 ( .A(n8898), .ZN(n5230) );
  NAND2_X1 U6717 ( .A1(n9050), .A2(n6590), .ZN(n5228) );
  NAND2_X1 U6718 ( .A1(n8094), .A2(n5098), .ZN(n5227) );
  NAND2_X1 U6719 ( .A1(n5228), .A2(n5227), .ZN(n8897) );
  NAND2_X1 U6720 ( .A1(n8898), .A2(n8897), .ZN(n5232) );
  INV_X1 U6721 ( .A(n7439), .ZN(n5262) );
  NAND2_X1 U6722 ( .A1(n7994), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6723 ( .A1(n5010), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6724 ( .A1(n5234), .A2(n10214), .ZN(n5235) );
  NAND2_X1 U6725 ( .A1(n5274), .A2(n5235), .ZN(n7443) );
  OR2_X1 U6726 ( .A1(n5581), .A2(n7443), .ZN(n5237) );
  NAND2_X1 U6727 ( .A1(n7995), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5236) );
  NAND4_X1 U6728 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n9049)
         );
  INV_X1 U6729 ( .A(n9049), .ZN(n7606) );
  AND2_X1 U6730 ( .A1(n5215), .A2(n5240), .ZN(n5244) );
  NOR2_X1 U6731 ( .A1(n5244), .A2(n4595), .ZN(n5241) );
  MUX2_X1 U6732 ( .A(n4595), .B(n5241), .S(P1_IR_REG_8__SCAN_IN), .Z(n5242) );
  INV_X1 U6733 ( .A(n5242), .ZN(n5246) );
  INV_X1 U6734 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5243) );
  INV_X1 U6735 ( .A(n5296), .ZN(n5245) );
  NAND2_X1 U6736 ( .A1(n5246), .A2(n5245), .ZN(n6902) );
  OR2_X1 U6737 ( .A1(n4405), .A2(n6650), .ZN(n5258) );
  NAND2_X1 U6738 ( .A1(n5248), .A2(n5247), .ZN(n5252) );
  INV_X1 U6739 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6740 ( .A1(n5250), .A2(SI_7_), .ZN(n5251) );
  INV_X1 U6741 ( .A(SI_8_), .ZN(n5253) );
  NAND2_X1 U6742 ( .A1(n5254), .A2(n5253), .ZN(n5265) );
  INV_X1 U6743 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6744 ( .A1(n5255), .A2(SI_8_), .ZN(n5256) );
  XNOR2_X1 U6745 ( .A(n5264), .B(n5004), .ZN(n6649) );
  OR2_X1 U6746 ( .A1(n5128), .A2(n6649), .ZN(n5257) );
  OAI211_X1 U6747 ( .C1(n5294), .C2(n6902), .A(n5258), .B(n5257), .ZN(n7445)
         );
  INV_X1 U6748 ( .A(n7445), .ZN(n9743) );
  OAI22_X1 U6749 ( .A1(n7606), .A2(n5613), .B1(n9743), .B2(n5187), .ZN(n5260)
         );
  INV_X1 U6750 ( .A(n5260), .ZN(n7436) );
  AOI22_X1 U6751 ( .A1(n9049), .A2(n5114), .B1(n7445), .B2(n6359), .ZN(n5259)
         );
  XOR2_X1 U6752 ( .A(n7169), .B(n5259), .Z(n7437) );
  OAI21_X1 U6753 ( .B1(n7439), .B2(n5260), .A(n7437), .ZN(n5261) );
  OAI21_X2 U6754 ( .B1(n5262), .B2(n7436), .A(n5261), .ZN(n7600) );
  OR2_X1 U6755 ( .A1(n5296), .A2(n4595), .ZN(n5263) );
  XNOR2_X1 U6756 ( .A(n5263), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9640) );
  INV_X1 U6757 ( .A(n9640), .ZN(n6652) );
  MUX2_X1 U6758 ( .A(n6654), .B(n10209), .S(n6628), .Z(n5267) );
  INV_X1 U6759 ( .A(SI_9_), .ZN(n5266) );
  NAND2_X1 U6760 ( .A1(n5267), .A2(n5266), .ZN(n5289) );
  INV_X1 U6761 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U6762 ( .A1(n5268), .A2(SI_9_), .ZN(n5269) );
  XNOR2_X1 U6763 ( .A(n5288), .B(n5005), .ZN(n6651) );
  NAND2_X1 U6764 ( .A1(n6651), .A2(n8035), .ZN(n5271) );
  OR2_X1 U6765 ( .A1(n4405), .A2(n10209), .ZN(n5270) );
  OAI211_X1 U6766 ( .C1(n5294), .C2(n6652), .A(n5271), .B(n5270), .ZN(n7393)
         );
  NAND2_X1 U6767 ( .A1(n7393), .A2(n6359), .ZN(n5281) );
  NAND2_X1 U6768 ( .A1(n5010), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5279) );
  INV_X1 U6769 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5272) );
  OR2_X1 U6770 ( .A1(n6388), .A2(n5272), .ZN(n5278) );
  AND2_X1 U6771 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  OR2_X1 U6772 ( .A1(n5275), .A2(n5300), .ZN(n7603) );
  OR2_X1 U6773 ( .A1(n5581), .A2(n7603), .ZN(n5277) );
  NAND2_X1 U6774 ( .A1(n7995), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5276) );
  NAND4_X1 U6775 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n9048)
         );
  NAND2_X1 U6776 ( .A1(n9048), .A2(n5114), .ZN(n5280) );
  NAND2_X1 U6777 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  XNOR2_X1 U6778 ( .A(n5282), .B(n6362), .ZN(n5286) );
  NAND2_X1 U6779 ( .A1(n7393), .A2(n6365), .ZN(n5284) );
  NAND2_X1 U6780 ( .A1(n9048), .A2(n6590), .ZN(n5283) );
  AND2_X1 U6781 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  NAND2_X1 U6782 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  OAI21_X1 U6783 ( .B1(n5286), .B2(n5285), .A(n5287), .ZN(n7601) );
  INV_X1 U6784 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5290) );
  MUX2_X1 U6785 ( .A(n6662), .B(n5290), .S(n4396), .Z(n5291) );
  NAND2_X1 U6786 ( .A1(n5291), .A2(n10120), .ZN(n5312) );
  INV_X1 U6787 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6788 ( .A1(n5292), .A2(SI_10_), .ZN(n5293) );
  XNOR2_X1 U6789 ( .A(n5311), .B(n4999), .ZN(n6655) );
  NAND2_X1 U6790 ( .A1(n6655), .A2(n8035), .ZN(n5299) );
  NAND2_X1 U6791 ( .A1(n5296), .A2(n5295), .ZN(n5313) );
  NAND2_X1 U6792 ( .A1(n5313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6793 ( .A(n5297), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U6794 ( .A1(n5513), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6613), .B2(
        n9655), .ZN(n5298) );
  NAND2_X1 U6795 ( .A1(n5299), .A2(n5298), .ZN(n7638) );
  NOR2_X1 U6796 ( .A1(n5300), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5301) );
  OR2_X1 U6797 ( .A1(n5318), .A2(n5301), .ZN(n7631) );
  OR2_X1 U6798 ( .A1(n5581), .A2(n7631), .ZN(n5305) );
  NAND2_X1 U6799 ( .A1(n5010), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6800 ( .A1(n7995), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6801 ( .A1(n7994), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5302) );
  NAND4_X1 U6802 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n9047)
         );
  AOI22_X1 U6803 ( .A1(n7638), .A2(n6359), .B1(n5114), .B2(n9047), .ZN(n5306)
         );
  XOR2_X1 U6804 ( .A(n7169), .B(n5306), .Z(n5307) );
  INV_X1 U6805 ( .A(n7638), .ZN(n9493) );
  INV_X1 U6806 ( .A(n9047), .ZN(n7734) );
  OAI22_X1 U6807 ( .A1(n9493), .A2(n5187), .B1(n7734), .B2(n5613), .ZN(n5308)
         );
  NAND2_X1 U6808 ( .A1(n5307), .A2(n5308), .ZN(n7629) );
  INV_X1 U6809 ( .A(n5307), .ZN(n5310) );
  INV_X1 U6810 ( .A(n5308), .ZN(n5309) );
  NAND2_X1 U6811 ( .A1(n5310), .A2(n5309), .ZN(n7628) );
  INV_X1 U6812 ( .A(n7728), .ZN(n5329) );
  MUX2_X1 U6813 ( .A(n10188), .B(n6679), .S(n4396), .Z(n5335) );
  XNOR2_X1 U6814 ( .A(n5335), .B(SI_11_), .ZN(n5334) );
  XNOR2_X1 U6815 ( .A(n5339), .B(n5334), .ZN(n6678) );
  NAND2_X1 U6816 ( .A1(n6678), .A2(n8035), .ZN(n5316) );
  OAI21_X1 U6817 ( .B1(n5313), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5314) );
  XNOR2_X1 U6818 ( .A(n5314), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U6819 ( .A1(n5513), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6613), .B2(
        n6991), .ZN(n5315) );
  INV_X1 U6820 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6821 ( .A1(n6388), .A2(n5317), .ZN(n5323) );
  OR2_X1 U6822 ( .A1(n5318), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6823 ( .A1(n5348), .A2(n5319), .ZN(n7731) );
  OR2_X1 U6824 ( .A1(n5581), .A2(n7731), .ZN(n5322) );
  INV_X1 U6825 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7460) );
  OR2_X1 U6826 ( .A1(n5690), .A2(n7460), .ZN(n5321) );
  NAND2_X1 U6827 ( .A1(n5010), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5320) );
  NAND4_X1 U6828 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n9046)
         );
  AND2_X1 U6829 ( .A1(n9046), .A2(n6590), .ZN(n5324) );
  AOI21_X1 U6830 ( .B1(n7476), .B2(n6365), .A(n5324), .ZN(n5331) );
  NAND2_X1 U6831 ( .A1(n7476), .A2(n6359), .ZN(n5326) );
  NAND2_X1 U6832 ( .A1(n9046), .A2(n5098), .ZN(n5325) );
  NAND2_X1 U6833 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  XNOR2_X1 U6834 ( .A(n5327), .B(n7169), .ZN(n5330) );
  XOR2_X1 U6835 ( .A(n5331), .B(n5330), .Z(n7727) );
  INV_X1 U6836 ( .A(n7727), .ZN(n5328) );
  INV_X1 U6837 ( .A(n5331), .ZN(n5332) );
  INV_X1 U6838 ( .A(n5334), .ZN(n5338) );
  INV_X1 U6839 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6840 ( .A1(n5336), .A2(SI_11_), .ZN(n5337) );
  MUX2_X1 U6841 ( .A(n6868), .B(n6870), .S(n4396), .Z(n5341) );
  INV_X1 U6842 ( .A(SI_12_), .ZN(n5340) );
  NAND2_X1 U6843 ( .A1(n5341), .A2(n5340), .ZN(n5361) );
  INV_X1 U6844 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6845 ( .A1(n5342), .A2(SI_12_), .ZN(n5343) );
  NAND2_X1 U6846 ( .A1(n5361), .A2(n5343), .ZN(n5362) );
  XNOR2_X1 U6847 ( .A(n5363), .B(n5362), .ZN(n6867) );
  NAND2_X1 U6848 ( .A1(n6867), .A2(n8035), .ZN(n5346) );
  NAND2_X1 U6849 ( .A1(n4477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6850 ( .A(n5344), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7186) );
  AOI22_X1 U6851 ( .A1(n5513), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6613), .B2(
        n7186), .ZN(n5345) );
  NAND2_X1 U6852 ( .A1(n5010), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5353) );
  INV_X1 U6853 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6985) );
  OR2_X1 U6854 ( .A1(n6388), .A2(n6985), .ZN(n5352) );
  NAND2_X1 U6855 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6856 ( .A1(n5373), .A2(n5349), .ZN(n9516) );
  OR2_X1 U6857 ( .A1(n5581), .A2(n9516), .ZN(n5351) );
  NAND2_X1 U6858 ( .A1(n7995), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5350) );
  NAND4_X1 U6859 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n9045)
         );
  AOI22_X1 U6860 ( .A1(n7563), .A2(n5098), .B1(n6590), .B2(n9045), .ZN(n5358)
         );
  NAND2_X1 U6861 ( .A1(n7563), .A2(n6359), .ZN(n5355) );
  NAND2_X1 U6862 ( .A1(n9045), .A2(n6365), .ZN(n5354) );
  NAND2_X1 U6863 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  XNOR2_X1 U6864 ( .A(n5356), .B(n7169), .ZN(n5357) );
  XOR2_X1 U6865 ( .A(n5358), .B(n5357), .Z(n9507) );
  INV_X1 U6866 ( .A(n5357), .ZN(n5359) );
  NAND2_X1 U6867 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X2 U6868 ( .A1(n9511), .A2(n5360), .ZN(n7894) );
  INV_X1 U6869 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5364) );
  MUX2_X1 U6870 ( .A(n6925), .B(n5364), .S(n4397), .Z(n5365) );
  NAND2_X1 U6871 ( .A1(n5365), .A2(n10219), .ZN(n5383) );
  INV_X1 U6872 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6873 ( .A1(n5366), .A2(SI_13_), .ZN(n5367) );
  XNOR2_X1 U6874 ( .A(n5382), .B(n5007), .ZN(n6913) );
  NAND2_X1 U6875 ( .A1(n6913), .A2(n8035), .ZN(n5371) );
  INV_X1 U6876 ( .A(n5368), .ZN(n5386) );
  NAND2_X1 U6877 ( .A1(n5386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U6878 ( .A(n5369), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7499) );
  AOI22_X1 U6879 ( .A1(n5513), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6613), .B2(
        n7499), .ZN(n5370) );
  INV_X1 U6880 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7179) );
  OR2_X1 U6881 ( .A1(n6388), .A2(n7179), .ZN(n5378) );
  NAND2_X1 U6882 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U6883 ( .A1(n5391), .A2(n5374), .ZN(n7901) );
  OR2_X1 U6884 ( .A1(n5581), .A2(n7901), .ZN(n5377) );
  INV_X1 U6885 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7574) );
  OR2_X1 U6886 ( .A1(n5690), .A2(n7574), .ZN(n5376) );
  NAND2_X1 U6887 ( .A1(n5010), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5375) );
  NAND4_X1 U6888 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(n9499)
         );
  AOI22_X1 U6889 ( .A1(n7662), .A2(n6359), .B1(n5114), .B2(n9499), .ZN(n5379)
         );
  XOR2_X1 U6890 ( .A(n7169), .B(n5379), .Z(n7892) );
  INV_X1 U6891 ( .A(n7662), .ZN(n7895) );
  INV_X1 U6892 ( .A(n9499), .ZN(n7976) );
  OAI22_X1 U6893 ( .A1(n7895), .A2(n5187), .B1(n7976), .B2(n5613), .ZN(n7891)
         );
  NOR2_X1 U6894 ( .A1(n7892), .A2(n7891), .ZN(n5381) );
  NAND2_X1 U6895 ( .A1(n7892), .A2(n7891), .ZN(n5380) );
  NAND2_X1 U6896 ( .A1(n5382), .A2(n5007), .ZN(n5384) );
  MUX2_X1 U6897 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4396), .Z(n5403) );
  XNOR2_X1 U6898 ( .A(n5403), .B(SI_14_), .ZN(n5405) );
  INV_X1 U6899 ( .A(n5405), .ZN(n5385) );
  XNOR2_X1 U6900 ( .A(n5406), .B(n5385), .ZN(n6933) );
  NAND2_X1 U6901 ( .A1(n6933), .A2(n8035), .ZN(n5390) );
  NOR2_X1 U6902 ( .A1(n5386), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5387) );
  OR2_X1 U6903 ( .A1(n5387), .A2(n4595), .ZN(n5388) );
  XNOR2_X1 U6904 ( .A(n5388), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7688) );
  AOI22_X1 U6905 ( .A1(n5513), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6613), .B2(
        n7688), .ZN(n5389) );
  NAND2_X1 U6906 ( .A1(n7982), .A2(n6359), .ZN(n5398) );
  INV_X1 U6907 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7491) );
  OR2_X1 U6908 ( .A1(n6388), .A2(n7491), .ZN(n5396) );
  INV_X1 U6909 ( .A(n5415), .ZN(n5417) );
  NAND2_X1 U6910 ( .A1(n5391), .A2(n7496), .ZN(n5392) );
  NAND2_X1 U6911 ( .A1(n5417), .A2(n5392), .ZN(n7980) );
  OR2_X1 U6912 ( .A1(n5581), .A2(n7980), .ZN(n5395) );
  INV_X1 U6913 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7673) );
  OR2_X1 U6914 ( .A1(n5690), .A2(n7673), .ZN(n5394) );
  NAND2_X1 U6915 ( .A1(n5010), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5393) );
  NAND4_X1 U6916 ( .A1(n5396), .A2(n5395), .A3(n5394), .A4(n5393), .ZN(n9044)
         );
  NAND2_X1 U6917 ( .A1(n9044), .A2(n5114), .ZN(n5397) );
  NAND2_X1 U6918 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  XNOR2_X1 U6919 ( .A(n5399), .B(n7169), .ZN(n7973) );
  INV_X1 U6920 ( .A(n7973), .ZN(n5402) );
  NAND2_X1 U6921 ( .A1(n7982), .A2(n5114), .ZN(n5401) );
  NAND2_X1 U6922 ( .A1(n9044), .A2(n6590), .ZN(n5400) );
  NAND2_X1 U6923 ( .A1(n5401), .A2(n5400), .ZN(n5426) );
  INV_X1 U6924 ( .A(n5426), .ZN(n7972) );
  NAND2_X1 U6925 ( .A1(n5402), .A2(n7972), .ZN(n5431) );
  NAND2_X1 U6926 ( .A1(n5403), .A2(SI_14_), .ZN(n5404) );
  MUX2_X1 U6927 ( .A(n7065), .B(n7063), .S(n4397), .Z(n5407) );
  NAND2_X1 U6928 ( .A1(n5407), .A2(n10088), .ZN(n5433) );
  INV_X1 U6929 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U6930 ( .A1(n5408), .A2(SI_15_), .ZN(n5409) );
  NAND2_X1 U6931 ( .A1(n5433), .A2(n5409), .ZN(n5434) );
  NAND2_X1 U6932 ( .A1(n7062), .A2(n8035), .ZN(n5414) );
  AND2_X1 U6933 ( .A1(n5368), .A2(n5410), .ZN(n5439) );
  OR2_X1 U6934 ( .A1(n5439), .A2(n4595), .ZN(n5411) );
  XNOR2_X1 U6935 ( .A(n5411), .B(n5438), .ZN(n7824) );
  INV_X1 U6936 ( .A(n7824), .ZN(n5412) );
  AOI22_X1 U6937 ( .A1(n5513), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6613), .B2(
        n5412), .ZN(n5413) );
  NAND2_X1 U6938 ( .A1(n9453), .A2(n6359), .ZN(n5424) );
  INV_X1 U6939 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7690) );
  OR2_X1 U6940 ( .A1(n6388), .A2(n7690), .ZN(n5422) );
  NAND2_X1 U6941 ( .A1(n5010), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5421) );
  INV_X1 U6942 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6943 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  NAND2_X1 U6944 ( .A1(n5443), .A2(n5418), .ZN(n9036) );
  OR2_X1 U6945 ( .A1(n5581), .A2(n9036), .ZN(n5420) );
  NAND2_X1 U6946 ( .A1(n7995), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5419) );
  NAND4_X1 U6947 ( .A1(n5422), .A2(n5421), .A3(n5420), .A4(n5419), .ZN(n9043)
         );
  NAND2_X1 U6948 ( .A1(n9043), .A2(n6365), .ZN(n5423) );
  NAND2_X1 U6949 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  XNOR2_X1 U6950 ( .A(n5425), .B(n7169), .ZN(n5430) );
  INV_X1 U6951 ( .A(n5430), .ZN(n5428) );
  AND2_X1 U6952 ( .A1(n7973), .A2(n5426), .ZN(n5432) );
  INV_X1 U6953 ( .A(n5432), .ZN(n5427) );
  NAND2_X1 U6954 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  AOI22_X1 U6955 ( .A1(n9453), .A2(n5114), .B1(n6590), .B2(n9043), .ZN(n9029)
         );
  MUX2_X1 U6956 ( .A(n7154), .B(n10112), .S(n4397), .Z(n5435) );
  NAND2_X1 U6957 ( .A1(n5435), .A2(n10216), .ZN(n5455) );
  INV_X1 U6958 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6959 ( .A1(n5436), .A2(SI_16_), .ZN(n5437) );
  NAND2_X1 U6960 ( .A1(n7081), .A2(n8035), .ZN(n5442) );
  NAND2_X1 U6961 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U6962 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5458) );
  XNOR2_X1 U6963 ( .A(n5458), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9080) );
  AOI22_X1 U6964 ( .A1(n5513), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6613), .B2(
        n9080), .ZN(n5441) );
  NAND2_X1 U6965 ( .A1(n7905), .A2(n6359), .ZN(n5450) );
  INV_X1 U6966 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10136) );
  OR2_X1 U6967 ( .A1(n6388), .A2(n10136), .ZN(n5448) );
  NAND2_X1 U6968 ( .A1(n5010), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5447) );
  OR2_X2 U6969 ( .A1(n5443), .A2(n7829), .ZN(n5464) );
  NAND2_X1 U6970 ( .A1(n5443), .A2(n7829), .ZN(n5444) );
  NAND2_X1 U6971 ( .A1(n5464), .A2(n5444), .ZN(n8956) );
  OR2_X1 U6972 ( .A1(n5581), .A2(n8956), .ZN(n5446) );
  NAND2_X1 U6973 ( .A1(n7995), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5445) );
  NAND4_X1 U6974 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n9364)
         );
  NAND2_X1 U6975 ( .A1(n9364), .A2(n6365), .ZN(n5449) );
  NAND2_X1 U6976 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  XNOR2_X1 U6977 ( .A(n5451), .B(n6362), .ZN(n5474) );
  AND2_X1 U6978 ( .A1(n9364), .A2(n6590), .ZN(n5452) );
  AOI21_X1 U6979 ( .B1(n7905), .B2(n5098), .A(n5452), .ZN(n5473) );
  NOR2_X1 U6980 ( .A1(n5474), .A2(n5473), .ZN(n8948) );
  MUX2_X1 U6981 ( .A(n7158), .B(n10235), .S(n4397), .Z(n5481) );
  XNOR2_X1 U6982 ( .A(n5481), .B(SI_17_), .ZN(n5480) );
  XNOR2_X1 U6983 ( .A(n5485), .B(n5480), .ZN(n7156) );
  NAND2_X1 U6984 ( .A1(n7156), .A2(n8035), .ZN(n5461) );
  NAND2_X1 U6985 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U6986 ( .A1(n5459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U6987 ( .A(n5487), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9098) );
  AOI22_X1 U6988 ( .A1(n5513), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6613), .B2(
        n9098), .ZN(n5460) );
  NAND2_X1 U6989 ( .A1(n9442), .A2(n6359), .ZN(n5471) );
  NAND2_X1 U6990 ( .A1(n5010), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6991 ( .A1(n7995), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5468) );
  INV_X1 U6992 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6993 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6994 ( .A1(n5492), .A2(n5465), .ZN(n9356) );
  OR2_X1 U6995 ( .A1(n5581), .A2(n9356), .ZN(n5467) );
  NAND2_X1 U6996 ( .A1(n7994), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5466) );
  NAND4_X1 U6997 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n9042)
         );
  NAND2_X1 U6998 ( .A1(n9042), .A2(n6365), .ZN(n5470) );
  NAND2_X1 U6999 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  XNOR2_X1 U7000 ( .A(n5472), .B(n7169), .ZN(n5477) );
  AOI22_X1 U7001 ( .A1(n9442), .A2(n5114), .B1(n6590), .B2(n9042), .ZN(n5478)
         );
  XNOR2_X1 U7002 ( .A(n5477), .B(n5478), .ZN(n8963) );
  INV_X1 U7003 ( .A(n8963), .ZN(n5475) );
  OR2_X1 U7004 ( .A1(n8948), .A2(n5475), .ZN(n5476) );
  NAND2_X1 U7005 ( .A1(n5474), .A2(n5473), .ZN(n8960) );
  INV_X1 U7006 ( .A(n5477), .ZN(n5479) );
  NAND2_X1 U7007 ( .A1(n5479), .A2(n5478), .ZN(n5499) );
  NAND2_X1 U7008 ( .A1(n4376), .A2(n5499), .ZN(n8998) );
  INV_X1 U7009 ( .A(n5480), .ZN(n5484) );
  INV_X1 U7010 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U7011 ( .A1(n5482), .A2(SI_17_), .ZN(n5483) );
  MUX2_X1 U7012 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4397), .Z(n5506) );
  XNOR2_X1 U7013 ( .A(n5506), .B(SI_18_), .ZN(n5503) );
  XNOR2_X1 U7014 ( .A(n5505), .B(n5503), .ZN(n7328) );
  NAND2_X1 U7015 ( .A1(n7328), .A2(n8035), .ZN(n5491) );
  NAND2_X1 U7016 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U7017 ( .A1(n5488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5489) );
  XNOR2_X1 U7018 ( .A(n5489), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9111) );
  AOI22_X1 U7019 ( .A1(n5513), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6613), .B2(
        n9111), .ZN(n5490) );
  INV_X1 U7020 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10185) );
  OR2_X1 U7021 ( .A1(n6388), .A2(n10185), .ZN(n5497) );
  NAND2_X1 U7022 ( .A1(n5492), .A2(n10149), .ZN(n5493) );
  NAND2_X1 U7023 ( .A1(n5518), .A2(n5493), .ZN(n9007) );
  OR2_X1 U7024 ( .A1(n5581), .A2(n9007), .ZN(n5496) );
  INV_X1 U7025 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7926) );
  OR2_X1 U7026 ( .A1(n5690), .A2(n7926), .ZN(n5495) );
  NAND2_X1 U7027 ( .A1(n5010), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5494) );
  NAND4_X1 U7028 ( .A1(n5497), .A2(n5496), .A3(n5495), .A4(n5494), .ZN(n9365)
         );
  AOI22_X1 U7029 ( .A1(n9437), .A2(n6359), .B1(n6365), .B2(n9365), .ZN(n5498)
         );
  XNOR2_X1 U7030 ( .A(n5498), .B(n7169), .ZN(n9000) );
  INV_X1 U7031 ( .A(n9000), .ZN(n5500) );
  AOI22_X1 U7032 ( .A1(n9437), .A2(n6365), .B1(n6590), .B2(n9365), .ZN(n8999)
         );
  INV_X1 U7033 ( .A(n5503), .ZN(n5504) );
  NAND2_X1 U7034 ( .A1(n5505), .A2(n5504), .ZN(n5508) );
  NAND2_X1 U7035 ( .A1(n5506), .A2(SI_18_), .ZN(n5507) );
  MUX2_X1 U7036 ( .A(n7433), .B(n7435), .S(n4396), .Z(n5510) );
  NAND2_X1 U7037 ( .A1(n5510), .A2(n5509), .ZN(n5531) );
  INV_X1 U7038 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U7039 ( .A1(n5511), .A2(SI_19_), .ZN(n5512) );
  NAND2_X1 U7040 ( .A1(n5531), .A2(n5512), .ZN(n5532) );
  XNOR2_X1 U7041 ( .A(n5533), .B(n5532), .ZN(n7432) );
  NAND2_X1 U7042 ( .A1(n7432), .A2(n8035), .ZN(n5515) );
  AOI22_X1 U7043 ( .A1(n5513), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9670), .B2(
        n6613), .ZN(n5514) );
  NAND2_X1 U7044 ( .A1(n9434), .A2(n6359), .ZN(n5525) );
  INV_X1 U7045 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7046 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  NAND2_X1 U7047 ( .A1(n5540), .A2(n5519), .ZN(n9341) );
  OR2_X1 U7048 ( .A1(n9341), .A2(n5581), .ZN(n5523) );
  NAND2_X1 U7049 ( .A1(n5010), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7050 ( .A1(n7994), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7051 ( .A1(n7995), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5520) );
  NAND4_X1 U7052 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9322)
         );
  NAND2_X1 U7053 ( .A1(n9322), .A2(n6365), .ZN(n5524) );
  NAND2_X1 U7054 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  XNOR2_X1 U7055 ( .A(n5526), .B(n7169), .ZN(n8918) );
  NAND2_X1 U7056 ( .A1(n9434), .A2(n5114), .ZN(n5528) );
  NAND2_X1 U7057 ( .A1(n9322), .A2(n6590), .ZN(n5527) );
  NAND2_X1 U7058 ( .A1(n5528), .A2(n5527), .ZN(n8919) );
  NAND2_X1 U7059 ( .A1(n8918), .A2(n8919), .ZN(n5530) );
  MUX2_X1 U7060 ( .A(n9970), .B(n7506), .S(n4397), .Z(n5535) );
  NAND2_X1 U7061 ( .A1(n5535), .A2(n5534), .ZN(n5551) );
  INV_X1 U7062 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U7063 ( .A1(n5536), .A2(SI_20_), .ZN(n5537) );
  XNOR2_X1 U7064 ( .A(n5550), .B(n5549), .ZN(n7505) );
  NAND2_X1 U7065 ( .A1(n7505), .A2(n8035), .ZN(n5539) );
  OR2_X1 U7066 ( .A1(n4405), .A2(n7506), .ZN(n5538) );
  NAND2_X1 U7067 ( .A1(n5540), .A2(n8983), .ZN(n5541) );
  NAND2_X1 U7068 ( .A1(n5579), .A2(n5541), .ZN(n9316) );
  NAND2_X1 U7069 ( .A1(n7994), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5543) );
  INV_X1 U7070 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10218) );
  OR2_X1 U7071 ( .A1(n5687), .A2(n10218), .ZN(n5542) );
  AND2_X1 U7072 ( .A1(n5543), .A2(n5542), .ZN(n5545) );
  NAND2_X1 U7073 ( .A1(n7995), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7074 ( .C1(n9316), .C2(n5581), .A(n5545), .B(n5544), .ZN(n9299)
         );
  AOI22_X1 U7075 ( .A1(n9427), .A2(n6359), .B1(n6365), .B2(n9299), .ZN(n5546)
         );
  XNOR2_X1 U7076 ( .A(n5546), .B(n7169), .ZN(n5548) );
  AOI22_X1 U7077 ( .A1(n9427), .A2(n6365), .B1(n6590), .B2(n9299), .ZN(n5547)
         );
  NAND2_X1 U7078 ( .A1(n5548), .A2(n5547), .ZN(n8927) );
  OAI21_X1 U7079 ( .B1(n5548), .B2(n5547), .A(n8927), .ZN(n8982) );
  MUX2_X1 U7080 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4396), .Z(n5566) );
  XNOR2_X1 U7081 ( .A(n5566), .B(n10076), .ZN(n5564) );
  XNOR2_X1 U7082 ( .A(n5563), .B(n5564), .ZN(n7580) );
  NAND2_X1 U7083 ( .A1(n7580), .A2(n8035), .ZN(n5553) );
  INV_X1 U7084 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7611) );
  OR2_X1 U7085 ( .A1(n4405), .A2(n7611), .ZN(n5552) );
  NAND2_X1 U7086 ( .A1(n9422), .A2(n6359), .ZN(n5561) );
  XNOR2_X1 U7087 ( .A(n5579), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U7088 ( .A1(n9304), .A2(n5686), .ZN(n5559) );
  INV_X1 U7089 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7090 ( .A1(n5010), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7091 ( .A1(n7995), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5554) );
  OAI211_X1 U7092 ( .C1(n6388), .C2(n5556), .A(n5555), .B(n5554), .ZN(n5557)
         );
  INV_X1 U7093 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7094 ( .A1(n5559), .A2(n5558), .ZN(n9323) );
  NAND2_X1 U7095 ( .A1(n9323), .A2(n6365), .ZN(n5560) );
  NAND2_X1 U7096 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  XNOR2_X1 U7097 ( .A(n5562), .B(n7169), .ZN(n5587) );
  AOI22_X1 U7098 ( .A1(n9422), .A2(n5114), .B1(n6590), .B2(n9323), .ZN(n5588)
         );
  XNOR2_X1 U7099 ( .A(n5587), .B(n5588), .ZN(n8932) );
  INV_X1 U7100 ( .A(n8932), .ZN(n5586) );
  OR2_X1 U7101 ( .A1(n8982), .A2(n5586), .ZN(n5593) );
  INV_X1 U7102 ( .A(n5563), .ZN(n5565) );
  NAND2_X1 U7103 ( .A1(n5565), .A2(n5564), .ZN(n5568) );
  NAND2_X1 U7104 ( .A1(n5566), .A2(SI_21_), .ZN(n5567) );
  NAND2_X1 U7105 ( .A1(n5568), .A2(n5567), .ZN(n5647) );
  INV_X1 U7106 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7645) );
  MUX2_X1 U7107 ( .A(n7645), .B(n7642), .S(n4396), .Z(n5570) );
  INV_X1 U7108 ( .A(SI_22_), .ZN(n5569) );
  NAND2_X1 U7109 ( .A1(n5570), .A2(n5569), .ZN(n5617) );
  INV_X1 U7110 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7111 ( .A1(n5571), .A2(SI_22_), .ZN(n5572) );
  NAND2_X1 U7112 ( .A1(n5617), .A2(n5572), .ZN(n5615) );
  XNOR2_X1 U7113 ( .A(n5647), .B(n5615), .ZN(n7641) );
  NAND2_X1 U7114 ( .A1(n7641), .A2(n8035), .ZN(n5574) );
  OR2_X1 U7115 ( .A1(n4405), .A2(n7642), .ZN(n5573) );
  INV_X1 U7116 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9287) );
  INV_X1 U7117 ( .A(n5579), .ZN(n5576) );
  AND2_X1 U7118 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5575) );
  INV_X1 U7119 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5578) );
  INV_X1 U7120 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U7121 ( .B1(n5579), .B2(n5578), .A(n5577), .ZN(n5580) );
  NAND2_X1 U7122 ( .A1(n5606), .A2(n5580), .ZN(n9286) );
  OR2_X1 U7123 ( .A1(n9286), .A2(n5581), .ZN(n5583) );
  AOI22_X1 U7124 ( .A1(n7994), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n5010), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5582) );
  OAI211_X1 U7125 ( .C1(n5690), .C2(n9287), .A(n5583), .B(n5582), .ZN(n9300)
         );
  AOI22_X1 U7126 ( .A1(n9417), .A2(n6365), .B1(n6590), .B2(n9300), .ZN(n5584)
         );
  INV_X1 U7127 ( .A(n5584), .ZN(n5594) );
  OR2_X1 U7128 ( .A1(n5593), .A2(n5594), .ZN(n5585) );
  NOR2_X1 U7129 ( .A1(n8926), .A2(n5585), .ZN(n5591) );
  OR2_X1 U7130 ( .A1(n5586), .A2(n8927), .ZN(n8928) );
  INV_X1 U7131 ( .A(n5587), .ZN(n5589) );
  NAND2_X1 U7132 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  AND2_X1 U7133 ( .A1(n8928), .A2(n5590), .ZN(n5595) );
  NOR2_X2 U7134 ( .A1(n5591), .A2(n4444), .ZN(n8989) );
  AOI22_X1 U7135 ( .A1(n9417), .A2(n6359), .B1(n5114), .B2(n9300), .ZN(n5592)
         );
  XOR2_X1 U7136 ( .A(n7169), .B(n5592), .Z(n8992) );
  NAND2_X1 U7137 ( .A1(n8989), .A2(n8992), .ZN(n5638) );
  AND2_X1 U7138 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NAND2_X1 U7139 ( .A1(n8929), .A2(n5596), .ZN(n8990) );
  OR2_X1 U7140 ( .A1(n5647), .A2(n5615), .ZN(n5597) );
  NAND2_X1 U7141 ( .A1(n5597), .A2(n5617), .ZN(n5603) );
  INV_X1 U7142 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5598) );
  MUX2_X1 U7143 ( .A(n5598), .B(n10022), .S(n4397), .Z(n5600) );
  INV_X1 U7144 ( .A(SI_23_), .ZN(n5599) );
  NAND2_X1 U7145 ( .A1(n5600), .A2(n5599), .ZN(n5616) );
  INV_X1 U7146 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7147 ( .A1(n5601), .A2(SI_23_), .ZN(n5614) );
  AND2_X1 U7148 ( .A1(n5616), .A2(n5614), .ZN(n5602) );
  NAND2_X1 U7149 ( .A1(n7721), .A2(n8035), .ZN(n5605) );
  OR2_X1 U7150 ( .A1(n4405), .A2(n10022), .ZN(n5604) );
  NAND2_X1 U7151 ( .A1(n9412), .A2(n6359), .ZN(n5611) );
  OR2_X2 U7152 ( .A1(n5606), .A2(n10099), .ZN(n5626) );
  NAND2_X1 U7153 ( .A1(n5606), .A2(n10099), .ZN(n5607) );
  NAND2_X1 U7154 ( .A1(n5626), .A2(n5607), .ZN(n9275) );
  AOI22_X1 U7155 ( .A1(n7995), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n5010), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7156 ( .A1(n7994), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5608) );
  OAI211_X1 U7157 ( .C1(n9275), .C2(n5581), .A(n5609), .B(n5608), .ZN(n9261)
         );
  NAND2_X1 U7158 ( .A1(n9261), .A2(n6365), .ZN(n5610) );
  NAND2_X1 U7159 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  XNOR2_X1 U7160 ( .A(n5612), .B(n6362), .ZN(n5639) );
  NAND3_X1 U7161 ( .A1(n5638), .A2(n8990), .A3(n5639), .ZN(n8909) );
  INV_X1 U7162 ( .A(n9412), .ZN(n9279) );
  INV_X1 U7163 ( .A(n9261), .ZN(n9294) );
  OAI22_X1 U7164 ( .A1(n9279), .A2(n5187), .B1(n9294), .B2(n5613), .ZN(n8911)
         );
  NAND2_X1 U7165 ( .A1(n8909), .A2(n8911), .ZN(n8969) );
  OR2_X1 U7166 ( .A1(n5647), .A2(n5645), .ZN(n5620) );
  AND2_X1 U7167 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  NAND2_X1 U7168 ( .A1(n5620), .A2(n5648), .ZN(n5621) );
  INV_X1 U7169 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7724) );
  MUX2_X1 U7170 ( .A(n7724), .B(n9958), .S(n4397), .Z(n5643) );
  XNOR2_X1 U7171 ( .A(n5643), .B(SI_24_), .ZN(n5649) );
  NAND2_X1 U7172 ( .A1(n7719), .A2(n8035), .ZN(n5623) );
  OR2_X1 U7173 ( .A1(n4405), .A2(n9958), .ZN(n5622) );
  INV_X1 U7174 ( .A(n5626), .ZN(n5624) );
  INV_X1 U7175 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7176 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U7177 ( .A1(n5658), .A2(n5627), .ZN(n9254) );
  INV_X1 U7178 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7179 ( .A1(n5010), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7180 ( .A1(n7995), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5628) );
  OAI211_X1 U7181 ( .C1(n5630), .C2(n6388), .A(n5629), .B(n5628), .ZN(n5631)
         );
  INV_X1 U7182 ( .A(n5631), .ZN(n5632) );
  AOI22_X1 U7183 ( .A1(n9406), .A2(n6359), .B1(n6365), .B2(n9245), .ZN(n5634)
         );
  XNOR2_X1 U7184 ( .A(n5634), .B(n7169), .ZN(n5636) );
  AOI22_X1 U7185 ( .A1(n9406), .A2(n6365), .B1(n6590), .B2(n9245), .ZN(n5635)
         );
  NAND2_X1 U7186 ( .A1(n5636), .A2(n5635), .ZN(n5642) );
  OAI21_X1 U7187 ( .B1(n5636), .B2(n5635), .A(n5642), .ZN(n8973) );
  INV_X1 U7188 ( .A(n8973), .ZN(n5637) );
  NAND2_X1 U7189 ( .A1(n5638), .A2(n8990), .ZN(n5641) );
  INV_X1 U7190 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7191 ( .A1(n5641), .A2(n5640), .ZN(n8970) );
  INV_X1 U7192 ( .A(n5643), .ZN(n5644) );
  MUX2_X1 U7193 ( .A(n10031), .B(n7944), .S(n4397), .Z(n5653) );
  INV_X1 U7194 ( .A(SI_25_), .ZN(n5652) );
  NAND2_X1 U7195 ( .A1(n5653), .A2(n5652), .ZN(n5676) );
  INV_X1 U7196 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7197 ( .A1(n5654), .A2(SI_25_), .ZN(n5655) );
  NAND2_X1 U7198 ( .A1(n5676), .A2(n5655), .ZN(n5672) );
  NAND2_X1 U7199 ( .A1(n7812), .A2(n8035), .ZN(n5657) );
  OR2_X1 U7200 ( .A1(n4405), .A2(n7944), .ZN(n5656) );
  INV_X1 U7201 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8942) );
  OR2_X2 U7202 ( .A1(n5658), .A2(n8942), .ZN(n5684) );
  NAND2_X1 U7203 ( .A1(n5658), .A2(n8942), .ZN(n5659) );
  NAND2_X1 U7204 ( .A1(n5684), .A2(n5659), .ZN(n9238) );
  INV_X1 U7205 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U7206 ( .A1(n5010), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7207 ( .A1(n7994), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U7208 ( .C1(n5690), .C2(n9973), .A(n5661), .B(n5660), .ZN(n5662)
         );
  INV_X1 U7209 ( .A(n5662), .ZN(n5663) );
  AND2_X1 U7210 ( .A1(n9262), .A2(n6590), .ZN(n5665) );
  AOI21_X1 U7211 ( .B1(n9400), .B2(n5114), .A(n5665), .ZN(n5668) );
  AOI22_X1 U7212 ( .A1(n9400), .A2(n6359), .B1(n6365), .B2(n9262), .ZN(n5666)
         );
  XNOR2_X1 U7213 ( .A(n5666), .B(n7169), .ZN(n5667) );
  XOR2_X1 U7214 ( .A(n5668), .B(n5667), .Z(n8940) );
  INV_X1 U7215 ( .A(n5667), .ZN(n5670) );
  INV_X1 U7216 ( .A(n5668), .ZN(n5669) );
  NOR2_X1 U7217 ( .A1(n5670), .A2(n5669), .ZN(n5700) );
  INV_X1 U7218 ( .A(n5700), .ZN(n5671) );
  INV_X1 U7219 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7814) );
  MUX2_X1 U7220 ( .A(n7814), .B(n7810), .S(n4397), .Z(n5678) );
  INV_X1 U7221 ( .A(SI_26_), .ZN(n5677) );
  NAND2_X1 U7222 ( .A1(n5678), .A2(n5677), .ZN(n6088) );
  INV_X1 U7223 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7224 ( .A1(n5679), .A2(SI_26_), .ZN(n5680) );
  XNOR2_X1 U7225 ( .A(n6087), .B(n6086), .ZN(n7809) );
  NAND2_X1 U7226 ( .A1(n7809), .A2(n8035), .ZN(n5682) );
  OR2_X1 U7227 ( .A1(n4405), .A2(n7810), .ZN(n5681) );
  NAND2_X1 U7228 ( .A1(n9397), .A2(n6359), .ZN(n5696) );
  INV_X1 U7229 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7230 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  NAND2_X1 U7231 ( .A1(n9229), .A2(n5686), .ZN(n5694) );
  INV_X1 U7232 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7233 ( .A1(n7994), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5689) );
  INV_X1 U7234 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10070) );
  OR2_X1 U7235 ( .A1(n5687), .A2(n10070), .ZN(n5688) );
  OAI211_X1 U7236 ( .C1(n5691), .C2(n5690), .A(n5689), .B(n5688), .ZN(n5692)
         );
  INV_X1 U7237 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7238 ( .A1(n9246), .A2(n5114), .ZN(n5695) );
  NAND2_X1 U7239 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  XNOR2_X1 U7240 ( .A(n5697), .B(n6362), .ZN(n6370) );
  AND2_X1 U7241 ( .A1(n9246), .A2(n6590), .ZN(n5698) );
  AOI21_X1 U7242 ( .B1(n9397), .B2(n6365), .A(n5698), .ZN(n6371) );
  XNOR2_X1 U7243 ( .A(n6370), .B(n6371), .ZN(n5701) );
  NOR2_X1 U7244 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  NAND2_X1 U7245 ( .A1(n5704), .A2(P1_B_REG_SCAN_IN), .ZN(n5705) );
  MUX2_X1 U7246 ( .A(n5705), .B(P1_B_REG_SCAN_IN), .S(n5717), .Z(n5706) );
  INV_X1 U7247 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6648) );
  INV_X1 U7248 ( .A(n5707), .ZN(n7811) );
  NOR4_X1 U7249 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5711) );
  NOR4_X1 U7250 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5710) );
  NOR4_X1 U7251 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5709) );
  NOR4_X1 U7252 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5708) );
  NAND4_X1 U7253 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n5716)
         );
  NOR2_X1 U7254 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .ZN(
        n10166) );
  NOR4_X1 U7255 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5714) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5713) );
  NOR4_X1 U7257 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5712) );
  NAND4_X1 U7258 ( .A1(n10166), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n5715)
         );
  NOR2_X1 U7259 ( .A1(n5716), .A2(n5715), .ZN(n6665) );
  NAND2_X1 U7260 ( .A1(n6665), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5718) );
  INV_X1 U7261 ( .A(n5717), .ZN(n7720) );
  NAND2_X1 U7262 ( .A1(n7107), .A2(n6693), .ZN(n5730) );
  NAND2_X1 U7263 ( .A1(n5720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5722) );
  XNOR2_X1 U7264 ( .A(n5722), .B(n5721), .ZN(n7722) );
  AND2_X1 U7265 ( .A1(n7722), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7266 ( .A1(n9742), .A2(n8198), .ZN(n5727) );
  NAND3_X1 U7267 ( .A1(n5730), .A2(n5008), .A3(n6647), .ZN(n5733) );
  NAND2_X1 U7268 ( .A1(n5733), .A2(n7108), .ZN(n6920) );
  AND3_X1 U7269 ( .A1(n5729), .A2(n5719), .A3(n7722), .ZN(n5731) );
  NAND2_X1 U7270 ( .A1(n5730), .A2(n9742), .ZN(n6921) );
  NAND2_X1 U7271 ( .A1(n5731), .A2(n6921), .ZN(n5732) );
  NAND2_X1 U7272 ( .A1(n5732), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5734) );
  INV_X1 U7273 ( .A(n9517), .ZN(n8936) );
  INV_X1 U7274 ( .A(n5736), .ZN(n5735) );
  NAND2_X1 U7275 ( .A1(n5735), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6383) );
  INV_X1 U7276 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U7277 ( .A1(n5736), .A2(n10228), .ZN(n5737) );
  NAND2_X1 U7278 ( .A1(n6383), .A2(n5737), .ZN(n9215) );
  INV_X1 U7279 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7280 ( .A1(n7995), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7281 ( .A1(n5010), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5738) );
  OAI211_X1 U7282 ( .C1(n6388), .C2(n5740), .A(n5739), .B(n5738), .ZN(n5741)
         );
  INV_X1 U7283 ( .A(n5741), .ZN(n5742) );
  NAND2_X2 U7284 ( .A1(n5743), .A2(n5742), .ZN(n9147) );
  INV_X1 U7285 ( .A(n5744), .ZN(n5746) );
  INV_X1 U7286 ( .A(n8260), .ZN(n5745) );
  NAND2_X1 U7287 ( .A1(n5746), .A2(n5745), .ZN(n5749) );
  INV_X1 U7288 ( .A(n5749), .ZN(n5748) );
  AOI22_X1 U7289 ( .A1(n9262), .A2(n9005), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n5750) );
  OAI21_X1 U7290 ( .B1(n9227), .B2(n9003), .A(n5750), .ZN(n5751) );
  AOI21_X1 U7291 ( .B1(n9229), .B2(n8936), .A(n5751), .ZN(n5752) );
  OAI21_X1 U7292 ( .B1(n9232), .B2(n9020), .A(n5752), .ZN(n5753) );
  OAI21_X1 U7293 ( .B1(n5013), .B2(n5755), .A(n5754), .ZN(P1_U3238) );
  INV_X1 U7294 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7295 ( .A1(n4458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  MUX2_X1 U7296 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5767), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5769) );
  NAND2_X1 U7297 ( .A1(n5770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7298 ( .A1(n7526), .A2(n4410), .ZN(n6576) );
  INV_X1 U7299 ( .A(n6576), .ZN(n6354) );
  NAND2_X2 U7300 ( .A1(n6399), .A2(n6354), .ZN(n6529) );
  INV_X1 U7301 ( .A(n7526), .ZN(n6555) );
  NAND2_X1 U7302 ( .A1(n6555), .A2(n6401), .ZN(n7031) );
  NOR2_X1 U7303 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5776) );
  NOR2_X1 U7304 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5775) );
  NOR2_X1 U7305 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5774) );
  NOR2_X1 U7306 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5773) );
  INV_X1 U7307 ( .A(n7019), .ZN(n5798) );
  OR2_X2 U7308 ( .A1(n5790), .A2(n10207), .ZN(n5788) );
  XNOR2_X2 U7309 ( .A(n5788), .B(n5787), .ZN(n6353) );
  INV_X1 U7310 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7311 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5793) );
  XNOR2_X1 U7312 ( .A(n5793), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U7313 ( .A1(n5821), .A2(n6792), .ZN(n5797) );
  INV_X1 U7314 ( .A(n6633), .ZN(n5794) );
  NAND2_X1 U7315 ( .A1(n5874), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7316 ( .A1(n5995), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7317 ( .A1(n4377), .A2(SI_0_), .ZN(n5799) );
  XNOR2_X1 U7318 ( .A(n5799), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U7319 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8895), .S(n4400), .Z(n9837) );
  INV_X1 U7320 ( .A(n9837), .ZN(n7041) );
  NAND2_X1 U7321 ( .A1(n4398), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7322 ( .A1(n4408), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7323 ( .A1(n5827), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7324 ( .A1(n4395), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7325 ( .A1(n6176), .A2(n7044), .ZN(n5805) );
  NAND2_X1 U7326 ( .A1(n5805), .A2(n6203), .ZN(n6205) );
  INV_X1 U7327 ( .A(n6205), .ZN(n7033) );
  NAND2_X1 U7328 ( .A1(n5815), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7329 ( .A1(n5827), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7330 ( .A1(n4395), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5806) );
  INV_X1 U7331 ( .A(n6629), .ZN(n5809) );
  NAND2_X1 U7332 ( .A1(n5874), .A2(n5809), .ZN(n5814) );
  XNOR2_X1 U7333 ( .A(n5811), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U7334 ( .A1(n5821), .A2(n6789), .ZN(n5812) );
  NAND2_X1 U7335 ( .A1(n8505), .A2(n9851), .ZN(n6208) );
  INV_X1 U7336 ( .A(n7021), .ZN(n7034) );
  NAND2_X1 U7337 ( .A1(n7033), .A2(n7034), .ZN(n7069) );
  NAND2_X1 U7338 ( .A1(n7069), .A2(n7068), .ZN(n5826) );
  NAND2_X1 U7339 ( .A1(n4407), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7340 ( .A1(n6079), .A2(n7050), .ZN(n5818) );
  NAND2_X1 U7341 ( .A1(n5827), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7342 ( .A1(n5828), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5816) );
  NAND4_X1 U7343 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n9788)
         );
  INV_X1 U7344 ( .A(n6631), .ZN(n5820) );
  NAND2_X1 U7345 ( .A1(n4382), .A2(n5820), .ZN(n5825) );
  NAND2_X1 U7346 ( .A1(n6093), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7347 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4438), .ZN(n5822) );
  XNOR2_X1 U7348 ( .A(n5822), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U7349 ( .A1(n6658), .A2(n6787), .ZN(n5823) );
  NAND2_X1 U7350 ( .A1(n9788), .A2(n7224), .ZN(n6217) );
  NAND2_X1 U7351 ( .A1(n6198), .A2(n6217), .ZN(n7222) );
  NAND2_X1 U7352 ( .A1(n4407), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5832) );
  XNOR2_X1 U7353 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9792) );
  INV_X1 U7354 ( .A(n9792), .ZN(n7087) );
  NAND2_X1 U7355 ( .A1(n6079), .A2(n7087), .ZN(n5831) );
  NAND2_X1 U7356 ( .A1(n6147), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7357 ( .A1(n5828), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5829) );
  NAND4_X1 U7358 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n8504)
         );
  INV_X1 U7359 ( .A(n6635), .ZN(n5833) );
  NAND2_X1 U7360 ( .A1(n4382), .A2(n5833), .ZN(n5840) );
  NAND2_X1 U7361 ( .A1(n6093), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5839) );
  NOR2_X1 U7362 ( .A1(n5835), .A2(n10207), .ZN(n5836) );
  MUX2_X1 U7363 ( .A(n10207), .B(n5836), .S(P2_IR_REG_4__SCAN_IN), .Z(n5837)
         );
  NOR2_X1 U7364 ( .A1(n5837), .A2(n5858), .ZN(n6795) );
  NAND2_X1 U7365 ( .A1(n6658), .A2(n6795), .ZN(n5838) );
  OR2_X1 U7366 ( .A1(n8504), .A2(n7230), .ZN(n6194) );
  INV_X1 U7367 ( .A(n6194), .ZN(n6199) );
  NAND2_X1 U7368 ( .A1(n8504), .A2(n7230), .ZN(n6218) );
  NAND2_X1 U7369 ( .A1(n6153), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7370 ( .A1(n4407), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5844) );
  AOI21_X1 U7371 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5841) );
  NOR2_X1 U7372 ( .A1(n5841), .A2(n5851), .ZN(n7238) );
  NAND2_X1 U7373 ( .A1(n6079), .A2(n7238), .ZN(n5843) );
  NAND2_X1 U7374 ( .A1(n6147), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5842) );
  NAND4_X1 U7375 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9786)
         );
  INV_X1 U7376 ( .A(n6638), .ZN(n5846) );
  NAND2_X1 U7377 ( .A1(n4382), .A2(n5846), .ZN(n5850) );
  NAND2_X1 U7378 ( .A1(n6093), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7379 ( .A1(n5858), .A2(n10207), .ZN(n5847) );
  XNOR2_X1 U7380 ( .A(n5847), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U7381 ( .A1(n6658), .A2(n6784), .ZN(n5848) );
  NAND2_X1 U7382 ( .A1(n4402), .A2(n7294), .ZN(n6195) );
  INV_X1 U7383 ( .A(n6195), .ZN(n6219) );
  OR2_X1 U7384 ( .A1(n4402), .A2(n7294), .ZN(n6200) );
  NAND2_X1 U7385 ( .A1(n6153), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7386 ( .A1(n4407), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5855) );
  NOR2_X1 U7387 ( .A1(n5851), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5852) );
  NOR2_X1 U7388 ( .A1(n5867), .A2(n5852), .ZN(n7337) );
  NAND2_X1 U7389 ( .A1(n6079), .A2(n7337), .ZN(n5854) );
  NAND2_X1 U7390 ( .A1(n6117), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5853) );
  NAND4_X1 U7391 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n8503)
         );
  INV_X1 U7392 ( .A(n8503), .ZN(n7236) );
  NAND2_X1 U7393 ( .A1(n5858), .A2(n5857), .ZN(n5863) );
  NAND2_X1 U7394 ( .A1(n5863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  INV_X1 U7395 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5859) );
  XNOR2_X1 U7396 ( .A(n5860), .B(n5859), .ZN(n6843) );
  OR2_X1 U7397 ( .A1(n5992), .A2(n6641), .ZN(n5862) );
  NAND2_X1 U7398 ( .A1(n6093), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7399 ( .A1(n7236), .A2(n7298), .ZN(n6223) );
  INV_X1 U7400 ( .A(n7298), .ZN(n9877) );
  NAND2_X1 U7401 ( .A1(n8503), .A2(n9877), .ZN(n6214) );
  AND2_X1 U7402 ( .A1(n6223), .A2(n6214), .ZN(n7341) );
  NAND2_X1 U7403 ( .A1(n7340), .A2(n7341), .ZN(n7339) );
  NAND2_X1 U7404 ( .A1(n7339), .A2(n6223), .ZN(n7301) );
  OR2_X1 U7405 ( .A1(n6644), .A2(n5992), .ZN(n5866) );
  NAND2_X1 U7406 ( .A1(n5875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U7407 ( .A(n5864), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6898) );
  AOI22_X1 U7408 ( .A1(n6093), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4406), .B2(
        n6898), .ZN(n5865) );
  NAND2_X1 U7409 ( .A1(n5866), .A2(n5865), .ZN(n8317) );
  INV_X1 U7410 ( .A(n8317), .ZN(n7964) );
  NAND2_X1 U7411 ( .A1(n6153), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7412 ( .A1(n5974), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5871) );
  NOR2_X1 U7413 ( .A1(n5867), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5868) );
  NOR2_X1 U7414 ( .A1(n5879), .A2(n5868), .ZN(n8316) );
  NAND2_X1 U7415 ( .A1(n6079), .A2(n8316), .ZN(n5870) );
  NAND2_X1 U7416 ( .A1(n6147), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5869) );
  INV_X1 U7417 ( .A(n7400), .ZN(n8502) );
  NAND2_X1 U7418 ( .A1(n7964), .A2(n8502), .ZN(n6228) );
  NAND2_X1 U7419 ( .A1(n7301), .A2(n6228), .ZN(n5873) );
  NAND2_X1 U7420 ( .A1(n7400), .A2(n8317), .ZN(n6227) );
  NAND2_X1 U7421 ( .A1(n5873), .A2(n6227), .ZN(n7949) );
  OR2_X1 U7422 ( .A1(n6649), .A2(n5992), .ZN(n5878) );
  NOR2_X1 U7423 ( .A1(n5875), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7424 ( .A1(n5886), .A2(n10207), .ZN(n5876) );
  XNOR2_X1 U7425 ( .A(n5876), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7426 ( .A1(n6093), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4406), .B2(
        n6961), .ZN(n5877) );
  NAND2_X1 U7427 ( .A1(n5878), .A2(n5877), .ZN(n9881) );
  NAND2_X1 U7428 ( .A1(n6153), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7429 ( .A1(n5974), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7430 ( .A1(n5879), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5901) );
  OAI21_X1 U7431 ( .B1(n5879), .B2(P2_REG3_REG_8__SCAN_IN), .A(n5901), .ZN(
        n7958) );
  INV_X1 U7432 ( .A(n7958), .ZN(n5880) );
  NAND2_X1 U7433 ( .A1(n6079), .A2(n5880), .ZN(n5882) );
  NAND2_X1 U7434 ( .A1(n6117), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5881) );
  OR2_X1 U7435 ( .A1(n9881), .A2(n7318), .ZN(n6232) );
  NAND2_X1 U7436 ( .A1(n9881), .A2(n7318), .ZN(n6233) );
  NAND2_X1 U7437 ( .A1(n6232), .A2(n6233), .ZN(n7948) );
  INV_X1 U7438 ( .A(n7948), .ZN(n7950) );
  NAND2_X1 U7439 ( .A1(n7949), .A2(n7950), .ZN(n5885) );
  NAND2_X1 U7440 ( .A1(n5885), .A2(n6233), .ZN(n7404) );
  NAND2_X1 U7441 ( .A1(n6651), .A2(n4403), .ZN(n5888) );
  NAND2_X1 U7442 ( .A1(n5886), .A2(n10208), .ZN(n5921) );
  NAND2_X1 U7443 ( .A1(n5921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5895) );
  XNOR2_X1 U7444 ( .A(n5895), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7130) );
  AOI22_X1 U7445 ( .A1(n6093), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4406), .B2(
        n7130), .ZN(n5887) );
  NAND2_X1 U7446 ( .A1(n5888), .A2(n5887), .ZN(n7528) );
  NAND2_X1 U7447 ( .A1(n6153), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7448 ( .A1(n5974), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U7449 ( .A(n5901), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U7450 ( .A1(n6079), .A2(n7411), .ZN(n5890) );
  NAND2_X1 U7451 ( .A1(n6147), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5889) );
  OR2_X1 U7452 ( .A1(n7528), .A2(n7533), .ZN(n6236) );
  NAND2_X1 U7453 ( .A1(n7404), .A2(n6236), .ZN(n5893) );
  NAND2_X1 U7454 ( .A1(n7528), .A2(n7533), .ZN(n6234) );
  NAND2_X1 U7455 ( .A1(n6655), .A2(n4403), .ZN(n5898) );
  INV_X1 U7456 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7457 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U7458 ( .A1(n5896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U7459 ( .A(n5908), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7355) );
  AOI22_X1 U7460 ( .A1(n6093), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4406), .B2(
        n7355), .ZN(n5897) );
  NAND2_X1 U7461 ( .A1(n5898), .A2(n5897), .ZN(n8351) );
  NAND2_X1 U7462 ( .A1(n6153), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7463 ( .A1(n5974), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5905) );
  INV_X1 U7464 ( .A(n5901), .ZN(n5899) );
  AOI21_X1 U7465 ( .B1(n5899), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7466 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5900) );
  NOR2_X1 U7467 ( .A1(n5901), .A2(n5900), .ZN(n5913) );
  OR2_X1 U7468 ( .A1(n5902), .A2(n5913), .ZN(n7538) );
  INV_X1 U7469 ( .A(n7538), .ZN(n8350) );
  NAND2_X1 U7470 ( .A1(n6079), .A2(n8350), .ZN(n5904) );
  NAND2_X1 U7471 ( .A1(n6117), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5903) );
  OR2_X1 U7472 ( .A1(n8351), .A2(n8444), .ZN(n6237) );
  NAND2_X1 U7473 ( .A1(n8351), .A2(n8444), .ZN(n7617) );
  NAND2_X1 U7474 ( .A1(n6237), .A2(n7617), .ZN(n7545) );
  INV_X1 U7475 ( .A(n7545), .ZN(n7532) );
  NAND2_X1 U7476 ( .A1(n6678), .A2(n4403), .ZN(n5912) );
  INV_X1 U7477 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7478 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  NAND2_X1 U7479 ( .A1(n5909), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U7480 ( .A(n5910), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U7481 ( .A1(n6093), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4406), .B2(
        n7418), .ZN(n5911) );
  NAND2_X1 U7482 ( .A1(n6153), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7483 ( .A1(n5974), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7484 ( .A1(n5913), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7485 ( .A1(n5913), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5914) );
  AND2_X1 U7486 ( .A1(n5926), .A2(n5914), .ZN(n8448) );
  NAND2_X1 U7487 ( .A1(n6079), .A2(n8448), .ZN(n5916) );
  NAND2_X1 U7488 ( .A1(n6147), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7489 ( .A1(n8449), .A2(n8381), .ZN(n6250) );
  AND2_X1 U7490 ( .A1(n6250), .A2(n7617), .ZN(n6245) );
  NAND2_X1 U7491 ( .A1(n6867), .A2(n4403), .ZN(n5924) );
  INV_X1 U7492 ( .A(n5919), .ZN(n5920) );
  NAND2_X1 U7493 ( .A1(n5932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7494 ( .A(n5922), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U7495 ( .A1(n6093), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4406), .B2(
        n7427), .ZN(n5923) );
  NAND2_X1 U7496 ( .A1(n6153), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7497 ( .A1(n5974), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7498 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  AND2_X1 U7499 ( .A1(n5936), .A2(n5927), .ZN(n8387) );
  NAND2_X1 U7500 ( .A1(n6079), .A2(n8387), .ZN(n5929) );
  NAND2_X1 U7501 ( .A1(n6117), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7502 ( .A1(n8388), .A2(n8432), .ZN(n6253) );
  AND2_X1 U7503 ( .A1(n6253), .A2(n7554), .ZN(n6248) );
  NAND2_X1 U7504 ( .A1(n8388), .A2(n8432), .ZN(n6251) );
  NAND2_X1 U7505 ( .A1(n6913), .A2(n4403), .ZN(n5934) );
  OAI21_X1 U7506 ( .B1(n5932), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5943) );
  XNOR2_X1 U7507 ( .A(n5943), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7589) );
  AOI22_X1 U7508 ( .A1(n6093), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4406), .B2(
        n7589), .ZN(n5933) );
  NAND2_X1 U7509 ( .A1(n6153), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7510 ( .A1(n5974), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5940) );
  AND2_X1 U7511 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NOR2_X1 U7512 ( .A1(n5959), .A2(n5937), .ZN(n8437) );
  NAND2_X1 U7513 ( .A1(n6079), .A2(n8437), .ZN(n5939) );
  NAND2_X1 U7514 ( .A1(n6147), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5938) );
  OR2_X1 U7515 ( .A1(n8866), .A2(n7709), .ZN(n6255) );
  NAND2_X1 U7516 ( .A1(n8866), .A2(n7709), .ZN(n6249) );
  NAND2_X1 U7517 ( .A1(n7782), .A2(n7783), .ZN(n7781) );
  NAND2_X1 U7518 ( .A1(n7781), .A2(n6249), .ZN(n7707) );
  NAND2_X1 U7519 ( .A1(n6933), .A2(n4403), .ZN(n5949) );
  INV_X1 U7520 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7521 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  NAND2_X1 U7522 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7523 ( .A1(n5946), .A2(n5945), .ZN(n5954) );
  OR2_X1 U7524 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  AOI22_X1 U7525 ( .A1(n6093), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4406), .B2(
        n7848), .ZN(n5948) );
  NAND2_X1 U7526 ( .A1(n5974), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5953) );
  INV_X1 U7527 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5960) );
  XNOR2_X1 U7528 ( .A(n5959), .B(n5960), .ZN(n7710) );
  NAND2_X1 U7529 ( .A1(n6079), .A2(n7710), .ZN(n5952) );
  NAND2_X1 U7530 ( .A1(n6117), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7531 ( .A1(n6153), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5950) );
  OR2_X1 U7532 ( .A1(n8277), .A2(n9532), .ZN(n6257) );
  NAND2_X1 U7533 ( .A1(n8277), .A2(n9532), .ZN(n6256) );
  INV_X1 U7534 ( .A(n8278), .ZN(n7706) );
  NAND2_X1 U7535 ( .A1(n7062), .A2(n4403), .ZN(n5957) );
  NAND2_X1 U7536 ( .A1(n5954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  XNOR2_X1 U7537 ( .A(n5955), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7864) );
  AOI22_X1 U7538 ( .A1(n7864), .A2(n4406), .B1(n6093), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7539 ( .A1(n5974), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5967) );
  AND2_X1 U7540 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5958) );
  NAND2_X1 U7541 ( .A1(n5959), .A2(n5958), .ZN(n5976) );
  INV_X1 U7542 ( .A(n5959), .ZN(n5961) );
  INV_X1 U7543 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8270) );
  OAI21_X1 U7544 ( .B1(n5961), .B2(n5960), .A(n8270), .ZN(n5962) );
  NAND2_X1 U7545 ( .A1(n5976), .A2(n5962), .ZN(n9541) );
  INV_X1 U7546 ( .A(n9541), .ZN(n5963) );
  NAND2_X1 U7547 ( .A1(n6079), .A2(n5963), .ZN(n5966) );
  NAND2_X1 U7548 ( .A1(n6147), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7549 ( .A1(n6153), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7550 ( .A1(n8294), .A2(n8280), .ZN(n6261) );
  OR2_X1 U7551 ( .A1(n8294), .A2(n8280), .ZN(n6260) );
  NAND2_X1 U7552 ( .A1(n7081), .A2(n4403), .ZN(n5973) );
  NAND2_X1 U7553 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  MUX2_X1 U7554 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5969), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5971) );
  INV_X1 U7555 ( .A(n5970), .ZN(n5982) );
  AOI22_X1 U7556 ( .A1(n6093), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4406), .B2(
        n8508), .ZN(n5972) );
  NAND2_X1 U7557 ( .A1(n6153), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7558 ( .A1(n5974), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5980) );
  INV_X1 U7559 ( .A(n5976), .ZN(n5975) );
  NAND2_X1 U7560 ( .A1(n5975), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5986) );
  INV_X1 U7561 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U7562 ( .A1(n5976), .A2(n7860), .ZN(n5977) );
  AND2_X1 U7563 ( .A1(n5986), .A2(n5977), .ZN(n8779) );
  NAND2_X1 U7564 ( .A1(n6079), .A2(n8779), .ZN(n5979) );
  NAND2_X1 U7565 ( .A1(n6117), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7566 ( .A1(n8861), .A2(n9534), .ZN(n6265) );
  NAND2_X1 U7567 ( .A1(n8861), .A2(n9534), .ZN(n6264) );
  NAND2_X1 U7568 ( .A1(n7156), .A2(n4403), .ZN(n5985) );
  NAND2_X1 U7569 ( .A1(n5982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7570 ( .A(n5983), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8529) );
  AOI22_X1 U7571 ( .A1(n6093), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4406), .B2(
        n8529), .ZN(n5984) );
  NAND2_X1 U7572 ( .A1(n6153), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7573 ( .A1(n5974), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7574 ( .A1(n5986), .A2(n8516), .ZN(n5987) );
  AND2_X1 U7575 ( .A1(n5999), .A2(n5987), .ZN(n8751) );
  NAND2_X1 U7576 ( .A1(n6079), .A2(n8751), .ZN(n5989) );
  NAND2_X1 U7577 ( .A1(n6117), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7578 ( .A1(n8295), .A2(n8471), .ZN(n6267) );
  NAND2_X1 U7579 ( .A1(n6266), .A2(n6267), .ZN(n8753) );
  NAND2_X1 U7580 ( .A1(n7328), .A2(n4403), .ZN(n5997) );
  NAND2_X1 U7581 ( .A1(n5993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5994) );
  XNOR2_X1 U7582 ( .A(n5994), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8540) );
  AOI22_X1 U7583 ( .A1(n6093), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4406), .B2(
        n8540), .ZN(n5996) );
  NAND2_X1 U7584 ( .A1(n6153), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7585 ( .A1(n5974), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6003) );
  INV_X1 U7586 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U7587 ( .A1(n5999), .A2(n10126), .ZN(n6000) );
  AND2_X1 U7588 ( .A1(n6007), .A2(n6000), .ZN(n8737) );
  NAND2_X1 U7589 ( .A1(n6079), .A2(n8737), .ZN(n6002) );
  NAND2_X1 U7590 ( .A1(n6147), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6001) );
  NAND4_X1 U7591 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n8493)
         );
  INV_X1 U7592 ( .A(n8493), .ZN(n8755) );
  NAND2_X1 U7593 ( .A1(n8852), .A2(n8755), .ZN(n6272) );
  OR2_X1 U7594 ( .A1(n8852), .A2(n8755), .ZN(n6273) );
  NAND2_X1 U7595 ( .A1(n7432), .A2(n4403), .ZN(n6006) );
  AOI22_X1 U7596 ( .A1(n6093), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4625), .B2(
        n4406), .ZN(n6005) );
  NAND2_X1 U7597 ( .A1(n6007), .A2(n8364), .ZN(n6008) );
  AND2_X1 U7598 ( .A1(n6016), .A2(n6008), .ZN(n8728) );
  NAND2_X1 U7599 ( .A1(n8728), .A2(n6079), .ZN(n6012) );
  NAND2_X1 U7600 ( .A1(n5974), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7601 ( .A1(n6153), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7602 ( .A1(n6117), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7603 ( .A1(n8849), .A2(n8425), .ZN(n6279) );
  NAND2_X1 U7604 ( .A1(n8849), .A2(n8425), .ZN(n8710) );
  NAND2_X1 U7605 ( .A1(n7505), .A2(n4403), .ZN(n6014) );
  NAND2_X1 U7606 ( .A1(n6093), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6013) );
  INV_X1 U7607 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U7608 ( .A1(n6016), .A2(n8423), .ZN(n6017) );
  NAND2_X1 U7609 ( .A1(n6026), .A2(n6017), .ZN(n8706) );
  OR2_X1 U7610 ( .A1(n8706), .A2(n6132), .ZN(n6020) );
  AOI22_X1 U7611 ( .A1(n6153), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n5974), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7612 ( .A1(n6147), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7613 ( .A1(n8842), .A2(n8373), .ZN(n6282) );
  NAND2_X1 U7614 ( .A1(n6284), .A2(n6282), .ZN(n8712) );
  INV_X1 U7615 ( .A(n8710), .ZN(n6021) );
  NOR2_X1 U7616 ( .A1(n8712), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U7617 ( .A1(n7580), .A2(n4403), .ZN(n6025) );
  NAND2_X1 U7618 ( .A1(n6093), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6024) );
  INV_X1 U7619 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U7620 ( .A1(n6026), .A2(n8371), .ZN(n6027) );
  NAND2_X1 U7621 ( .A1(n6034), .A2(n6027), .ZN(n8691) );
  AOI22_X1 U7622 ( .A1(n6153), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5974), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7623 ( .A1(n6117), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6028) );
  OAI211_X1 U7624 ( .C1(n8691), .C2(n6132), .A(n6029), .B(n6028), .ZN(n8713)
         );
  INV_X1 U7625 ( .A(n8713), .ZN(n8680) );
  XNOR2_X1 U7626 ( .A(n8837), .B(n8680), .ZN(n8695) );
  NAND2_X1 U7627 ( .A1(n7641), .A2(n4403), .ZN(n6032) );
  NAND2_X1 U7628 ( .A1(n6093), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6031) );
  INV_X1 U7629 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U7630 ( .A1(n6034), .A2(n10196), .ZN(n6035) );
  NAND2_X1 U7631 ( .A1(n6046), .A2(n6035), .ZN(n8672) );
  OR2_X1 U7632 ( .A1(n8672), .A2(n6132), .ZN(n6041) );
  INV_X1 U7633 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7634 ( .A1(n5974), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7635 ( .A1(n6153), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7636 ( .C1(n6135), .C2(n6038), .A(n6037), .B(n6036), .ZN(n6039)
         );
  INV_X1 U7637 ( .A(n6039), .ZN(n6040) );
  OR2_X1 U7638 ( .A1(n8832), .A2(n8372), .ZN(n6053) );
  NAND2_X1 U7639 ( .A1(n8832), .A2(n8372), .ZN(n6288) );
  AND2_X1 U7640 ( .A1(n8837), .A2(n8680), .ZN(n8676) );
  NOR2_X1 U7641 ( .A1(n8669), .A2(n8676), .ZN(n6042) );
  NAND2_X1 U7642 ( .A1(n7721), .A2(n4403), .ZN(n6044) );
  NAND2_X1 U7643 ( .A1(n6093), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6043) );
  INV_X1 U7644 ( .A(n6046), .ZN(n6045) );
  NAND2_X1 U7645 ( .A1(n6045), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6057) );
  INV_X1 U7646 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U7647 ( .A1(n6046), .A2(n10234), .ZN(n6047) );
  NAND2_X1 U7648 ( .A1(n6057), .A2(n6047), .ZN(n8655) );
  OR2_X1 U7649 ( .A1(n8655), .A2(n6132), .ZN(n6052) );
  INV_X1 U7650 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U7651 ( .A1(n6153), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7652 ( .A1(n6147), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U7653 ( .C1(n4409), .C2(n10233), .A(n6049), .B(n6048), .ZN(n6050)
         );
  INV_X1 U7654 ( .A(n6050), .ZN(n6051) );
  OR2_X1 U7655 ( .A1(n8827), .A2(n8681), .ZN(n6295) );
  NAND2_X1 U7656 ( .A1(n8827), .A2(n8681), .ZN(n8643) );
  NAND2_X1 U7657 ( .A1(n6295), .A2(n8643), .ZN(n8659) );
  INV_X1 U7658 ( .A(n6053), .ZN(n8660) );
  NOR2_X1 U7659 ( .A1(n8659), .A2(n8660), .ZN(n6054) );
  NAND2_X1 U7660 ( .A1(n7719), .A2(n4403), .ZN(n6056) );
  NAND2_X1 U7661 ( .A1(n6093), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7662 ( .A1(n6057), .A2(n10225), .ZN(n6058) );
  NAND2_X1 U7663 ( .A1(n6077), .A2(n6058), .ZN(n8638) );
  OR2_X1 U7664 ( .A1(n8638), .A2(n6132), .ZN(n6065) );
  INV_X1 U7665 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7666 ( .A1(n5974), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7667 ( .A1(n6147), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7668 ( .C1(n6062), .C2(n6061), .A(n6060), .B(n6059), .ZN(n6063)
         );
  INV_X1 U7669 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7670 ( .A1(n8822), .A2(n8398), .ZN(n6297) );
  INV_X1 U7671 ( .A(n8643), .ZN(n6290) );
  NOR2_X1 U7672 ( .A1(n8633), .A2(n6290), .ZN(n6066) );
  NAND2_X1 U7673 ( .A1(n8661), .A2(n6066), .ZN(n8647) );
  NAND2_X1 U7674 ( .A1(n8647), .A2(n6296), .ZN(n8623) );
  NAND2_X1 U7675 ( .A1(n7812), .A2(n4403), .ZN(n6068) );
  NAND2_X1 U7676 ( .A1(n6093), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7677 ( .A(n6077), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8627) );
  INV_X1 U7678 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7679 ( .A1(n5828), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7680 ( .A1(n5974), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6069) );
  OAI211_X1 U7681 ( .C1(n6071), .C2(n6135), .A(n6070), .B(n6069), .ZN(n6072)
         );
  AOI21_X1 U7682 ( .B1(n8627), .B2(n6079), .A(n6072), .ZN(n8645) );
  XNOR2_X1 U7683 ( .A(n8818), .B(n8645), .ZN(n8622) );
  INV_X1 U7684 ( .A(n8622), .ZN(n6298) );
  NOR2_X1 U7685 ( .A1(n8818), .A2(n8645), .ZN(n6301) );
  NAND2_X1 U7686 ( .A1(n7809), .A2(n4403), .ZN(n6074) );
  NAND2_X1 U7687 ( .A1(n6093), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6073) );
  INV_X1 U7688 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8397) );
  INV_X1 U7689 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6075) );
  OAI21_X1 U7690 ( .B1(n6077), .B2(n8397), .A(n6075), .ZN(n6078) );
  NAND2_X1 U7691 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n6076) );
  NAND2_X1 U7692 ( .A1(n8611), .A2(n6079), .ZN(n6085) );
  INV_X1 U7693 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7694 ( .A1(n5828), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7695 ( .A1(n5974), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6080) );
  OAI211_X1 U7696 ( .C1(n6082), .C2(n6135), .A(n6081), .B(n6080), .ZN(n6083)
         );
  INV_X1 U7697 ( .A(n6083), .ZN(n6084) );
  OR2_X1 U7698 ( .A1(n8810), .A2(n8400), .ZN(n6304) );
  NAND2_X1 U7699 ( .A1(n8810), .A2(n8400), .ZN(n8585) );
  NAND2_X1 U7700 ( .A1(n6304), .A2(n8585), .ZN(n8595) );
  INV_X1 U7701 ( .A(n8595), .ZN(n8599) );
  INV_X1 U7702 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7842) );
  INV_X1 U7703 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7838) );
  MUX2_X1 U7704 ( .A(n7842), .B(n7838), .S(n4396), .Z(n6090) );
  INV_X1 U7705 ( .A(SI_27_), .ZN(n6089) );
  NAND2_X1 U7706 ( .A1(n6090), .A2(n6089), .ZN(n6108) );
  INV_X1 U7707 ( .A(n6090), .ZN(n6091) );
  NAND2_X1 U7708 ( .A1(n6091), .A2(SI_27_), .ZN(n6092) );
  NAND2_X1 U7709 ( .A1(n7839), .A2(n4403), .ZN(n6095) );
  NAND2_X1 U7710 ( .A1(n6093), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6094) );
  INV_X1 U7711 ( .A(n6097), .ZN(n6096) );
  NAND2_X1 U7712 ( .A1(n6096), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6115) );
  INV_X1 U7713 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U7714 ( .A1(n6097), .A2(n10110), .ZN(n6098) );
  NAND2_X1 U7715 ( .A1(n6115), .A2(n6098), .ZN(n8581) );
  INV_X1 U7716 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7717 ( .A1(n5828), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7718 ( .A1(n5974), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6099) );
  OAI211_X1 U7719 ( .C1(n6101), .C2(n6135), .A(n6100), .B(n6099), .ZN(n6102)
         );
  INV_X1 U7720 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7721 ( .A1(n8804), .A2(n8604), .ZN(n6307) );
  NAND2_X1 U7722 ( .A1(n6308), .A2(n6307), .ZN(n8587) );
  INV_X1 U7723 ( .A(n8587), .ZN(n6306) );
  NAND2_X1 U7724 ( .A1(n6306), .A2(n8585), .ZN(n6105) );
  INV_X1 U7725 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7882) );
  INV_X1 U7726 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U7727 ( .A(n7882), .B(n6110), .S(n4377), .Z(n6127) );
  XNOR2_X1 U7728 ( .A(n6127), .B(SI_28_), .ZN(n6124) );
  NAND2_X1 U7729 ( .A1(n7879), .A2(n4403), .ZN(n6112) );
  NAND2_X1 U7730 ( .A1(n6093), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6111) );
  INV_X1 U7731 ( .A(n6115), .ZN(n6113) );
  NAND2_X1 U7732 ( .A1(n6113), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8296) );
  INV_X1 U7733 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7734 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  NAND2_X1 U7735 ( .A1(n8296), .A2(n6116), .ZN(n6580) );
  INV_X1 U7736 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U7737 ( .A1(n5828), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7738 ( .A1(n6117), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7739 ( .C1(n4409), .C2(n10198), .A(n6119), .B(n6118), .ZN(n6120)
         );
  INV_X1 U7740 ( .A(n6120), .ZN(n6121) );
  NAND2_X1 U7741 ( .A1(n8799), .A2(n8328), .ZN(n6314) );
  INV_X1 U7742 ( .A(n8569), .ZN(n6310) );
  INV_X1 U7743 ( .A(n6313), .ZN(n6123) );
  INV_X1 U7744 ( .A(SI_28_), .ZN(n6126) );
  NAND2_X1 U7745 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  INV_X1 U7746 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8002) );
  INV_X1 U7747 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7934) );
  MUX2_X1 U7748 ( .A(n8002), .B(n7934), .S(n4377), .Z(n6139) );
  XNOR2_X1 U7749 ( .A(n6139), .B(SI_29_), .ZN(n6129) );
  NAND2_X1 U7750 ( .A1(n8001), .A2(n4403), .ZN(n6131) );
  NAND2_X1 U7751 ( .A1(n6093), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6130) );
  OR2_X1 U7752 ( .A1(n8296), .A2(n6132), .ZN(n6138) );
  INV_X1 U7753 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U7754 ( .A1(n5974), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7755 ( .A1(n5828), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6133) );
  OAI211_X1 U7756 ( .C1(n9971), .C2(n6135), .A(n6134), .B(n6133), .ZN(n6136)
         );
  INV_X1 U7757 ( .A(n6136), .ZN(n6137) );
  OR2_X1 U7758 ( .A1(n8794), .A2(n6573), .ZN(n6318) );
  NAND2_X1 U7759 ( .A1(n8794), .A2(n6573), .ZN(n6317) );
  NAND2_X1 U7760 ( .A1(n8301), .A2(n4423), .ZN(n8300) );
  INV_X1 U7761 ( .A(n6139), .ZN(n6140) );
  NOR2_X1 U7762 ( .A1(n6140), .A2(SI_29_), .ZN(n6142) );
  NAND2_X1 U7763 ( .A1(n6140), .A2(SI_29_), .ZN(n6141) );
  INV_X1 U7764 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10227) );
  INV_X1 U7765 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10251) );
  MUX2_X1 U7766 ( .A(n10227), .B(n10251), .S(n4377), .Z(n6161) );
  INV_X1 U7767 ( .A(SI_30_), .ZN(n6144) );
  NAND2_X1 U7768 ( .A1(n8310), .A2(n4403), .ZN(n6146) );
  NAND2_X1 U7769 ( .A1(n6093), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7770 ( .A1(n5974), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7771 ( .A1(n6147), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7772 ( .A1(n5828), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7773 ( .A1(n6681), .A2(n6401), .ZN(n6156) );
  INV_X1 U7774 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U7775 ( .A1(n5974), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7776 ( .A1(n5828), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6154) );
  OAI211_X1 U7777 ( .C1(n6135), .C2(n10007), .A(n6155), .B(n6154), .ZN(n8489)
         );
  NAND2_X1 U7778 ( .A1(n8556), .A2(n8489), .ZN(n6319) );
  INV_X1 U7779 ( .A(n6319), .ZN(n6157) );
  NAND2_X1 U7780 ( .A1(n6159), .A2(n6158), .ZN(n6173) );
  NAND2_X1 U7781 ( .A1(n6160), .A2(SI_30_), .ZN(n6165) );
  INV_X1 U7782 ( .A(n6161), .ZN(n6162) );
  NAND2_X1 U7783 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  NAND2_X1 U7784 ( .A1(n6165), .A2(n6164), .ZN(n6168) );
  MUX2_X1 U7785 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4377), .Z(n6166) );
  XNOR2_X1 U7786 ( .A(n6166), .B(SI_31_), .ZN(n6167) );
  NAND2_X1 U7787 ( .A1(n8888), .A2(n4403), .ZN(n6170) );
  NAND2_X1 U7788 ( .A1(n6093), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6169) );
  OR2_X1 U7789 ( .A1(n8787), .A2(n6681), .ZN(n6328) );
  INV_X1 U7790 ( .A(n8556), .ZN(n8790) );
  INV_X1 U7791 ( .A(n8489), .ZN(n6171) );
  NAND2_X1 U7792 ( .A1(n8790), .A2(n6171), .ZN(n6321) );
  NAND2_X1 U7793 ( .A1(n8787), .A2(n6681), .ZN(n6326) );
  INV_X1 U7794 ( .A(n6326), .ZN(n6172) );
  AOI21_X1 U7795 ( .B1(n6173), .B2(n6322), .A(n6172), .ZN(n6174) );
  XNOR2_X1 U7796 ( .A(n6174), .B(n4625), .ZN(n6175) );
  AOI21_X1 U7797 ( .B1(n6529), .B2(n7031), .A(n6175), .ZN(n6342) );
  NAND2_X1 U7798 ( .A1(n6326), .A2(n6319), .ZN(n6325) );
  INV_X1 U7799 ( .A(n6325), .ZN(n6188) );
  INV_X1 U7800 ( .A(n8659), .ZN(n6291) );
  NAND2_X1 U7801 ( .A1(n6260), .A2(n6261), .ZN(n9524) );
  INV_X1 U7802 ( .A(n7018), .ZN(n6177) );
  NAND3_X1 U7803 ( .A1(n6177), .A2(n4695), .A3(n6555), .ZN(n6178) );
  NAND2_X1 U7804 ( .A1(n6403), .A2(n7041), .ZN(n6202) );
  NAND2_X1 U7805 ( .A1(n7044), .A2(n6202), .ZN(n9838) );
  NOR4_X1 U7806 ( .A1(n6178), .A2(n9803), .A3(n7021), .A4(n9838), .ZN(n6179)
         );
  NAND2_X1 U7807 ( .A1(n6200), .A2(n6195), .ZN(n7292) );
  INV_X1 U7808 ( .A(n7292), .ZN(n7233) );
  NAND4_X1 U7809 ( .A1(n6179), .A2(n7399), .A3(n7341), .A4(n7233), .ZN(n6180)
         );
  NAND2_X1 U7810 ( .A1(n6236), .A2(n6234), .ZN(n7405) );
  NOR4_X1 U7811 ( .A1(n6180), .A2(n7545), .A3(n7405), .A4(n7948), .ZN(n6181)
         );
  NAND4_X1 U7812 ( .A1(n7783), .A2(n7702), .A3(n4899), .A4(n6181), .ZN(n6182)
         );
  NOR4_X1 U7813 ( .A1(n8772), .A2(n9524), .A3(n7706), .A4(n6182), .ZN(n6183)
         );
  NAND4_X1 U7814 ( .A1(n8284), .A2(n8740), .A3(n4744), .A4(n6183), .ZN(n6184)
         );
  NOR4_X1 U7815 ( .A1(n8669), .A2(n8695), .A3(n8712), .A4(n6184), .ZN(n6185)
         );
  NAND4_X1 U7816 ( .A1(n8599), .A2(n8642), .A3(n6291), .A4(n6185), .ZN(n6186)
         );
  NOR4_X1 U7817 ( .A1(n8569), .A2(n8622), .A3(n8587), .A4(n6186), .ZN(n6187)
         );
  NAND4_X1 U7818 ( .A1(n6188), .A2(n6322), .A3(n4423), .A4(n6187), .ZN(n6189)
         );
  XNOR2_X1 U7819 ( .A(n6189), .B(n4410), .ZN(n6190) );
  OAI22_X1 U7820 ( .A1(n6190), .A2(n6401), .B1(n6555), .B2(n7032), .ZN(n6331)
         );
  NAND2_X1 U7821 ( .A1(n6401), .A2(n4625), .ZN(n6192) );
  OR2_X1 U7822 ( .A1(n6191), .A2(n6192), .ZN(n6324) );
  NOR2_X1 U7823 ( .A1(n8622), .A2(n6297), .ZN(n6193) );
  AOI211_X1 U7824 ( .C1(n8645), .C2(n8818), .A(n6193), .B(n8595), .ZN(n6300)
         );
  NOR2_X1 U7825 ( .A1(n8660), .A2(n6324), .ZN(n6294) );
  INV_X1 U7826 ( .A(n6324), .ZN(n6327) );
  NAND2_X1 U7827 ( .A1(n6200), .A2(n6194), .ZN(n6197) );
  NAND2_X1 U7828 ( .A1(n6195), .A2(n6218), .ZN(n6196) );
  NOR2_X1 U7829 ( .A1(n6199), .A2(n4749), .ZN(n6201) );
  OAI211_X1 U7830 ( .C1(n6216), .C2(n6201), .A(n6223), .B(n6200), .ZN(n6213)
         );
  NAND2_X1 U7831 ( .A1(n6203), .A2(n6202), .ZN(n6206) );
  NAND3_X1 U7832 ( .A1(n6206), .A2(n7068), .A3(n6176), .ZN(n6204) );
  AND2_X1 U7833 ( .A1(n6204), .A2(n6208), .ZN(n6211) );
  OAI21_X1 U7834 ( .B1(n6206), .B2(n7581), .A(n6205), .ZN(n6209) );
  INV_X1 U7835 ( .A(n7068), .ZN(n6207) );
  AOI21_X1 U7836 ( .B1(n6209), .B2(n6208), .A(n6207), .ZN(n6210) );
  MUX2_X1 U7837 ( .A(n6211), .B(n6210), .S(n6316), .Z(n6212) );
  INV_X1 U7838 ( .A(n6214), .ZN(n6220) );
  NOR2_X1 U7839 ( .A1(n6215), .A2(n6220), .ZN(n6226) );
  AOI21_X1 U7840 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6221) );
  NOR3_X1 U7841 ( .A1(n6221), .A2(n6220), .A3(n6219), .ZN(n6222) );
  NOR2_X1 U7842 ( .A1(n6222), .A2(n6316), .ZN(n6225) );
  MUX2_X1 U7843 ( .A(n6228), .B(n6227), .S(n6316), .Z(n6229) );
  NAND3_X1 U7844 ( .A1(n6230), .A2(n7950), .A3(n6229), .ZN(n6231) );
  OAI21_X1 U7845 ( .B1(n6327), .B2(n6232), .A(n6231), .ZN(n6240) );
  NAND2_X1 U7846 ( .A1(n6234), .A2(n6233), .ZN(n6239) );
  NAND3_X1 U7847 ( .A1(n6240), .A2(n7617), .A3(n6234), .ZN(n6235) );
  NAND2_X1 U7848 ( .A1(n6235), .A2(n6324), .ZN(n6238) );
  AND2_X1 U7849 ( .A1(n6237), .A2(n6236), .ZN(n6241) );
  OAI211_X1 U7850 ( .C1(n6240), .C2(n6239), .A(n6238), .B(n6241), .ZN(n6247)
         );
  INV_X1 U7851 ( .A(n6241), .ZN(n6243) );
  INV_X1 U7852 ( .A(n7554), .ZN(n6242) );
  AOI21_X1 U7853 ( .B1(n7617), .B2(n6243), .A(n6242), .ZN(n6244) );
  MUX2_X1 U7854 ( .A(n6245), .B(n6244), .S(n6316), .Z(n6246) );
  NAND2_X1 U7855 ( .A1(n6247), .A2(n6246), .ZN(n6252) );
  NAND3_X1 U7856 ( .A1(n6252), .A2(n6251), .A3(n6250), .ZN(n6254) );
  INV_X1 U7857 ( .A(n9524), .ZN(n9529) );
  MUX2_X1 U7858 ( .A(n6257), .B(n6256), .S(n6316), .Z(n6258) );
  NAND3_X1 U7859 ( .A1(n6259), .A2(n9529), .A3(n6258), .ZN(n6263) );
  MUX2_X1 U7860 ( .A(n6261), .B(n6260), .S(n6316), .Z(n6262) );
  MUX2_X1 U7861 ( .A(n6265), .B(n6264), .S(n6316), .Z(n6271) );
  NAND2_X1 U7862 ( .A1(n6273), .A2(n6266), .ZN(n6269) );
  INV_X1 U7863 ( .A(n6267), .ZN(n6268) );
  MUX2_X1 U7864 ( .A(n6269), .B(n6268), .S(n6327), .Z(n6270) );
  INV_X1 U7865 ( .A(n6272), .ZN(n6280) );
  OAI211_X1 U7866 ( .C1(n6274), .C2(n6280), .A(n6279), .B(n6273), .ZN(n6275)
         );
  NAND2_X1 U7867 ( .A1(n6275), .A2(n8710), .ZN(n6277) );
  INV_X1 U7868 ( .A(n6282), .ZN(n6276) );
  AOI211_X1 U7869 ( .C1(n6277), .C2(n6284), .A(n8676), .B(n6276), .ZN(n6278)
         );
  NOR2_X1 U7870 ( .A1(n8837), .A2(n8680), .ZN(n6285) );
  INV_X1 U7871 ( .A(n6296), .ZN(n6293) );
  OAI21_X1 U7872 ( .B1(n6281), .B2(n6280), .A(n6279), .ZN(n6283) );
  NAND3_X1 U7873 ( .A1(n6283), .A2(n6282), .A3(n8710), .ZN(n6287) );
  NOR2_X1 U7874 ( .A1(n6285), .A2(n4761), .ZN(n6286) );
  AOI21_X1 U7875 ( .B1(n6287), .B2(n6286), .A(n8676), .ZN(n6289) );
  OAI211_X1 U7876 ( .C1(n6289), .C2(n8660), .A(n6324), .B(n6288), .ZN(n6292)
         );
  AOI21_X1 U7877 ( .B1(n6296), .B2(n6295), .A(n6324), .ZN(n6299) );
  INV_X1 U7878 ( .A(n6301), .ZN(n6302) );
  AOI21_X1 U7879 ( .B1(n6304), .B2(n6302), .A(n6316), .ZN(n6303) );
  AOI21_X1 U7880 ( .B1(n6305), .B2(n6304), .A(n6303), .ZN(n6312) );
  OAI21_X1 U7881 ( .B1(n8585), .B2(n6324), .A(n6306), .ZN(n6311) );
  MUX2_X1 U7882 ( .A(n6308), .B(n6307), .S(n6316), .Z(n6309) );
  MUX2_X1 U7883 ( .A(n6314), .B(n6313), .S(n6316), .Z(n6315) );
  MUX2_X1 U7884 ( .A(n6318), .B(n6317), .S(n6316), .Z(n6320) );
  NAND3_X1 U7885 ( .A1(n6321), .A2(n6320), .A3(n6319), .ZN(n6323) );
  NOR2_X1 U7886 ( .A1(n6328), .A2(n6327), .ZN(n6329) );
  OAI21_X1 U7887 ( .B1(n6330), .B2(n6329), .A(n7526), .ZN(n6333) );
  INV_X1 U7888 ( .A(n7032), .ZN(n6332) );
  NOR3_X1 U7889 ( .A1(n6333), .A2(n6332), .A3(n6399), .ZN(n6334) );
  OR2_X1 U7890 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  NAND2_X1 U7891 ( .A1(n6343), .A2(n6340), .ZN(n6610) );
  OR2_X1 U7892 ( .A1(n6610), .A2(P2_U3152), .ZN(n6761) );
  NAND2_X1 U7893 ( .A1(n4389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6347) );
  MUX2_X1 U7894 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6347), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6349) );
  NAND2_X1 U7895 ( .A1(n6350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6351) );
  MUX2_X1 U7896 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6351), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6352) );
  NAND2_X1 U7897 ( .A1(n6352), .A2(n4389), .ZN(n7813) );
  NAND2_X1 U7898 ( .A1(n6762), .A2(n6610), .ZN(n6578) );
  INV_X1 U7899 ( .A(n7840), .ZN(n8302) );
  INV_X1 U7900 ( .A(n6353), .ZN(n6571) );
  NAND4_X1 U7901 ( .A1(n7023), .A2(n8302), .A3(n6354), .A4(n9787), .ZN(n6355)
         );
  OAI211_X1 U7902 ( .C1(n6191), .C2(n6761), .A(n6355), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6356) );
  NAND2_X1 U7903 ( .A1(n7839), .A2(n8035), .ZN(n6358) );
  OR2_X1 U7904 ( .A1(n4405), .A2(n7838), .ZN(n6357) );
  NAND2_X1 U7905 ( .A1(n9392), .A2(n6359), .ZN(n6361) );
  NAND2_X1 U7906 ( .A1(n9147), .A2(n5098), .ZN(n6360) );
  NAND2_X1 U7907 ( .A1(n6361), .A2(n6360), .ZN(n6363) );
  XNOR2_X1 U7908 ( .A(n6363), .B(n6362), .ZN(n6367) );
  INV_X1 U7909 ( .A(n6367), .ZN(n6369) );
  AND2_X1 U7910 ( .A1(n9147), .A2(n6590), .ZN(n6364) );
  AOI21_X1 U7911 ( .B1(n9392), .B2(n6365), .A(n6364), .ZN(n6366) );
  INV_X1 U7912 ( .A(n6366), .ZN(n6368) );
  AOI21_X1 U7913 ( .B1(n6369), .B2(n6368), .A(n6593), .ZN(n6377) );
  INV_X1 U7914 ( .A(n6377), .ZN(n6375) );
  INV_X1 U7915 ( .A(n6370), .ZN(n6373) );
  INV_X1 U7916 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U7917 ( .A1(n6373), .A2(n6372), .ZN(n6378) );
  INV_X1 U7918 ( .A(n6378), .ZN(n6374) );
  NOR2_X1 U7919 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  AND2_X2 U7920 ( .A1(n6379), .A2(n6376), .ZN(n6607) );
  AOI21_X1 U7921 ( .B1(n6379), .B2(n6378), .A(n6377), .ZN(n6380) );
  INV_X1 U7922 ( .A(n6383), .ZN(n6381) );
  NAND2_X1 U7923 ( .A1(n6381), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9177) );
  INV_X1 U7924 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7925 ( .A1(n6383), .A2(n6382), .ZN(n6384) );
  NAND2_X1 U7926 ( .A1(n9177), .A2(n6384), .ZN(n9198) );
  INV_X1 U7927 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U7928 ( .A1(n5010), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7929 ( .A1(n7995), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6385) );
  OAI211_X1 U7930 ( .C1(n6388), .C2(n6387), .A(n6386), .B(n6385), .ZN(n6389)
         );
  INV_X1 U7931 ( .A(n6389), .ZN(n6390) );
  NOR2_X1 U7932 ( .A1(n9215), .A2(n9517), .ZN(n6393) );
  OAI22_X1 U7933 ( .A1(n9213), .A2(n9503), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10228), .ZN(n6392) );
  AOI211_X1 U7934 ( .C1(n9500), .C2(n9210), .A(n6393), .B(n6392), .ZN(n6394)
         );
  INV_X1 U7935 ( .A(n6395), .ZN(n6396) );
  NAND2_X1 U7936 ( .A1(n6397), .A2(n6396), .ZN(P1_U3212) );
  INV_X1 U7937 ( .A(n6399), .ZN(n6400) );
  NAND3_X1 U7938 ( .A1(n6400), .A2(n7032), .A3(n7581), .ZN(n6402) );
  NAND2_X1 U7939 ( .A1(n6401), .A2(n7526), .ZN(n7027) );
  INV_X1 U7940 ( .A(n6973), .ZN(n6406) );
  AND2_X1 U7941 ( .A1(n6403), .A2(n9837), .ZN(n7040) );
  NAND2_X1 U7942 ( .A1(n7040), .A2(n6529), .ZN(n6980) );
  NAND2_X1 U7943 ( .A1(n4401), .A2(n7041), .ZN(n6404) );
  NAND2_X1 U7944 ( .A1(n6980), .A2(n6404), .ZN(n6974) );
  NAND2_X1 U7945 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  AND2_X1 U7946 ( .A1(n8505), .A2(n6529), .ZN(n6411) );
  NAND2_X1 U7947 ( .A1(n6410), .A2(n6411), .ZN(n6414) );
  INV_X1 U7948 ( .A(n6410), .ZN(n7053) );
  INV_X1 U7949 ( .A(n6411), .ZN(n6412) );
  NAND2_X1 U7950 ( .A1(n7053), .A2(n6412), .ZN(n6413) );
  AND2_X1 U7951 ( .A1(n6414), .A2(n6413), .ZN(n8457) );
  AND2_X1 U7952 ( .A1(n9788), .A2(n6529), .ZN(n6416) );
  NAND2_X1 U7953 ( .A1(n7084), .A2(n6416), .ZN(n6422) );
  INV_X1 U7954 ( .A(n7084), .ZN(n6418) );
  INV_X1 U7955 ( .A(n6416), .ZN(n6417) );
  NAND2_X1 U7956 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  AND2_X1 U7957 ( .A1(n6422), .A2(n6419), .ZN(n7055) );
  AND2_X1 U7958 ( .A1(n8504), .A2(n6529), .ZN(n6424) );
  XNOR2_X1 U7959 ( .A(n6426), .B(n6424), .ZN(n7083) );
  AND2_X1 U7960 ( .A1(n7083), .A2(n6422), .ZN(n6423) );
  INV_X1 U7961 ( .A(n6424), .ZN(n6425) );
  NAND2_X1 U7962 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  XNOR2_X1 U7963 ( .A(n7294), .B(n4401), .ZN(n7097) );
  AND2_X1 U7964 ( .A1(n9786), .A2(n6529), .ZN(n6428) );
  NAND2_X1 U7965 ( .A1(n7097), .A2(n6428), .ZN(n6433) );
  INV_X1 U7966 ( .A(n7097), .ZN(n6430) );
  INV_X1 U7967 ( .A(n6428), .ZN(n6429) );
  NAND2_X1 U7968 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U7969 ( .A1(n6433), .A2(n6431), .ZN(n7139) );
  XNOR2_X1 U7970 ( .A(n7298), .B(n6538), .ZN(n6435) );
  NAND2_X1 U7971 ( .A1(n8503), .A2(n6529), .ZN(n6436) );
  XNOR2_X1 U7972 ( .A(n6435), .B(n6436), .ZN(n7096) );
  AND2_X1 U7973 ( .A1(n7096), .A2(n6433), .ZN(n6434) );
  INV_X1 U7974 ( .A(n6435), .ZN(n6437) );
  NAND2_X1 U7975 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  AND2_X1 U7976 ( .A1(n7095), .A2(n6438), .ZN(n8313) );
  NOR2_X1 U7977 ( .A1(n7400), .A2(n6979), .ZN(n6440) );
  XNOR2_X1 U7978 ( .A(n8317), .B(n4380), .ZN(n6439) );
  NAND2_X1 U7979 ( .A1(n6440), .A2(n6439), .ZN(n6443) );
  INV_X1 U7980 ( .A(n6439), .ZN(n7278) );
  INV_X1 U7981 ( .A(n6440), .ZN(n6441) );
  NAND2_X1 U7982 ( .A1(n7278), .A2(n6441), .ZN(n6442) );
  AND2_X1 U7983 ( .A1(n6443), .A2(n6442), .ZN(n8312) );
  XNOR2_X1 U7984 ( .A(n9881), .B(n4380), .ZN(n6444) );
  NOR2_X1 U7985 ( .A1(n7318), .A2(n6979), .ZN(n6445) );
  NAND2_X1 U7986 ( .A1(n6444), .A2(n6445), .ZN(n6449) );
  INV_X1 U7987 ( .A(n6444), .ZN(n7314) );
  INV_X1 U7988 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U7989 ( .A1(n7314), .A2(n6446), .ZN(n6447) );
  AND2_X1 U7990 ( .A1(n6449), .A2(n6447), .ZN(n7276) );
  XNOR2_X1 U7991 ( .A(n7528), .B(n4401), .ZN(n6453) );
  NOR2_X1 U7992 ( .A1(n7533), .A2(n6979), .ZN(n6451) );
  XNOR2_X1 U7993 ( .A(n6453), .B(n6451), .ZN(n7326) );
  AND2_X1 U7994 ( .A1(n7326), .A2(n6449), .ZN(n6450) );
  INV_X1 U7995 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U7996 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  XNOR2_X1 U7997 ( .A(n8351), .B(n4380), .ZN(n6455) );
  NOR2_X1 U7998 ( .A1(n8444), .A2(n6979), .ZN(n6456) );
  NAND2_X1 U7999 ( .A1(n6455), .A2(n6456), .ZN(n6460) );
  INV_X1 U8000 ( .A(n6455), .ZN(n8445) );
  INV_X1 U8001 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U8002 ( .A1(n8445), .A2(n6457), .ZN(n6458) );
  NAND2_X1 U8003 ( .A1(n6460), .A2(n6458), .ZN(n8345) );
  XNOR2_X1 U8004 ( .A(n8449), .B(n4380), .ZN(n6461) );
  NOR2_X1 U8005 ( .A1(n8381), .A2(n6979), .ZN(n6462) );
  NAND2_X1 U8006 ( .A1(n6461), .A2(n6462), .ZN(n6466) );
  INV_X1 U8007 ( .A(n6461), .ZN(n8382) );
  INV_X1 U8008 ( .A(n6462), .ZN(n6463) );
  NAND2_X1 U8009 ( .A1(n8382), .A2(n6463), .ZN(n6464) );
  AND2_X1 U8010 ( .A1(n6466), .A2(n6464), .ZN(n8442) );
  NAND2_X1 U8011 ( .A1(n6465), .A2(n8442), .ZN(n8378) );
  NAND2_X1 U8012 ( .A1(n8378), .A2(n6466), .ZN(n6471) );
  XNOR2_X1 U8013 ( .A(n8388), .B(n4380), .ZN(n6467) );
  NOR2_X1 U8014 ( .A1(n8432), .A2(n6979), .ZN(n6468) );
  NAND2_X1 U8015 ( .A1(n6467), .A2(n6468), .ZN(n6472) );
  INV_X1 U8016 ( .A(n6467), .ZN(n8433) );
  INV_X1 U8017 ( .A(n6468), .ZN(n6469) );
  NAND2_X1 U8018 ( .A1(n8433), .A2(n6469), .ZN(n6470) );
  AND2_X1 U8019 ( .A1(n6472), .A2(n6470), .ZN(n8379) );
  NAND2_X1 U8020 ( .A1(n6471), .A2(n8379), .ZN(n8383) );
  NAND2_X1 U8021 ( .A1(n8383), .A2(n6472), .ZN(n6477) );
  XNOR2_X1 U8022 ( .A(n8866), .B(n4380), .ZN(n6473) );
  NOR2_X1 U8023 ( .A1(n7709), .A2(n6979), .ZN(n6474) );
  NAND2_X1 U8024 ( .A1(n6473), .A2(n6474), .ZN(n6478) );
  INV_X1 U8025 ( .A(n6473), .ZN(n7647) );
  INV_X1 U8026 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8027 ( .A1(n7647), .A2(n6475), .ZN(n6476) );
  AND2_X1 U8028 ( .A1(n6478), .A2(n6476), .ZN(n8430) );
  XNOR2_X1 U8029 ( .A(n8277), .B(n4401), .ZN(n6482) );
  NOR2_X1 U8030 ( .A1(n9532), .A2(n6979), .ZN(n6480) );
  XNOR2_X1 U8031 ( .A(n6482), .B(n6480), .ZN(n7658) );
  AND2_X1 U8032 ( .A1(n7658), .A2(n6478), .ZN(n6479) );
  INV_X1 U8033 ( .A(n6480), .ZN(n6481) );
  NAND2_X1 U8034 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  XNOR2_X1 U8035 ( .A(n8294), .B(n4401), .ZN(n6486) );
  NOR2_X1 U8036 ( .A1(n8280), .A2(n6979), .ZN(n6484) );
  INV_X1 U8037 ( .A(n6486), .ZN(n6487) );
  XNOR2_X1 U8038 ( .A(n8861), .B(n4380), .ZN(n6490) );
  NOR2_X1 U8039 ( .A1(n9534), .A2(n6979), .ZN(n6491) );
  XNOR2_X1 U8040 ( .A(n6490), .B(n6491), .ZN(n7885) );
  INV_X1 U8041 ( .A(n6490), .ZN(n6493) );
  INV_X1 U8042 ( .A(n6491), .ZN(n6492) );
  NAND2_X1 U8043 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  XNOR2_X1 U8044 ( .A(n8295), .B(n4380), .ZN(n6495) );
  NOR2_X1 U8045 ( .A1(n8471), .A2(n6979), .ZN(n6496) );
  NAND2_X1 U8046 ( .A1(n6495), .A2(n6496), .ZN(n6499) );
  INV_X1 U8047 ( .A(n6495), .ZN(n8465) );
  INV_X1 U8048 ( .A(n6496), .ZN(n6497) );
  NAND2_X1 U8049 ( .A1(n8465), .A2(n6497), .ZN(n6498) );
  NAND2_X1 U8050 ( .A1(n6499), .A2(n6498), .ZN(n8406) );
  XNOR2_X1 U8051 ( .A(n8852), .B(n4380), .ZN(n6504) );
  NAND2_X1 U8052 ( .A1(n8493), .A2(n6529), .ZN(n6502) );
  XOR2_X1 U8053 ( .A(n6504), .B(n6502), .Z(n8462) );
  OR2_X1 U8054 ( .A1(n8462), .A2(n6499), .ZN(n6500) );
  OAI21_X1 U8055 ( .B1(n8407), .B2(n5016), .A(n6500), .ZN(n6501) );
  INV_X1 U8056 ( .A(n6502), .ZN(n6503) );
  NAND2_X1 U8057 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  XNOR2_X1 U8058 ( .A(n8849), .B(n4380), .ZN(n8357) );
  NOR2_X1 U8059 ( .A1(n8425), .A2(n6979), .ZN(n6506) );
  AND2_X1 U8060 ( .A1(n8357), .A2(n6506), .ZN(n8356) );
  INV_X1 U8061 ( .A(n8357), .ZN(n6508) );
  INV_X1 U8062 ( .A(n6506), .ZN(n6507) );
  NAND2_X1 U8063 ( .A1(n6508), .A2(n6507), .ZN(n8359) );
  XNOR2_X1 U8064 ( .A(n8842), .B(n4401), .ZN(n6509) );
  NAND2_X1 U8065 ( .A1(n8697), .A2(n6529), .ZN(n6510) );
  XNOR2_X1 U8066 ( .A(n6509), .B(n6510), .ZN(n8421) );
  INV_X1 U8067 ( .A(n6509), .ZN(n6512) );
  INV_X1 U8068 ( .A(n6510), .ZN(n6511) );
  NAND2_X1 U8069 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  NAND2_X1 U8070 ( .A1(n6514), .A2(n6513), .ZN(n8370) );
  XNOR2_X1 U8071 ( .A(n8837), .B(n4380), .ZN(n6517) );
  NAND2_X1 U8072 ( .A1(n8713), .A2(n6529), .ZN(n6515) );
  XNOR2_X1 U8073 ( .A(n6517), .B(n6515), .ZN(n8369) );
  INV_X1 U8074 ( .A(n6515), .ZN(n6516) );
  AND2_X1 U8075 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  AOI21_X2 U8076 ( .B1(n8370), .B2(n8369), .A(n6518), .ZN(n6522) );
  XNOR2_X1 U8077 ( .A(n8832), .B(n4401), .ZN(n6521) );
  XNOR2_X2 U8078 ( .A(n6519), .B(n6521), .ZN(n7940) );
  NAND2_X1 U8079 ( .A1(n8698), .A2(n6529), .ZN(n6520) );
  NAND2_X2 U8080 ( .A1(n7940), .A2(n6520), .ZN(n7937) );
  XNOR2_X1 U8081 ( .A(n8827), .B(n4401), .ZN(n8335) );
  OR2_X1 U8082 ( .A1(n8681), .A2(n6979), .ZN(n8338) );
  AND2_X1 U8083 ( .A1(n6522), .A2(n6521), .ZN(n8333) );
  INV_X1 U8084 ( .A(n8335), .ZN(n6524) );
  INV_X1 U8085 ( .A(n8338), .ZN(n6523) );
  AOI21_X2 U8086 ( .B1(n7937), .B2(n6525), .A(n5002), .ZN(n6526) );
  XNOR2_X1 U8087 ( .A(n8822), .B(n4380), .ZN(n6527) );
  XNOR2_X1 U8088 ( .A(n6526), .B(n6527), .ZN(n8414) );
  NOR2_X1 U8089 ( .A1(n8398), .A2(n6979), .ZN(n8413) );
  INV_X1 U8090 ( .A(n6526), .ZN(n6528) );
  XOR2_X1 U8091 ( .A(n4380), .B(n8818), .Z(n8395) );
  INV_X1 U8092 ( .A(n8645), .ZN(n8490) );
  NAND2_X1 U8093 ( .A1(n8490), .A2(n6529), .ZN(n8394) );
  XNOR2_X1 U8094 ( .A(n8810), .B(n4380), .ZN(n8323) );
  NOR2_X1 U8095 ( .A1(n8400), .A2(n6979), .ZN(n6530) );
  NAND2_X1 U8096 ( .A1(n8323), .A2(n6530), .ZN(n6531) );
  OAI21_X1 U8097 ( .B1(n8323), .B2(n6530), .A(n6531), .ZN(n8479) );
  XNOR2_X1 U8098 ( .A(n8804), .B(n4380), .ZN(n6532) );
  NOR2_X1 U8099 ( .A1(n8604), .A2(n6979), .ZN(n6533) );
  NAND2_X1 U8100 ( .A1(n6532), .A2(n6533), .ZN(n6537) );
  INV_X1 U8101 ( .A(n6532), .ZN(n6535) );
  INV_X1 U8102 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U8103 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND2_X1 U8104 ( .A1(n8326), .A2(n6537), .ZN(n6568) );
  INV_X1 U8105 ( .A(n8799), .ZN(n8568) );
  NOR2_X1 U8106 ( .A1(n8328), .A2(n6979), .ZN(n6539) );
  XNOR2_X1 U8107 ( .A(n6539), .B(n4380), .ZN(n6560) );
  INV_X1 U8108 ( .A(n6560), .ZN(n6561) );
  XNOR2_X1 U8109 ( .A(n7726), .B(P2_B_REG_SCAN_IN), .ZN(n6540) );
  INV_X1 U8110 ( .A(n9810), .ZN(n6542) );
  NAND2_X1 U8111 ( .A1(n7813), .A2(n7816), .ZN(n9834) );
  NOR4_X1 U8112 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6549) );
  INV_X1 U8113 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9968) );
  INV_X1 U8114 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10039) );
  INV_X1 U8115 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10138) );
  INV_X1 U8116 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10144) );
  NAND4_X1 U8117 ( .A1(n9968), .A2(n10039), .A3(n10138), .A4(n10144), .ZN(
        n10175) );
  NOR4_X1 U8118 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6546) );
  NOR4_X1 U8119 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6545) );
  NOR4_X1 U8120 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6544) );
  NOR4_X1 U8121 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6543) );
  NAND4_X1 U8122 ( .A1(n6546), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(n6547)
         );
  NOR4_X1 U8123 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        n10175), .A4(n6547), .ZN(n6548) );
  NOR4_X1 U8124 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n10167) );
  NAND3_X1 U8125 ( .A1(n6549), .A2(n6548), .A3(n10167), .ZN(n6550) );
  INV_X1 U8126 ( .A(n7025), .ZN(n6553) );
  NAND2_X1 U8127 ( .A1(n7726), .A2(n7816), .ZN(n9831) );
  INV_X1 U8128 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8129 ( .A1(n9810), .A2(n6551), .ZN(n6552) );
  NAND2_X1 U8130 ( .A1(n6553), .A2(n7309), .ZN(n6554) );
  NOR2_X1 U8131 ( .A1(n7289), .A2(n6554), .ZN(n6574) );
  AND2_X1 U8132 ( .A1(n6399), .A2(n6555), .ZN(n9526) );
  NAND2_X1 U8133 ( .A1(n6569), .A2(n9526), .ZN(n6557) );
  INV_X1 U8134 ( .A(n7288), .ZN(n6556) );
  NOR3_X1 U8135 ( .A1(n8568), .A2(n8455), .A3(n6561), .ZN(n6558) );
  AOI21_X1 U8136 ( .B1(n8568), .B2(n6561), .A(n6558), .ZN(n6567) );
  AND2_X2 U8137 ( .A1(n6399), .A2(n6576), .ZN(n9882) );
  NOR2_X1 U8138 ( .A1(n9882), .A2(n6765), .ZN(n6559) );
  OAI21_X1 U8139 ( .B1(n8568), .B2(n8485), .A(n8478), .ZN(n6566) );
  NOR3_X1 U8140 ( .A1(n8568), .A2(n6560), .A3(n8455), .ZN(n6563) );
  NOR2_X1 U8141 ( .A1(n8799), .A2(n6561), .ZN(n6562) );
  OR2_X1 U8142 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  NAND2_X1 U8143 ( .A1(n6568), .A2(n6564), .ZN(n6565) );
  OAI211_X1 U8144 ( .C1(n6568), .C2(n6567), .A(n6566), .B(n6565), .ZN(n6584)
         );
  INV_X1 U8145 ( .A(n6569), .ZN(n6570) );
  INV_X1 U8146 ( .A(n6765), .ZN(n6572) );
  INV_X1 U8147 ( .A(n6574), .ZN(n6575) );
  NAND2_X1 U8148 ( .A1(n6575), .A2(n7288), .ZN(n6577) );
  NAND2_X1 U8149 ( .A1(n6765), .A2(n6576), .ZN(n7022) );
  NAND2_X1 U8150 ( .A1(n6577), .A2(n7022), .ZN(n6971) );
  OR2_X1 U8151 ( .A1(n6971), .A2(n6578), .ZN(n6579) );
  INV_X1 U8152 ( .A(n6580), .ZN(n8566) );
  AOI22_X1 U8153 ( .A1(n8480), .A2(n8571), .B1(n8481), .B2(n8566), .ZN(n6582)
         );
  AOI22_X1 U8154 ( .A1(n8482), .A2(n8572), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6581) );
  NAND2_X1 U8155 ( .A1(n6584), .A2(n6583), .ZN(P2_U3222) );
  NAND2_X1 U8156 ( .A1(n7879), .A2(n8035), .ZN(n6586) );
  OR2_X1 U8157 ( .A1(n4405), .A2(n7882), .ZN(n6585) );
  NAND2_X1 U8158 ( .A1(n9388), .A2(n6359), .ZN(n6588) );
  NAND2_X1 U8159 ( .A1(n9210), .A2(n5098), .ZN(n6587) );
  NAND2_X1 U8160 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  XNOR2_X1 U8161 ( .A(n6589), .B(n7169), .ZN(n6592) );
  AOI22_X1 U8162 ( .A1(n9388), .A2(n5114), .B1(n6590), .B2(n9210), .ZN(n6591)
         );
  XNOR2_X1 U8163 ( .A(n6592), .B(n6591), .ZN(n6594) );
  OR4_X2 U8164 ( .A1(n6607), .A2(n6593), .A3(n6594), .A4(n9509), .ZN(n6609) );
  AND2_X1 U8165 ( .A1(n6594), .A2(n9016), .ZN(n6606) );
  NAND3_X1 U8166 ( .A1(n6594), .A2(n9016), .A3(n6593), .ZN(n6604) );
  OR2_X1 U8167 ( .A1(n9177), .A2(n5581), .ZN(n6599) );
  NAND2_X1 U8168 ( .A1(n7995), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8169 ( .A1(n7994), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8170 ( .A1(n5010), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6595) );
  AND3_X1 U8171 ( .A1(n6597), .A2(n6596), .A3(n6595), .ZN(n6598) );
  NAND2_X1 U8172 ( .A1(n6599), .A2(n6598), .ZN(n9041) );
  AOI22_X1 U8173 ( .A1(n9041), .A2(n9500), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6601) );
  NAND2_X1 U8174 ( .A1(n9147), .A2(n9005), .ZN(n6600) );
  OAI211_X1 U8175 ( .C1(n9517), .C2(n9198), .A(n6601), .B(n6600), .ZN(n6602)
         );
  AOI21_X1 U8176 ( .B1(n9388), .B2(n9038), .A(n6602), .ZN(n6603) );
  AOI21_X1 U8177 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6608) );
  NAND2_X1 U8178 ( .A1(n6609), .A2(n6608), .ZN(P1_U3218) );
  NAND2_X1 U8179 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6610), .ZN(n9833) );
  INV_X1 U8180 ( .A(n7722), .ZN(n6611) );
  NOR2_X4 U8181 ( .A1(n6683), .A2(P1_U3084), .ZN(P1_U4006) );
  OR2_X1 U8182 ( .A1(n8198), .A2(n6611), .ZN(n6612) );
  NAND2_X1 U8183 ( .A1(n6612), .A2(n6683), .ZN(n6705) );
  OR2_X1 U8184 ( .A1(n6705), .A2(n6613), .ZN(n6614) );
  NAND2_X1 U8185 ( .A1(n6614), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8186 ( .A1(n6615), .A2(n6616), .ZN(n6617) );
  AOI21_X1 U8187 ( .B1(n6618), .B2(n6617), .A(n9509), .ZN(n6623) );
  NOR2_X1 U8188 ( .A1(n9517), .A2(n9666), .ZN(n6622) );
  NAND2_X1 U8189 ( .A1(n9500), .A2(n9665), .ZN(n6619) );
  NAND2_X1 U8190 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U8191 ( .A1(n6619), .A2(n6735), .ZN(n6621) );
  INV_X1 U8192 ( .A(n9052), .ZN(n9684) );
  OAI22_X1 U8193 ( .A1(n9684), .A2(n9503), .B1(n9020), .B2(n9722), .ZN(n6620)
         );
  OR4_X1 U8194 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(P1_U3225)
         );
  NOR2_X1 U8195 ( .A1(n4377), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8892) );
  INV_X2 U8196 ( .A(n8892), .ZN(n8311) );
  NAND2_X1 U8197 ( .A1(n4377), .A2(P2_U3152), .ZN(n8894) );
  INV_X1 U8198 ( .A(n6789), .ZN(n9481) );
  OAI222_X1 U8199 ( .A1(n8311), .A2(n6624), .B1(n8894), .B2(n6629), .C1(
        P2_U3152), .C2(n9481), .ZN(P2_U3356) );
  INV_X1 U8200 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6625) );
  INV_X1 U8201 ( .A(n6792), .ZN(n6866) );
  OAI222_X1 U8202 ( .A1(n8311), .A2(n6625), .B1(n7582), .B2(n6633), .C1(
        P2_U3152), .C2(n6866), .ZN(P2_U3357) );
  INV_X1 U8203 ( .A(n6787), .ZN(n6821) );
  OAI222_X1 U8204 ( .A1(n8311), .A2(n6626), .B1(n8894), .B2(n6631), .C1(
        P2_U3152), .C2(n6821), .ZN(P2_U3355) );
  INV_X1 U8205 ( .A(n6795), .ZN(n6832) );
  OAI222_X1 U8206 ( .A1(n8311), .A2(n6627), .B1(n8894), .B2(n6635), .C1(
        P2_U3152), .C2(n6832), .ZN(P2_U3354) );
  INV_X2 U8207 ( .A(n7878), .ZN(n9479) );
  OAI222_X1 U8208 ( .A1(n7945), .A2(n6630), .B1(n9479), .B2(n6629), .C1(
        P1_U3084), .C2(n9587), .ZN(P1_U3351) );
  OAI222_X1 U8209 ( .A1(n7945), .A2(n6632), .B1(n9479), .B2(n6631), .C1(
        P1_U3084), .C2(n6714), .ZN(P1_U3350) );
  OAI222_X1 U8210 ( .A1(n7945), .A2(n6634), .B1(n9479), .B2(n6633), .C1(
        P1_U3084), .C2(n6710), .ZN(P1_U3352) );
  OAI222_X1 U8211 ( .A1(n7945), .A2(n6636), .B1(P1_U3084), .B2(n9620), .C1(
        n9479), .C2(n6635), .ZN(P1_U3349) );
  INV_X1 U8212 ( .A(n6784), .ZN(n6854) );
  OAI222_X1 U8213 ( .A1(n8311), .A2(n6637), .B1(n7582), .B2(n6638), .C1(
        P2_U3152), .C2(n6854), .ZN(P2_U3353) );
  OAI222_X1 U8214 ( .A1(n7945), .A2(n6639), .B1(n9479), .B2(n6638), .C1(
        P1_U3084), .C2(n6737), .ZN(P1_U3348) );
  OAI222_X1 U8215 ( .A1(n7945), .A2(n6640), .B1(n9479), .B2(n6641), .C1(
        P1_U3084), .C2(n6747), .ZN(P1_U3347) );
  OAI222_X1 U8216 ( .A1(n8311), .A2(n6642), .B1(n7582), .B2(n6641), .C1(
        P2_U3152), .C2(n6843), .ZN(P2_U3352) );
  INV_X1 U8217 ( .A(n6898), .ZN(n6643) );
  OAI222_X1 U8218 ( .A1(n8311), .A2(n10204), .B1(n7582), .B2(n6644), .C1(
        P2_U3152), .C2(n6643), .ZN(P2_U3351) );
  OAI222_X1 U8219 ( .A1(n7945), .A2(n10226), .B1(n9479), .B2(n6644), .C1(
        P1_U3084), .C2(n6748), .ZN(P1_U3346) );
  INV_X1 U8220 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U8221 ( .A1(n9700), .A2(n6645), .B1(n6647), .B2(n6668), .ZN(
        P1_U3440) );
  AOI22_X1 U8222 ( .A1(n9700), .A2(n6648), .B1(n6647), .B2(n6646), .ZN(
        P1_U3441) );
  INV_X1 U8223 ( .A(n6961), .ZN(n6810) );
  OAI222_X1 U8224 ( .A1(n8311), .A2(n10011), .B1(n7582), .B2(n6649), .C1(
        P2_U3152), .C2(n6810), .ZN(P2_U3350) );
  OAI222_X1 U8225 ( .A1(n7945), .A2(n6650), .B1(n9479), .B2(n6649), .C1(
        P1_U3084), .C2(n6902), .ZN(P1_U3345) );
  INV_X1 U8226 ( .A(n6651), .ZN(n6653) );
  OAI222_X1 U8227 ( .A1(n9479), .A2(n6653), .B1(n6652), .B2(P1_U3084), .C1(
        n10209), .C2(n7945), .ZN(P1_U3344) );
  INV_X1 U8228 ( .A(n7130), .ZN(n6970) );
  OAI222_X1 U8229 ( .A1(n8311), .A2(n6654), .B1(n7582), .B2(n6653), .C1(n6970), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8230 ( .A(n6655), .ZN(n6661) );
  INV_X1 U8231 ( .A(n7945), .ZN(n9474) );
  AOI22_X1 U8232 ( .A1(n9655), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9474), .ZN(n6656) );
  OAI21_X1 U8233 ( .B1(n6661), .B2(n9479), .A(n6656), .ZN(P1_U3343) );
  NAND2_X1 U8234 ( .A1(n6341), .A2(n4406), .ZN(n6657) );
  NAND2_X1 U8235 ( .A1(n9809), .A2(n6657), .ZN(n6660) );
  OR2_X1 U8236 ( .A1(n4406), .A2(n6765), .ZN(n6659) );
  NOR2_X1 U8237 ( .A1(n9775), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8238 ( .A(n7355), .ZN(n7137) );
  OAI222_X1 U8239 ( .A1(n8311), .A2(n6662), .B1(n7582), .B2(n6661), .C1(n7137), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8240 ( .A(n7107), .ZN(n6663) );
  NAND2_X1 U8241 ( .A1(n5728), .A2(n9670), .ZN(n9374) );
  AND2_X1 U8242 ( .A1(n6663), .A2(n7109), .ZN(n6664) );
  INV_X1 U8243 ( .A(n6665), .ZN(n6666) );
  NAND2_X1 U8244 ( .A1(n6667), .A2(n6666), .ZN(n6672) );
  INV_X1 U8245 ( .A(n6668), .ZN(n6669) );
  OAI21_X1 U8246 ( .B1(n6670), .B2(P1_D_REG_0__SCAN_IN), .A(n6669), .ZN(n6671)
         );
  INV_X1 U8247 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6677) );
  INV_X1 U8248 ( .A(n7150), .ZN(n7111) );
  AND2_X1 U8249 ( .A1(n7111), .A2(n7117), .ZN(n8208) );
  NOR2_X1 U8250 ( .A1(n7118), .A2(n8208), .ZN(n8011) );
  NAND2_X1 U8251 ( .A1(n8260), .A2(n6936), .ZN(n6673) );
  OR2_X1 U8252 ( .A1(n8011), .A2(n6673), .ZN(n6675) );
  INV_X1 U8253 ( .A(n4378), .ZN(n9606) );
  NAND2_X1 U8254 ( .A1(n9055), .A2(n9664), .ZN(n6674) );
  AND2_X1 U8255 ( .A1(n6675), .A2(n6674), .ZN(n7153) );
  OAI21_X1 U8256 ( .B1(n7111), .B2(n6936), .A(n7153), .ZN(n6695) );
  NAND2_X1 U8257 ( .A1(n6695), .A2(n9759), .ZN(n6676) );
  OAI21_X1 U8258 ( .B1(n9759), .B2(n6677), .A(n6676), .ZN(P1_U3454) );
  INV_X1 U8259 ( .A(n6678), .ZN(n6680) );
  INV_X1 U8260 ( .A(n6991), .ZN(n6885) );
  OAI222_X1 U8261 ( .A1(n9479), .A2(n6680), .B1(n6885), .B2(P1_U3084), .C1(
        n6679), .C2(n7945), .ZN(P1_U3342) );
  INV_X1 U8262 ( .A(n7418), .ZN(n7425) );
  OAI222_X1 U8263 ( .A1(n8311), .A2(n10188), .B1(n7582), .B2(n6680), .C1(n7425), .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8264 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10121) );
  INV_X1 U8265 ( .A(n6681), .ZN(n8551) );
  NAND2_X1 U8266 ( .A1(P2_U3966), .A2(n8551), .ZN(n6682) );
  OAI21_X1 U8267 ( .B1(P2_U3966), .B2(n10121), .A(n6682), .ZN(P2_U3583) );
  INV_X1 U8268 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6692) );
  INV_X1 U8269 ( .A(n6683), .ZN(n6684) );
  INV_X1 U8270 ( .A(n9603), .ZN(n6720) );
  INV_X1 U8271 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6685) );
  AOI21_X1 U8272 ( .B1(n6720), .B2(n6685), .A(n4378), .ZN(n9609) );
  XNOR2_X1 U8273 ( .A(n9609), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6688) );
  OR2_X1 U8274 ( .A1(n4378), .A2(P1_U3084), .ZN(n7880) );
  INV_X1 U8275 ( .A(n7880), .ZN(n6686) );
  INV_X1 U8276 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6697) );
  OR2_X1 U8277 ( .A1(n9603), .A2(P1_U3084), .ZN(n7836) );
  INV_X1 U8278 ( .A(n7836), .ZN(n9108) );
  AOI21_X1 U8279 ( .B1(n6686), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9108), .ZN(
        n6687) );
  NOR3_X1 U8280 ( .A1(n6688), .A2(n6687), .A3(n6705), .ZN(n6689) );
  AOI21_X1 U8281 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6689), .ZN(
        n6691) );
  NOR2_X2 U8282 ( .A1(n6719), .A2(n6720), .ZN(n9653) );
  NAND3_X1 U8283 ( .A1(n9653), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6697), .ZN(
        n6690) );
  OAI211_X1 U8284 ( .C1(n6692), .C2(n9629), .A(n6691), .B(n6690), .ZN(P1_U3241) );
  NAND2_X1 U8285 ( .A1(n6695), .A2(n9772), .ZN(n6696) );
  OAI21_X1 U8286 ( .B1(n9772), .B2(n6697), .A(n6696), .ZN(P1_U3523) );
  INV_X1 U8287 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10012) );
  MUX2_X1 U8288 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10012), .S(n6747), .Z(n6704)
         );
  INV_X1 U8289 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6702) );
  XNOR2_X1 U8290 ( .A(n9587), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9596) );
  XNOR2_X1 U8291 ( .A(n6710), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9060) );
  AND2_X1 U8292 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9059) );
  NAND2_X1 U8293 ( .A1(n9060), .A2(n9059), .ZN(n9058) );
  INV_X1 U8294 ( .A(n6710), .ZN(n9057) );
  NAND2_X1 U8295 ( .A1(n9057), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8296 ( .A1(n9058), .A2(n6698), .ZN(n9595) );
  NAND2_X1 U8297 ( .A1(n9596), .A2(n9595), .ZN(n9594) );
  INV_X1 U8298 ( .A(n9587), .ZN(n9597) );
  NAND2_X1 U8299 ( .A1(n9597), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8300 ( .A1(n9594), .A2(n6699), .ZN(n9070) );
  XNOR2_X1 U8301 ( .A(n6714), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U8302 ( .A1(n9070), .A2(n9071), .ZN(n9069) );
  INV_X1 U8303 ( .A(n6714), .ZN(n9068) );
  NAND2_X1 U8304 ( .A1(n9068), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U8305 ( .A1(n9069), .A2(n6700), .ZN(n9617) );
  XNOR2_X1 U8306 ( .A(n9620), .B(n6701), .ZN(n9616) );
  NOR2_X1 U8307 ( .A1(n9617), .A2(n9616), .ZN(n9619) );
  AOI21_X1 U8308 ( .B1(n9620), .B2(n6701), .A(n9619), .ZN(n6733) );
  XNOR2_X1 U8309 ( .A(n6737), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8310 ( .A1(n6733), .A2(n6734), .ZN(n6732) );
  OAI21_X1 U8311 ( .B1(n6702), .B2(n6737), .A(n6732), .ZN(n6703) );
  NOR2_X1 U8312 ( .A1(n6703), .A2(n6704), .ZN(n6746) );
  AOI21_X1 U8313 ( .B1(n6704), .B2(n6703), .A(n6746), .ZN(n6727) );
  INV_X1 U8314 ( .A(n9653), .ZN(n9115) );
  INV_X1 U8315 ( .A(n6705), .ZN(n9109) );
  NOR2_X1 U8316 ( .A1(n9606), .A2(n7836), .ZN(n6706) );
  INV_X1 U8317 ( .A(n6747), .ZN(n6742) );
  NOR2_X1 U8318 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6707), .ZN(n9018) );
  INV_X1 U8319 ( .A(n6737), .ZN(n6717) );
  INV_X1 U8320 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6708) );
  MUX2_X1 U8321 ( .A(n6708), .B(P1_REG2_REG_2__SCAN_IN), .S(n9587), .Z(n6712)
         );
  INV_X1 U8322 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6709) );
  MUX2_X1 U8323 ( .A(n6709), .B(P1_REG2_REG_1__SCAN_IN), .S(n6710), .Z(n9056)
         );
  AND2_X1 U8324 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9605) );
  NAND2_X1 U8325 ( .A1(n9056), .A2(n9605), .ZN(n9589) );
  OR2_X1 U8326 ( .A1(n6710), .A2(n6709), .ZN(n9588) );
  NAND2_X1 U8327 ( .A1(n9589), .A2(n9588), .ZN(n6711) );
  NAND2_X1 U8328 ( .A1(n6712), .A2(n6711), .ZN(n9592) );
  NAND2_X1 U8329 ( .A1(n9597), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6713) );
  INV_X1 U8330 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6715) );
  MUX2_X1 U8331 ( .A(n6715), .B(P1_REG2_REG_3__SCAN_IN), .S(n6714), .Z(n9067)
         );
  NAND2_X1 U8332 ( .A1(n9068), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6716) );
  INV_X1 U8333 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10205) );
  MUX2_X1 U8334 ( .A(n10205), .B(P1_REG2_REG_4__SCAN_IN), .S(n9620), .Z(n9612)
         );
  AND2_X1 U8335 ( .A1(n9620), .A2(n10205), .ZN(n6728) );
  MUX2_X1 U8336 ( .A(n5166), .B(P1_REG2_REG_5__SCAN_IN), .S(n6737), .Z(n6729)
         );
  OAI21_X1 U8337 ( .B1(n9615), .B2(n6728), .A(n6729), .ZN(n6731) );
  INV_X1 U8338 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6718) );
  MUX2_X1 U8339 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6718), .S(n6747), .Z(n6722)
         );
  INV_X1 U8340 ( .A(n6719), .ZN(n6721) );
  AOI211_X1 U8341 ( .C1(n6723), .C2(n6722), .A(n6741), .B(n9647), .ZN(n6724)
         );
  AOI211_X1 U8342 ( .C1(n9654), .C2(n6742), .A(n9018), .B(n6724), .ZN(n6726)
         );
  NAND2_X1 U8343 ( .A1(n9656), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6725) );
  OAI211_X1 U8344 ( .C1(n6727), .C2(n9115), .A(n6726), .B(n6725), .ZN(P1_U3247) );
  OR3_X1 U8345 ( .A1(n9615), .A2(n6729), .A3(n6728), .ZN(n6730) );
  AOI21_X1 U8346 ( .B1(n6731), .B2(n6730), .A(n9647), .ZN(n6739) );
  INV_X1 U8347 ( .A(n9654), .ZN(n9096) );
  OAI211_X1 U8348 ( .C1(n6734), .C2(n6733), .A(n9653), .B(n6732), .ZN(n6736)
         );
  OAI211_X1 U8349 ( .C1(n9096), .C2(n6737), .A(n6736), .B(n6735), .ZN(n6738)
         );
  AOI211_X1 U8350 ( .C1(P1_ADDR_REG_5__SCAN_IN), .C2(n9656), .A(n6739), .B(
        n6738), .ZN(n6740) );
  INV_X1 U8351 ( .A(n6740), .ZN(P1_U3246) );
  INV_X1 U8352 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6754) );
  INV_X1 U8353 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7216) );
  MUX2_X1 U8354 ( .A(n7216), .B(P1_REG2_REG_7__SCAN_IN), .S(n6748), .Z(n6743)
         );
  OAI21_X1 U8355 ( .B1(n6744), .B2(n6743), .A(n6871), .ZN(n6752) );
  XNOR2_X1 U8356 ( .A(n6748), .B(n6745), .ZN(n6880) );
  AOI21_X1 U8357 ( .B1(n10012), .B2(n6747), .A(n6746), .ZN(n6881) );
  XOR2_X1 U8358 ( .A(n6880), .B(n6881), .Z(n6750) );
  INV_X1 U8359 ( .A(n6748), .ZN(n6879) );
  AND2_X1 U8360 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8901) );
  AOI21_X1 U8361 ( .B1(n9654), .B2(n6879), .A(n8901), .ZN(n6749) );
  OAI21_X1 U8362 ( .B1(n9115), .B2(n6750), .A(n6749), .ZN(n6751) );
  AOI21_X1 U8363 ( .B1(n9593), .B2(n6752), .A(n6751), .ZN(n6753) );
  OAI21_X1 U8364 ( .B1(n9629), .B2(n6754), .A(n6753), .ZN(P1_U3248) );
  INV_X1 U8365 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U8366 ( .A1(n7994), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8367 ( .A1(n7995), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U8368 ( .A1(n5010), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6755) );
  INV_X1 U8369 ( .A(n9127), .ZN(n6758) );
  NAND2_X1 U8370 ( .A1(n6758), .A2(P1_U4006), .ZN(n6759) );
  OAI21_X1 U8371 ( .B1(P1_U4006), .B2(n10151), .A(n6759), .ZN(P1_U3586) );
  INV_X1 U8372 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U8373 ( .A1(n7117), .A2(P1_U4006), .ZN(n6760) );
  OAI21_X1 U8374 ( .B1(P1_U4006), .B2(n10124), .A(n6760), .ZN(P1_U3555) );
  OR2_X1 U8375 ( .A1(n6353), .A2(P2_U3152), .ZN(n7876) );
  OAI21_X1 U8376 ( .B1(n6762), .B2(n7876), .A(n6761), .ZN(n6763) );
  INV_X1 U8377 ( .A(n6763), .ZN(n6764) );
  OAI21_X1 U8378 ( .B1(n9809), .B2(n6765), .A(n6764), .ZN(n6779) );
  NAND2_X1 U8379 ( .A1(n6779), .A2(n4399), .ZN(n6766) );
  NAND2_X1 U8380 ( .A1(n6766), .A2(n8491), .ZN(n6805) );
  INV_X1 U8381 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7284) );
  NOR2_X1 U8382 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7284), .ZN(n6783) );
  INV_X1 U8383 ( .A(n6843), .ZN(n6775) );
  XNOR2_X1 U8384 ( .A(n6795), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8385 ( .A1(n6789), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U8386 ( .B1(n6789), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6767), .ZN(
        n6768) );
  INV_X1 U8387 ( .A(n6768), .ZN(n9483) );
  INV_X1 U8388 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6769) );
  XNOR2_X1 U8389 ( .A(n6792), .B(n6769), .ZN(n6855) );
  NAND2_X1 U8390 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6858) );
  INV_X1 U8391 ( .A(n6858), .ZN(n6770) );
  AND2_X1 U8392 ( .A1(n6855), .A2(n6770), .ZN(n6856) );
  AND2_X1 U8393 ( .A1(n6792), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6771) );
  OR2_X1 U8394 ( .A1(n6856), .A2(n6771), .ZN(n9482) );
  NAND2_X1 U8395 ( .A1(n6787), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6772) );
  OAI21_X1 U8396 ( .B1(n6787), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6772), .ZN(
        n6812) );
  NOR2_X1 U8397 ( .A1(n6823), .A2(n6824), .ZN(n6822) );
  AOI21_X1 U8398 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6795), .A(n6822), .ZN(
        n6846) );
  NAND2_X1 U8399 ( .A1(n6784), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6773) );
  OAI21_X1 U8400 ( .B1(n6784), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6773), .ZN(
        n6845) );
  INV_X1 U8401 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6774) );
  MUX2_X1 U8402 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6774), .S(n6843), .Z(n6834)
         );
  NAND2_X1 U8403 ( .A1(n6898), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6776) );
  OAI21_X1 U8404 ( .B1(n6898), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6776), .ZN(
        n6894) );
  NOR2_X1 U8405 ( .A1(n6895), .A2(n6894), .ZN(n6893) );
  INV_X1 U8406 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6777) );
  MUX2_X1 U8407 ( .A(n6777), .B(P2_REG1_REG_8__SCAN_IN), .S(n6961), .Z(n6780)
         );
  AND2_X1 U8408 ( .A1(n4399), .A2(n7840), .ZN(n6778) );
  AOI211_X1 U8409 ( .C1(n6781), .C2(n6780), .A(n6955), .B(n9778), .ZN(n6782)
         );
  AOI211_X1 U8410 ( .C1(n9775), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6783), .B(
        n6782), .ZN(n6809) );
  NAND2_X1 U8411 ( .A1(n6898), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6801) );
  INV_X1 U8412 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8413 ( .A1(n6784), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6797) );
  INV_X1 U8414 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6785) );
  MUX2_X1 U8415 ( .A(n6785), .B(P2_REG2_REG_5__SCAN_IN), .S(n6784), .Z(n6786)
         );
  INV_X1 U8416 ( .A(n6786), .ZN(n6850) );
  INV_X1 U8417 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U8418 ( .A1(n6787), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6794) );
  INV_X1 U8419 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6788) );
  MUX2_X1 U8420 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6788), .S(n6787), .Z(n6817)
         );
  NAND2_X1 U8421 ( .A1(n6789), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6793) );
  INV_X1 U8422 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6790) );
  MUX2_X1 U8423 ( .A(n6790), .B(P2_REG2_REG_2__SCAN_IN), .S(n6789), .Z(n6791)
         );
  INV_X1 U8424 ( .A(n6791), .ZN(n9487) );
  INV_X1 U8425 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7046) );
  MUX2_X1 U8426 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7046), .S(n6792), .Z(n6862)
         );
  NAND3_X1 U8427 ( .A1(n6862), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6861) );
  OAI21_X1 U8428 ( .B1(n7046), .B2(n6866), .A(n6861), .ZN(n9488) );
  NAND2_X1 U8429 ( .A1(n9487), .A2(n9488), .ZN(n9486) );
  NAND2_X1 U8430 ( .A1(n6793), .A2(n9486), .ZN(n6818) );
  NAND2_X1 U8431 ( .A1(n6817), .A2(n6818), .ZN(n6816) );
  NAND2_X1 U8432 ( .A1(n6794), .A2(n6816), .ZN(n6829) );
  MUX2_X1 U8433 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6796), .S(n6795), .Z(n6828)
         );
  NAND2_X1 U8434 ( .A1(n6829), .A2(n6828), .ZN(n6827) );
  OAI21_X1 U8435 ( .B1(n6796), .B2(n6832), .A(n6827), .ZN(n6851) );
  NAND2_X1 U8436 ( .A1(n6850), .A2(n6851), .ZN(n6849) );
  NAND2_X1 U8437 ( .A1(n6797), .A2(n6849), .ZN(n6840) );
  MUX2_X1 U8438 ( .A(n6798), .B(P2_REG2_REG_6__SCAN_IN), .S(n6843), .Z(n6839)
         );
  NAND2_X1 U8439 ( .A1(n6840), .A2(n6839), .ZN(n6838) );
  OAI21_X1 U8440 ( .B1(n6798), .B2(n6843), .A(n6838), .ZN(n6891) );
  INV_X1 U8441 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10083) );
  MUX2_X1 U8442 ( .A(n10083), .B(P2_REG2_REG_7__SCAN_IN), .S(n6898), .Z(n6892)
         );
  INV_X1 U8443 ( .A(n6892), .ZN(n6799) );
  NAND2_X1 U8444 ( .A1(n6891), .A2(n6799), .ZN(n6800) );
  NAND2_X1 U8445 ( .A1(n6801), .A2(n6800), .ZN(n6807) );
  INV_X1 U8446 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U8447 ( .A(n6802), .B(P2_REG2_REG_8__SCAN_IN), .S(n6961), .Z(n6803)
         );
  INV_X1 U8448 ( .A(n6803), .ZN(n6806) );
  NOR2_X1 U8449 ( .A1(n6353), .A2(n7840), .ZN(n6804) );
  NAND2_X1 U8450 ( .A1(n6806), .A2(n6807), .ZN(n6962) );
  OAI211_X1 U8451 ( .C1(n6807), .C2(n6806), .A(n9774), .B(n6962), .ZN(n6808)
         );
  OAI211_X1 U8452 ( .C1(n9777), .C2(n6810), .A(n6809), .B(n6808), .ZN(P2_U3253) );
  INV_X1 U8453 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7050) );
  NOR2_X1 U8454 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7050), .ZN(n6815) );
  AOI211_X1 U8455 ( .C1(n6813), .C2(n6812), .A(n6811), .B(n9778), .ZN(n6814)
         );
  AOI211_X1 U8456 ( .C1(n9775), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6815), .B(
        n6814), .ZN(n6820) );
  OAI211_X1 U8457 ( .C1(n6818), .C2(n6817), .A(n9774), .B(n6816), .ZN(n6819)
         );
  OAI211_X1 U8458 ( .C1(n9777), .C2(n6821), .A(n6820), .B(n6819), .ZN(P2_U3248) );
  NAND2_X1 U8459 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7088) );
  INV_X1 U8460 ( .A(n7088), .ZN(n6826) );
  AOI211_X1 U8461 ( .C1(n6824), .C2(n6823), .A(n6822), .B(n9778), .ZN(n6825)
         );
  AOI211_X1 U8462 ( .C1(n9775), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6826), .B(
        n6825), .ZN(n6831) );
  OAI211_X1 U8463 ( .C1(n6829), .C2(n6828), .A(n9774), .B(n6827), .ZN(n6830)
         );
  OAI211_X1 U8464 ( .C1(n9777), .C2(n6832), .A(n6831), .B(n6830), .ZN(P2_U3249) );
  NAND2_X1 U8465 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7100) );
  INV_X1 U8466 ( .A(n7100), .ZN(n6837) );
  AOI211_X1 U8467 ( .C1(n6835), .C2(n6834), .A(n6833), .B(n9778), .ZN(n6836)
         );
  AOI211_X1 U8468 ( .C1(n9775), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6837), .B(
        n6836), .ZN(n6842) );
  OAI211_X1 U8469 ( .C1(n6840), .C2(n6839), .A(n9774), .B(n6838), .ZN(n6841)
         );
  OAI211_X1 U8470 ( .C1(n9777), .C2(n6843), .A(n6842), .B(n6841), .ZN(P2_U3251) );
  INV_X1 U8471 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7143) );
  NOR2_X1 U8472 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7143), .ZN(n6848) );
  AOI211_X1 U8473 ( .C1(n6846), .C2(n6845), .A(n6844), .B(n9778), .ZN(n6847)
         );
  AOI211_X1 U8474 ( .C1(n9775), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6848), .B(
        n6847), .ZN(n6853) );
  OAI211_X1 U8475 ( .C1(n6851), .C2(n6850), .A(n9774), .B(n6849), .ZN(n6852)
         );
  OAI211_X1 U8476 ( .C1(n9777), .C2(n6854), .A(n6853), .B(n6852), .ZN(P2_U3250) );
  NOR2_X1 U8477 ( .A1(n4988), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6860) );
  INV_X1 U8478 ( .A(n6855), .ZN(n6857) );
  AOI211_X1 U8479 ( .C1(n6858), .C2(n6857), .A(n6856), .B(n9778), .ZN(n6859)
         );
  AOI211_X1 U8480 ( .C1(n9775), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6860), .B(
        n6859), .ZN(n6865) );
  AND2_X1 U8481 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6863) );
  OAI211_X1 U8482 ( .C1(n6863), .C2(n6862), .A(n9774), .B(n6861), .ZN(n6864)
         );
  OAI211_X1 U8483 ( .C1(n9777), .C2(n6866), .A(n6865), .B(n6864), .ZN(P2_U3246) );
  INV_X1 U8484 ( .A(n6867), .ZN(n6869) );
  INV_X1 U8485 ( .A(n7427), .ZN(n7513) );
  OAI222_X1 U8486 ( .A1(n8311), .A2(n6868), .B1(n7582), .B2(n6869), .C1(
        P2_U3152), .C2(n7513), .ZN(P2_U3346) );
  INV_X1 U8487 ( .A(n7186), .ZN(n6989) );
  OAI222_X1 U8488 ( .A1(n7945), .A2(n6870), .B1(n9479), .B2(n6869), .C1(
        P1_U3084), .C2(n6989), .ZN(P1_U3341) );
  INV_X1 U8489 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6890) );
  OAI21_X1 U8490 ( .B1(n6879), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6871), .ZN(
        n6904) );
  INV_X1 U8491 ( .A(n6902), .ZN(n6909) );
  NAND2_X1 U8492 ( .A1(n6909), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6872) );
  INV_X1 U8493 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U8494 ( .A1(n6904), .A2(n6872), .B1(n10152), .B2(n6902), .ZN(n6873)
         );
  INV_X1 U8495 ( .A(n6873), .ZN(n9635) );
  NAND2_X1 U8496 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9640), .ZN(n6874) );
  OAI21_X1 U8497 ( .B1(n9640), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6874), .ZN(
        n9636) );
  NOR2_X1 U8498 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  AOI21_X1 U8499 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9640), .A(n9634), .ZN(
        n9649) );
  XNOR2_X1 U8500 ( .A(n9655), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9648) );
  NOR2_X1 U8501 ( .A1(n9649), .A2(n9648), .ZN(n9646) );
  AOI22_X1 U8502 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6991), .B1(n6885), .B2(
        n7460), .ZN(n6875) );
  OAI21_X1 U8503 ( .B1(n6876), .B2(n6875), .A(n6990), .ZN(n6877) );
  NAND2_X1 U8504 ( .A1(n6877), .A2(n9593), .ZN(n6889) );
  AOI22_X1 U8505 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6991), .B1(n6885), .B2(
        n5317), .ZN(n6884) );
  INV_X1 U8506 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6878) );
  MUX2_X1 U8507 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6878), .S(n9655), .Z(n9644)
         );
  OAI22_X1 U8508 ( .A1(n6881), .A2(n6880), .B1(n6879), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6906) );
  XNOR2_X1 U8509 ( .A(n6909), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6907) );
  NOR2_X1 U8510 ( .A1(n6906), .A2(n6907), .ZN(n6905) );
  AOI21_X1 U8511 ( .B1(n6909), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6905), .ZN(
        n9633) );
  NOR2_X1 U8512 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9640), .ZN(n6882) );
  AOI21_X1 U8513 ( .B1(n9640), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6882), .ZN(
        n9632) );
  NAND2_X1 U8514 ( .A1(n9633), .A2(n9632), .ZN(n9631) );
  OAI21_X1 U8515 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9640), .A(n9631), .ZN(
        n9645) );
  NAND2_X1 U8516 ( .A1(n9644), .A2(n9645), .ZN(n9643) );
  OAI21_X1 U8517 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9655), .A(n9643), .ZN(
        n6883) );
  NAND2_X1 U8518 ( .A1(n6884), .A2(n6883), .ZN(n6984) );
  OAI21_X1 U8519 ( .B1(n6884), .B2(n6883), .A(n6984), .ZN(n6887) );
  AND2_X1 U8520 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7732) );
  NOR2_X1 U8521 ( .A1(n9096), .A2(n6885), .ZN(n6886) );
  AOI211_X1 U8522 ( .C1(n9653), .C2(n6887), .A(n7732), .B(n6886), .ZN(n6888)
         );
  OAI211_X1 U8523 ( .C1(n9629), .C2(n6890), .A(n6889), .B(n6888), .ZN(P1_U3252) );
  XOR2_X1 U8524 ( .A(n6892), .B(n6891), .Z(n6901) );
  AND2_X1 U8525 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6897) );
  AOI211_X1 U8526 ( .C1(n6895), .C2(n6894), .A(n6893), .B(n9778), .ZN(n6896)
         );
  AOI211_X1 U8527 ( .C1(n9775), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6897), .B(
        n6896), .ZN(n6900) );
  INV_X1 U8528 ( .A(n9777), .ZN(n8534) );
  NAND2_X1 U8529 ( .A1(n8534), .A2(n6898), .ZN(n6899) );
  OAI211_X1 U8530 ( .C1(n6901), .C2(n9776), .A(n6900), .B(n6899), .ZN(P2_U3252) );
  MUX2_X1 U8531 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10152), .S(n6902), .Z(n6903)
         );
  XNOR2_X1 U8532 ( .A(n6904), .B(n6903), .ZN(n6912) );
  NOR2_X1 U8533 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10214), .ZN(n7441) );
  AOI211_X1 U8534 ( .C1(n6907), .C2(n6906), .A(n6905), .B(n9115), .ZN(n6908)
         );
  AOI211_X1 U8535 ( .C1(n9654), .C2(n6909), .A(n7441), .B(n6908), .ZN(n6911)
         );
  NAND2_X1 U8536 ( .A1(n9656), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6910) );
  OAI211_X1 U8537 ( .C1(n6912), .C2(n9647), .A(n6911), .B(n6910), .ZN(P1_U3249) );
  INV_X1 U8538 ( .A(n6913), .ZN(n6924) );
  AOI22_X1 U8539 ( .A1(n7499), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9474), .ZN(n6914) );
  OAI21_X1 U8540 ( .B1(n6924), .B2(n9479), .A(n6914), .ZN(P1_U3340) );
  INV_X1 U8541 ( .A(n6915), .ZN(n6918) );
  INV_X1 U8542 ( .A(n6916), .ZN(n6917) );
  AOI21_X1 U8543 ( .B1(n6919), .B2(n6918), .A(n6917), .ZN(n9604) );
  INV_X1 U8544 ( .A(n6920), .ZN(n9513) );
  NAND2_X1 U8545 ( .A1(n9513), .A2(n6921), .ZN(n7987) );
  AOI22_X1 U8546 ( .A1(n9500), .A2(n9055), .B1(n7987), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8547 ( .A1(n9038), .A2(n7150), .ZN(n6922) );
  OAI211_X1 U8548 ( .C1(n9604), .C2(n9509), .A(n6923), .B(n6922), .ZN(P1_U3230) );
  INV_X1 U8549 ( .A(n7589), .ZN(n7516) );
  OAI222_X1 U8550 ( .A1(n8311), .A2(n6925), .B1(n7582), .B2(n6924), .C1(n7516), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XNOR2_X1 U8551 ( .A(n5014), .B(n6926), .ZN(n6927) );
  XNOR2_X1 U8552 ( .A(n6928), .B(n6927), .ZN(n6932) );
  AOI22_X1 U8553 ( .A1(n9005), .A2(n7117), .B1(n9500), .B2(n9054), .ZN(n6931)
         );
  NAND2_X1 U8554 ( .A1(n7122), .A2(n9727), .ZN(n9701) );
  NOR2_X1 U8555 ( .A1(n7987), .A2(n9701), .ZN(n6929) );
  AOI21_X1 U8556 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7987), .A(n6929), .ZN(
        n6930) );
  OAI211_X1 U8557 ( .C1(n6932), .C2(n9509), .A(n6931), .B(n6930), .ZN(P1_U3220) );
  INV_X1 U8558 ( .A(n6933), .ZN(n6953) );
  INV_X1 U8559 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10206) );
  OAI222_X1 U8560 ( .A1(n9479), .A2(n6953), .B1(n7694), .B2(P1_U3084), .C1(
        n10206), .C2(n7945), .ZN(P1_U3339) );
  OR2_X1 U8561 ( .A1(n7122), .A2(n7150), .ZN(n7110) );
  AND2_X1 U8562 ( .A1(n7110), .A2(n7988), .ZN(n6934) );
  OR2_X1 U8563 ( .A1(n6934), .A2(n9678), .ZN(n7196) );
  INV_X1 U8564 ( .A(n5728), .ZN(n6935) );
  INV_X1 U8565 ( .A(n7988), .ZN(n6937) );
  OAI22_X1 U8566 ( .A1(n7196), .A2(n9753), .B1(n6937), .B2(n9742), .ZN(n6951)
         );
  NAND2_X1 U8567 ( .A1(n9686), .A2(n7988), .ZN(n8212) );
  NAND2_X1 U8568 ( .A1(n6937), .A2(n9054), .ZN(n8214) );
  NAND2_X1 U8569 ( .A1(n6942), .A2(n7118), .ZN(n6939) );
  INV_X1 U8570 ( .A(n7122), .ZN(n8209) );
  OR2_X1 U8571 ( .A1(n9055), .A2(n8209), .ZN(n6938) );
  XNOR2_X1 U8572 ( .A(n4568), .B(n8216), .ZN(n6950) );
  OR2_X1 U8573 ( .A1(n9376), .A2(n9305), .ZN(n6941) );
  OR2_X1 U8574 ( .A1(n5725), .A2(n5728), .ZN(n6940) );
  INV_X1 U8575 ( .A(n6942), .ZN(n6944) );
  NAND2_X1 U8576 ( .A1(n7117), .A2(n7150), .ZN(n7114) );
  NAND2_X1 U8577 ( .A1(n6944), .A2(n6943), .ZN(n7112) );
  NAND2_X1 U8578 ( .A1(n9055), .A2(n7122), .ZN(n6945) );
  XNOR2_X1 U8579 ( .A(n7159), .B(n8010), .ZN(n6947) );
  MUX2_X1 U8580 ( .A(n5726), .B(n6946), .S(n5080), .Z(n9690) );
  INV_X1 U8581 ( .A(n9690), .ZN(n7242) );
  NAND2_X1 U8582 ( .A1(n6947), .A2(n7242), .ZN(n6949) );
  AOI22_X1 U8583 ( .A1(n9363), .A2(n9055), .B1(n9053), .B2(n9664), .ZN(n6948)
         );
  OAI211_X1 U8584 ( .C1(n6950), .C2(n9672), .A(n6949), .B(n6948), .ZN(n7197)
         );
  NOR2_X1 U8585 ( .A1(n6951), .A2(n7197), .ZN(n9708) );
  NAND2_X1 U8586 ( .A1(n9770), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6952) );
  OAI21_X1 U8587 ( .B1(n9708), .B2(n9770), .A(n6952), .ZN(P1_U3525) );
  INV_X1 U8588 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6954) );
  OAI222_X1 U8589 ( .A1(n8311), .A2(n6954), .B1(n7582), .B2(n6953), .C1(n7845), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8590 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7321) );
  INV_X1 U8591 ( .A(n7321), .ZN(n6960) );
  INV_X1 U8592 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6956) );
  MUX2_X1 U8593 ( .A(n6956), .B(P2_REG1_REG_9__SCAN_IN), .S(n7130), .Z(n6957)
         );
  AOI211_X1 U8594 ( .C1(n6958), .C2(n6957), .A(n7125), .B(n9778), .ZN(n6959)
         );
  AOI211_X1 U8595 ( .C1(n9775), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6960), .B(
        n6959), .ZN(n6969) );
  NAND2_X1 U8596 ( .A1(n6961), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8597 ( .A1(n6963), .A2(n6962), .ZN(n6967) );
  INV_X1 U8598 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6964) );
  MUX2_X1 U8599 ( .A(n6964), .B(P2_REG2_REG_9__SCAN_IN), .S(n7130), .Z(n6965)
         );
  INV_X1 U8600 ( .A(n6965), .ZN(n6966) );
  NAND2_X1 U8601 ( .A1(n6966), .A2(n6967), .ZN(n7131) );
  OAI211_X1 U8602 ( .C1(n6967), .C2(n6966), .A(n9774), .B(n7131), .ZN(n6968)
         );
  OAI211_X1 U8603 ( .C1(n9777), .C2(n6970), .A(n6969), .B(n6968), .ZN(P2_U3254) );
  OR2_X1 U8604 ( .A1(n6971), .A2(n9809), .ZN(n8454) );
  NAND2_X1 U8605 ( .A1(n6973), .A2(n6974), .ZN(n6975) );
  AOI21_X1 U8606 ( .B1(n6972), .B2(n6975), .A(n8478), .ZN(n6976) );
  AOI21_X1 U8607 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8454), .A(n6976), .ZN(
        n6978) );
  AOI22_X1 U8608 ( .A1(n8480), .A2(n8505), .B1(n9844), .B2(n8455), .ZN(n6977)
         );
  OAI211_X1 U8609 ( .C1(n5804), .C2(n8472), .A(n6978), .B(n6977), .ZN(P2_U3224) );
  OAI22_X1 U8610 ( .A1(n8464), .A2(n5804), .B1(n7041), .B2(n8478), .ZN(n6981)
         );
  NAND2_X1 U8611 ( .A1(n6981), .A2(n6980), .ZN(n6983) );
  AOI22_X1 U8612 ( .A1(n8455), .A2(n9837), .B1(n8454), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6982) );
  OAI211_X1 U8613 ( .C1(n8424), .C2(n5798), .A(n6983), .B(n6982), .ZN(P2_U3234) );
  INV_X1 U8614 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6999) );
  OAI21_X1 U8615 ( .B1(n6991), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6984), .ZN(
        n6988) );
  NOR2_X1 U8616 ( .A1(n6989), .A2(n6985), .ZN(n6986) );
  AOI21_X1 U8617 ( .B1(n6985), .B2(n6989), .A(n6986), .ZN(n6987) );
  NAND2_X1 U8618 ( .A1(n6987), .A2(n6988), .ZN(n7181) );
  OAI21_X1 U8619 ( .B1(n6988), .B2(n6987), .A(n7181), .ZN(n6997) );
  NAND2_X1 U8620 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9501) );
  OAI21_X1 U8621 ( .B1(n9096), .B2(n6989), .A(n9501), .ZN(n6996) );
  NAND2_X1 U8622 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7186), .ZN(n6992) );
  OAI21_X1 U8623 ( .B1(n7186), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6992), .ZN(
        n6993) );
  AOI211_X1 U8624 ( .C1(n6994), .C2(n6993), .A(n7185), .B(n9647), .ZN(n6995)
         );
  AOI211_X1 U8625 ( .C1(n9653), .C2(n6997), .A(n6996), .B(n6995), .ZN(n6998)
         );
  OAI21_X1 U8626 ( .B1(n9629), .B2(n6999), .A(n6998), .ZN(P1_U3253) );
  INV_X1 U8627 ( .A(n7254), .ZN(n7007) );
  OAI21_X1 U8628 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  NAND2_X1 U8629 ( .A1(n7003), .A2(n9016), .ZN(n7006) );
  AND2_X1 U8630 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9621) );
  INV_X1 U8631 ( .A(n7255), .ZN(n9714) );
  OAI22_X1 U8632 ( .A1(n9003), .A2(n9021), .B1(n9714), .B2(n9020), .ZN(n7004)
         );
  AOI211_X1 U8633 ( .C1(n9005), .C2(n9053), .A(n9621), .B(n7004), .ZN(n7005)
         );
  OAI211_X1 U8634 ( .C1(n9517), .C2(n7007), .A(n7006), .B(n7005), .ZN(P1_U3228) );
  INV_X1 U8635 ( .A(n7008), .ZN(n7013) );
  NOR3_X1 U8636 ( .A1(n7009), .A2(n7011), .A3(n7010), .ZN(n7012) );
  OAI21_X1 U8637 ( .B1(n7013), .B2(n7012), .A(n9016), .ZN(n7017) );
  OAI22_X1 U8638 ( .A1(n9003), .A2(n9684), .B1(n9686), .B2(n9503), .ZN(n7015)
         );
  MUX2_X1 U8639 ( .A(n8936), .B(P1_U3084), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n7014) );
  AOI211_X1 U8640 ( .C1(n9038), .C2(n7160), .A(n7015), .B(n7014), .ZN(n7016)
         );
  NAND2_X1 U8641 ( .A1(n7017), .A2(n7016), .ZN(P1_U3216) );
  NAND2_X1 U8642 ( .A1(n7018), .A2(n7040), .ZN(n7039) );
  NAND2_X1 U8643 ( .A1(n7019), .A2(n9844), .ZN(n7020) );
  OAI21_X1 U8644 ( .B1(n4480), .B2(n7021), .A(n7067), .ZN(n9853) );
  INV_X1 U8645 ( .A(n9853), .ZN(n7038) );
  NAND2_X1 U8646 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8647 ( .A1(n7290), .A2(n7291), .ZN(n7026) );
  XNOR2_X1 U8648 ( .A(n6191), .B(n7027), .ZN(n8762) );
  NAND2_X1 U8649 ( .A1(n8762), .A2(n4410), .ZN(n8774) );
  INV_X1 U8650 ( .A(n7027), .ZN(n7028) );
  NAND2_X1 U8651 ( .A1(n7028), .A2(n4625), .ZN(n7076) );
  NAND2_X1 U8652 ( .A1(n8774), .A2(n7076), .ZN(n9537) );
  NOR2_X1 U8653 ( .A1(n7029), .A2(n4625), .ZN(n7968) );
  INV_X1 U8654 ( .A(n7968), .ZN(n7713) );
  NAND2_X1 U8655 ( .A1(n9841), .A2(n9851), .ZN(n7075) );
  OAI211_X1 U8656 ( .C1(n9841), .C2(n9851), .A(n7075), .B(n9883), .ZN(n9849)
         );
  OAI22_X1 U8657 ( .A1(n7713), .A2(n9849), .B1(n4754), .B2(n9793), .ZN(n7030)
         );
  AOI21_X1 U8658 ( .B1(n8598), .B2(n4751), .A(n7030), .ZN(n7037) );
  OAI21_X1 U8659 ( .B1(n7034), .B2(n7033), .A(n7069), .ZN(n7035) );
  AOI222_X1 U8660 ( .A1(n9790), .A2(n7035), .B1(n8506), .B2(n9787), .C1(n9788), 
        .C2(n9785), .ZN(n9850) );
  MUX2_X1 U8661 ( .A(n6790), .B(n9850), .S(n9791), .Z(n7036) );
  OAI211_X1 U8662 ( .C1(n7038), .C2(n8748), .A(n7037), .B(n7036), .ZN(P2_U3294) );
  OAI21_X1 U8663 ( .B1(n7018), .B2(n7040), .A(n7039), .ZN(n9847) );
  INV_X1 U8664 ( .A(n9521), .ZN(n8560) );
  NOR3_X1 U8665 ( .A1(n8560), .A2(n9841), .A3(n9842), .ZN(n7042) );
  AOI211_X1 U8666 ( .C1(n8778), .C2(P2_REG3_REG_1__SCAN_IN), .A(n7043), .B(
        n7042), .ZN(n7048) );
  XNOR2_X1 U8667 ( .A(n7018), .B(n7044), .ZN(n7045) );
  AOI222_X1 U8668 ( .A1(n9790), .A2(n7045), .B1(n8505), .B2(n9785), .C1(n6403), 
        .C2(n9787), .ZN(n9846) );
  MUX2_X1 U8669 ( .A(n7046), .B(n9846), .S(n9791), .Z(n7047) );
  NAND2_X1 U8670 ( .A1(n7048), .A2(n7047), .ZN(P2_U3295) );
  INV_X1 U8671 ( .A(n7224), .ZN(n9855) );
  NAND2_X1 U8672 ( .A1(n8455), .A2(n9855), .ZN(n7049) );
  OAI21_X1 U8673 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7050), .A(n7049), .ZN(n7052) );
  INV_X1 U8674 ( .A(n8504), .ZN(n7235) );
  OAI22_X1 U8675 ( .A1(n4752), .A2(n8472), .B1(n8424), .B2(n7235), .ZN(n7051)
         );
  AOI211_X1 U8676 ( .C1(n8481), .C2(n7050), .A(n7052), .B(n7051), .ZN(n7061)
         );
  NOR3_X1 U8677 ( .A1(n8464), .A2(n7053), .A3(n4752), .ZN(n7059) );
  INV_X1 U8678 ( .A(n7055), .ZN(n7056) );
  AOI21_X1 U8679 ( .B1(n7054), .B2(n7056), .A(n8478), .ZN(n7058) );
  OAI21_X1 U8680 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7060) );
  NAND2_X1 U8681 ( .A1(n7061), .A2(n7060), .ZN(P2_U3220) );
  INV_X1 U8682 ( .A(n7062), .ZN(n7064) );
  OAI222_X1 U8683 ( .A1(n7945), .A2(n7063), .B1(n9479), .B2(n7064), .C1(
        P1_U3084), .C2(n7824), .ZN(P1_U3338) );
  INV_X1 U8684 ( .A(n7864), .ZN(n7857) );
  OAI222_X1 U8685 ( .A1(n8311), .A2(n7065), .B1(n7582), .B2(n7064), .C1(
        P2_U3152), .C2(n7857), .ZN(P2_U3343) );
  INV_X1 U8686 ( .A(n8774), .ZN(n7409) );
  NAND2_X1 U8687 ( .A1(n4752), .A2(n9851), .ZN(n7066) );
  XNOR2_X1 U8688 ( .A(n7223), .B(n4695), .ZN(n9859) );
  INV_X1 U8689 ( .A(n9859), .ZN(n7074) );
  OAI22_X1 U8690 ( .A1(n4752), .A2(n9533), .B1(n7235), .B2(n9535), .ZN(n7073)
         );
  NAND3_X1 U8691 ( .A1(n7069), .A2(n7068), .A3(n7222), .ZN(n7070) );
  AOI21_X1 U8692 ( .B1(n7071), .B2(n7070), .A(n9531), .ZN(n7072) );
  AOI211_X1 U8693 ( .C1(n7409), .C2(n7074), .A(n7073), .B(n7072), .ZN(n9858)
         );
  OR2_X1 U8694 ( .A1(n7075), .A2(n9855), .ZN(n9795) );
  AOI21_X1 U8695 ( .B1(n9855), .B2(n7075), .A(n4819), .ZN(n9856) );
  OAI22_X1 U8696 ( .A1(n9791), .A2(n6788), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9793), .ZN(n7079) );
  INV_X1 U8697 ( .A(n7076), .ZN(n7077) );
  OAI22_X1 U8698 ( .A1(n8783), .A2(n9859), .B1(n7224), .B2(n8781), .ZN(n7078)
         );
  AOI211_X1 U8699 ( .C1(n9521), .C2(n9856), .A(n7079), .B(n7078), .ZN(n7080)
         );
  OAI21_X1 U8700 ( .B1(n9808), .B2(n9858), .A(n7080), .ZN(P2_U3293) );
  INV_X1 U8701 ( .A(n7081), .ZN(n7155) );
  INV_X1 U8702 ( .A(n9080), .ZN(n7832) );
  OAI222_X1 U8703 ( .A1(n9479), .A2(n7155), .B1(n7832), .B2(P1_U3084), .C1(
        n10112), .C2(n7945), .ZN(P1_U3337) );
  OAI21_X1 U8704 ( .B1(n7083), .B2(n7057), .A(n4383), .ZN(n7092) );
  INV_X1 U8705 ( .A(n7083), .ZN(n7085) );
  NAND3_X1 U8706 ( .A1(n8412), .A2(n7085), .A3(n7084), .ZN(n7086) );
  INV_X1 U8707 ( .A(n9788), .ZN(n7225) );
  AOI21_X1 U8708 ( .B1(n7086), .B2(n8472), .A(n7225), .ZN(n7091) );
  AOI22_X1 U8709 ( .A1(n8480), .A2(n4402), .B1(n8481), .B2(n7087), .ZN(n7089)
         );
  OAI211_X1 U8710 ( .C1(n7230), .C2(n8485), .A(n7089), .B(n7088), .ZN(n7090)
         );
  AOI211_X1 U8711 ( .C1(n8456), .C2(n7092), .A(n7091), .B(n7090), .ZN(n7093)
         );
  INV_X1 U8712 ( .A(n7093), .ZN(P2_U3232) );
  OAI21_X1 U8713 ( .B1(n7096), .B2(n7094), .A(n7095), .ZN(n7104) );
  INV_X1 U8714 ( .A(n7096), .ZN(n7098) );
  NAND3_X1 U8715 ( .A1(n8412), .A2(n7098), .A3(n7097), .ZN(n7099) );
  INV_X1 U8716 ( .A(n4402), .ZN(n7295) );
  AOI21_X1 U8717 ( .B1(n7099), .B2(n8472), .A(n7295), .ZN(n7103) );
  AOI22_X1 U8718 ( .A1(n8480), .A2(n8502), .B1(n8481), .B2(n7337), .ZN(n7101)
         );
  OAI211_X1 U8719 ( .C1(n9877), .C2(n8485), .A(n7101), .B(n7100), .ZN(n7102)
         );
  AOI211_X1 U8720 ( .C1(n8456), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7105)
         );
  INV_X1 U8721 ( .A(n7105), .ZN(P2_U3241) );
  NAND3_X1 U8722 ( .A1(n7108), .A2(n7107), .A3(n7106), .ZN(n7149) );
  NAND2_X2 U8723 ( .A1(n7149), .A2(n9693), .ZN(n9692) );
  OAI211_X1 U8724 ( .C1(n8209), .C2(n7111), .A(n9728), .B(n7110), .ZN(n9702)
         );
  INV_X1 U8725 ( .A(n7112), .ZN(n7113) );
  AOI21_X1 U8726 ( .B1(n6942), .B2(n7114), .A(n7113), .ZN(n9705) );
  NAND2_X1 U8727 ( .A1(n9705), .A2(n7242), .ZN(n7116) );
  INV_X1 U8728 ( .A(n9693), .ZN(n9357) );
  NAND2_X1 U8729 ( .A1(n9357), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7115) );
  OAI211_X1 U8730 ( .C1(n9670), .C2(n9702), .A(n7116), .B(n7115), .ZN(n7121)
         );
  INV_X1 U8731 ( .A(n7117), .ZN(n7120) );
  XOR2_X1 U8732 ( .A(n6942), .B(n7118), .Z(n7119) );
  OAI222_X1 U8733 ( .A1(n9683), .A2(n9686), .B1(n9685), .B2(n7120), .C1(n7119), 
        .C2(n9672), .ZN(n9703) );
  OAI21_X1 U8734 ( .B1(n7121), .B2(n9703), .A(n9692), .ZN(n7124) );
  NAND2_X1 U8735 ( .A1(n9309), .A2(n7122), .ZN(n7123) );
  OAI211_X1 U8736 ( .C1(n6709), .C2(n9692), .A(n7124), .B(n7123), .ZN(P1_U3290) );
  AND2_X1 U8737 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8349) );
  AOI21_X1 U8738 ( .B1(n7130), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7125), .ZN(
        n7128) );
  INV_X1 U8739 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7126) );
  MUX2_X1 U8740 ( .A(n7126), .B(P2_REG1_REG_10__SCAN_IN), .S(n7355), .Z(n7127)
         );
  NOR2_X1 U8741 ( .A1(n7128), .A2(n7127), .ZN(n7354) );
  AOI211_X1 U8742 ( .C1(n7128), .C2(n7127), .A(n7354), .B(n9778), .ZN(n7129)
         );
  AOI211_X1 U8743 ( .C1(n9775), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8349), .B(
        n7129), .ZN(n7136) );
  NAND2_X1 U8744 ( .A1(n7130), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8745 ( .A1(n7132), .A2(n7131), .ZN(n7134) );
  INV_X1 U8746 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7539) );
  MUX2_X1 U8747 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7539), .S(n7355), .Z(n7133)
         );
  NAND2_X1 U8748 ( .A1(n7133), .A2(n7134), .ZN(n7348) );
  OAI211_X1 U8749 ( .C1(n7134), .C2(n7133), .A(n9774), .B(n7348), .ZN(n7135)
         );
  OAI211_X1 U8750 ( .C1(n9777), .C2(n7137), .A(n7136), .B(n7135), .ZN(P2_U3255) );
  INV_X1 U8751 ( .A(n7094), .ZN(n7138) );
  AOI211_X1 U8752 ( .C1(n7140), .C2(n7139), .A(n8478), .B(n7138), .ZN(n7146)
         );
  OAI22_X1 U8753 ( .A1(n7235), .A2(n8472), .B1(n8424), .B2(n7236), .ZN(n7145)
         );
  NAND2_X1 U8754 ( .A1(n8481), .A2(n7238), .ZN(n7142) );
  NAND2_X1 U8755 ( .A1(n8455), .A2(n4821), .ZN(n7141) );
  OAI211_X1 U8756 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7143), .A(n7142), .B(n7141), .ZN(n7144) );
  OR3_X1 U8757 ( .A1(n7146), .A2(n7145), .A3(n7144), .ZN(P2_U3229) );
  INV_X1 U8758 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7147) );
  OAI22_X1 U8759 ( .A1(n9692), .A2(n6685), .B1(n7147), .B2(n9693), .ZN(n7148)
         );
  INV_X1 U8760 ( .A(n7148), .ZN(n7152) );
  OR2_X1 U8761 ( .A1(n7149), .A2(n9670), .ZN(n7676) );
  INV_X1 U8762 ( .A(n9176), .ZN(n9679) );
  OAI21_X1 U8763 ( .B1(n9679), .B2(n9309), .A(n7150), .ZN(n7151) );
  OAI211_X1 U8764 ( .C1(n7153), .C2(n4381), .A(n7152), .B(n7151), .ZN(P1_U3291) );
  INV_X1 U8765 ( .A(n8508), .ZN(n8513) );
  OAI222_X1 U8766 ( .A1(P2_U3152), .A2(n8513), .B1(n7582), .B2(n7155), .C1(
        n7154), .C2(n8311), .ZN(P2_U3342) );
  INV_X1 U8767 ( .A(n7156), .ZN(n7157) );
  INV_X1 U8768 ( .A(n9098), .ZN(n9085) );
  OAI222_X1 U8769 ( .A1(n9479), .A2(n7157), .B1(n9085), .B2(P1_U3084), .C1(
        n10235), .C2(n7945), .ZN(P1_U3336) );
  INV_X1 U8770 ( .A(n8529), .ZN(n8520) );
  OAI222_X1 U8771 ( .A1(n8311), .A2(n7158), .B1(n7582), .B2(n7157), .C1(n8520), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8772 ( .A(n9665), .ZN(n8902) );
  NAND2_X1 U8773 ( .A1(n8902), .A2(n9726), .ZN(n8097) );
  INV_X1 U8774 ( .A(n9726), .ZN(n9019) );
  NAND2_X1 U8775 ( .A1(n9019), .A2(n9665), .ZN(n8100) );
  INV_X1 U8776 ( .A(n9053), .ZN(n7161) );
  NAND2_X1 U8777 ( .A1(n7161), .A2(n7160), .ZN(n8217) );
  NAND2_X1 U8778 ( .A1(n9709), .A2(n9053), .ZN(n8007) );
  NAND2_X1 U8779 ( .A1(n8217), .A2(n8007), .ZN(n7171) );
  NAND2_X1 U8780 ( .A1(n7161), .A2(n9709), .ZN(n7162) );
  NAND2_X1 U8781 ( .A1(n9684), .A2(n7255), .ZN(n8222) );
  NAND2_X1 U8782 ( .A1(n9714), .A2(n9052), .ZN(n8012) );
  NAND2_X1 U8783 ( .A1(n8222), .A2(n8012), .ZN(n7244) );
  NAND2_X1 U8784 ( .A1(n7241), .A2(n7244), .ZN(n7164) );
  NAND2_X1 U8785 ( .A1(n9684), .A2(n9714), .ZN(n7163) );
  NAND2_X1 U8786 ( .A1(n7164), .A2(n7163), .ZN(n9660) );
  NAND2_X1 U8787 ( .A1(n9021), .A2(n9668), .ZN(n7207) );
  NAND2_X1 U8788 ( .A1(n9051), .A2(n9668), .ZN(n7165) );
  INV_X1 U8789 ( .A(n7206), .ZN(n7167) );
  AOI21_X1 U8790 ( .B1(n8101), .B2(n7168), .A(n7167), .ZN(n9732) );
  NAND2_X1 U8791 ( .A1(n8216), .A2(n8010), .ZN(n7170) );
  NAND2_X1 U8792 ( .A1(n9682), .A2(n4566), .ZN(n7172) );
  INV_X1 U8793 ( .A(n8222), .ZN(n7173) );
  INV_X1 U8794 ( .A(n7208), .ZN(n7174) );
  INV_X1 U8795 ( .A(n9671), .ZN(n9659) );
  INV_X1 U8796 ( .A(n8102), .ZN(n8099) );
  XNOR2_X1 U8797 ( .A(n8099), .B(n8101), .ZN(n7175) );
  AOI222_X1 U8798 ( .A1(n9189), .A2(n7175), .B1(n9051), .B2(n9363), .C1(n9050), 
        .C2(n9664), .ZN(n9731) );
  MUX2_X1 U8799 ( .A(n6718), .B(n9731), .S(n9692), .Z(n7178) );
  NAND2_X1 U8800 ( .A1(n9678), .A2(n9709), .ZN(n9677) );
  OR2_X1 U8801 ( .A1(n9677), .A2(n7255), .ZN(n9661) );
  AOI21_X1 U8802 ( .B1(n9726), .B2(n9662), .A(n7215), .ZN(n9729) );
  OAI22_X1 U8803 ( .A1(n9694), .A2(n9019), .B1(n9023), .B2(n9693), .ZN(n7176)
         );
  AOI21_X1 U8804 ( .B1(n9729), .B2(n9679), .A(n7176), .ZN(n7177) );
  OAI211_X1 U8805 ( .C1(n9732), .C2(n9370), .A(n7178), .B(n7177), .ZN(P1_U3285) );
  INV_X1 U8806 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7194) );
  INV_X1 U8807 ( .A(n7499), .ZN(n7184) );
  NOR2_X1 U8808 ( .A1(n7184), .A2(n7179), .ZN(n7180) );
  AOI21_X1 U8809 ( .B1(n7179), .B2(n7184), .A(n7180), .ZN(n7183) );
  OAI21_X1 U8810 ( .B1(n7186), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7181), .ZN(
        n7182) );
  NAND2_X1 U8811 ( .A1(n7183), .A2(n7182), .ZN(n7493) );
  OAI21_X1 U8812 ( .B1(n7183), .B2(n7182), .A(n7493), .ZN(n7192) );
  NAND2_X1 U8813 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7896) );
  OAI21_X1 U8814 ( .B1(n9096), .B2(n7184), .A(n7896), .ZN(n7191) );
  AOI21_X1 U8815 ( .B1(n7186), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7185), .ZN(
        n7189) );
  NAND2_X1 U8816 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7499), .ZN(n7187) );
  OAI21_X1 U8817 ( .B1(n7499), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7187), .ZN(
        n7188) );
  NOR2_X1 U8818 ( .A1(n7189), .A2(n7188), .ZN(n7498) );
  AOI211_X1 U8819 ( .C1(n7189), .C2(n7188), .A(n7498), .B(n9647), .ZN(n7190)
         );
  AOI211_X1 U8820 ( .C1(n9653), .C2(n7192), .A(n7191), .B(n7190), .ZN(n7193)
         );
  OAI21_X1 U8821 ( .B1(n9629), .B2(n7194), .A(n7193), .ZN(P1_U3254) );
  AOI22_X1 U8822 ( .A1(n9309), .A2(n7988), .B1(n9357), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7195) );
  OAI21_X1 U8823 ( .B1(n9176), .B2(n7196), .A(n7195), .ZN(n7199) );
  MUX2_X1 U8824 ( .A(n7197), .B(P1_REG2_REG_2__SCAN_IN), .S(n4381), .Z(n7198)
         );
  INV_X1 U8825 ( .A(n9838), .ZN(n7204) );
  NAND2_X1 U8826 ( .A1(n8560), .A2(n8781), .ZN(n9805) );
  NAND2_X1 U8827 ( .A1(n9805), .A2(n9837), .ZN(n7203) );
  AOI22_X1 U8828 ( .A1(n9838), .A2(n9790), .B1(n9785), .B2(n8506), .ZN(n9840)
         );
  INV_X1 U8829 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7200) );
  OAI22_X1 U8830 ( .A1(n9808), .A2(n9840), .B1(n7200), .B2(n9793), .ZN(n7201)
         );
  AOI21_X1 U8831 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9808), .A(n7201), .ZN(
        n7202) );
  OAI211_X1 U8832 ( .C1(n7204), .C2(n8748), .A(n7203), .B(n7202), .ZN(P2_U3296) );
  NAND2_X1 U8833 ( .A1(n8902), .A2(n9019), .ZN(n7205) );
  INV_X1 U8834 ( .A(n9050), .ZN(n8095) );
  NAND2_X1 U8835 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  NAND2_X1 U8836 ( .A1(n9736), .A2(n9050), .ZN(n8219) );
  XNOR2_X1 U8837 ( .A(n7266), .B(n8016), .ZN(n9739) );
  INV_X1 U8838 ( .A(n9739), .ZN(n7221) );
  AND2_X1 U8839 ( .A1(n8097), .A2(n7207), .ZN(n8223) );
  INV_X1 U8840 ( .A(n8013), .ZN(n7209) );
  NAND2_X1 U8841 ( .A1(n7209), .A2(n8097), .ZN(n8225) );
  AND2_X1 U8842 ( .A1(n8225), .A2(n8100), .ZN(n8009) );
  INV_X1 U8843 ( .A(n7260), .ZN(n7212) );
  AOI21_X1 U8844 ( .B1(n8016), .B2(n7213), .A(n7212), .ZN(n7214) );
  OAI222_X1 U8845 ( .A1(n9683), .A2(n7606), .B1(n9685), .B2(n8902), .C1(n9672), 
        .C2(n7214), .ZN(n9737) );
  NAND2_X1 U8846 ( .A1(n7215), .A2(n9736), .ZN(n7262) );
  OAI211_X1 U8847 ( .C1(n7215), .C2(n9736), .A(n7262), .B(n9728), .ZN(n9735)
         );
  OAI22_X1 U8848 ( .A1(n9692), .A2(n7216), .B1(n8904), .B2(n9693), .ZN(n7217)
         );
  AOI21_X1 U8849 ( .B1(n9309), .B2(n8094), .A(n7217), .ZN(n7218) );
  OAI21_X1 U8850 ( .B1(n9735), .B2(n7676), .A(n7218), .ZN(n7219) );
  AOI21_X1 U8851 ( .B1(n9737), .B2(n9692), .A(n7219), .ZN(n7220) );
  OAI21_X1 U8852 ( .B1(n7221), .B2(n9370), .A(n7220), .ZN(P1_U3284) );
  NAND2_X1 U8853 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  NAND2_X1 U8854 ( .A1(n7227), .A2(n7226), .ZN(n9802) );
  NAND2_X1 U8855 ( .A1(n9802), .A2(n9803), .ZN(n7229) );
  NAND2_X1 U8856 ( .A1(n7235), .A2(n7230), .ZN(n7228) );
  NAND2_X1 U8857 ( .A1(n7229), .A2(n7228), .ZN(n7293) );
  XNOR2_X1 U8858 ( .A(n7293), .B(n7233), .ZN(n9870) );
  INV_X1 U8859 ( .A(n7230), .ZN(n9799) );
  INV_X1 U8860 ( .A(n9797), .ZN(n7231) );
  AOI211_X1 U8861 ( .C1(n4821), .C2(n7231), .A(n9900), .B(n7334), .ZN(n9868)
         );
  XNOR2_X1 U8862 ( .A(n7232), .B(n7233), .ZN(n7234) );
  OAI222_X1 U8863 ( .A1(n9535), .A2(n7236), .B1(n9533), .B2(n7235), .C1(n9531), 
        .C2(n7234), .ZN(n9867) );
  AOI21_X1 U8864 ( .B1(n9868), .B2(n4410), .A(n9867), .ZN(n7237) );
  MUX2_X1 U8865 ( .A(n6785), .B(n7237), .S(n9791), .Z(n7240) );
  AOI22_X1 U8866 ( .A1(n8598), .A2(n4821), .B1(n8778), .B2(n7238), .ZN(n7239)
         );
  OAI211_X1 U8867 ( .C1(n9870), .C2(n8748), .A(n7240), .B(n7239), .ZN(P2_U3291) );
  XNOR2_X1 U8868 ( .A(n7241), .B(n7244), .ZN(n7243) );
  NAND2_X1 U8869 ( .A1(n7243), .A2(n7242), .ZN(n7252) );
  INV_X1 U8870 ( .A(n7244), .ZN(n7245) );
  XNOR2_X1 U8871 ( .A(n7246), .B(n7245), .ZN(n7250) );
  NAND2_X1 U8872 ( .A1(n9051), .A2(n9664), .ZN(n7248) );
  NAND2_X1 U8873 ( .A1(n9053), .A2(n9363), .ZN(n7247) );
  NAND2_X1 U8874 ( .A1(n7248), .A2(n7247), .ZN(n7249) );
  AOI21_X1 U8875 ( .B1(n7250), .B2(n9189), .A(n7249), .ZN(n7251) );
  AND2_X1 U8876 ( .A1(n7252), .A2(n7251), .ZN(n9718) );
  NAND2_X1 U8877 ( .A1(n9677), .A2(n7255), .ZN(n7253) );
  NAND2_X1 U8878 ( .A1(n9661), .A2(n7253), .ZN(n9715) );
  AOI22_X1 U8879 ( .A1(n4381), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7254), .B2(
        n9357), .ZN(n7257) );
  NAND2_X1 U8880 ( .A1(n9309), .A2(n7255), .ZN(n7256) );
  OAI211_X1 U8881 ( .C1(n9715), .C2(n9176), .A(n7257), .B(n7256), .ZN(n7258)
         );
  INV_X1 U8882 ( .A(n7258), .ZN(n7259) );
  OAI21_X1 U8883 ( .B1(n9718), .B2(n4381), .A(n7259), .ZN(P1_U3287) );
  INV_X1 U8884 ( .A(n9048), .ZN(n7635) );
  NAND2_X1 U8885 ( .A1(n7606), .A2(n7445), .ZN(n8107) );
  NAND2_X1 U8886 ( .A1(n9743), .A2(n9049), .ZN(n7381) );
  XNOR2_X1 U8887 ( .A(n7368), .B(n8018), .ZN(n7261) );
  OAI222_X1 U8888 ( .A1(n9683), .A2(n7635), .B1(n9685), .B2(n8095), .C1(n7261), 
        .C2(n9672), .ZN(n9745) );
  OR2_X1 U8889 ( .A1(n7262), .A2(n7445), .ZN(n7387) );
  NAND2_X1 U8890 ( .A1(n7262), .A2(n7445), .ZN(n7263) );
  NAND2_X1 U8891 ( .A1(n7387), .A2(n7263), .ZN(n9744) );
  OAI22_X1 U8892 ( .A1(n9692), .A2(n10152), .B1(n7443), .B2(n9693), .ZN(n7264)
         );
  AOI21_X1 U8893 ( .B1(n9309), .B2(n7445), .A(n7264), .ZN(n7265) );
  OAI21_X1 U8894 ( .B1(n9744), .B2(n9176), .A(n7265), .ZN(n7273) );
  NAND2_X1 U8895 ( .A1(n8095), .A2(n9736), .ZN(n7267) );
  NAND2_X1 U8896 ( .A1(n7268), .A2(n7267), .ZN(n7270) );
  INV_X1 U8897 ( .A(n9747), .ZN(n7271) );
  AND2_X1 U8898 ( .A1(n7270), .A2(n8018), .ZN(n9741) );
  NOR3_X1 U8899 ( .A1(n7271), .A2(n9741), .A3(n9370), .ZN(n7272) );
  AOI211_X1 U8900 ( .C1(n9692), .C2(n9745), .A(n7273), .B(n7272), .ZN(n7274)
         );
  INV_X1 U8901 ( .A(n7274), .ZN(P1_U3283) );
  INV_X1 U8902 ( .A(n7276), .ZN(n7277) );
  AOI21_X1 U8903 ( .B1(n7275), .B2(n7277), .A(n8478), .ZN(n7281) );
  NOR3_X1 U8904 ( .A1(n8464), .A2(n7278), .A3(n7400), .ZN(n7280) );
  OAI21_X1 U8905 ( .B1(n7281), .B2(n7280), .A(n7279), .ZN(n7287) );
  INV_X1 U8906 ( .A(n8315), .ZN(n8365) );
  OR2_X1 U8907 ( .A1(n7533), .A2(n9535), .ZN(n7283) );
  OR2_X1 U8908 ( .A1(n7400), .A2(n9533), .ZN(n7282) );
  AND2_X1 U8909 ( .A1(n7283), .A2(n7282), .ZN(n7953) );
  OAI22_X1 U8910 ( .A1(n8365), .A2(n7953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7284), .ZN(n7285) );
  AOI21_X1 U8911 ( .B1(n9881), .B2(n8455), .A(n7285), .ZN(n7286) );
  OAI211_X1 U8912 ( .C1(n8470), .C2(n7958), .A(n7287), .B(n7286), .ZN(P2_U3223) );
  NAND3_X1 U8913 ( .A1(n7290), .A2(n7289), .A3(n7288), .ZN(n7310) );
  INV_X1 U8914 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U8915 ( .A1(n7293), .A2(n7292), .ZN(n7297) );
  NAND2_X1 U8916 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  NAND2_X1 U8917 ( .A1(n7297), .A2(n7296), .ZN(n7332) );
  NAND2_X1 U8918 ( .A1(n8503), .A2(n7298), .ZN(n7299) );
  XOR2_X1 U8919 ( .A(n7398), .B(n7399), .Z(n7971) );
  AND2_X1 U8920 ( .A1(n7526), .A2(n4625), .ZN(n7300) );
  NAND2_X1 U8921 ( .A1(n7643), .A2(n7300), .ZN(n9890) );
  XNOR2_X1 U8922 ( .A(n7301), .B(n7399), .ZN(n7304) );
  OR2_X1 U8923 ( .A1(n7318), .A2(n9535), .ZN(n7303) );
  NAND2_X1 U8924 ( .A1(n8503), .A2(n9787), .ZN(n7302) );
  NAND2_X1 U8925 ( .A1(n7303), .A2(n7302), .ZN(n8314) );
  AOI21_X1 U8926 ( .B1(n7304), .B2(n9790), .A(n8314), .ZN(n7965) );
  AOI21_X1 U8927 ( .B1(n7336), .B2(n8317), .A(n9900), .ZN(n7305) );
  AND2_X1 U8928 ( .A1(n7305), .A2(n7955), .ZN(n7969) );
  AOI21_X1 U8929 ( .B1(n9882), .B2(n8317), .A(n7969), .ZN(n7306) );
  OAI211_X1 U8930 ( .C1(n7971), .C2(n9871), .A(n7965), .B(n7306), .ZN(n7311)
         );
  NAND2_X1 U8931 ( .A1(n7311), .A2(n9924), .ZN(n7307) );
  OAI21_X1 U8932 ( .B1(n9924), .B2(n7308), .A(n7307), .ZN(P2_U3527) );
  INV_X1 U8933 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U8934 ( .A1(n7311), .A2(n9908), .ZN(n7312) );
  OAI21_X1 U8935 ( .B1(n9908), .B2(n7313), .A(n7312), .ZN(P2_U3472) );
  INV_X1 U8936 ( .A(n7279), .ZN(n7316) );
  NOR3_X1 U8937 ( .A1(n8464), .A2(n7314), .A3(n7318), .ZN(n7315) );
  AOI21_X1 U8938 ( .B1(n7316), .B2(n8456), .A(n7315), .ZN(n7327) );
  INV_X1 U8939 ( .A(n7317), .ZN(n7324) );
  INV_X1 U8940 ( .A(n8444), .ZN(n8499) );
  AOI22_X1 U8941 ( .A1(n8480), .A2(n8499), .B1(n8481), .B2(n7411), .ZN(n7322)
         );
  INV_X1 U8942 ( .A(n7318), .ZN(n8501) );
  NAND2_X1 U8943 ( .A1(n8482), .A2(n8501), .ZN(n7320) );
  NAND2_X1 U8944 ( .A1(n8455), .A2(n7528), .ZN(n7319) );
  NAND4_X1 U8945 ( .A1(n7322), .A2(n7321), .A3(n7320), .A4(n7319), .ZN(n7323)
         );
  AOI21_X1 U8946 ( .B1(n7324), .B2(n8456), .A(n7323), .ZN(n7325) );
  OAI21_X1 U8947 ( .B1(n7327), .B2(n7326), .A(n7325), .ZN(P2_U3233) );
  INV_X1 U8948 ( .A(n7328), .ZN(n7331) );
  AOI22_X1 U8949 ( .A1(n9111), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9474), .ZN(n7329) );
  OAI21_X1 U8950 ( .B1(n7331), .B2(n9479), .A(n7329), .ZN(P1_U3335) );
  AOI22_X1 U8951 ( .A1(n8540), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8892), .ZN(n7330) );
  OAI21_X1 U8952 ( .B1(n7331), .B2(n8894), .A(n7330), .ZN(P2_U3340) );
  INV_X1 U8953 ( .A(n8748), .ZN(n9804) );
  INV_X1 U8954 ( .A(n7341), .ZN(n7333) );
  XNOR2_X1 U8955 ( .A(n7332), .B(n7333), .ZN(n9874) );
  OR2_X1 U8956 ( .A1(n7334), .A2(n9877), .ZN(n7335) );
  AND2_X1 U8957 ( .A1(n7336), .A2(n7335), .ZN(n9875) );
  AOI22_X1 U8958 ( .A1(n9521), .A2(n9875), .B1(n7337), .B2(n8778), .ZN(n7338)
         );
  OAI21_X1 U8959 ( .B1(n9877), .B2(n8781), .A(n7338), .ZN(n7346) );
  OAI21_X1 U8960 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(n7342) );
  NAND2_X1 U8961 ( .A1(n7342), .A2(n9790), .ZN(n7344) );
  AOI22_X1 U8962 ( .A1(n8502), .A2(n9785), .B1(n9787), .B2(n4402), .ZN(n7343)
         );
  NAND2_X1 U8963 ( .A1(n7344), .A2(n7343), .ZN(n9879) );
  MUX2_X1 U8964 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9879), .S(n9791), .Z(n7345)
         );
  AOI211_X1 U8965 ( .C1(n9804), .C2(n9874), .A(n7346), .B(n7345), .ZN(n7347)
         );
  INV_X1 U8966 ( .A(n7347), .ZN(P2_U3290) );
  NAND2_X1 U8967 ( .A1(n7355), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U8968 ( .A1(n7349), .A2(n7348), .ZN(n7352) );
  INV_X1 U8969 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7350) );
  MUX2_X1 U8970 ( .A(n7350), .B(P2_REG2_REG_11__SCAN_IN), .S(n7418), .Z(n7351)
         );
  NOR2_X1 U8971 ( .A1(n7352), .A2(n7351), .ZN(n7424) );
  AOI21_X1 U8972 ( .B1(n7352), .B2(n7351), .A(n7424), .ZN(n7363) );
  INV_X1 U8973 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7353) );
  NOR2_X1 U8974 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7353), .ZN(n7360) );
  INV_X1 U8975 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7356) );
  MUX2_X1 U8976 ( .A(n7356), .B(P2_REG1_REG_11__SCAN_IN), .S(n7418), .Z(n7357)
         );
  AOI211_X1 U8977 ( .C1(n7358), .C2(n7357), .A(n7417), .B(n9778), .ZN(n7359)
         );
  AOI211_X1 U8978 ( .C1(n9775), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7360), .B(
        n7359), .ZN(n7362) );
  NAND2_X1 U8979 ( .A1(n8534), .A2(n7418), .ZN(n7361) );
  OAI211_X1 U8980 ( .C1(n7363), .C2(n9776), .A(n7362), .B(n7361), .ZN(P2_U3256) );
  NAND2_X1 U8981 ( .A1(n9049), .A2(n7445), .ZN(n7364) );
  INV_X1 U8982 ( .A(n7393), .ZN(n7602) );
  NAND2_X1 U8983 ( .A1(n7602), .A2(n7635), .ZN(n7366) );
  AND2_X1 U8984 ( .A1(n7393), .A2(n9048), .ZN(n7365) );
  OR2_X1 U8985 ( .A1(n7734), .A2(n7638), .ZN(n8111) );
  NAND2_X1 U8986 ( .A1(n7638), .A2(n7734), .ZN(n7451) );
  NAND2_X1 U8987 ( .A1(n8111), .A2(n7451), .ZN(n8020) );
  NAND2_X1 U8988 ( .A1(n7367), .A2(n8020), .ZN(n7449) );
  OAI21_X1 U8989 ( .B1(n7367), .B2(n8020), .A(n7449), .ZN(n9496) );
  INV_X1 U8990 ( .A(n9496), .ZN(n7380) );
  NAND2_X1 U8991 ( .A1(n7602), .A2(n9048), .ZN(n7383) );
  AND2_X1 U8992 ( .A1(n7383), .A2(n7381), .ZN(n8108) );
  NAND2_X1 U8993 ( .A1(n7635), .A2(n7393), .ZN(n7450) );
  NAND2_X1 U8994 ( .A1(n7452), .A2(n7450), .ZN(n7370) );
  INV_X1 U8995 ( .A(n8020), .ZN(n7369) );
  XNOR2_X1 U8996 ( .A(n7370), .B(n7369), .ZN(n7371) );
  NAND2_X1 U8997 ( .A1(n7371), .A2(n9189), .ZN(n7373) );
  AOI22_X1 U8998 ( .A1(n9363), .A2(n9048), .B1(n9046), .B2(n9664), .ZN(n7372)
         );
  NAND2_X1 U8999 ( .A1(n7373), .A2(n7372), .ZN(n9495) );
  NOR2_X2 U9000 ( .A1(n7387), .A2(n7393), .ZN(n7388) );
  AND2_X1 U9001 ( .A1(n7388), .A2(n9493), .ZN(n7458) );
  INV_X1 U9002 ( .A(n7458), .ZN(n7374) );
  OAI211_X1 U9003 ( .C1(n9493), .C2(n7388), .A(n7374), .B(n9728), .ZN(n9492)
         );
  INV_X1 U9004 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7375) );
  OAI22_X1 U9005 ( .A1(n9692), .A2(n7375), .B1(n7631), .B2(n9693), .ZN(n7376)
         );
  AOI21_X1 U9006 ( .B1(n9309), .B2(n7638), .A(n7376), .ZN(n7377) );
  OAI21_X1 U9007 ( .B1(n9492), .B2(n7676), .A(n7377), .ZN(n7378) );
  AOI21_X1 U9008 ( .B1(n9495), .B2(n9692), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9009 ( .B1(n7380), .B2(n9370), .A(n7379), .ZN(P1_U3281) );
  NAND2_X1 U9010 ( .A1(n7382), .A2(n7381), .ZN(n7384) );
  NAND2_X1 U9011 ( .A1(n7383), .A2(n7450), .ZN(n8019) );
  XNOR2_X1 U9012 ( .A(n7384), .B(n8019), .ZN(n7385) );
  AOI222_X1 U9013 ( .A1(n9189), .A2(n7385), .B1(n9047), .B2(n9664), .C1(n9049), 
        .C2(n9363), .ZN(n9751) );
  INV_X1 U9014 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7386) );
  OAI22_X1 U9015 ( .A1(n9692), .A2(n7386), .B1(n7603), .B2(n9693), .ZN(n7392)
         );
  INV_X1 U9016 ( .A(n7387), .ZN(n7390) );
  INV_X1 U9017 ( .A(n7388), .ZN(n7389) );
  OAI21_X1 U9018 ( .B1(n7602), .B2(n7390), .A(n7389), .ZN(n9752) );
  NOR2_X1 U9019 ( .A1(n9752), .A2(n9176), .ZN(n7391) );
  AOI211_X1 U9020 ( .C1(n9309), .C2(n7393), .A(n7392), .B(n7391), .ZN(n7397)
         );
  XOR2_X1 U9021 ( .A(n8019), .B(n7394), .Z(n9756) );
  INV_X1 U9022 ( .A(n9370), .ZN(n7395) );
  NAND2_X1 U9023 ( .A1(n9756), .A2(n7395), .ZN(n7396) );
  OAI211_X1 U9024 ( .C1(n9751), .C2(n4381), .A(n7397), .B(n7396), .ZN(P1_U3282) );
  NAND2_X1 U9025 ( .A1(n9881), .A2(n8501), .ZN(n7402) );
  NAND2_X1 U9026 ( .A1(n7403), .A2(n7405), .ZN(n7530) );
  OAI21_X1 U9027 ( .B1(n7403), .B2(n7405), .A(n7530), .ZN(n7482) );
  XNOR2_X1 U9028 ( .A(n7404), .B(n7405), .ZN(n7407) );
  AOI22_X1 U9029 ( .A1(n9787), .A2(n8501), .B1(n8499), .B2(n9785), .ZN(n7406)
         );
  OAI21_X1 U9030 ( .B1(n7407), .B2(n9531), .A(n7406), .ZN(n7408) );
  AOI21_X1 U9031 ( .B1(n7409), .B2(n7482), .A(n7408), .ZN(n7485) );
  INV_X1 U9032 ( .A(n7528), .ZN(n7414) );
  INV_X1 U9033 ( .A(n7957), .ZN(n7410) );
  AOI21_X1 U9034 ( .B1(n7528), .B2(n7410), .A(n7540), .ZN(n7483) );
  NAND2_X1 U9035 ( .A1(n7483), .A2(n9521), .ZN(n7413) );
  AOI22_X1 U9036 ( .A1(n9808), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7411), .B2(
        n8778), .ZN(n7412) );
  OAI211_X1 U9037 ( .C1(n7414), .C2(n8781), .A(n7413), .B(n7412), .ZN(n7415)
         );
  AOI21_X1 U9038 ( .B1(n7482), .B2(n8767), .A(n7415), .ZN(n7416) );
  OAI21_X1 U9039 ( .B1(n7485), .B2(n9808), .A(n7416), .ZN(P2_U3287) );
  INV_X1 U9040 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7512) );
  MUX2_X1 U9041 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7512), .S(n7427), .Z(n7419)
         );
  OAI21_X1 U9042 ( .B1(n7420), .B2(n7419), .A(n7515), .ZN(n7423) );
  AND2_X1 U9043 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8386) );
  INV_X1 U9044 ( .A(n9775), .ZN(n7592) );
  INV_X1 U9045 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7421) );
  NOR2_X1 U9046 ( .A1(n7592), .A2(n7421), .ZN(n7422) );
  AOI211_X1 U9047 ( .C1(n9773), .C2(n7423), .A(n8386), .B(n7422), .ZN(n7431)
         );
  AOI21_X1 U9048 ( .B1(n7425), .B2(n7350), .A(n7424), .ZN(n7429) );
  INV_X1 U9049 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7426) );
  MUX2_X1 U9050 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7426), .S(n7427), .Z(n7428)
         );
  NAND2_X1 U9051 ( .A1(n7427), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7508) );
  OAI211_X1 U9052 ( .C1(n7427), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7429), .B(
        n7508), .ZN(n7507) );
  OAI211_X1 U9053 ( .C1(n7429), .C2(n7428), .A(n9774), .B(n7507), .ZN(n7430)
         );
  OAI211_X1 U9054 ( .C1(n9777), .C2(n7513), .A(n7431), .B(n7430), .ZN(P2_U3257) );
  INV_X1 U9055 ( .A(n7432), .ZN(n7434) );
  OAI222_X1 U9056 ( .A1(n8311), .A2(n7433), .B1(n7582), .B2(n7434), .C1(
        P2_U3152), .C2(n4410), .ZN(P2_U3339) );
  OAI222_X1 U9057 ( .A1(n7945), .A2(n7435), .B1(n9479), .B2(n7434), .C1(n9305), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  XNOR2_X1 U9058 ( .A(n7437), .B(n7436), .ZN(n7438) );
  XNOR2_X1 U9059 ( .A(n7439), .B(n7438), .ZN(n7447) );
  NOR2_X1 U9060 ( .A1(n9503), .A2(n8095), .ZN(n7440) );
  AOI211_X1 U9061 ( .C1(n9500), .C2(n9048), .A(n7441), .B(n7440), .ZN(n7442)
         );
  OAI21_X1 U9062 ( .B1(n9517), .B2(n7443), .A(n7442), .ZN(n7444) );
  AOI21_X1 U9063 ( .B1(n9038), .B2(n7445), .A(n7444), .ZN(n7446) );
  OAI21_X1 U9064 ( .B1(n7447), .B2(n9509), .A(n7446), .ZN(P1_U3219) );
  OR2_X1 U9065 ( .A1(n7638), .A2(n9047), .ZN(n7448) );
  NAND2_X1 U9066 ( .A1(n7449), .A2(n7448), .ZN(n7467) );
  XNOR2_X1 U9067 ( .A(n7476), .B(n9046), .ZN(n8122) );
  XOR2_X1 U9068 ( .A(n7467), .B(n8122), .Z(n9580) );
  INV_X1 U9069 ( .A(n9580), .ZN(n7465) );
  AND2_X1 U9070 ( .A1(n7451), .A2(n7450), .ZN(n8109) );
  NAND2_X1 U9071 ( .A1(n7453), .A2(n8111), .ZN(n7475) );
  INV_X1 U9072 ( .A(n8122), .ZN(n7454) );
  XNOR2_X1 U9073 ( .A(n7475), .B(n7454), .ZN(n7455) );
  NAND2_X1 U9074 ( .A1(n7455), .A2(n9189), .ZN(n7457) );
  AOI22_X1 U9075 ( .A1(n9363), .A2(n9047), .B1(n9045), .B2(n9664), .ZN(n7456)
         );
  NAND2_X1 U9076 ( .A1(n7457), .A2(n7456), .ZN(n9579) );
  NAND2_X1 U9077 ( .A1(n7458), .A2(n9576), .ZN(n7471) );
  OR2_X1 U9078 ( .A1(n7458), .A2(n9576), .ZN(n7459) );
  NAND2_X1 U9079 ( .A1(n7471), .A2(n7459), .ZN(n9577) );
  OAI22_X1 U9080 ( .A1(n9692), .A2(n7460), .B1(n7731), .B2(n9693), .ZN(n7461)
         );
  AOI21_X1 U9081 ( .B1(n9309), .B2(n7476), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9082 ( .B1(n9577), .B2(n9176), .A(n7462), .ZN(n7463) );
  AOI21_X1 U9083 ( .B1(n9579), .B2(n9692), .A(n7463), .ZN(n7464) );
  OAI21_X1 U9084 ( .B1(n7465), .B2(n9370), .A(n7464), .ZN(P1_U3280) );
  NAND2_X1 U9085 ( .A1(n7476), .A2(n9046), .ZN(n7466) );
  INV_X1 U9086 ( .A(n9045), .ZN(n7897) );
  OR2_X1 U9087 ( .A1(n7563), .A2(n7897), .ZN(n8125) );
  NAND2_X1 U9088 ( .A1(n7563), .A2(n7897), .ZN(n8121) );
  NAND2_X1 U9089 ( .A1(n7469), .A2(n7468), .ZN(n7565) );
  OAI21_X1 U9090 ( .B1(n7469), .B2(n7468), .A(n7565), .ZN(n9571) );
  OR2_X2 U9091 ( .A1(n7471), .A2(n7563), .ZN(n7572) );
  INV_X1 U9092 ( .A(n7572), .ZN(n7470) );
  AOI211_X1 U9093 ( .C1(n7563), .C2(n7471), .A(n9753), .B(n7470), .ZN(n9573)
         );
  INV_X1 U9094 ( .A(n7563), .ZN(n9506) );
  NOR2_X1 U9095 ( .A1(n9506), .A2(n9694), .ZN(n7474) );
  INV_X1 U9096 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7472) );
  OAI22_X1 U9097 ( .A1(n9692), .A2(n7472), .B1(n9516), .B2(n9693), .ZN(n7473)
         );
  AOI211_X1 U9098 ( .C1(n9573), .C2(n9340), .A(n7474), .B(n7473), .ZN(n7481)
         );
  INV_X1 U9099 ( .A(n9046), .ZN(n9504) );
  NAND2_X1 U9100 ( .A1(n7476), .A2(n9504), .ZN(n8044) );
  OR2_X1 U9101 ( .A1(n7476), .A2(n9504), .ZN(n8057) );
  XNOR2_X1 U9102 ( .A(n7566), .B(n7468), .ZN(n7477) );
  NAND2_X1 U9103 ( .A1(n7477), .A2(n9189), .ZN(n7479) );
  AOI22_X1 U9104 ( .A1(n9363), .A2(n9046), .B1(n9499), .B2(n9664), .ZN(n7478)
         );
  NAND2_X1 U9105 ( .A1(n7479), .A2(n7478), .ZN(n9572) );
  NAND2_X1 U9106 ( .A1(n9572), .A2(n9692), .ZN(n7480) );
  OAI211_X1 U9107 ( .C1(n9571), .C2(n9370), .A(n7481), .B(n7480), .ZN(P1_U3279) );
  INV_X1 U9108 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7488) );
  INV_X1 U9109 ( .A(n7482), .ZN(n7486) );
  AOI22_X1 U9110 ( .A1(n7483), .A2(n9883), .B1(n9882), .B2(n7528), .ZN(n7484)
         );
  OAI211_X1 U9111 ( .C1(n7486), .C2(n9890), .A(n7485), .B(n7484), .ZN(n7489)
         );
  NAND2_X1 U9112 ( .A1(n7489), .A2(n9908), .ZN(n7487) );
  OAI21_X1 U9113 ( .B1(n9908), .B2(n7488), .A(n7487), .ZN(P2_U3478) );
  NAND2_X1 U9114 ( .A1(n7489), .A2(n9924), .ZN(n7490) );
  OAI21_X1 U9115 ( .B1(n9924), .B2(n6956), .A(n7490), .ZN(P2_U3529) );
  NOR2_X1 U9116 ( .A1(n7694), .A2(n7491), .ZN(n7492) );
  AOI21_X1 U9117 ( .B1(n7491), .B2(n7694), .A(n7492), .ZN(n7495) );
  OAI21_X1 U9118 ( .B1(n7499), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7493), .ZN(
        n7494) );
  NAND2_X1 U9119 ( .A1(n7495), .A2(n7494), .ZN(n7687) );
  OAI21_X1 U9120 ( .B1(n7495), .B2(n7494), .A(n7687), .ZN(n7503) );
  NOR2_X1 U9121 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7496), .ZN(n7978) );
  INV_X1 U9122 ( .A(n7978), .ZN(n7497) );
  OAI21_X1 U9123 ( .B1(n9096), .B2(n7694), .A(n7497), .ZN(n7502) );
  AOI211_X1 U9124 ( .C1(n7500), .C2(n7673), .A(n7696), .B(n9647), .ZN(n7501)
         );
  AOI211_X1 U9125 ( .C1(n9653), .C2(n7503), .A(n7502), .B(n7501), .ZN(n7504)
         );
  OAI21_X1 U9126 ( .B1(n9629), .B2(n10173), .A(n7504), .ZN(P1_U3255) );
  INV_X1 U9127 ( .A(n7505), .ZN(n7527) );
  OAI222_X1 U9128 ( .A1(n9479), .A2(n7527), .B1(P1_U3084), .B2(n5728), .C1(
        n7506), .C2(n7945), .ZN(P1_U3333) );
  NAND2_X1 U9129 ( .A1(n7508), .A2(n7507), .ZN(n7511) );
  INV_X1 U9130 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7509) );
  AOI22_X1 U9131 ( .A1(n7589), .A2(n7509), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7516), .ZN(n7510) );
  NOR2_X1 U9132 ( .A1(n7511), .A2(n7510), .ZN(n7584) );
  AOI21_X1 U9133 ( .B1(n7511), .B2(n7510), .A(n7584), .ZN(n7525) );
  NAND2_X1 U9134 ( .A1(n7513), .A2(n7512), .ZN(n7514) );
  NAND2_X1 U9135 ( .A1(n7515), .A2(n7514), .ZN(n7519) );
  INV_X1 U9136 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7517) );
  AOI22_X1 U9137 ( .A1(n7589), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7517), .B2(
        n7516), .ZN(n7518) );
  NAND2_X1 U9138 ( .A1(n7518), .A2(n7519), .ZN(n7588) );
  OAI21_X1 U9139 ( .B1(n7519), .B2(n7518), .A(n7588), .ZN(n7522) );
  AND2_X1 U9140 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8436) );
  INV_X1 U9141 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7520) );
  NOR2_X1 U9142 ( .A1(n7592), .A2(n7520), .ZN(n7521) );
  AOI211_X1 U9143 ( .C1(n9773), .C2(n7522), .A(n8436), .B(n7521), .ZN(n7524)
         );
  NAND2_X1 U9144 ( .A1(n8534), .A2(n7589), .ZN(n7523) );
  OAI211_X1 U9145 ( .C1(n7525), .C2(n9776), .A(n7524), .B(n7523), .ZN(P2_U3258) );
  OAI222_X1 U9146 ( .A1(n8311), .A2(n9970), .B1(n7582), .B2(n7527), .C1(n7526), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U9147 ( .A(n7533), .ZN(n8500) );
  OR2_X1 U9148 ( .A1(n7528), .A2(n8500), .ZN(n7529) );
  NAND2_X1 U9149 ( .A1(n7547), .A2(n7545), .ZN(n7614) );
  OAI21_X1 U9150 ( .B1(n7547), .B2(n7545), .A(n7614), .ZN(n9891) );
  OR2_X1 U9151 ( .A1(n9891), .A2(n8774), .ZN(n7537) );
  OAI21_X1 U9152 ( .B1(n7532), .B2(n7531), .A(n7618), .ZN(n7535) );
  OAI22_X1 U9153 ( .A1(n7533), .A2(n9533), .B1(n8381), .B2(n9535), .ZN(n7534)
         );
  AOI21_X1 U9154 ( .B1(n7535), .B2(n9790), .A(n7534), .ZN(n7536) );
  NAND2_X1 U9155 ( .A1(n7537), .A2(n7536), .ZN(n9894) );
  NAND2_X1 U9156 ( .A1(n9894), .A2(n9791), .ZN(n7544) );
  OAI22_X1 U9157 ( .A1(n9791), .A2(n7539), .B1(n7538), .B2(n9793), .ZN(n7542)
         );
  INV_X1 U9158 ( .A(n8351), .ZN(n9892) );
  NAND2_X1 U9159 ( .A1(n7540), .A2(n9892), .ZN(n7621) );
  OAI21_X1 U9160 ( .B1(n7540), .B2(n9892), .A(n7621), .ZN(n9893) );
  NOR2_X1 U9161 ( .A1(n9893), .A2(n8560), .ZN(n7541) );
  AOI211_X1 U9162 ( .C1(n8598), .C2(n8351), .A(n7542), .B(n7541), .ZN(n7543)
         );
  OAI211_X1 U9163 ( .C1(n9891), .C2(n8783), .A(n7544), .B(n7543), .ZN(P2_U3286) );
  NAND2_X1 U9164 ( .A1(n8449), .A2(n4900), .ZN(n7549) );
  AND2_X1 U9165 ( .A1(n7545), .A2(n7548), .ZN(n7546) );
  NAND2_X1 U9166 ( .A1(n7547), .A2(n7546), .ZN(n7553) );
  INV_X1 U9167 ( .A(n7548), .ZN(n7551) );
  NAND2_X1 U9168 ( .A1(n8351), .A2(n8499), .ZN(n7613) );
  AND2_X1 U9169 ( .A1(n7613), .A2(n7549), .ZN(n7550) );
  OR2_X1 U9170 ( .A1(n7551), .A2(n7550), .ZN(n7552) );
  NAND2_X1 U9171 ( .A1(n7553), .A2(n7552), .ZN(n7703) );
  XNOR2_X1 U9172 ( .A(n7703), .B(n7702), .ZN(n9905) );
  INV_X1 U9173 ( .A(n9905), .ZN(n7562) );
  NAND2_X1 U9174 ( .A1(n7555), .A2(n7554), .ZN(n7556) );
  XNOR2_X1 U9175 ( .A(n7556), .B(n7702), .ZN(n7557) );
  OAI222_X1 U9176 ( .A1(n9533), .A2(n8381), .B1(n9535), .B2(n7709), .C1(n9531), 
        .C2(n7557), .ZN(n9902) );
  OAI21_X1 U9177 ( .B1(n4807), .B2(n4806), .A(n7791), .ZN(n9901) );
  AOI22_X1 U9178 ( .A1(n9808), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8387), .B2(
        n8778), .ZN(n7559) );
  NAND2_X1 U9179 ( .A1(n8598), .A2(n8388), .ZN(n7558) );
  OAI211_X1 U9180 ( .C1(n9901), .C2(n8560), .A(n7559), .B(n7558), .ZN(n7560)
         );
  AOI21_X1 U9181 ( .B1(n9902), .B2(n9791), .A(n7560), .ZN(n7561) );
  OAI21_X1 U9182 ( .B1(n8748), .B2(n7562), .A(n7561), .ZN(P2_U3284) );
  NAND2_X1 U9183 ( .A1(n7563), .A2(n9045), .ZN(n7564) );
  NAND2_X1 U9184 ( .A1(n7565), .A2(n7564), .ZN(n7661) );
  OR2_X1 U9185 ( .A1(n7662), .A2(n7976), .ZN(n8056) );
  NAND2_X1 U9186 ( .A1(n7662), .A2(n7976), .ZN(n8043) );
  XNOR2_X1 U9187 ( .A(n7661), .B(n8023), .ZN(n9570) );
  INV_X1 U9188 ( .A(n9570), .ZN(n7579) );
  OAI21_X1 U9189 ( .B1(n8023), .B2(n7568), .A(n7668), .ZN(n7569) );
  NAND2_X1 U9190 ( .A1(n7569), .A2(n9189), .ZN(n7571) );
  AOI22_X1 U9191 ( .A1(n9363), .A2(n9045), .B1(n9044), .B2(n9664), .ZN(n7570)
         );
  NAND2_X1 U9192 ( .A1(n7571), .A2(n7570), .ZN(n9569) );
  AND2_X1 U9193 ( .A1(n7572), .A2(n7662), .ZN(n7573) );
  OR2_X1 U9194 ( .A1(n7573), .A2(n7672), .ZN(n9567) );
  OAI22_X1 U9195 ( .A1(n9692), .A2(n7574), .B1(n7901), .B2(n9693), .ZN(n7575)
         );
  AOI21_X1 U9196 ( .B1(n7662), .B2(n9309), .A(n7575), .ZN(n7576) );
  OAI21_X1 U9197 ( .B1(n9567), .B2(n9176), .A(n7576), .ZN(n7577) );
  AOI21_X1 U9198 ( .B1(n9569), .B2(n9692), .A(n7577), .ZN(n7578) );
  OAI21_X1 U9199 ( .B1(n7579), .B2(n9370), .A(n7578), .ZN(P1_U3278) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7583) );
  INV_X1 U9201 ( .A(n7580), .ZN(n7612) );
  OAI222_X1 U9202 ( .A1(n8311), .A2(n7583), .B1(n7582), .B2(n7612), .C1(n7581), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NOR2_X1 U9203 ( .A1(n7589), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7585) );
  NOR2_X1 U9204 ( .A1(n7585), .A2(n7584), .ZN(n7587) );
  INV_X1 U9205 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7844) );
  AOI22_X1 U9206 ( .A1(n7848), .A2(n7844), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7845), .ZN(n7586) );
  NOR2_X1 U9207 ( .A1(n7587), .A2(n7586), .ZN(n7843) );
  AOI21_X1 U9208 ( .B1(n7587), .B2(n7586), .A(n7843), .ZN(n7597) );
  INV_X1 U9209 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U9210 ( .A1(n7848), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9552), .B2(
        n7845), .ZN(n7591) );
  OAI21_X1 U9211 ( .B1(n7589), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7588), .ZN(
        n7590) );
  NAND2_X1 U9212 ( .A1(n7591), .A2(n7590), .ZN(n7847) );
  OAI21_X1 U9213 ( .B1(n7591), .B2(n7590), .A(n7847), .ZN(n7595) );
  NOR2_X1 U9214 ( .A1(n9777), .A2(n7845), .ZN(n7594) );
  INV_X1 U9215 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U9216 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7653) );
  OAI21_X1 U9217 ( .B1(n7592), .B2(n10172), .A(n7653), .ZN(n7593) );
  AOI211_X1 U9218 ( .C1(n7595), .C2(n9773), .A(n7594), .B(n7593), .ZN(n7596)
         );
  OAI21_X1 U9219 ( .B1(n7597), .B2(n9776), .A(n7596), .ZN(P2_U3259) );
  INV_X1 U9220 ( .A(n7598), .ZN(n7599) );
  AOI21_X1 U9221 ( .B1(n7601), .B2(n7600), .A(n7599), .ZN(n7610) );
  NOR2_X1 U9222 ( .A1(n7602), .A2(n9742), .ZN(n9749) );
  NOR2_X1 U9223 ( .A1(n9517), .A2(n7603), .ZN(n7608) );
  NAND2_X1 U9224 ( .A1(n9500), .A2(n9047), .ZN(n7605) );
  AND2_X1 U9225 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9638) );
  INV_X1 U9226 ( .A(n9638), .ZN(n7604) );
  OAI211_X1 U9227 ( .C1(n7606), .C2(n9503), .A(n7605), .B(n7604), .ZN(n7607)
         );
  AOI211_X1 U9228 ( .C1(n9749), .C2(n9513), .A(n7608), .B(n7607), .ZN(n7609)
         );
  OAI21_X1 U9229 ( .B1(n7610), .B2(n9509), .A(n7609), .ZN(P1_U3229) );
  OAI222_X1 U9230 ( .A1(n9479), .A2(n7612), .B1(P1_U3084), .B2(n5725), .C1(
        n7611), .C2(n7945), .ZN(P1_U3332) );
  INV_X1 U9231 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9232 ( .A1(n7614), .A2(n7613), .ZN(n7616) );
  XNOR2_X1 U9233 ( .A(n7616), .B(n7615), .ZN(n7686) );
  NAND2_X1 U9234 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  XNOR2_X1 U9235 ( .A(n7619), .B(n4899), .ZN(n7620) );
  INV_X1 U9236 ( .A(n8432), .ZN(n8498) );
  AOI222_X1 U9237 ( .A1(n9790), .A2(n7620), .B1(n8498), .B2(n9785), .C1(n8499), 
        .C2(n9787), .ZN(n7681) );
  AOI21_X1 U9238 ( .B1(n8449), .B2(n7621), .A(n4807), .ZN(n7684) );
  AOI22_X1 U9239 ( .A1(n7684), .A2(n9883), .B1(n9882), .B2(n8449), .ZN(n7622)
         );
  OAI211_X1 U9240 ( .C1(n9871), .C2(n7686), .A(n7681), .B(n7622), .ZN(n7625)
         );
  NAND2_X1 U9241 ( .A1(n7625), .A2(n9908), .ZN(n7623) );
  OAI21_X1 U9242 ( .B1(n9908), .B2(n7624), .A(n7623), .ZN(P2_U3484) );
  NAND2_X1 U9243 ( .A1(n7625), .A2(n9924), .ZN(n7626) );
  OAI21_X1 U9244 ( .B1(n9924), .B2(n7356), .A(n7626), .ZN(P2_U3531) );
  NAND2_X1 U9245 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  XNOR2_X1 U9246 ( .A(n7627), .B(n7630), .ZN(n7640) );
  NOR2_X1 U9247 ( .A1(n9517), .A2(n7631), .ZN(n7637) );
  NAND2_X1 U9248 ( .A1(n9500), .A2(n9046), .ZN(n7634) );
  INV_X1 U9249 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7632) );
  NOR2_X1 U9250 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7632), .ZN(n9651) );
  INV_X1 U9251 ( .A(n9651), .ZN(n7633) );
  OAI211_X1 U9252 ( .C1(n7635), .C2(n9503), .A(n7634), .B(n7633), .ZN(n7636)
         );
  AOI211_X1 U9253 ( .C1(n9038), .C2(n7638), .A(n7637), .B(n7636), .ZN(n7639)
         );
  OAI21_X1 U9254 ( .B1(n7640), .B2(n9509), .A(n7639), .ZN(P1_U3215) );
  INV_X1 U9255 ( .A(n7641), .ZN(n7644) );
  OAI222_X1 U9256 ( .A1(n7945), .A2(n7642), .B1(n9479), .B2(n7644), .C1(n9376), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U9257 ( .A1(n8311), .A2(n7645), .B1(n8894), .B2(n7644), .C1(
        P2_U3152), .C2(n7643), .ZN(P2_U3336) );
  INV_X1 U9258 ( .A(n7646), .ZN(n7649) );
  NOR3_X1 U9259 ( .A1(n7647), .A2(n7709), .A3(n8464), .ZN(n7648) );
  AOI21_X1 U9260 ( .B1(n7649), .B2(n8456), .A(n7648), .ZN(n7659) );
  INV_X1 U9261 ( .A(n7650), .ZN(n7656) );
  INV_X1 U9262 ( .A(n8280), .ZN(n8495) );
  AOI22_X1 U9263 ( .A1(n8480), .A2(n8495), .B1(n8481), .B2(n7710), .ZN(n7654)
         );
  NAND2_X1 U9264 ( .A1(n8277), .A2(n8455), .ZN(n7652) );
  INV_X1 U9265 ( .A(n7709), .ZN(n8497) );
  NAND2_X1 U9266 ( .A1(n8482), .A2(n8497), .ZN(n7651) );
  NAND4_X1 U9267 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n7655)
         );
  AOI21_X1 U9268 ( .B1(n7656), .B2(n8456), .A(n7655), .ZN(n7657) );
  OAI21_X1 U9269 ( .B1(n7659), .B2(n7658), .A(n7657), .ZN(P2_U3217) );
  OR2_X1 U9270 ( .A1(n7662), .A2(n9499), .ZN(n7660) );
  NAND2_X1 U9271 ( .A1(n7661), .A2(n7660), .ZN(n7664) );
  NAND2_X1 U9272 ( .A1(n7662), .A2(n9499), .ZN(n7663) );
  INV_X1 U9273 ( .A(n9044), .ZN(n9032) );
  OR2_X1 U9274 ( .A1(n7982), .A2(n9032), .ZN(n8062) );
  NAND2_X1 U9275 ( .A1(n7982), .A2(n9032), .ZN(n8128) );
  NAND2_X1 U9276 ( .A1(n8062), .A2(n8128), .ZN(n8026) );
  XOR2_X1 U9277 ( .A(n7741), .B(n8026), .Z(n9564) );
  INV_X1 U9278 ( .A(n9564), .ZN(n7679) );
  INV_X1 U9279 ( .A(n8043), .ZN(n7665) );
  NOR2_X1 U9280 ( .A1(n8026), .A2(n7665), .ZN(n7666) );
  NAND2_X1 U9281 ( .A1(n7746), .A2(n9189), .ZN(n7671) );
  INV_X1 U9282 ( .A(n8026), .ZN(n7667) );
  AOI21_X1 U9283 ( .B1(n7668), .B2(n8043), .A(n7667), .ZN(n7670) );
  AOI22_X1 U9284 ( .A1(n9363), .A2(n9499), .B1(n9043), .B2(n9664), .ZN(n7669)
         );
  OAI21_X1 U9285 ( .B1(n7671), .B2(n7670), .A(n7669), .ZN(n9563) );
  INV_X1 U9286 ( .A(n7982), .ZN(n9561) );
  OAI211_X1 U9287 ( .C1(n9561), .C2(n7672), .A(n4424), .B(n9728), .ZN(n9560)
         );
  OAI22_X1 U9288 ( .A1(n9692), .A2(n7673), .B1(n7980), .B2(n9693), .ZN(n7674)
         );
  AOI21_X1 U9289 ( .B1(n7982), .B2(n9309), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9290 ( .B1(n9560), .B2(n7676), .A(n7675), .ZN(n7677) );
  AOI21_X1 U9291 ( .B1(n9563), .B2(n9692), .A(n7677), .ZN(n7678) );
  OAI21_X1 U9292 ( .B1(n7679), .B2(n9370), .A(n7678), .ZN(P1_U3277) );
  AOI22_X1 U9293 ( .A1(n9808), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8448), .B2(
        n8778), .ZN(n7680) );
  OAI21_X1 U9294 ( .B1(n4901), .B2(n8781), .A(n7680), .ZN(n7683) );
  NOR2_X1 U9295 ( .A1(n7681), .A2(n9808), .ZN(n7682) );
  AOI211_X1 U9296 ( .C1(n7684), .C2(n9521), .A(n7683), .B(n7682), .ZN(n7685)
         );
  OAI21_X1 U9297 ( .B1(n8748), .B2(n7686), .A(n7685), .ZN(P2_U3285) );
  OAI21_X1 U9298 ( .B1(n7688), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7687), .ZN(
        n7823) );
  XNOR2_X1 U9299 ( .A(n7824), .B(n7823), .ZN(n7689) );
  INV_X1 U9300 ( .A(n7689), .ZN(n7692) );
  NOR2_X1 U9301 ( .A1(n7690), .A2(n7689), .ZN(n7825) );
  INV_X1 U9302 ( .A(n7825), .ZN(n7691) );
  OAI211_X1 U9303 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7692), .A(n9653), .B(
        n7691), .ZN(n7693) );
  NAND2_X1 U9304 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U9305 ( .C1(n9096), .C2(n7824), .A(n7693), .B(n9031), .ZN(n7700)
         );
  NOR2_X1 U9306 ( .A1(n7695), .A2(n7694), .ZN(n7697) );
  XNOR2_X1 U9307 ( .A(n7817), .B(n7824), .ZN(n7698) );
  INV_X1 U9308 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9309 ( .A1(n7743), .A2(n7698), .ZN(n7818) );
  AOI211_X1 U9310 ( .C1(n7698), .C2(n7743), .A(n7818), .B(n9647), .ZN(n7699)
         );
  AOI211_X1 U9311 ( .C1(n9656), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7700), .B(
        n7699), .ZN(n7701) );
  INV_X1 U9312 ( .A(n7701), .ZN(P1_U3256) );
  NAND2_X1 U9313 ( .A1(n8866), .A2(n8497), .ZN(n7705) );
  XNOR2_X1 U9314 ( .A(n8279), .B(n8278), .ZN(n9551) );
  INV_X1 U9315 ( .A(n9551), .ZN(n7716) );
  XNOR2_X1 U9316 ( .A(n7707), .B(n7706), .ZN(n7708) );
  OAI222_X1 U9317 ( .A1(n9533), .A2(n7709), .B1(n9535), .B2(n8280), .C1(n7708), 
        .C2(n9531), .ZN(n9549) );
  INV_X1 U9318 ( .A(n8277), .ZN(n9548) );
  OAI211_X1 U9319 ( .C1(n7790), .C2(n9548), .A(n9518), .B(n9883), .ZN(n9547)
         );
  AOI22_X1 U9320 ( .A1(n9808), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7710), .B2(
        n8778), .ZN(n7712) );
  NAND2_X1 U9321 ( .A1(n8277), .A2(n8598), .ZN(n7711) );
  OAI211_X1 U9322 ( .C1(n9547), .C2(n7713), .A(n7712), .B(n7711), .ZN(n7714)
         );
  AOI21_X1 U9323 ( .B1(n9549), .B2(n9791), .A(n7714), .ZN(n7715) );
  OAI21_X1 U9324 ( .B1(n7716), .B2(n8748), .A(n7715), .ZN(P2_U3282) );
  INV_X1 U9325 ( .A(n7721), .ZN(n7718) );
  AOI21_X1 U9326 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8892), .A(n6341), .ZN(
        n7717) );
  OAI21_X1 U9327 ( .B1(n7718), .B2(n8894), .A(n7717), .ZN(P2_U3335) );
  INV_X1 U9328 ( .A(n7719), .ZN(n7725) );
  OAI222_X1 U9329 ( .A1(n9479), .A2(n7725), .B1(P1_U3084), .B2(n7720), .C1(
        n9958), .C2(n7945), .ZN(P1_U3329) );
  NAND2_X1 U9330 ( .A1(n7721), .A2(n7878), .ZN(n7723) );
  OR2_X1 U9331 ( .A1(n7722), .A2(P1_U3084), .ZN(n8261) );
  OAI211_X1 U9332 ( .C1(n10022), .C2(n7945), .A(n7723), .B(n8261), .ZN(
        P1_U3330) );
  OAI222_X1 U9333 ( .A1(n7726), .A2(P2_U3152), .B1(n8894), .B2(n7725), .C1(
        n7724), .C2(n8311), .ZN(P2_U3334) );
  AOI21_X1 U9334 ( .B1(n7728), .B2(n7727), .A(n9509), .ZN(n7730) );
  NAND2_X1 U9335 ( .A1(n7730), .A2(n7729), .ZN(n7738) );
  INV_X1 U9336 ( .A(n7731), .ZN(n7736) );
  AOI21_X1 U9337 ( .B1(n9500), .B2(n9045), .A(n7732), .ZN(n7733) );
  OAI21_X1 U9338 ( .B1(n7734), .B2(n9503), .A(n7733), .ZN(n7735) );
  AOI21_X1 U9339 ( .B1(n7736), .B2(n8936), .A(n7735), .ZN(n7737) );
  OAI211_X1 U9340 ( .C1(n9576), .C2(n9020), .A(n7738), .B(n7737), .ZN(P1_U3234) );
  AND2_X1 U9341 ( .A1(n7982), .A2(n9044), .ZN(n7740) );
  INV_X1 U9342 ( .A(n9043), .ZN(n8952) );
  NOR2_X1 U9343 ( .A1(n9453), .A2(n8952), .ZN(n8133) );
  NAND2_X1 U9344 ( .A1(n9453), .A2(n8952), .ZN(n8068) );
  INV_X1 U9345 ( .A(n8068), .ZN(n8134) );
  XOR2_X1 U9346 ( .A(n7912), .B(n8131), .Z(n9455) );
  INV_X1 U9347 ( .A(n9453), .ZN(n7742) );
  AOI211_X1 U9348 ( .C1(n9453), .C2(n4424), .A(n9753), .B(n4605), .ZN(n9452)
         );
  NOR2_X1 U9349 ( .A1(n7742), .A2(n9694), .ZN(n7745) );
  OAI22_X1 U9350 ( .A1(n9692), .A2(n7743), .B1(n9036), .B2(n9693), .ZN(n7744)
         );
  AOI211_X1 U9351 ( .C1(n9452), .C2(n9340), .A(n7745), .B(n7744), .ZN(n7749)
         );
  INV_X1 U9352 ( .A(n9364), .ZN(n7798) );
  XOR2_X1 U9353 ( .A(n8131), .B(n7805), .Z(n7747) );
  OAI222_X1 U9354 ( .A1(n9683), .A2(n7798), .B1(n9685), .B2(n9032), .C1(n9672), 
        .C2(n7747), .ZN(n9451) );
  NAND2_X1 U9355 ( .A1(n9451), .A2(n9692), .ZN(n7748) );
  OAI211_X1 U9356 ( .C1(n9455), .C2(n9370), .A(n7749), .B(n7748), .ZN(P1_U3276) );
  INV_X1 U9357 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U9358 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7750) );
  AOI21_X1 U9359 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7750), .ZN(n9931) );
  NOR2_X1 U9360 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7751) );
  AOI21_X1 U9361 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7751), .ZN(n9934) );
  NAND2_X1 U9362 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7752) );
  OAI21_X1 U9363 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7752), .ZN(n9940) );
  NOR2_X1 U9364 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7753) );
  AOI21_X1 U9365 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7753), .ZN(n9943) );
  NOR2_X1 U9366 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7760) );
  XNOR2_X1 U9367 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10273) );
  NAND2_X1 U9368 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7758) );
  XOR2_X1 U9369 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10271) );
  NAND2_X1 U9370 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7756) );
  XOR2_X1 U9371 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10269) );
  AOI21_X1 U9372 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9925) );
  INV_X1 U9373 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7754) );
  NAND3_X1 U9374 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9927) );
  OAI21_X1 U9375 ( .B1(n9925), .B2(n7754), .A(n9927), .ZN(n10268) );
  NAND2_X1 U9376 ( .A1(n10269), .A2(n10268), .ZN(n7755) );
  NAND2_X1 U9377 ( .A1(n7756), .A2(n7755), .ZN(n10270) );
  NAND2_X1 U9378 ( .A1(n10271), .A2(n10270), .ZN(n7757) );
  NAND2_X1 U9379 ( .A1(n7758), .A2(n7757), .ZN(n10272) );
  NOR2_X1 U9380 ( .A1(n10273), .A2(n10272), .ZN(n7759) );
  NOR2_X1 U9381 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  NOR2_X1 U9382 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7761), .ZN(n10257) );
  AND2_X1 U9383 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7761), .ZN(n10256) );
  NOR2_X1 U9384 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10256), .ZN(n7762) );
  NAND2_X1 U9385 ( .A1(n7763), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7765) );
  XOR2_X1 U9386 ( .A(n7763), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10255) );
  NAND2_X1 U9387 ( .A1(n10255), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U9388 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  NAND2_X1 U9389 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7766), .ZN(n7768) );
  XOR2_X1 U9390 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7766), .Z(n10254) );
  NAND2_X1 U9391 ( .A1(n10254), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U9392 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  NAND2_X1 U9393 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7769), .ZN(n7771) );
  XOR2_X1 U9394 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7769), .Z(n10267) );
  NAND2_X1 U9395 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10267), .ZN(n7770) );
  NAND2_X1 U9396 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  AND2_X1 U9397 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7772), .ZN(n7773) );
  INV_X1 U9398 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10265) );
  XNOR2_X1 U9399 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7772), .ZN(n10264) );
  NOR2_X1 U9400 ( .A1(n10265), .A2(n10264), .ZN(n10263) );
  NAND2_X1 U9401 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7774) );
  OAI21_X1 U9402 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7774), .ZN(n9951) );
  NAND2_X1 U9403 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7775) );
  OAI21_X1 U9404 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7775), .ZN(n9948) );
  NOR2_X1 U9405 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7776) );
  AOI21_X1 U9406 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7776), .ZN(n9945) );
  NAND2_X1 U9407 ( .A1(n9946), .A2(n9945), .ZN(n9944) );
  NAND2_X1 U9408 ( .A1(n9943), .A2(n9942), .ZN(n9941) );
  AOI21_X1 U9409 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9938), .ZN(n9937) );
  NOR2_X1 U9410 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7777) );
  AOI21_X1 U9411 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7777), .ZN(n9936) );
  NAND2_X1 U9412 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  OAI21_X1 U9413 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9935), .ZN(n9933) );
  NAND2_X1 U9414 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  OAI21_X1 U9415 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9932), .ZN(n9930) );
  NAND2_X1 U9416 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  NOR2_X1 U9417 ( .A1(n10261), .A2(n10260), .ZN(n7778) );
  NAND2_X1 U9418 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  OAI21_X1 U9419 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7778), .A(n10259), .ZN(
        n7780) );
  XNOR2_X1 U9420 ( .A(n4803), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7779) );
  XNOR2_X1 U9421 ( .A(n7780), .B(n7779), .ZN(ADD_1071_U4) );
  OAI21_X1 U9422 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7789) );
  OAI22_X1 U9423 ( .A1(n9532), .A2(n9535), .B1(n8432), .B2(n9533), .ZN(n7788)
         );
  NAND2_X1 U9424 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U9425 ( .A1(n7786), .A2(n7785), .ZN(n8870) );
  NOR2_X1 U9426 ( .A1(n8870), .A2(n8774), .ZN(n7787) );
  AOI211_X1 U9427 ( .C1(n9790), .C2(n7789), .A(n7788), .B(n7787), .ZN(n8869)
         );
  AOI21_X1 U9428 ( .B1(n8866), .B2(n7791), .A(n7790), .ZN(n8867) );
  INV_X1 U9429 ( .A(n8866), .ZN(n7793) );
  AOI22_X1 U9430 ( .A1(n9808), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8437), .B2(
        n8778), .ZN(n7792) );
  OAI21_X1 U9431 ( .B1(n7793), .B2(n8781), .A(n7792), .ZN(n7795) );
  NOR2_X1 U9432 ( .A1(n8870), .A2(n8783), .ZN(n7794) );
  AOI211_X1 U9433 ( .C1(n8867), .C2(n9521), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI21_X1 U9434 ( .B1(n8869), .B2(n9808), .A(n7796), .ZN(P2_U3283) );
  NOR2_X1 U9435 ( .A1(n9453), .A2(n9043), .ZN(n7906) );
  OR2_X1 U9436 ( .A1(n7912), .A2(n7906), .ZN(n7797) );
  NAND2_X1 U9437 ( .A1(n9453), .A2(n9043), .ZN(n7908) );
  NAND2_X1 U9438 ( .A1(n7797), .A2(n7908), .ZN(n7799) );
  NAND2_X1 U9439 ( .A1(n7905), .A2(n7798), .ZN(n8069) );
  XNOR2_X1 U9440 ( .A(n7799), .B(n8135), .ZN(n9450) );
  INV_X1 U9441 ( .A(n7928), .ZN(n9355) );
  AOI211_X1 U9442 ( .C1(n7905), .C2(n7800), .A(n9753), .B(n7928), .ZN(n9448)
         );
  INV_X1 U9443 ( .A(n7905), .ZN(n7801) );
  NOR2_X1 U9444 ( .A1(n7801), .A2(n9694), .ZN(n7804) );
  INV_X1 U9445 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7802) );
  OAI22_X1 U9446 ( .A1(n9692), .A2(n7802), .B1(n8956), .B2(n9693), .ZN(n7803)
         );
  AOI211_X1 U9447 ( .C1(n9448), .C2(n9340), .A(n7804), .B(n7803), .ZN(n7808)
         );
  INV_X1 U9448 ( .A(n9042), .ZN(n7920) );
  XNOR2_X1 U9449 ( .A(n7916), .B(n8135), .ZN(n7806) );
  OAI222_X1 U9450 ( .A1(n9683), .A2(n7920), .B1(n9685), .B2(n8952), .C1(n7806), 
        .C2(n9672), .ZN(n9447) );
  NAND2_X1 U9451 ( .A1(n9447), .A2(n9692), .ZN(n7807) );
  OAI211_X1 U9452 ( .C1(n9450), .C2(n9370), .A(n7808), .B(n7807), .ZN(P1_U3275) );
  INV_X1 U9453 ( .A(n7809), .ZN(n7815) );
  OAI222_X1 U9454 ( .A1(n9479), .A2(n7815), .B1(P1_U3084), .B2(n7811), .C1(
        n7810), .C2(n7945), .ZN(P1_U3327) );
  INV_X1 U9455 ( .A(n7812), .ZN(n7943) );
  OAI222_X1 U9456 ( .A1(n8311), .A2(n10031), .B1(n8894), .B2(n7943), .C1(n7813), .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9457 ( .A1(n7816), .A2(P2_U3152), .B1(n8894), .B2(n7815), .C1(
        n7814), .C2(n8311), .ZN(P2_U3332) );
  NOR2_X1 U9458 ( .A1(n7817), .A2(n7824), .ZN(n7819) );
  NOR2_X1 U9459 ( .A1(n7819), .A2(n7818), .ZN(n7822) );
  NAND2_X1 U9460 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9080), .ZN(n7820) );
  OAI21_X1 U9461 ( .B1(n9080), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7820), .ZN(
        n7821) );
  NOR2_X1 U9462 ( .A1(n7822), .A2(n7821), .ZN(n9079) );
  AOI211_X1 U9463 ( .C1(n7822), .C2(n7821), .A(n9079), .B(n9647), .ZN(n7835)
         );
  NOR2_X1 U9464 ( .A1(n7824), .A2(n7823), .ZN(n7826) );
  NOR2_X1 U9465 ( .A1(n7826), .A2(n7825), .ZN(n7828) );
  XNOR2_X1 U9466 ( .A(n9080), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7827) );
  NOR2_X1 U9467 ( .A1(n7828), .A2(n7827), .ZN(n9076) );
  AOI211_X1 U9468 ( .C1(n7828), .C2(n7827), .A(n9076), .B(n9115), .ZN(n7834)
         );
  NAND2_X1 U9469 ( .A1(n9656), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7831) );
  NOR2_X1 U9470 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7829), .ZN(n8954) );
  INV_X1 U9471 ( .A(n8954), .ZN(n7830) );
  OAI211_X1 U9472 ( .C1(n9096), .C2(n7832), .A(n7831), .B(n7830), .ZN(n7833)
         );
  OR3_X1 U9473 ( .A1(n7835), .A2(n7834), .A3(n7833), .ZN(P1_U3257) );
  NAND2_X1 U9474 ( .A1(n7839), .A2(n7878), .ZN(n7837) );
  OAI211_X1 U9475 ( .C1(n7945), .C2(n7838), .A(n7837), .B(n7836), .ZN(P1_U3326) );
  INV_X1 U9476 ( .A(n7839), .ZN(n7841) );
  OAI222_X1 U9477 ( .A1(n8311), .A2(n7842), .B1(n8894), .B2(n7841), .C1(n7840), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  AOI21_X1 U9478 ( .B1(n7845), .B2(n7844), .A(n7843), .ZN(n7863) );
  XNOR2_X1 U9479 ( .A(n7863), .B(n7864), .ZN(n7846) );
  NOR2_X1 U9480 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7846), .ZN(n7865) );
  AOI21_X1 U9481 ( .B1(n7846), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7865), .ZN(
        n7855) );
  OAI21_X1 U9482 ( .B1(n7848), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7847), .ZN(
        n7856) );
  XNOR2_X1 U9483 ( .A(n7856), .B(n7857), .ZN(n7849) );
  INV_X1 U9484 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U9485 ( .A1(n10145), .A2(n7849), .ZN(n7858) );
  AOI211_X1 U9486 ( .C1(n7849), .C2(n10145), .A(n7858), .B(n9778), .ZN(n7853)
         );
  NOR2_X1 U9487 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8270), .ZN(n7850) );
  AOI21_X1 U9488 ( .B1(n9775), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7850), .ZN(
        n7851) );
  OAI21_X1 U9489 ( .B1(n9777), .B2(n7857), .A(n7851), .ZN(n7852) );
  NOR2_X1 U9490 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  OAI21_X1 U9491 ( .B1(n7855), .B2(n9776), .A(n7854), .ZN(P2_U3260) );
  NOR2_X1 U9492 ( .A1(n7857), .A2(n7856), .ZN(n7859) );
  XNOR2_X1 U9493 ( .A(n8508), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8509) );
  XNOR2_X1 U9494 ( .A(n8507), .B(n8509), .ZN(n7874) );
  NOR2_X1 U9495 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7860), .ZN(n7862) );
  NOR2_X1 U9496 ( .A1(n9777), .A2(n8513), .ZN(n7861) );
  AOI211_X1 U9497 ( .C1(n9775), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7862), .B(
        n7861), .ZN(n7873) );
  NOR2_X1 U9498 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  NOR2_X1 U9499 ( .A1(n7866), .A2(n7865), .ZN(n7871) );
  INV_X1 U9500 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9501 ( .A1(n8508), .A2(n7868), .ZN(n7867) );
  OAI21_X1 U9502 ( .B1(n8508), .B2(n7868), .A(n7867), .ZN(n7870) );
  NAND2_X1 U9503 ( .A1(n8513), .A2(n7868), .ZN(n7869) );
  OAI211_X1 U9504 ( .C1(n7868), .C2(n8513), .A(n7871), .B(n7869), .ZN(n8512)
         );
  OAI211_X1 U9505 ( .C1(n7871), .C2(n7870), .A(n8512), .B(n9774), .ZN(n7872)
         );
  OAI211_X1 U9506 ( .C1(n7874), .C2(n9778), .A(n7873), .B(n7872), .ZN(P2_U3261) );
  INV_X1 U9507 ( .A(n7879), .ZN(n7877) );
  NAND2_X1 U9508 ( .A1(n8892), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7875) );
  OAI211_X1 U9509 ( .C1(n7877), .C2(n8894), .A(n7876), .B(n7875), .ZN(P2_U3330) );
  NAND2_X1 U9510 ( .A1(n7879), .A2(n7878), .ZN(n7881) );
  OAI211_X1 U9511 ( .C1(n7945), .C2(n7882), .A(n7881), .B(n7880), .ZN(P1_U3325) );
  INV_X1 U9512 ( .A(n7883), .ZN(n7884) );
  AOI21_X1 U9513 ( .B1(n7885), .B2(n8275), .A(n7884), .ZN(n7890) );
  INV_X1 U9514 ( .A(n8779), .ZN(n7887) );
  OAI22_X1 U9515 ( .A1(n8280), .A2(n9533), .B1(n8471), .B2(n9535), .ZN(n8776)
         );
  AOI22_X1 U9516 ( .A1(n8315), .A2(n8776), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7886) );
  OAI21_X1 U9517 ( .B1(n8470), .B2(n7887), .A(n7886), .ZN(n7888) );
  AOI21_X1 U9518 ( .B1(n8861), .B2(n8455), .A(n7888), .ZN(n7889) );
  OAI21_X1 U9519 ( .B1(n7890), .B2(n8478), .A(n7889), .ZN(P2_U3228) );
  XNOR2_X1 U9520 ( .A(n7892), .B(n7891), .ZN(n7893) );
  XNOR2_X1 U9521 ( .A(n7894), .B(n7893), .ZN(n7904) );
  NOR2_X1 U9522 ( .A1(n7895), .A2(n9742), .ZN(n9565) );
  INV_X1 U9523 ( .A(n7896), .ZN(n7899) );
  NOR2_X1 U9524 ( .A1(n9503), .A2(n7897), .ZN(n7898) );
  AOI211_X1 U9525 ( .C1(n9500), .C2(n9044), .A(n7899), .B(n7898), .ZN(n7900)
         );
  OAI21_X1 U9526 ( .B1(n9517), .B2(n7901), .A(n7900), .ZN(n7902) );
  AOI21_X1 U9527 ( .B1(n9565), .B2(n9513), .A(n7902), .ZN(n7903) );
  OAI21_X1 U9528 ( .B1(n7904), .B2(n9509), .A(n7903), .ZN(P1_U3232) );
  OR2_X1 U9529 ( .A1(n7906), .A2(n7909), .ZN(n9348) );
  OR2_X1 U9530 ( .A1(n9442), .A2(n9042), .ZN(n7907) );
  INV_X1 U9531 ( .A(n7907), .ZN(n7910) );
  OR2_X1 U9532 ( .A1(n7912), .A2(n7913), .ZN(n7911) );
  NAND2_X1 U9533 ( .A1(n7911), .A2(n7914), .ZN(n7915) );
  INV_X1 U9534 ( .A(n9365), .ZN(n9335) );
  NAND2_X1 U9535 ( .A1(n9437), .A2(n9335), .ZN(n9330) );
  INV_X1 U9536 ( .A(n8028), .ZN(n7921) );
  OAI21_X1 U9537 ( .B1(n7915), .B2(n7921), .A(n9136), .ZN(n9441) );
  INV_X1 U9538 ( .A(n9362), .ZN(n7919) );
  AND2_X1 U9539 ( .A1(n9442), .A2(n7920), .ZN(n8042) );
  NAND2_X1 U9540 ( .A1(n7919), .A2(n7918), .ZN(n9150) );
  OR2_X1 U9541 ( .A1(n9442), .A2(n7920), .ZN(n8075) );
  NAND2_X1 U9542 ( .A1(n9150), .A2(n8075), .ZN(n7922) );
  XNOR2_X1 U9543 ( .A(n7922), .B(n7921), .ZN(n7923) );
  NAND2_X1 U9544 ( .A1(n7923), .A2(n9189), .ZN(n7925) );
  AOI22_X1 U9545 ( .A1(n9363), .A2(n9042), .B1(n9322), .B2(n9664), .ZN(n7924)
         );
  OAI22_X1 U9546 ( .A1(n9692), .A2(n7926), .B1(n9007), .B2(n9693), .ZN(n7927)
         );
  AOI21_X1 U9547 ( .B1(n9437), .B2(n9309), .A(n7927), .ZN(n7931) );
  AND2_X1 U9548 ( .A1(n9353), .A2(n9437), .ZN(n7929) );
  NOR2_X1 U9549 ( .A1(n9337), .A2(n7929), .ZN(n9438) );
  NAND2_X1 U9550 ( .A1(n9438), .A2(n9679), .ZN(n7930) );
  OAI211_X1 U9551 ( .C1(n9440), .C2(n4381), .A(n7931), .B(n7930), .ZN(n7932)
         );
  INV_X1 U9552 ( .A(n7932), .ZN(n7933) );
  OAI21_X1 U9553 ( .B1(n9441), .B2(n9370), .A(n7933), .ZN(P1_U3273) );
  INV_X1 U9554 ( .A(n8001), .ZN(n7936) );
  OAI22_X1 U9555 ( .A1(n8424), .A2(n8681), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10196), .ZN(n7939) );
  OAI22_X1 U9556 ( .A1(n8472), .A2(n8680), .B1(n8470), .B2(n8672), .ZN(n7938)
         );
  AOI211_X1 U9557 ( .C1(n8832), .C2(n8455), .A(n7939), .B(n7938), .ZN(n7942)
         );
  OR3_X1 U9558 ( .A1(n7940), .A2(n8372), .A3(n8464), .ZN(n7941) );
  OAI211_X1 U9559 ( .C1(n7937), .C2(n8478), .A(n7942), .B(n7941), .ZN(P2_U3237) );
  OAI222_X1 U9560 ( .A1(n7945), .A2(n7944), .B1(n9479), .B2(n7943), .C1(n5704), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI21_X1 U9561 ( .B1(n7946), .B2(n7948), .A(n7947), .ZN(n9886) );
  XNOR2_X1 U9562 ( .A(n7949), .B(n7950), .ZN(n7951) );
  NAND2_X1 U9563 ( .A1(n7951), .A2(n9790), .ZN(n7952) );
  OAI211_X1 U9564 ( .C1(n9886), .C2(n8774), .A(n7953), .B(n7952), .ZN(n9888)
         );
  MUX2_X1 U9565 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9888), .S(n9791), .Z(n7954)
         );
  INV_X1 U9566 ( .A(n7954), .ZN(n7962) );
  AND2_X1 U9567 ( .A1(n7955), .A2(n9881), .ZN(n7956) );
  NOR2_X1 U9568 ( .A1(n7957), .A2(n7956), .ZN(n9884) );
  INV_X1 U9569 ( .A(n9881), .ZN(n7959) );
  OAI22_X1 U9570 ( .A1(n8781), .A2(n7959), .B1(n9793), .B2(n7958), .ZN(n7960)
         );
  AOI21_X1 U9571 ( .B1(n9884), .B2(n9521), .A(n7960), .ZN(n7961) );
  OAI211_X1 U9572 ( .C1(n9886), .C2(n8783), .A(n7962), .B(n7961), .ZN(P2_U3288) );
  AOI22_X1 U9573 ( .A1(n9808), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8316), .B2(
        n8778), .ZN(n7963) );
  OAI21_X1 U9574 ( .B1(n7964), .B2(n8781), .A(n7963), .ZN(n7967) );
  NOR2_X1 U9575 ( .A1(n7965), .A2(n9808), .ZN(n7966) );
  AOI211_X1 U9576 ( .C1(n7969), .C2(n7968), .A(n7967), .B(n7966), .ZN(n7970)
         );
  OAI21_X1 U9577 ( .B1(n8748), .B2(n7971), .A(n7970), .ZN(P2_U3289) );
  XNOR2_X1 U9578 ( .A(n7973), .B(n7972), .ZN(n7974) );
  XNOR2_X1 U9579 ( .A(n7975), .B(n7974), .ZN(n7984) );
  NOR2_X1 U9580 ( .A1(n9503), .A2(n7976), .ZN(n7977) );
  AOI211_X1 U9581 ( .C1(n9500), .C2(n9043), .A(n7978), .B(n7977), .ZN(n7979)
         );
  OAI21_X1 U9582 ( .B1(n9517), .B2(n7980), .A(n7979), .ZN(n7981) );
  AOI21_X1 U9583 ( .B1(n9038), .B2(n7982), .A(n7981), .ZN(n7983) );
  OAI21_X1 U9584 ( .B1(n7984), .B2(n9509), .A(n7983), .ZN(P1_U3213) );
  AOI21_X1 U9585 ( .B1(n7986), .B2(n7985), .A(n7009), .ZN(n7991) );
  AOI22_X1 U9586 ( .A1(n9005), .A2(n9055), .B1(n9500), .B2(n9053), .ZN(n7990)
         );
  AOI22_X1 U9587 ( .A1(n9038), .A2(n7988), .B1(n7987), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7989) );
  OAI211_X1 U9588 ( .C1(n7991), .C2(n9509), .A(n7990), .B(n7989), .ZN(P1_U3235) );
  NAND2_X1 U9589 ( .A1(n8310), .A2(n8035), .ZN(n7993) );
  OR2_X1 U9590 ( .A1(n4405), .A2(n10227), .ZN(n7992) );
  NAND2_X1 U9591 ( .A1(n7994), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U9592 ( .A1(n5010), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U9593 ( .A1(n7995), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7996) );
  AND3_X1 U9594 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n10250) );
  NAND2_X1 U9595 ( .A1(n8001), .A2(n8035), .ZN(n8004) );
  OR2_X1 U9596 ( .A1(n4405), .A2(n8002), .ZN(n8003) );
  OR2_X1 U9597 ( .A1(n9380), .A2(n9191), .ZN(n8040) );
  NAND2_X1 U9598 ( .A1(n9380), .A2(n9191), .ZN(n8192) );
  NAND2_X1 U9599 ( .A1(n8040), .A2(n8192), .ZN(n9166) );
  INV_X1 U9600 ( .A(n9210), .ZN(n9171) );
  OR2_X2 U9601 ( .A1(n9388), .A2(n9171), .ZN(n9163) );
  NAND2_X1 U9602 ( .A1(n9388), .A2(n9171), .ZN(n9164) );
  INV_X1 U9603 ( .A(n9187), .ZN(n8033) );
  OR2_X2 U9604 ( .A1(n9392), .A2(n9227), .ZN(n9162) );
  NAND2_X1 U9605 ( .A1(n9392), .A2(n9227), .ZN(n8178) );
  AND2_X1 U9606 ( .A1(n9397), .A2(n9213), .ZN(n9160) );
  INV_X1 U9607 ( .A(n9160), .ZN(n8005) );
  OR2_X1 U9608 ( .A1(n9397), .A2(n9213), .ZN(n8173) );
  INV_X1 U9609 ( .A(n9262), .ZN(n9226) );
  NAND2_X1 U9610 ( .A1(n9400), .A2(n9226), .ZN(n8171) );
  OR2_X1 U9611 ( .A1(n9406), .A2(n9273), .ZN(n8241) );
  NAND2_X1 U9612 ( .A1(n9406), .A2(n9273), .ZN(n9242) );
  NOR2_X1 U9613 ( .A1(n9412), .A2(n9294), .ZN(n9158) );
  NAND2_X1 U9614 ( .A1(n9412), .A2(n9294), .ZN(n9157) );
  INV_X1 U9615 ( .A(n9267), .ZN(n9269) );
  INV_X1 U9616 ( .A(n9300), .ZN(n9272) );
  AND2_X1 U9617 ( .A1(n9417), .A2(n9272), .ZN(n9156) );
  INV_X1 U9618 ( .A(n9156), .ZN(n8157) );
  NAND2_X1 U9619 ( .A1(n9155), .A2(n8157), .ZN(n9290) );
  INV_X1 U9620 ( .A(n9323), .ZN(n9293) );
  OR2_X1 U9621 ( .A1(n9422), .A2(n9293), .ZN(n8155) );
  NAND2_X1 U9622 ( .A1(n9422), .A2(n9293), .ZN(n9154) );
  INV_X1 U9623 ( .A(n9307), .ZN(n8030) );
  INV_X1 U9624 ( .A(n9299), .ZN(n9336) );
  NOR2_X1 U9625 ( .A1(n9427), .A2(n9336), .ZN(n9152) );
  NAND2_X1 U9626 ( .A1(n9427), .A2(n9336), .ZN(n9153) );
  NAND2_X1 U9627 ( .A1(n4715), .A2(n9153), .ZN(n9320) );
  INV_X1 U9628 ( .A(n9322), .ZN(n9002) );
  OR2_X1 U9629 ( .A1(n9434), .A2(n9002), .ZN(n8147) );
  NAND2_X1 U9630 ( .A1(n9434), .A2(n9002), .ZN(n9151) );
  NAND2_X1 U9631 ( .A1(n8147), .A2(n9151), .ZN(n9329) );
  INV_X1 U9632 ( .A(n8075), .ZN(n8006) );
  INV_X1 U9633 ( .A(n9351), .ZN(n9361) );
  AND2_X1 U9634 ( .A1(n8012), .A2(n8007), .ZN(n8008) );
  NAND2_X1 U9635 ( .A1(n8009), .A2(n8008), .ZN(n8051) );
  NAND3_X1 U9636 ( .A1(n8011), .A2(n8010), .A3(n6942), .ZN(n8017) );
  NAND2_X1 U9637 ( .A1(n8222), .A2(n8217), .ZN(n8014) );
  NAND3_X1 U9638 ( .A1(n8014), .A2(n8013), .A3(n8012), .ZN(n8015) );
  NAND2_X1 U9639 ( .A1(n8015), .A2(n8223), .ZN(n8052) );
  OR4_X1 U9640 ( .A1(n8051), .A2(n8017), .A3(n8052), .A4(n8016), .ZN(n8021) );
  NOR4_X1 U9641 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n7269), .ZN(n8024)
         );
  NAND4_X1 U9642 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8122), .ZN(n8025)
         );
  NOR4_X1 U9643 ( .A1(n8135), .A2(n8131), .A3(n8026), .A4(n8025), .ZN(n8027)
         );
  NAND4_X1 U9644 ( .A1(n4720), .A2(n8028), .A3(n9361), .A4(n8027), .ZN(n8029)
         );
  NOR4_X1 U9645 ( .A1(n9290), .A2(n8030), .A3(n9320), .A4(n8029), .ZN(n8031)
         );
  NAND4_X1 U9646 ( .A1(n9223), .A2(n9243), .A3(n8164), .A4(n8031), .ZN(n8032)
         );
  NOR4_X1 U9647 ( .A1(n9166), .A2(n8033), .A3(n4510), .A4(n8032), .ZN(n8036)
         );
  NOR2_X1 U9648 ( .A1(n4405), .A2(n10121), .ZN(n8034) );
  INV_X1 U9649 ( .A(n9129), .ZN(n9371) );
  NAND3_X1 U9650 ( .A1(n8248), .A2(n8036), .A3(n8253), .ZN(n8038) );
  OR2_X1 U9651 ( .A1(n9371), .A2(n9127), .ZN(n8200) );
  NAND2_X1 U9652 ( .A1(n9558), .A2(n10250), .ZN(n8037) );
  NAND2_X1 U9653 ( .A1(n8200), .A2(n8037), .ZN(n8206) );
  OAI21_X1 U9654 ( .B1(n8038), .B2(n8206), .A(n5725), .ZN(n8201) );
  INV_X1 U9655 ( .A(n8201), .ZN(n8093) );
  OR2_X1 U9656 ( .A1(n9129), .A2(n8248), .ZN(n8039) );
  NAND2_X1 U9657 ( .A1(n8039), .A2(n8253), .ZN(n8182) );
  INV_X1 U9658 ( .A(n8182), .ZN(n8184) );
  AND2_X1 U9659 ( .A1(n8040), .A2(n9163), .ZN(n8089) );
  INV_X1 U9660 ( .A(n8089), .ZN(n8246) );
  AND2_X1 U9661 ( .A1(n8173), .A2(n9221), .ZN(n9161) );
  AND2_X1 U9662 ( .A1(n8171), .A2(n9242), .ZN(n9159) );
  NAND2_X1 U9663 ( .A1(n8241), .A2(n4704), .ZN(n8041) );
  NAND2_X1 U9664 ( .A1(n9159), .A2(n8041), .ZN(n8162) );
  INV_X1 U9665 ( .A(n8162), .ZN(n8083) );
  NOR2_X1 U9666 ( .A1(n9158), .A2(n4708), .ZN(n8207) );
  NAND2_X1 U9667 ( .A1(n9330), .A2(n7918), .ZN(n8142) );
  INV_X1 U9668 ( .A(n8069), .ZN(n8138) );
  NAND2_X1 U9669 ( .A1(n8128), .A2(n8043), .ZN(n8123) );
  INV_X1 U9670 ( .A(n8123), .ZN(n8049) );
  NAND2_X1 U9671 ( .A1(n8121), .A2(n8044), .ZN(n8124) );
  INV_X1 U9672 ( .A(n8111), .ZN(n8045) );
  NOR2_X1 U9673 ( .A1(n8109), .A2(n8045), .ZN(n8046) );
  OR2_X1 U9674 ( .A1(n8124), .A2(n8046), .ZN(n8061) );
  INV_X1 U9675 ( .A(n8061), .ZN(n8048) );
  AND2_X1 U9676 ( .A1(n8096), .A2(n8107), .ZN(n8047) );
  NAND4_X1 U9677 ( .A1(n8068), .A2(n8049), .A3(n8048), .A4(n8047), .ZN(n8050)
         );
  OR3_X1 U9678 ( .A1(n8142), .A2(n8138), .A3(n8050), .ZN(n8232) );
  INV_X1 U9679 ( .A(n8051), .ZN(n8220) );
  NAND2_X1 U9680 ( .A1(n8220), .A2(n9682), .ZN(n8055) );
  NAND2_X1 U9681 ( .A1(n8052), .A2(n8100), .ZN(n8054) );
  INV_X1 U9682 ( .A(n8219), .ZN(n8053) );
  AOI21_X1 U9683 ( .B1(n8055), .B2(n8054), .A(n8053), .ZN(n8073) );
  INV_X1 U9684 ( .A(n8133), .ZN(n8067) );
  NAND2_X1 U9685 ( .A1(n8062), .A2(n8056), .ZN(n8129) );
  NAND2_X1 U9686 ( .A1(n8125), .A2(n8057), .ZN(n8058) );
  AND2_X1 U9687 ( .A1(n8058), .A2(n8121), .ZN(n8059) );
  NOR2_X1 U9688 ( .A1(n8129), .A2(n8059), .ZN(n8126) );
  INV_X1 U9689 ( .A(n8126), .ZN(n8065) );
  AND2_X1 U9690 ( .A1(n8108), .A2(n8111), .ZN(n8060) );
  NOR2_X1 U9691 ( .A1(n8061), .A2(n8060), .ZN(n8064) );
  AND2_X1 U9692 ( .A1(n8123), .A2(n8062), .ZN(n8130) );
  INV_X1 U9693 ( .A(n8130), .ZN(n8063) );
  OAI21_X1 U9694 ( .B1(n8065), .B2(n8064), .A(n8063), .ZN(n8066) );
  NAND2_X1 U9695 ( .A1(n8067), .A2(n8066), .ZN(n8070) );
  NAND3_X1 U9696 ( .A1(n8070), .A2(n8069), .A3(n8068), .ZN(n8071) );
  AND2_X1 U9697 ( .A1(n8071), .A2(n8137), .ZN(n8072) );
  OR2_X1 U9698 ( .A1(n8142), .A2(n8072), .ZN(n8230) );
  OAI21_X1 U9699 ( .B1(n8232), .B2(n8073), .A(n8230), .ZN(n8074) );
  AND2_X1 U9700 ( .A1(n8074), .A2(n9151), .ZN(n8080) );
  AND2_X1 U9701 ( .A1(n8146), .A2(n8075), .ZN(n9149) );
  NAND2_X1 U9702 ( .A1(n9151), .A2(n9330), .ZN(n8151) );
  INV_X1 U9703 ( .A(n8147), .ZN(n8076) );
  NOR2_X1 U9704 ( .A1(n9152), .A2(n8076), .ZN(n8150) );
  OAI211_X1 U9705 ( .C1(n9149), .C2(n8151), .A(n8150), .B(n8155), .ZN(n8235)
         );
  INV_X1 U9706 ( .A(n9153), .ZN(n8077) );
  NAND2_X1 U9707 ( .A1(n8155), .A2(n8077), .ZN(n8078) );
  NAND2_X1 U9708 ( .A1(n8078), .A2(n9154), .ZN(n8079) );
  NOR2_X1 U9709 ( .A1(n9156), .A2(n8079), .ZN(n8236) );
  OAI21_X1 U9710 ( .B1(n8080), .B2(n8235), .A(n8236), .ZN(n8081) );
  NAND3_X1 U9711 ( .A1(n8207), .A2(n8241), .A3(n8081), .ZN(n8082) );
  NAND2_X1 U9712 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  NAND3_X1 U9713 ( .A1(n9162), .A2(n9161), .A3(n8084), .ZN(n8090) );
  OR2_X1 U9714 ( .A1(n9127), .A2(n10250), .ZN(n8085) );
  NAND2_X1 U9715 ( .A1(n9558), .A2(n8085), .ZN(n8186) );
  NAND2_X1 U9716 ( .A1(n9162), .A2(n9160), .ZN(n8086) );
  NAND3_X1 U9717 ( .A1(n9164), .A2(n8178), .A3(n8086), .ZN(n8088) );
  INV_X1 U9718 ( .A(n8192), .ZN(n8087) );
  AOI21_X1 U9719 ( .B1(n8089), .B2(n8088), .A(n8087), .ZN(n8247) );
  OAI211_X1 U9720 ( .C1(n8246), .C2(n8090), .A(n8186), .B(n8247), .ZN(n8091)
         );
  NAND2_X1 U9721 ( .A1(n8200), .A2(n5049), .ZN(n8203) );
  AOI21_X1 U9722 ( .B1(n8184), .B2(n8091), .A(n8203), .ZN(n8092) );
  NOR2_X1 U9723 ( .A1(n8093), .A2(n8092), .ZN(n8202) );
  NAND2_X1 U9724 ( .A1(n9376), .A2(n9670), .ZN(n8188) );
  OAI21_X1 U9725 ( .B1(n9050), .B2(n8188), .A(n8094), .ZN(n8106) );
  OAI21_X1 U9726 ( .B1(n8095), .B2(n4535), .A(n9736), .ZN(n8105) );
  NAND3_X1 U9727 ( .A1(n8097), .A2(n8096), .A3(n8188), .ZN(n8098) );
  AOI21_X1 U9728 ( .B1(n8099), .B2(n8101), .A(n8098), .ZN(n8104) );
  NAND2_X1 U9729 ( .A1(n8100), .A2(n8219), .ZN(n8224) );
  AOI211_X1 U9730 ( .C1(n8102), .C2(n8101), .A(n8188), .B(n8224), .ZN(n8103)
         );
  AND2_X1 U9731 ( .A1(n8109), .A2(n8107), .ZN(n8114) );
  INV_X1 U9732 ( .A(n8125), .ZN(n8113) );
  INV_X1 U9733 ( .A(n8108), .ZN(n8110) );
  NAND2_X1 U9734 ( .A1(n8110), .A2(n8109), .ZN(n8112) );
  NAND2_X1 U9735 ( .A1(n8112), .A2(n8111), .ZN(n8115) );
  AOI211_X1 U9736 ( .C1(n8118), .C2(n8114), .A(n8113), .B(n8115), .ZN(n8120)
         );
  INV_X1 U9737 ( .A(n8114), .ZN(n8117) );
  INV_X1 U9738 ( .A(n8115), .ZN(n8116) );
  OAI21_X1 U9739 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n8119) );
  AOI21_X1 U9740 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8127) );
  MUX2_X1 U9741 ( .A(n8127), .B(n8126), .S(n8188), .Z(n8132) );
  MUX2_X1 U9742 ( .A(n8134), .B(n8133), .S(n8188), .Z(n8136) );
  INV_X1 U9743 ( .A(n8137), .ZN(n8139) );
  MUX2_X1 U9744 ( .A(n8139), .B(n8138), .S(n8188), .Z(n8140) );
  NOR3_X1 U9745 ( .A1(n8141), .A2(n8140), .A3(n9351), .ZN(n8145) );
  INV_X1 U9746 ( .A(n9149), .ZN(n8143) );
  MUX2_X1 U9747 ( .A(n8143), .B(n8142), .S(n4535), .Z(n8144) );
  INV_X1 U9748 ( .A(n8152), .ZN(n8148) );
  NAND3_X1 U9749 ( .A1(n8148), .A2(n8147), .A3(n8146), .ZN(n8149) );
  NAND3_X1 U9750 ( .A1(n8149), .A2(n9153), .A3(n9151), .ZN(n8154) );
  OAI21_X1 U9751 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8153) );
  INV_X1 U9752 ( .A(n8155), .ZN(n8158) );
  INV_X1 U9753 ( .A(n9154), .ZN(n8156) );
  INV_X1 U9754 ( .A(n8241), .ZN(n8159) );
  OAI21_X1 U9755 ( .B1(n8159), .B2(n9158), .A(n9242), .ZN(n8160) );
  NAND2_X1 U9756 ( .A1(n8160), .A2(n9221), .ZN(n8161) );
  MUX2_X1 U9757 ( .A(n8162), .B(n8161), .S(n8188), .Z(n8163) );
  INV_X1 U9758 ( .A(n8178), .ZN(n8166) );
  AOI21_X1 U9759 ( .B1(n9397), .B2(n9221), .A(n8166), .ZN(n8169) );
  INV_X1 U9760 ( .A(n9162), .ZN(n8167) );
  AOI21_X1 U9761 ( .B1(n9246), .B2(n8171), .A(n8167), .ZN(n8168) );
  MUX2_X1 U9762 ( .A(n8169), .B(n8168), .S(n8188), .Z(n8170) );
  NOR2_X1 U9763 ( .A1(n9397), .A2(n9246), .ZN(n9146) );
  OAI21_X1 U9764 ( .B1(n9397), .B2(n9221), .A(n9213), .ZN(n8175) );
  INV_X1 U9765 ( .A(n8171), .ZN(n8172) );
  NAND2_X1 U9766 ( .A1(n8173), .A2(n8172), .ZN(n8242) );
  NAND2_X1 U9767 ( .A1(n8242), .A2(n9232), .ZN(n8174) );
  MUX2_X1 U9768 ( .A(n8175), .B(n8174), .S(n8188), .Z(n8176) );
  MUX2_X1 U9769 ( .A(n9162), .B(n8178), .S(n8188), .Z(n8179) );
  MUX2_X1 U9770 ( .A(n9164), .B(n9163), .S(n8188), .Z(n8180) );
  OAI21_X1 U9771 ( .B1(n9180), .B2(n8188), .A(n8186), .ZN(n8181) );
  OAI21_X1 U9772 ( .B1(n8183), .B2(n9191), .A(n8184), .ZN(n8190) );
  INV_X1 U9773 ( .A(n8253), .ZN(n8185) );
  AOI21_X1 U9774 ( .B1(n8187), .B2(n8186), .A(n8185), .ZN(n8189) );
  INV_X1 U9775 ( .A(n8191), .ZN(n8193) );
  OAI21_X1 U9776 ( .B1(n8193), .B2(n9041), .A(n8192), .ZN(n8194) );
  AND2_X1 U9777 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  INV_X1 U9778 ( .A(n8198), .ZN(n8199) );
  NOR3_X1 U9779 ( .A1(n8204), .A2(n5726), .A3(n8203), .ZN(n8205) );
  INV_X1 U9780 ( .A(n8206), .ZN(n8252) );
  INV_X1 U9781 ( .A(n8208), .ZN(n8211) );
  NAND2_X1 U9782 ( .A1(n8209), .A2(n9055), .ZN(n8210) );
  NAND3_X1 U9783 ( .A1(n8211), .A2(n8210), .A3(n5049), .ZN(n8213) );
  NAND2_X1 U9784 ( .A1(n8213), .A2(n8212), .ZN(n8215) );
  OAI21_X1 U9785 ( .B1(n8216), .B2(n8215), .A(n8214), .ZN(n8218) );
  NAND2_X1 U9786 ( .A1(n8218), .A2(n8217), .ZN(n8221) );
  NAND3_X1 U9787 ( .A1(n8221), .A2(n8220), .A3(n8219), .ZN(n8229) );
  NAND2_X1 U9788 ( .A1(n8223), .A2(n8222), .ZN(n8227) );
  INV_X1 U9789 ( .A(n8224), .ZN(n8226) );
  NAND3_X1 U9790 ( .A1(n8227), .A2(n8226), .A3(n8225), .ZN(n8228) );
  NAND2_X1 U9791 ( .A1(n8229), .A2(n8228), .ZN(n8231) );
  OAI21_X1 U9792 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8233) );
  AND2_X1 U9793 ( .A1(n8233), .A2(n9151), .ZN(n8234) );
  NOR2_X1 U9794 ( .A1(n8235), .A2(n8234), .ZN(n8238) );
  INV_X1 U9795 ( .A(n8236), .ZN(n8237) );
  NOR2_X1 U9796 ( .A1(n8238), .A2(n8237), .ZN(n8239) );
  OAI211_X1 U9797 ( .C1(n4706), .C2(n8239), .A(n9242), .B(n9157), .ZN(n8240)
         );
  NAND3_X1 U9798 ( .A1(n9161), .A2(n8241), .A3(n8240), .ZN(n8243) );
  NAND2_X1 U9799 ( .A1(n8243), .A2(n8242), .ZN(n8244) );
  NAND2_X1 U9800 ( .A1(n9208), .A2(n8244), .ZN(n8245) );
  NOR2_X1 U9801 ( .A1(n8246), .A2(n8245), .ZN(n8250) );
  INV_X1 U9802 ( .A(n8247), .ZN(n8249) );
  OAI21_X1 U9803 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8251) );
  NAND2_X1 U9804 ( .A1(n8252), .A2(n8251), .ZN(n8254) );
  NAND2_X1 U9805 ( .A1(n8254), .A2(n8253), .ZN(n8258) );
  NAND2_X1 U9806 ( .A1(n8258), .A2(n8255), .ZN(n8257) );
  INV_X1 U9807 ( .A(n8261), .ZN(n8256) );
  OAI211_X1 U9808 ( .C1(n8258), .C2(n9374), .A(n8257), .B(n8256), .ZN(n8264)
         );
  NOR4_X1 U9809 ( .A1(n8260), .A2(n8259), .A3(n4378), .A4(n9603), .ZN(n8263)
         );
  OAI21_X1 U9810 ( .B1(n5726), .B2(n8261), .A(P1_B_REG_SCAN_IN), .ZN(n8262) );
  OAI22_X1 U9811 ( .A1(n8265), .A2(n8264), .B1(n8263), .B2(n8262), .ZN(
        P1_U3240) );
  NAND2_X1 U9812 ( .A1(n8266), .A2(n8456), .ZN(n8276) );
  INV_X1 U9813 ( .A(n8267), .ZN(n8269) );
  OAI211_X1 U9814 ( .C1(n8269), .C2(n8268), .A(n8412), .B(n8495), .ZN(n8274)
         );
  OAI22_X1 U9815 ( .A1(n8472), .A2(n9532), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8270), .ZN(n8272) );
  OAI22_X1 U9816 ( .A1(n8424), .A2(n9534), .B1(n8470), .B2(n9541), .ZN(n8271)
         );
  AOI211_X1 U9817 ( .C1(n8294), .C2(n8455), .A(n8272), .B(n8271), .ZN(n8273)
         );
  OAI211_X1 U9818 ( .C1(n8276), .C2(n8275), .A(n8274), .B(n8273), .ZN(P2_U3243) );
  INV_X1 U9819 ( .A(n9532), .ZN(n8496) );
  NAND2_X1 U9820 ( .A1(n9525), .A2(n9524), .ZN(n9523) );
  NAND2_X1 U9821 ( .A1(n9542), .A2(n8280), .ZN(n8281) );
  INV_X1 U9822 ( .A(n9534), .ZN(n8494) );
  INV_X1 U9823 ( .A(n8471), .ZN(n8742) );
  NAND2_X1 U9824 ( .A1(n8852), .A2(n8493), .ZN(n8283) );
  AOI21_X1 U9825 ( .B1(n8735), .B2(n8283), .A(n4472), .ZN(n8725) );
  NAND2_X1 U9826 ( .A1(n8725), .A2(n4771), .ZN(n8724) );
  NAND2_X1 U9827 ( .A1(n8849), .A2(n8743), .ZN(n8285) );
  NAND2_X1 U9828 ( .A1(n8724), .A2(n8285), .ZN(n8704) );
  NAND2_X1 U9829 ( .A1(n8842), .A2(n8697), .ZN(n8286) );
  NAND2_X1 U9830 ( .A1(n8703), .A2(n8286), .ZN(n8687) );
  OR2_X1 U9831 ( .A1(n8837), .A2(n8713), .ZN(n8287) );
  NAND2_X1 U9832 ( .A1(n8687), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U9833 ( .A1(n8837), .A2(n8713), .ZN(n8288) );
  INV_X1 U9834 ( .A(n8681), .ZN(n8492) );
  NAND2_X1 U9835 ( .A1(n8618), .A2(n8622), .ZN(n8617) );
  OR2_X1 U9836 ( .A1(n8818), .A2(n8490), .ZN(n8292) );
  NAND2_X1 U9837 ( .A1(n8576), .A2(n8293), .ZN(n8561) );
  NAND2_X1 U9838 ( .A1(n8561), .A2(n8569), .ZN(n8562) );
  INV_X1 U9839 ( .A(n8852), .ZN(n8739) );
  INV_X1 U9840 ( .A(n8837), .ZN(n8694) );
  INV_X1 U9841 ( .A(n8822), .ZN(n8641) );
  INV_X1 U9842 ( .A(n8794), .ZN(n8299) );
  INV_X1 U9843 ( .A(n8296), .ZN(n8297) );
  AOI22_X1 U9844 ( .A1(n9808), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8778), .B2(
        n8297), .ZN(n8298) );
  OAI21_X1 U9845 ( .B1(n8299), .B2(n8781), .A(n8298), .ZN(n8308) );
  OAI21_X1 U9846 ( .B1(n4423), .B2(n8301), .A(n8300), .ZN(n8306) );
  AOI21_X1 U9847 ( .B1(n8302), .B2(P2_B_REG_SCAN_IN), .A(n9535), .ZN(n8550) );
  NAND2_X1 U9848 ( .A1(n8489), .A2(n8550), .ZN(n8303) );
  NOR2_X1 U9849 ( .A1(n8797), .A2(n9808), .ZN(n8307) );
  OAI21_X1 U9850 ( .B1(n8798), .B2(n8748), .A(n8309), .ZN(P2_U3267) );
  INV_X1 U9851 ( .A(n8310), .ZN(n9478) );
  OAI222_X1 U9852 ( .A1(P2_U3152), .A2(n5784), .B1(n8894), .B2(n9478), .C1(
        n10251), .C2(n8311), .ZN(P2_U3328) );
  OAI211_X1 U9853 ( .C1(n8313), .C2(n8312), .A(n7275), .B(n8456), .ZN(n8321)
         );
  AOI22_X1 U9854 ( .A1(n8315), .A2(n8314), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n8320) );
  NAND2_X1 U9855 ( .A1(n8481), .A2(n8316), .ZN(n8319) );
  NAND2_X1 U9856 ( .A1(n8455), .A2(n8317), .ZN(n8318) );
  NAND4_X1 U9857 ( .A1(n8321), .A2(n8320), .A3(n8319), .A4(n8318), .ZN(
        P2_U3215) );
  NOR2_X1 U9858 ( .A1(n8477), .A2(n8322), .ZN(n8325) );
  NAND3_X1 U9859 ( .A1(n8323), .A2(n8412), .A3(n8624), .ZN(n8324) );
  NAND2_X1 U9860 ( .A1(n8327), .A2(n8326), .ZN(n8332) );
  NOR2_X1 U9861 ( .A1(n8470), .A2(n8581), .ZN(n8330) );
  OAI22_X1 U9862 ( .A1(n8424), .A2(n8328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10110), .ZN(n8329) );
  AOI211_X1 U9863 ( .C1(n8482), .C2(n8624), .A(n8330), .B(n8329), .ZN(n8331)
         );
  OAI211_X1 U9864 ( .C1(n8584), .C2(n8485), .A(n8332), .B(n8331), .ZN(P2_U3216) );
  INV_X1 U9865 ( .A(n8333), .ZN(n8334) );
  NAND2_X1 U9866 ( .A1(n7937), .A2(n8334), .ZN(n8336) );
  XNOR2_X1 U9867 ( .A(n8336), .B(n8335), .ZN(n8337) );
  NAND3_X1 U9868 ( .A1(n8337), .A2(n8412), .A3(n8492), .ZN(n8344) );
  INV_X1 U9869 ( .A(n8337), .ZN(n8339) );
  NAND3_X1 U9870 ( .A1(n8339), .A2(n8456), .A3(n8338), .ZN(n8343) );
  OAI22_X1 U9871 ( .A1(n8472), .A2(n8372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10234), .ZN(n8341) );
  OAI22_X1 U9872 ( .A1(n8424), .A2(n8398), .B1(n8470), .B2(n8655), .ZN(n8340)
         );
  AOI211_X1 U9873 ( .C1(n8827), .C2(n8455), .A(n8341), .B(n8340), .ZN(n8342)
         );
  NAND3_X1 U9874 ( .A1(n8344), .A2(n8343), .A3(n8342), .ZN(P2_U3218) );
  AOI21_X1 U9875 ( .B1(n8346), .B2(n8345), .A(n8478), .ZN(n8348) );
  NAND2_X1 U9876 ( .A1(n8348), .A2(n8347), .ZN(n8355) );
  AOI21_X1 U9877 ( .B1(n8480), .B2(n4900), .A(n8349), .ZN(n8354) );
  AOI22_X1 U9878 ( .A1(n8482), .A2(n8500), .B1(n8481), .B2(n8350), .ZN(n8353)
         );
  NAND2_X1 U9879 ( .A1(n8455), .A2(n8351), .ZN(n8352) );
  NAND4_X1 U9880 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(
        P2_U3219) );
  INV_X1 U9881 ( .A(n8849), .ZN(n8730) );
  NOR3_X1 U9882 ( .A1(n4978), .A2(n8356), .A3(n8478), .ZN(n8362) );
  NAND3_X1 U9883 ( .A1(n8357), .A2(n8412), .A3(n8743), .ZN(n8358) );
  OAI21_X1 U9884 ( .B1(n8359), .B2(n8478), .A(n8358), .ZN(n8361) );
  MUX2_X1 U9885 ( .A(n8362), .B(n8361), .S(n8360), .Z(n8363) );
  INV_X1 U9886 ( .A(n8363), .ZN(n8368) );
  AOI22_X1 U9887 ( .A1(n8697), .A2(n9785), .B1(n9787), .B2(n8493), .ZN(n8722)
         );
  OAI22_X1 U9888 ( .A1(n8365), .A2(n8722), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8364), .ZN(n8366) );
  AOI21_X1 U9889 ( .B1(n8728), .B2(n8481), .A(n8366), .ZN(n8367) );
  OAI211_X1 U9890 ( .C1(n8730), .C2(n8485), .A(n8368), .B(n8367), .ZN(P2_U3221) );
  XNOR2_X1 U9891 ( .A(n8370), .B(n8369), .ZN(n8377) );
  OAI22_X1 U9892 ( .A1(n8424), .A2(n8372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8371), .ZN(n8375) );
  OAI22_X1 U9893 ( .A1(n8472), .A2(n8373), .B1(n8470), .B2(n8691), .ZN(n8374)
         );
  AOI211_X1 U9894 ( .C1(n8837), .C2(n8455), .A(n8375), .B(n8374), .ZN(n8376)
         );
  OAI21_X1 U9895 ( .B1(n8377), .B2(n8478), .A(n8376), .ZN(P2_U3225) );
  INV_X1 U9896 ( .A(n8379), .ZN(n8380) );
  AOI21_X1 U9897 ( .B1(n8378), .B2(n8380), .A(n8478), .ZN(n8385) );
  NOR3_X1 U9898 ( .A1(n8464), .A2(n8382), .A3(n8381), .ZN(n8384) );
  OAI21_X1 U9899 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8392) );
  AOI21_X1 U9900 ( .B1(n8480), .B2(n8497), .A(n8386), .ZN(n8391) );
  AOI22_X1 U9901 ( .A1(n8482), .A2(n4900), .B1(n8481), .B2(n8387), .ZN(n8390)
         );
  NAND2_X1 U9902 ( .A1(n8455), .A2(n8388), .ZN(n8389) );
  NAND4_X1 U9903 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(
        P2_U3226) );
  XNOR2_X1 U9904 ( .A(n8395), .B(n8394), .ZN(n8396) );
  XNOR2_X1 U9905 ( .A(n4390), .B(n8396), .ZN(n8404) );
  OAI22_X1 U9906 ( .A1(n8472), .A2(n8398), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8397), .ZN(n8402) );
  INV_X1 U9907 ( .A(n8627), .ZN(n8399) );
  OAI22_X1 U9908 ( .A1(n8424), .A2(n8400), .B1(n8470), .B2(n8399), .ZN(n8401)
         );
  AOI211_X1 U9909 ( .C1(n8818), .C2(n8455), .A(n8402), .B(n8401), .ZN(n8403)
         );
  OAI21_X1 U9910 ( .B1(n8404), .B2(n8478), .A(n8403), .ZN(P2_U3227) );
  OR2_X1 U9911 ( .A1(n8407), .A2(n8406), .ZN(n8463) );
  INV_X1 U9912 ( .A(n8463), .ZN(n8405) );
  AOI22_X1 U9913 ( .A1(n8480), .A2(n8493), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8409) );
  AOI22_X1 U9914 ( .A1(n8482), .A2(n8494), .B1(n8481), .B2(n8751), .ZN(n8408)
         );
  OAI211_X1 U9915 ( .C1(n8860), .C2(n8485), .A(n8409), .B(n8408), .ZN(n8410)
         );
  OR2_X1 U9916 ( .A1(n8411), .A2(n8410), .ZN(P2_U3230) );
  NAND2_X1 U9917 ( .A1(n8412), .A2(n8663), .ZN(n8416) );
  OR2_X1 U9918 ( .A1(n8478), .A2(n8413), .ZN(n8415) );
  MUX2_X1 U9919 ( .A(n8416), .B(n8415), .S(n8414), .Z(n8420) );
  OAI22_X1 U9920 ( .A1(n8472), .A2(n8681), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10225), .ZN(n8418) );
  OAI22_X1 U9921 ( .A1(n8424), .A2(n8645), .B1(n8470), .B2(n8638), .ZN(n8417)
         );
  AOI211_X1 U9922 ( .C1(n8822), .C2(n8455), .A(n8418), .B(n8417), .ZN(n8419)
         );
  NAND2_X1 U9923 ( .A1(n8420), .A2(n8419), .ZN(P2_U3231) );
  XNOR2_X1 U9924 ( .A(n8422), .B(n8421), .ZN(n8429) );
  OAI22_X1 U9925 ( .A1(n8424), .A2(n8680), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8423), .ZN(n8427) );
  OAI22_X1 U9926 ( .A1(n8472), .A2(n8425), .B1(n8470), .B2(n8706), .ZN(n8426)
         );
  AOI211_X1 U9927 ( .C1(n8842), .C2(n8455), .A(n8427), .B(n8426), .ZN(n8428)
         );
  OAI21_X1 U9928 ( .B1(n8429), .B2(n8478), .A(n8428), .ZN(P2_U3235) );
  INV_X1 U9929 ( .A(n8430), .ZN(n8431) );
  AOI21_X1 U9930 ( .B1(n8383), .B2(n8431), .A(n8478), .ZN(n8435) );
  NOR3_X1 U9931 ( .A1(n8433), .A2(n8464), .A3(n8432), .ZN(n8434) );
  OAI21_X1 U9932 ( .B1(n8435), .B2(n8434), .A(n7646), .ZN(n8441) );
  AOI21_X1 U9933 ( .B1(n8480), .B2(n8496), .A(n8436), .ZN(n8440) );
  AOI22_X1 U9934 ( .A1(n8482), .A2(n8498), .B1(n8481), .B2(n8437), .ZN(n8439)
         );
  NAND2_X1 U9935 ( .A1(n8455), .A2(n8866), .ZN(n8438) );
  NAND4_X1 U9936 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(
        P2_U3236) );
  INV_X1 U9937 ( .A(n8442), .ZN(n8443) );
  AOI21_X1 U9938 ( .B1(n8347), .B2(n8443), .A(n8478), .ZN(n8447) );
  NOR3_X1 U9939 ( .A1(n8464), .A2(n8445), .A3(n8444), .ZN(n8446) );
  OAI21_X1 U9940 ( .B1(n8447), .B2(n8446), .A(n8378), .ZN(n8453) );
  AOI22_X1 U9941 ( .A1(n8480), .A2(n8498), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n8452) );
  AOI22_X1 U9942 ( .A1(n8482), .A2(n8499), .B1(n8481), .B2(n8448), .ZN(n8451)
         );
  NAND2_X1 U9943 ( .A1(n8455), .A2(n8449), .ZN(n8450) );
  NAND4_X1 U9944 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(
        P2_U3238) );
  AOI22_X1 U9945 ( .A1(n8480), .A2(n9788), .B1(n8482), .B2(n8506), .ZN(n8461)
         );
  AOI22_X1 U9946 ( .A1(n8455), .A2(n4751), .B1(n8454), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8460) );
  OAI211_X1 U9947 ( .C1(n8458), .C2(n8457), .A(n8456), .B(n7054), .ZN(n8459)
         );
  NAND3_X1 U9948 ( .A1(n8461), .A2(n8460), .A3(n8459), .ZN(P2_U3239) );
  AOI21_X1 U9949 ( .B1(n8463), .B2(n8462), .A(n8478), .ZN(n8468) );
  NOR3_X1 U9950 ( .A1(n8465), .A2(n8471), .A3(n8464), .ZN(n8467) );
  OAI21_X1 U9951 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8475) );
  AND2_X1 U9952 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8530) );
  INV_X1 U9953 ( .A(n8737), .ZN(n8469) );
  OAI22_X1 U9954 ( .A1(n8472), .A2(n8471), .B1(n8470), .B2(n8469), .ZN(n8473)
         );
  AOI211_X1 U9955 ( .C1(n8480), .C2(n8743), .A(n8530), .B(n8473), .ZN(n8474)
         );
  OAI211_X1 U9956 ( .C1(n8739), .C2(n8485), .A(n8475), .B(n8474), .ZN(P2_U3240) );
  AOI211_X1 U9957 ( .C1(n8479), .C2(n8476), .A(n8478), .B(n8477), .ZN(n8488)
         );
  INV_X1 U9958 ( .A(n8810), .ZN(n8486) );
  AOI22_X1 U9959 ( .A1(n8480), .A2(n8572), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8484) );
  AOI22_X1 U9960 ( .A1(n8482), .A2(n8490), .B1(n8481), .B2(n8611), .ZN(n8483)
         );
  OAI211_X1 U9961 ( .C1(n8486), .C2(n8485), .A(n8484), .B(n8483), .ZN(n8487)
         );
  OR2_X1 U9962 ( .A1(n8488), .A2(n8487), .ZN(P2_U3242) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8489), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9964 ( .A(n8571), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8491), .Z(
        P2_U3581) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8589), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9966 ( .A(n8572), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8491), .Z(
        P2_U3579) );
  MUX2_X1 U9967 ( .A(n8624), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8491), .Z(
        P2_U3578) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8490), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9969 ( .A(n8663), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8491), .Z(
        P2_U3576) );
  MUX2_X1 U9970 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8492), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8698), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8713), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8697), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9974 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8743), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9975 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8493), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8742), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9977 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8494), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9978 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8495), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9979 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8496), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8497), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9981 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8498), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9982 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n4900), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8499), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9984 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8500), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8501), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8502), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8503), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n4402), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9989 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8504), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9788), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8505), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8506), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6403), .S(P2_U3966), .Z(
        P2_U3552) );
  XNOR2_X1 U9994 ( .A(n8529), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8511) );
  AOI211_X1 U9995 ( .C1(n8511), .C2(n8510), .A(n9778), .B(n8528), .ZN(n8522)
         );
  OAI21_X1 U9996 ( .B1(n7868), .B2(n8513), .A(n8512), .ZN(n8515) );
  XOR2_X1 U9997 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8529), .Z(n8514) );
  NAND2_X1 U9998 ( .A1(n8514), .A2(n8515), .ZN(n8523) );
  OAI211_X1 U9999 ( .C1(n8515), .C2(n8514), .A(n9774), .B(n8523), .ZN(n8519)
         );
  NOR2_X1 U10000 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8516), .ZN(n8517) );
  AOI21_X1 U10001 ( .B1(n9775), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8517), .ZN(
        n8518) );
  OAI211_X1 U10002 ( .C1(n9777), .C2(n8520), .A(n8519), .B(n8518), .ZN(n8521)
         );
  OR2_X1 U10003 ( .A1(n8522), .A2(n8521), .ZN(P2_U3262) );
  NAND2_X1 U10004 ( .A1(n8529), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10005 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  NOR2_X1 U10006 ( .A1(n8525), .A2(n8540), .ZN(n8538) );
  AOI21_X1 U10007 ( .B1(n8540), .B2(n8525), .A(n8538), .ZN(n8526) );
  INV_X1 U10008 ( .A(n8526), .ZN(n8527) );
  NOR2_X1 U10009 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8527), .ZN(n8537) );
  AOI21_X1 U10010 ( .B1(n8527), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8537), .ZN(
        n8536) );
  AOI21_X1 U10011 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8529), .A(n8528), .ZN(
        n8542) );
  INV_X1 U10012 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10095) );
  XNOR2_X1 U10013 ( .A(n8540), .B(n10095), .ZN(n8543) );
  XOR2_X1 U10014 ( .A(n8542), .B(n8543), .Z(n8532) );
  AOI21_X1 U10015 ( .B1(n9775), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8530), .ZN(
        n8531) );
  OAI21_X1 U10016 ( .B1(n9778), .B2(n8532), .A(n8531), .ZN(n8533) );
  AOI21_X1 U10017 ( .B1(n8540), .B2(n8534), .A(n8533), .ZN(n8535) );
  OAI21_X1 U10018 ( .B1(n8536), .B2(n9776), .A(n8535), .ZN(P2_U3263) );
  NOR2_X1 U10019 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  XOR2_X1 U10020 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8539), .Z(n8547) );
  NOR2_X1 U10021 ( .A1(n8540), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8541) );
  AOI21_X1 U10022 ( .B1(n8543), .B2(n8542), .A(n8541), .ZN(n8544) );
  XNOR2_X1 U10023 ( .A(n8544), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10024 ( .A1(n9773), .A2(n8546), .ZN(n8545) );
  AND2_X1 U10025 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8548) );
  AOI21_X1 U10026 ( .B1(n9775), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8548), .ZN(
        n8549) );
  NAND2_X1 U10027 ( .A1(n8556), .A2(n8555), .ZN(n8554) );
  XNOR2_X1 U10028 ( .A(n8554), .B(n8787), .ZN(n8789) );
  NAND2_X1 U10029 ( .A1(n8551), .A2(n8550), .ZN(n8792) );
  NOR2_X1 U10030 ( .A1(n9808), .A2(n8792), .ZN(n8558) );
  AOI21_X1 U10031 ( .B1(n9808), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8558), .ZN(
        n8553) );
  NAND2_X1 U10032 ( .A1(n8787), .A2(n8598), .ZN(n8552) );
  OAI211_X1 U10033 ( .C1(n8789), .C2(n8560), .A(n8553), .B(n8552), .ZN(
        P2_U3265) );
  OAI21_X1 U10034 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8793) );
  NOR2_X1 U10035 ( .A1(n8556), .A2(n8781), .ZN(n8557) );
  AOI211_X1 U10036 ( .C1(n9808), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8558), .B(
        n8557), .ZN(n8559) );
  OAI21_X1 U10037 ( .B1(n8560), .B2(n8793), .A(n8559), .ZN(P2_U3266) );
  OAI21_X1 U10038 ( .B1(n8561), .B2(n8569), .A(n8562), .ZN(n8563) );
  INV_X1 U10039 ( .A(n8563), .ZN(n8803) );
  INV_X1 U10040 ( .A(n8564), .ZN(n8565) );
  AOI21_X1 U10041 ( .B1(n8799), .B2(n8578), .A(n8565), .ZN(n8800) );
  AOI22_X1 U10042 ( .A1(n9808), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8566), .B2(
        n8778), .ZN(n8567) );
  OAI21_X1 U10043 ( .B1(n8568), .B2(n8781), .A(n8567), .ZN(n8573) );
  OAI21_X1 U10044 ( .B1(n8803), .B2(n8748), .A(n8574), .ZN(P2_U3268) );
  OAI21_X1 U10045 ( .B1(n8575), .B2(n8587), .A(n8576), .ZN(n8577) );
  INV_X1 U10046 ( .A(n8577), .ZN(n8808) );
  INV_X1 U10047 ( .A(n8610), .ZN(n8580) );
  INV_X1 U10048 ( .A(n8578), .ZN(n8579) );
  AOI21_X1 U10049 ( .B1(n8804), .B2(n8580), .A(n8579), .ZN(n8805) );
  INV_X1 U10050 ( .A(n8581), .ZN(n8582) );
  AOI22_X1 U10051 ( .A1(n9808), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8582), .B2(
        n8778), .ZN(n8583) );
  OAI21_X1 U10052 ( .B1(n8584), .B2(n8781), .A(n8583), .ZN(n8592) );
  INV_X1 U10053 ( .A(n8585), .ZN(n8586) );
  NOR2_X1 U10054 ( .A1(n8602), .A2(n8586), .ZN(n8588) );
  XNOR2_X1 U10055 ( .A(n8588), .B(n8587), .ZN(n8590) );
  AOI222_X1 U10056 ( .A1(n9790), .A2(n8590), .B1(n8624), .B2(n9787), .C1(n8589), .C2(n9785), .ZN(n8807) );
  NOR2_X1 U10057 ( .A1(n8807), .A2(n9808), .ZN(n8591) );
  AOI211_X1 U10058 ( .C1(n8805), .C2(n9521), .A(n8592), .B(n8591), .ZN(n8593)
         );
  OAI21_X1 U10059 ( .B1(n8808), .B2(n8748), .A(n8593), .ZN(P2_U3269) );
  OR2_X1 U10060 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  NAND2_X1 U10061 ( .A1(n8594), .A2(n8597), .ZN(n8809) );
  INV_X1 U10062 ( .A(n8809), .ZN(n8616) );
  AOI22_X1 U10063 ( .A1(n8810), .A2(n8598), .B1(n9808), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8615) );
  NOR2_X1 U10064 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  OR2_X1 U10065 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  NAND2_X1 U10066 ( .A1(n8603), .A2(n9790), .ZN(n8607) );
  OAI22_X1 U10067 ( .A1(n8604), .A2(n9535), .B1(n8645), .B2(n9533), .ZN(n8605)
         );
  INV_X1 U10068 ( .A(n8605), .ZN(n8606) );
  NAND2_X1 U10069 ( .A1(n8607), .A2(n8606), .ZN(n8814) );
  NAND2_X1 U10070 ( .A1(n8810), .A2(n8620), .ZN(n8608) );
  NAND2_X1 U10071 ( .A1(n8608), .A2(n9883), .ZN(n8609) );
  OR2_X1 U10072 ( .A1(n8610), .A2(n8609), .ZN(n8812) );
  INV_X1 U10073 ( .A(n8611), .ZN(n8612) );
  OAI22_X1 U10074 ( .A1(n8812), .A2(n4625), .B1(n9793), .B2(n8612), .ZN(n8613)
         );
  OAI21_X1 U10075 ( .B1(n8814), .B2(n8613), .A(n9791), .ZN(n8614) );
  OAI211_X1 U10076 ( .C1(n8616), .C2(n8748), .A(n8615), .B(n8614), .ZN(
        P2_U3270) );
  OAI21_X1 U10077 ( .B1(n8618), .B2(n8622), .A(n8617), .ZN(n8619) );
  INV_X1 U10078 ( .A(n8619), .ZN(n8821) );
  INV_X1 U10079 ( .A(n8620), .ZN(n8621) );
  AOI211_X1 U10080 ( .C1(n8818), .C2(n8635), .A(n9900), .B(n8621), .ZN(n8817)
         );
  INV_X1 U10081 ( .A(n8817), .ZN(n8626) );
  XNOR2_X1 U10082 ( .A(n8623), .B(n8622), .ZN(n8625) );
  AOI222_X1 U10083 ( .A1(n9790), .A2(n8625), .B1(n8624), .B2(n9785), .C1(n8663), .C2(n9787), .ZN(n8820) );
  OAI21_X1 U10084 ( .B1(n4625), .B2(n8626), .A(n8820), .ZN(n8631) );
  INV_X1 U10085 ( .A(n8818), .ZN(n8629) );
  AOI22_X1 U10086 ( .A1(n9808), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8627), .B2(
        n8778), .ZN(n8628) );
  OAI21_X1 U10087 ( .B1(n8629), .B2(n8781), .A(n8628), .ZN(n8630) );
  AOI21_X1 U10088 ( .B1(n8631), .B2(n9791), .A(n8630), .ZN(n8632) );
  OAI21_X1 U10089 ( .B1(n8821), .B2(n8748), .A(n8632), .ZN(P2_U3271) );
  XNOR2_X1 U10090 ( .A(n8634), .B(n8633), .ZN(n8826) );
  INV_X1 U10091 ( .A(n8654), .ZN(n8637) );
  INV_X1 U10092 ( .A(n8635), .ZN(n8636) );
  AOI21_X1 U10093 ( .B1(n8822), .B2(n8637), .A(n8636), .ZN(n8823) );
  INV_X1 U10094 ( .A(n8638), .ZN(n8639) );
  AOI22_X1 U10095 ( .A1(n9808), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8639), .B2(
        n8778), .ZN(n8640) );
  OAI21_X1 U10096 ( .B1(n8641), .B2(n8781), .A(n8640), .ZN(n8650) );
  AOI21_X1 U10097 ( .B1(n8661), .B2(n8643), .A(n8642), .ZN(n8644) );
  NOR2_X1 U10098 ( .A1(n8644), .A2(n9531), .ZN(n8648) );
  OAI22_X1 U10099 ( .A1(n8645), .A2(n9535), .B1(n8681), .B2(n9533), .ZN(n8646)
         );
  AOI21_X1 U10100 ( .B1(n8648), .B2(n8647), .A(n8646), .ZN(n8825) );
  NOR2_X1 U10101 ( .A1(n8825), .A2(n9808), .ZN(n8649) );
  AOI211_X1 U10102 ( .C1(n8823), .C2(n9521), .A(n8650), .B(n8649), .ZN(n8651)
         );
  OAI21_X1 U10103 ( .B1(n8826), .B2(n8748), .A(n8651), .ZN(P2_U3272) );
  OAI21_X1 U10104 ( .B1(n8653), .B2(n8659), .A(n8652), .ZN(n8831) );
  AOI21_X1 U10105 ( .B1(n8827), .B2(n8670), .A(n8654), .ZN(n8828) );
  INV_X1 U10106 ( .A(n8827), .ZN(n8658) );
  INV_X1 U10107 ( .A(n8655), .ZN(n8656) );
  AOI22_X1 U10108 ( .A1(n9808), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8656), .B2(
        n8778), .ZN(n8657) );
  OAI21_X1 U10109 ( .B1(n8658), .B2(n8781), .A(n8657), .ZN(n8666) );
  OAI21_X1 U10110 ( .B1(n4428), .B2(n8660), .A(n8659), .ZN(n8662) );
  NAND2_X1 U10111 ( .A1(n8662), .A2(n8661), .ZN(n8664) );
  AOI222_X1 U10112 ( .A1(n9790), .A2(n8664), .B1(n8698), .B2(n9787), .C1(n8663), .C2(n9785), .ZN(n8830) );
  NOR2_X1 U10113 ( .A1(n8830), .A2(n9808), .ZN(n8665) );
  AOI211_X1 U10114 ( .C1(n8828), .C2(n9521), .A(n8666), .B(n8665), .ZN(n8667)
         );
  OAI21_X1 U10115 ( .B1(n8748), .B2(n8831), .A(n8667), .ZN(P2_U3273) );
  XNOR2_X1 U10116 ( .A(n8668), .B(n8669), .ZN(n8836) );
  INV_X1 U10117 ( .A(n8670), .ZN(n8671) );
  AOI21_X1 U10118 ( .B1(n8832), .B2(n8688), .A(n8671), .ZN(n8833) );
  INV_X1 U10119 ( .A(n8832), .ZN(n8675) );
  INV_X1 U10120 ( .A(n8672), .ZN(n8673) );
  AOI22_X1 U10121 ( .A1(n9808), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8673), .B2(
        n8778), .ZN(n8674) );
  OAI21_X1 U10122 ( .B1(n8675), .B2(n8781), .A(n8674), .ZN(n8685) );
  INV_X1 U10123 ( .A(n8676), .ZN(n8678) );
  AOI21_X1 U10124 ( .B1(n8696), .B2(n8678), .A(n8677), .ZN(n8679) );
  NOR3_X1 U10125 ( .A1(n4428), .A2(n8679), .A3(n9531), .ZN(n8683) );
  OAI22_X1 U10126 ( .A1(n8681), .A2(n9535), .B1(n8680), .B2(n9533), .ZN(n8682)
         );
  NOR2_X1 U10127 ( .A1(n8683), .A2(n8682), .ZN(n8835) );
  NOR2_X1 U10128 ( .A1(n8835), .A2(n9808), .ZN(n8684) );
  AOI211_X1 U10129 ( .C1(n8833), .C2(n9521), .A(n8685), .B(n8684), .ZN(n8686)
         );
  OAI21_X1 U10130 ( .B1(n8748), .B2(n8836), .A(n8686), .ZN(P2_U3274) );
  XNOR2_X1 U10131 ( .A(n8687), .B(n8695), .ZN(n8841) );
  INV_X1 U10132 ( .A(n8705), .ZN(n8690) );
  INV_X1 U10133 ( .A(n8688), .ZN(n8689) );
  AOI21_X1 U10134 ( .B1(n8837), .B2(n8690), .A(n8689), .ZN(n8838) );
  INV_X1 U10135 ( .A(n8691), .ZN(n8692) );
  AOI22_X1 U10136 ( .A1(n9808), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8692), .B2(
        n8778), .ZN(n8693) );
  OAI21_X1 U10137 ( .B1(n8694), .B2(n8781), .A(n8693), .ZN(n8701) );
  OAI21_X1 U10138 ( .B1(n4998), .B2(n6030), .A(n8696), .ZN(n8699) );
  AOI222_X1 U10139 ( .A1(n9790), .A2(n8699), .B1(n8698), .B2(n9785), .C1(n8697), .C2(n9787), .ZN(n8840) );
  NOR2_X1 U10140 ( .A1(n8840), .A2(n9808), .ZN(n8700) );
  AOI211_X1 U10141 ( .C1(n8838), .C2(n9521), .A(n8701), .B(n8700), .ZN(n8702)
         );
  OAI21_X1 U10142 ( .B1(n8841), .B2(n8748), .A(n8702), .ZN(P2_U3275) );
  OAI21_X1 U10143 ( .B1(n8704), .B2(n8712), .A(n8703), .ZN(n8846) );
  AOI21_X1 U10144 ( .B1(n8842), .B2(n8718), .A(n8705), .ZN(n8843) );
  INV_X1 U10145 ( .A(n8842), .ZN(n8709) );
  INV_X1 U10146 ( .A(n8706), .ZN(n8707) );
  AOI22_X1 U10147 ( .A1(n9808), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8707), .B2(
        n8778), .ZN(n8708) );
  OAI21_X1 U10148 ( .B1(n8709), .B2(n8781), .A(n8708), .ZN(n8716) );
  NAND2_X1 U10149 ( .A1(n8719), .A2(n8710), .ZN(n8711) );
  XOR2_X1 U10150 ( .A(n8712), .B(n8711), .Z(n8714) );
  AOI222_X1 U10151 ( .A1(n9790), .A2(n8714), .B1(n8713), .B2(n9785), .C1(n8743), .C2(n9787), .ZN(n8845) );
  NOR2_X1 U10152 ( .A1(n8845), .A2(n9808), .ZN(n8715) );
  AOI211_X1 U10153 ( .C1(n8843), .C2(n9521), .A(n8716), .B(n8715), .ZN(n8717)
         );
  OAI21_X1 U10154 ( .B1(n8748), .B2(n8846), .A(n8717), .ZN(P2_U3276) );
  AOI211_X1 U10155 ( .C1(n8849), .C2(n8736), .A(n9900), .B(n4808), .ZN(n8848)
         );
  INV_X1 U10156 ( .A(n8719), .ZN(n8720) );
  AOI21_X1 U10157 ( .B1(n4771), .B2(n8721), .A(n8720), .ZN(n8723) );
  OAI21_X1 U10158 ( .B1(n8723), .B2(n9531), .A(n8722), .ZN(n8847) );
  OAI21_X1 U10159 ( .B1(n8725), .B2(n4771), .A(n8724), .ZN(n8851) );
  NOR2_X1 U10160 ( .A1(n8851), .A2(n8774), .ZN(n8726) );
  AOI211_X1 U10161 ( .C1(n8848), .C2(n4410), .A(n8847), .B(n8726), .ZN(n8734)
         );
  INV_X1 U10162 ( .A(n8851), .ZN(n8732) );
  AOI22_X1 U10163 ( .A1(n9808), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8728), .B2(
        n8778), .ZN(n8729) );
  OAI21_X1 U10164 ( .B1(n8730), .B2(n8781), .A(n8729), .ZN(n8731) );
  AOI21_X1 U10165 ( .B1(n8732), .B2(n8767), .A(n8731), .ZN(n8733) );
  OAI21_X1 U10166 ( .B1(n8734), .B2(n9808), .A(n8733), .ZN(P2_U3277) );
  XNOR2_X1 U10167 ( .A(n8735), .B(n8740), .ZN(n8856) );
  AOI21_X1 U10168 ( .B1(n8852), .B2(n4425), .A(n4809), .ZN(n8853) );
  AOI22_X1 U10169 ( .A1(n9808), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8737), .B2(
        n8778), .ZN(n8738) );
  OAI21_X1 U10170 ( .B1(n8739), .B2(n8781), .A(n8738), .ZN(n8746) );
  XOR2_X1 U10171 ( .A(n8741), .B(n8740), .Z(n8744) );
  AOI222_X1 U10172 ( .A1(n9790), .A2(n8744), .B1(n8743), .B2(n9785), .C1(n8742), .C2(n9787), .ZN(n8855) );
  NOR2_X1 U10173 ( .A1(n8855), .A2(n9808), .ZN(n8745) );
  AOI211_X1 U10174 ( .C1(n8853), .C2(n9521), .A(n8746), .B(n8745), .ZN(n8747)
         );
  OAI21_X1 U10175 ( .B1(n8856), .B2(n8748), .A(n8747), .ZN(P2_U3278) );
  OAI21_X1 U10176 ( .B1(n8749), .B2(n8753), .A(n8750), .ZN(n8857) );
  AOI22_X1 U10177 ( .A1(n9808), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8751), .B2(
        n8778), .ZN(n8752) );
  OAI21_X1 U10178 ( .B1(n8860), .B2(n8781), .A(n8752), .ZN(n8766) );
  AOI21_X1 U10179 ( .B1(n8754), .B2(n8753), .A(n9531), .ZN(n8758) );
  OAI22_X1 U10180 ( .A1(n8755), .A2(n9535), .B1(n9534), .B2(n9533), .ZN(n8756)
         );
  AOI21_X1 U10181 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8764) );
  OAI211_X1 U10182 ( .C1(n8860), .C2(n8759), .A(n4425), .B(n9883), .ZN(n8760)
         );
  INV_X1 U10183 ( .A(n8858), .ZN(n8761) );
  AOI21_X1 U10184 ( .B1(n8857), .B2(n8762), .A(n8761), .ZN(n8763) );
  AOI211_X1 U10185 ( .C1(n8767), .C2(n8857), .A(n8766), .B(n8765), .ZN(n8768)
         );
  INV_X1 U10186 ( .A(n8768), .ZN(P2_U3279) );
  XNOR2_X1 U10187 ( .A(n8769), .B(n8772), .ZN(n8777) );
  INV_X1 U10188 ( .A(n8770), .ZN(n8773) );
  OAI21_X1 U10189 ( .B1(n8773), .B2(n8772), .A(n4543), .ZN(n8865) );
  NOR2_X1 U10190 ( .A1(n8865), .A2(n8774), .ZN(n8775) );
  AOI211_X1 U10191 ( .C1(n9790), .C2(n8777), .A(n8776), .B(n8775), .ZN(n8864)
         );
  XOR2_X1 U10192 ( .A(n9519), .B(n8861), .Z(n8862) );
  INV_X1 U10193 ( .A(n8861), .ZN(n8782) );
  AOI22_X1 U10194 ( .A1(n9808), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8779), .B2(
        n8778), .ZN(n8780) );
  OAI21_X1 U10195 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8785) );
  NOR2_X1 U10196 ( .A1(n8865), .A2(n8783), .ZN(n8784) );
  AOI211_X1 U10197 ( .C1(n8862), .C2(n9521), .A(n8785), .B(n8784), .ZN(n8786)
         );
  OAI21_X1 U10198 ( .B1(n8864), .B2(n9808), .A(n8786), .ZN(P2_U3280) );
  NAND2_X1 U10199 ( .A1(n8787), .A2(n9882), .ZN(n8788) );
  OAI211_X1 U10200 ( .C1(n8789), .C2(n9900), .A(n8792), .B(n8788), .ZN(n8871)
         );
  MUX2_X1 U10201 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8871), .S(n9924), .Z(
        P2_U3551) );
  NAND2_X1 U10202 ( .A1(n8790), .A2(n9882), .ZN(n8791) );
  OAI211_X1 U10203 ( .C1(n8793), .C2(n9900), .A(n8792), .B(n8791), .ZN(n8872)
         );
  MUX2_X1 U10204 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8872), .S(n9924), .Z(
        P2_U3550) );
  AOI22_X1 U10205 ( .A1(n8795), .A2(n9883), .B1(n9882), .B2(n8794), .ZN(n8796)
         );
  AOI22_X1 U10206 ( .A1(n8800), .A2(n9883), .B1(n9882), .B2(n8799), .ZN(n8801)
         );
  OAI211_X1 U10207 ( .C1(n8803), .C2(n9871), .A(n8802), .B(n8801), .ZN(n8874)
         );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8874), .S(n9924), .Z(
        P2_U3548) );
  AOI22_X1 U10209 ( .A1(n8805), .A2(n9883), .B1(n9882), .B2(n8804), .ZN(n8806)
         );
  OAI211_X1 U10210 ( .C1(n8808), .C2(n9871), .A(n8807), .B(n8806), .ZN(n8875)
         );
  MUX2_X1 U10211 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8875), .S(n9924), .Z(
        P2_U3547) );
  NAND2_X1 U10212 ( .A1(n8809), .A2(n9904), .ZN(n8816) );
  NAND2_X1 U10213 ( .A1(n8810), .A2(n9882), .ZN(n8811) );
  NAND2_X1 U10214 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NOR2_X1 U10215 ( .A1(n8814), .A2(n8813), .ZN(n8815) );
  NAND2_X1 U10216 ( .A1(n8816), .A2(n8815), .ZN(n8876) );
  MUX2_X1 U10217 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8876), .S(n9924), .Z(
        P2_U3546) );
  AOI21_X1 U10218 ( .B1(n9882), .B2(n8818), .A(n8817), .ZN(n8819) );
  OAI211_X1 U10219 ( .C1(n8821), .C2(n9871), .A(n8820), .B(n8819), .ZN(n8877)
         );
  MUX2_X1 U10220 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8877), .S(n9924), .Z(
        P2_U3545) );
  AOI22_X1 U10221 ( .A1(n8823), .A2(n9883), .B1(n9882), .B2(n8822), .ZN(n8824)
         );
  OAI211_X1 U10222 ( .C1(n8826), .C2(n9871), .A(n8825), .B(n8824), .ZN(n8878)
         );
  MUX2_X1 U10223 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8878), .S(n9924), .Z(
        P2_U3544) );
  AOI22_X1 U10224 ( .A1(n8828), .A2(n9883), .B1(n9882), .B2(n8827), .ZN(n8829)
         );
  OAI211_X1 U10225 ( .C1(n8831), .C2(n9871), .A(n8830), .B(n8829), .ZN(n8879)
         );
  MUX2_X1 U10226 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8879), .S(n9924), .Z(
        P2_U3543) );
  AOI22_X1 U10227 ( .A1(n8833), .A2(n9883), .B1(n9882), .B2(n8832), .ZN(n8834)
         );
  OAI211_X1 U10228 ( .C1(n8836), .C2(n9871), .A(n8835), .B(n8834), .ZN(n8880)
         );
  MUX2_X1 U10229 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8880), .S(n9924), .Z(
        P2_U3542) );
  AOI22_X1 U10230 ( .A1(n8838), .A2(n9883), .B1(n9882), .B2(n8837), .ZN(n8839)
         );
  OAI211_X1 U10231 ( .C1(n8841), .C2(n9871), .A(n8840), .B(n8839), .ZN(n8881)
         );
  MUX2_X1 U10232 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8881), .S(n9924), .Z(
        P2_U3541) );
  AOI22_X1 U10233 ( .A1(n8843), .A2(n9883), .B1(n9882), .B2(n8842), .ZN(n8844)
         );
  OAI211_X1 U10234 ( .C1(n8846), .C2(n9871), .A(n8845), .B(n8844), .ZN(n8882)
         );
  MUX2_X1 U10235 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8882), .S(n9924), .Z(
        P2_U3540) );
  AOI211_X1 U10236 ( .C1(n9882), .C2(n8849), .A(n8848), .B(n8847), .ZN(n8850)
         );
  OAI21_X1 U10237 ( .B1(n9871), .B2(n8851), .A(n8850), .ZN(n8883) );
  MUX2_X1 U10238 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8883), .S(n9924), .Z(
        P2_U3539) );
  AOI22_X1 U10239 ( .A1(n8853), .A2(n9883), .B1(n9882), .B2(n8852), .ZN(n8854)
         );
  OAI211_X1 U10240 ( .C1(n8856), .C2(n9871), .A(n8855), .B(n8854), .ZN(n8884)
         );
  MUX2_X1 U10241 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8884), .S(n9924), .Z(
        P2_U3538) );
  NAND2_X1 U10242 ( .A1(n8857), .A2(n9904), .ZN(n8859) );
  OAI211_X1 U10243 ( .C1(n8860), .C2(n9899), .A(n8859), .B(n8858), .ZN(n8885)
         );
  MUX2_X1 U10244 ( .A(n8885), .B(P2_REG1_REG_17__SCAN_IN), .S(n9922), .Z(
        P2_U3537) );
  AOI22_X1 U10245 ( .A1(n8862), .A2(n9883), .B1(n9882), .B2(n8861), .ZN(n8863)
         );
  OAI211_X1 U10246 ( .C1(n9890), .C2(n8865), .A(n8864), .B(n8863), .ZN(n8886)
         );
  MUX2_X1 U10247 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8886), .S(n9924), .Z(
        P2_U3536) );
  AOI22_X1 U10248 ( .A1(n8867), .A2(n9883), .B1(n9882), .B2(n8866), .ZN(n8868)
         );
  OAI211_X1 U10249 ( .C1(n9890), .C2(n8870), .A(n8869), .B(n8868), .ZN(n8887)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8887), .S(n9924), .Z(
        P2_U3533) );
  MUX2_X1 U10251 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8871), .S(n9908), .Z(
        P2_U3519) );
  MUX2_X1 U10252 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8872), .S(n9908), .Z(
        P2_U3518) );
  MUX2_X1 U10253 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8874), .S(n9908), .Z(
        P2_U3516) );
  MUX2_X1 U10254 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8875), .S(n9908), .Z(
        P2_U3515) );
  MUX2_X1 U10255 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8876), .S(n9908), .Z(
        P2_U3514) );
  MUX2_X1 U10256 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8877), .S(n9908), .Z(
        P2_U3513) );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8878), .S(n9908), .Z(
        P2_U3512) );
  MUX2_X1 U10258 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8879), .S(n9908), .Z(
        P2_U3511) );
  MUX2_X1 U10259 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8880), .S(n9908), .Z(
        P2_U3510) );
  MUX2_X1 U10260 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8881), .S(n9908), .Z(
        P2_U3509) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8882), .S(n9908), .Z(
        P2_U3508) );
  MUX2_X1 U10262 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8883), .S(n9908), .Z(
        P2_U3507) );
  MUX2_X1 U10263 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8884), .S(n9908), .Z(
        P2_U3505) );
  MUX2_X1 U10264 ( .A(n8885), .B(P2_REG0_REG_17__SCAN_IN), .S(n9906), .Z(
        P2_U3502) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8886), .S(n9908), .Z(
        P2_U3499) );
  MUX2_X1 U10266 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8887), .S(n9908), .Z(
        P2_U3490) );
  INV_X1 U10267 ( .A(n8888), .ZN(n9476) );
  INV_X1 U10268 ( .A(n8889), .ZN(n8890) );
  NOR4_X1 U10269 ( .A1(n8890), .A2(P2_IR_REG_30__SCAN_IN), .A3(n10207), .A4(
        P2_U3152), .ZN(n8891) );
  AOI21_X1 U10270 ( .B1(n8892), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8891), .ZN(
        n8893) );
  OAI21_X1 U10271 ( .B1(n9476), .B2(n8894), .A(n8893), .ZN(P2_U3327) );
  MUX2_X1 U10272 ( .A(n8895), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10273 ( .A(n8898), .B(n8897), .ZN(n8899) );
  XNOR2_X1 U10274 ( .A(n8896), .B(n8899), .ZN(n8900) );
  NAND2_X1 U10275 ( .A1(n8900), .A2(n9016), .ZN(n8908) );
  AOI21_X1 U10276 ( .B1(n9500), .B2(n9049), .A(n8901), .ZN(n8907) );
  OAI22_X1 U10277 ( .A1(n8902), .A2(n9503), .B1(n9020), .B2(n9736), .ZN(n8903)
         );
  INV_X1 U10278 ( .A(n8903), .ZN(n8906) );
  OR2_X1 U10279 ( .A1(n9517), .A2(n8904), .ZN(n8905) );
  NAND4_X1 U10280 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(
        P1_U3211) );
  NAND2_X1 U10281 ( .A1(n8970), .A2(n8909), .ZN(n8910) );
  XOR2_X1 U10282 ( .A(n8911), .B(n8910), .Z(n8916) );
  OAI22_X1 U10283 ( .A1(n9273), .A2(n9003), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10099), .ZN(n8912) );
  AOI21_X1 U10284 ( .B1(n9005), .B2(n9300), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10285 ( .B1(n9517), .B2(n9275), .A(n8913), .ZN(n8914) );
  AOI21_X1 U10286 ( .B1(n9412), .B2(n9038), .A(n8914), .ZN(n8915) );
  OAI21_X1 U10287 ( .B1(n8916), .B2(n9509), .A(n8915), .ZN(P1_U3214) );
  XOR2_X1 U10288 ( .A(n8919), .B(n8918), .Z(n8920) );
  XNOR2_X1 U10289 ( .A(n8917), .B(n8920), .ZN(n8925) );
  NAND2_X1 U10290 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9120) );
  OAI21_X1 U10291 ( .B1(n9003), .B2(n9336), .A(n9120), .ZN(n8921) );
  AOI21_X1 U10292 ( .B1(n9005), .B2(n9365), .A(n8921), .ZN(n8922) );
  OAI21_X1 U10293 ( .B1(n9517), .B2(n9341), .A(n8922), .ZN(n8923) );
  AOI21_X1 U10294 ( .B1(n9434), .B2(n9038), .A(n8923), .ZN(n8924) );
  OAI21_X1 U10295 ( .B1(n8925), .B2(n9509), .A(n8924), .ZN(P1_U3217) );
  INV_X1 U10296 ( .A(n9422), .ZN(n9123) );
  OR2_X1 U10297 ( .A1(n8926), .A2(n8982), .ZN(n8980) );
  NAND2_X1 U10298 ( .A1(n8980), .A2(n8927), .ZN(n8931) );
  AND2_X1 U10299 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  OAI21_X1 U10300 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8933) );
  NAND2_X1 U10301 ( .A1(n8933), .A2(n9016), .ZN(n8938) );
  AOI22_X1 U10302 ( .A1(n9005), .A2(n9299), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8934) );
  OAI21_X1 U10303 ( .B1(n9272), .B2(n9003), .A(n8934), .ZN(n8935) );
  AOI21_X1 U10304 ( .B1(n9304), .B2(n8936), .A(n8935), .ZN(n8937) );
  OAI211_X1 U10305 ( .C1(n9123), .C2(n9020), .A(n8938), .B(n8937), .ZN(
        P1_U3221) );
  INV_X1 U10306 ( .A(n9400), .ZN(n9241) );
  OAI21_X1 U10307 ( .B1(n8940), .B2(n8939), .A(n5703), .ZN(n8941) );
  NAND2_X1 U10308 ( .A1(n8941), .A2(n9016), .ZN(n8946) );
  NOR2_X1 U10309 ( .A1(n9238), .A2(n9517), .ZN(n8944) );
  OAI22_X1 U10310 ( .A1(n9213), .A2(n9003), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8942), .ZN(n8943) );
  AOI211_X1 U10311 ( .C1(n9005), .C2(n9245), .A(n8944), .B(n8943), .ZN(n8945)
         );
  OAI211_X1 U10312 ( .C1(n9241), .C2(n9020), .A(n8946), .B(n8945), .ZN(
        P1_U3223) );
  OR2_X1 U10313 ( .A1(n8947), .A2(n8948), .ZN(n8961) );
  INV_X1 U10314 ( .A(n8961), .ZN(n8951) );
  INV_X1 U10315 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U10316 ( .A1(n8949), .A2(n8960), .ZN(n8950) );
  AOI22_X1 U10317 ( .A1(n8951), .A2(n8960), .B1(n8947), .B2(n8950), .ZN(n8959)
         );
  NOR2_X1 U10318 ( .A1(n9503), .A2(n8952), .ZN(n8953) );
  AOI211_X1 U10319 ( .C1(n9500), .C2(n9042), .A(n8954), .B(n8953), .ZN(n8955)
         );
  OAI21_X1 U10320 ( .B1(n9517), .B2(n8956), .A(n8955), .ZN(n8957) );
  AOI21_X1 U10321 ( .B1(n7905), .B2(n9038), .A(n8957), .ZN(n8958) );
  OAI21_X1 U10322 ( .B1(n8959), .B2(n9509), .A(n8958), .ZN(P1_U3224) );
  INV_X1 U10323 ( .A(n9442), .ZN(n9360) );
  NAND2_X1 U10324 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  OAI21_X1 U10325 ( .B1(n8963), .B2(n8962), .A(n4376), .ZN(n8964) );
  NAND2_X1 U10326 ( .A1(n8964), .A2(n9016), .ZN(n8968) );
  NOR2_X1 U10327 ( .A1(n9517), .A2(n9356), .ZN(n8966) );
  NAND2_X1 U10328 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9084) );
  OAI21_X1 U10329 ( .B1(n9003), .B2(n9335), .A(n9084), .ZN(n8965) );
  AOI211_X1 U10330 ( .C1(n9005), .C2(n9364), .A(n8966), .B(n8965), .ZN(n8967)
         );
  OAI211_X1 U10331 ( .C1(n9360), .C2(n9020), .A(n8968), .B(n8967), .ZN(
        P1_U3226) );
  NAND2_X1 U10332 ( .A1(n8970), .A2(n8969), .ZN(n8974) );
  AND2_X1 U10333 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  AOI21_X1 U10334 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8979) );
  AOI22_X1 U10335 ( .A1(n9262), .A2(n9500), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8976) );
  NAND2_X1 U10336 ( .A1(n9261), .A2(n9005), .ZN(n8975) );
  OAI211_X1 U10337 ( .C1(n9517), .C2(n9254), .A(n8976), .B(n8975), .ZN(n8977)
         );
  AOI21_X1 U10338 ( .B1(n9406), .B2(n9038), .A(n8977), .ZN(n8978) );
  OAI21_X1 U10339 ( .B1(n8979), .B2(n9509), .A(n8978), .ZN(P1_U3227) );
  INV_X1 U10340 ( .A(n8980), .ZN(n8981) );
  AOI21_X1 U10341 ( .B1(n8982), .B2(n8926), .A(n8981), .ZN(n8988) );
  OAI22_X1 U10342 ( .A1(n9003), .A2(n9293), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8983), .ZN(n8984) );
  AOI21_X1 U10343 ( .B1(n9005), .B2(n9322), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10344 ( .B1(n9517), .B2(n9316), .A(n8985), .ZN(n8986) );
  AOI21_X1 U10345 ( .B1(n9427), .B2(n9038), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10346 ( .B1(n8988), .B2(n9509), .A(n8987), .ZN(P1_U3231) );
  NAND2_X1 U10347 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  XOR2_X1 U10348 ( .A(n8992), .B(n8991), .Z(n8997) );
  AOI22_X1 U10349 ( .A1(n9005), .A2(n9323), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8994) );
  NAND2_X1 U10350 ( .A1(n9261), .A2(n9500), .ZN(n8993) );
  OAI211_X1 U10351 ( .C1(n9517), .C2(n9286), .A(n8994), .B(n8993), .ZN(n8995)
         );
  AOI21_X1 U10352 ( .B1(n9417), .B2(n9038), .A(n8995), .ZN(n8996) );
  OAI21_X1 U10353 ( .B1(n8997), .B2(n9509), .A(n8996), .ZN(P1_U3233) );
  XNOR2_X1 U10354 ( .A(n9000), .B(n8999), .ZN(n9001) );
  XNOR2_X1 U10355 ( .A(n8998), .B(n9001), .ZN(n9010) );
  NAND2_X1 U10356 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9094) );
  OAI21_X1 U10357 ( .B1(n9003), .B2(n9002), .A(n9094), .ZN(n9004) );
  AOI21_X1 U10358 ( .B1(n9005), .B2(n9042), .A(n9004), .ZN(n9006) );
  OAI21_X1 U10359 ( .B1(n9517), .B2(n9007), .A(n9006), .ZN(n9008) );
  AOI21_X1 U10360 ( .B1(n9437), .B2(n9038), .A(n9008), .ZN(n9009) );
  OAI21_X1 U10361 ( .B1(n9010), .B2(n9509), .A(n9009), .ZN(P1_U3236) );
  INV_X1 U10362 ( .A(n9012), .ZN(n9014) );
  NOR2_X1 U10363 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  XNOR2_X1 U10364 ( .A(n9011), .B(n9015), .ZN(n9017) );
  NAND2_X1 U10365 ( .A1(n9017), .A2(n9016), .ZN(n9027) );
  AOI21_X1 U10366 ( .B1(n9500), .B2(n9050), .A(n9018), .ZN(n9026) );
  OAI22_X1 U10367 ( .A1(n9021), .A2(n9503), .B1(n9020), .B2(n9019), .ZN(n9022)
         );
  INV_X1 U10368 ( .A(n9022), .ZN(n9025) );
  OR2_X1 U10369 ( .A1(n9517), .A2(n9023), .ZN(n9024) );
  NAND4_X1 U10370 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(
        P1_U3237) );
  NAND2_X1 U10371 ( .A1(n4476), .A2(n9028), .ZN(n9030) );
  XNOR2_X1 U10372 ( .A(n9030), .B(n9029), .ZN(n9040) );
  INV_X1 U10373 ( .A(n9031), .ZN(n9034) );
  NOR2_X1 U10374 ( .A1(n9503), .A2(n9032), .ZN(n9033) );
  AOI211_X1 U10375 ( .C1(n9500), .C2(n9364), .A(n9034), .B(n9033), .ZN(n9035)
         );
  OAI21_X1 U10376 ( .B1(n9517), .B2(n9036), .A(n9035), .ZN(n9037) );
  AOI21_X1 U10377 ( .B1(n9453), .B2(n9038), .A(n9037), .ZN(n9039) );
  OAI21_X1 U10378 ( .B1(n9040), .B2(n9509), .A(n9039), .ZN(P1_U3239) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9041), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9210), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9147), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9246), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9262), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9245), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9261), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9300), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9323), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9299), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9322), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9365), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9042), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9364), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9043), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9044), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9499), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9045), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9046), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9047), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9048), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9049), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9050), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9665), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9051), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9052), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9053), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9054), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9055), .S(P1_U4006), .Z(
        P1_U3556) );
  OAI211_X1 U10408 ( .C1(n9605), .C2(n9056), .A(n9593), .B(n9589), .ZN(n9064)
         );
  NAND2_X1 U10409 ( .A1(n9656), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n9063) );
  AOI22_X1 U10410 ( .A1(n9654), .A2(n9057), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9062) );
  OAI211_X1 U10411 ( .C1(n9060), .C2(n9059), .A(n9653), .B(n9058), .ZN(n9061)
         );
  NAND4_X1 U10412 ( .A1(n9064), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(
        P1_U3242) );
  OAI211_X1 U10413 ( .C1(n9067), .C2(n9066), .A(n9593), .B(n9065), .ZN(n9075)
         );
  NAND2_X1 U10414 ( .A1(n9656), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9074) );
  AOI22_X1 U10415 ( .A1(n9654), .A2(n9068), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n9073) );
  OAI211_X1 U10416 ( .C1(n9071), .C2(n9070), .A(n9653), .B(n9069), .ZN(n9072)
         );
  NAND4_X1 U10417 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(
        P1_U3244) );
  INV_X1 U10418 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9090) );
  AOI21_X1 U10419 ( .B1(n9080), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9076), .ZN(
        n9078) );
  XNOR2_X1 U10420 ( .A(n9098), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U10421 ( .A1(n9078), .A2(n9077), .ZN(n9091) );
  AOI211_X1 U10422 ( .C1(n9078), .C2(n9077), .A(n9091), .B(n9115), .ZN(n9088)
         );
  AOI21_X1 U10423 ( .B1(n9080), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9079), .ZN(
        n9083) );
  NAND2_X1 U10424 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9098), .ZN(n9081) );
  OAI21_X1 U10425 ( .B1(n9098), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9081), .ZN(
        n9082) );
  NOR2_X1 U10426 ( .A1(n9083), .A2(n9082), .ZN(n9097) );
  AOI211_X1 U10427 ( .C1(n9083), .C2(n9082), .A(n9097), .B(n9647), .ZN(n9087)
         );
  OAI21_X1 U10428 ( .B1(n9096), .B2(n9085), .A(n9084), .ZN(n9086) );
  NOR3_X1 U10429 ( .A1(n9088), .A2(n9087), .A3(n9086), .ZN(n9089) );
  OAI21_X1 U10430 ( .B1(n9629), .B2(n9090), .A(n9089), .ZN(P1_U3258) );
  INV_X1 U10431 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9106) );
  XOR2_X1 U10432 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9111), .Z(n9093) );
  AOI21_X1 U10433 ( .B1(n9098), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9091), .ZN(
        n9092) );
  NAND2_X1 U10434 ( .A1(n9093), .A2(n9092), .ZN(n9110) );
  OAI21_X1 U10435 ( .B1(n9093), .B2(n9092), .A(n9110), .ZN(n9104) );
  INV_X1 U10436 ( .A(n9111), .ZN(n9095) );
  OAI21_X1 U10437 ( .B1(n9096), .B2(n9095), .A(n9094), .ZN(n9103) );
  NAND2_X1 U10438 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9111), .ZN(n9099) );
  OAI21_X1 U10439 ( .B1(n9111), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9099), .ZN(
        n9100) );
  AOI211_X1 U10440 ( .C1(n9101), .C2(n9100), .A(n9107), .B(n9647), .ZN(n9102)
         );
  AOI211_X1 U10441 ( .C1(n9653), .C2(n9104), .A(n9103), .B(n9102), .ZN(n9105)
         );
  OAI21_X1 U10442 ( .B1(n9629), .B2(n9106), .A(n9105), .ZN(P1_U3259) );
  NAND3_X1 U10443 ( .A1(n9117), .A2(n9109), .A3(n9108), .ZN(n9114) );
  OAI21_X1 U10444 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9111), .A(n9110), .ZN(
        n9112) );
  XOR2_X1 U10445 ( .A(n9112), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9116) );
  AOI21_X1 U10446 ( .B1(n9116), .B2(n9653), .A(n9654), .ZN(n9113) );
  NAND2_X1 U10447 ( .A1(n9114), .A2(n9113), .ZN(n9119) );
  OAI22_X1 U10448 ( .A1(n9117), .A2(n9647), .B1(n9116), .B2(n9115), .ZN(n9118)
         );
  MUX2_X1 U10449 ( .A(n9119), .B(n9118), .S(n9305), .Z(n9122) );
  OAI21_X1 U10450 ( .B1(n9629), .B2(n5058), .A(n9120), .ZN(n9121) );
  INV_X1 U10451 ( .A(n9434), .ZN(n9345) );
  INV_X1 U10452 ( .A(n9427), .ZN(n9319) );
  OR2_X2 U10453 ( .A1(n9302), .A2(n9417), .ZN(n9283) );
  INV_X1 U10454 ( .A(n9406), .ZN(n9257) );
  NOR2_X2 U10455 ( .A1(n9228), .A2(n9392), .ZN(n9214) );
  INV_X1 U10456 ( .A(n9388), .ZN(n9202) );
  NAND2_X1 U10457 ( .A1(n9196), .A2(n9180), .ZN(n9175) );
  NOR2_X1 U10458 ( .A1(n9558), .A2(n9175), .ZN(n9124) );
  XNOR2_X1 U10459 ( .A(n9129), .B(n9124), .ZN(n9373) );
  INV_X1 U10460 ( .A(P1_B_REG_SCAN_IN), .ZN(n9125) );
  NOR2_X1 U10461 ( .A1(n9603), .A2(n9125), .ZN(n9126) );
  OR2_X1 U10462 ( .A1(n9683), .A2(n9126), .ZN(n9170) );
  NOR2_X1 U10463 ( .A1(n9127), .A2(n9170), .ZN(n9557) );
  INV_X1 U10464 ( .A(n9557), .ZN(n9128) );
  NOR2_X1 U10465 ( .A1(n9128), .A2(n4381), .ZN(n9132) );
  NOR2_X1 U10466 ( .A1(n9129), .A2(n9694), .ZN(n9130) );
  AOI211_X1 U10467 ( .C1(n4381), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9132), .B(
        n9130), .ZN(n9131) );
  OAI21_X1 U10468 ( .B1(n9176), .B2(n9373), .A(n9131), .ZN(P1_U3261) );
  XNOR2_X1 U10469 ( .A(n9175), .B(n9558), .ZN(n9555) );
  AOI21_X1 U10470 ( .B1(n4381), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9132), .ZN(
        n9134) );
  NAND2_X1 U10471 ( .A1(n9558), .A2(n9309), .ZN(n9133) );
  OAI211_X1 U10472 ( .C1(n9555), .C2(n9176), .A(n9134), .B(n9133), .ZN(
        P1_U3262) );
  NAND2_X1 U10473 ( .A1(n9437), .A2(n9365), .ZN(n9135) );
  NAND2_X1 U10474 ( .A1(n9136), .A2(n9135), .ZN(n9328) );
  OR2_X1 U10475 ( .A1(n9434), .A2(n9322), .ZN(n9137) );
  NAND2_X1 U10476 ( .A1(n9328), .A2(n9137), .ZN(n9139) );
  NAND2_X1 U10477 ( .A1(n9434), .A2(n9322), .ZN(n9138) );
  NAND2_X1 U10478 ( .A1(n9139), .A2(n9138), .ZN(n9313) );
  AND2_X1 U10479 ( .A1(n9427), .A2(n9299), .ZN(n9141) );
  NOR2_X1 U10480 ( .A1(n9417), .A2(n9300), .ZN(n9142) );
  INV_X1 U10481 ( .A(n9417), .ZN(n9285) );
  NOR2_X1 U10482 ( .A1(n9251), .A2(n9144), .ZN(n9145) );
  AOI21_X1 U10483 ( .B1(n9257), .B2(n9273), .A(n9145), .ZN(n9235) );
  OAI22_X1 U10484 ( .A1(n9235), .A2(n9243), .B1(n9262), .B2(n9400), .ZN(n9220)
         );
  XNOR2_X1 U10485 ( .A(n9148), .B(n9166), .ZN(n9378) );
  INV_X1 U10486 ( .A(n9378), .ZN(n9184) );
  NAND2_X1 U10487 ( .A1(n9298), .A2(n9307), .ZN(n9297) );
  NAND2_X1 U10488 ( .A1(n9209), .A2(n9208), .ZN(n9207) );
  INV_X1 U10489 ( .A(n9163), .ZN(n9165) );
  INV_X1 U10490 ( .A(n9166), .ZN(n9167) );
  OAI22_X1 U10491 ( .A1(n9171), .A2(n9685), .B1(n9170), .B2(n10250), .ZN(n9172) );
  INV_X1 U10492 ( .A(n9172), .ZN(n9173) );
  OAI21_X1 U10493 ( .B1(n9196), .B2(n9180), .A(n9175), .ZN(n9379) );
  NOR2_X1 U10494 ( .A1(n9379), .A2(n9176), .ZN(n9182) );
  INV_X1 U10495 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U10496 ( .A1(n9178), .A2(n9357), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n4381), .ZN(n9179) );
  OAI21_X1 U10497 ( .B1(n9180), .B2(n9694), .A(n9179), .ZN(n9181) );
  AOI211_X1 U10498 ( .C1(n9382), .C2(n9692), .A(n9182), .B(n9181), .ZN(n9183)
         );
  OAI21_X1 U10499 ( .B1(n9184), .B2(n9370), .A(n9183), .ZN(P1_U3355) );
  AOI21_X1 U10500 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9385) );
  INV_X1 U10501 ( .A(n9385), .ZN(n9205) );
  XNOR2_X1 U10502 ( .A(n9188), .B(n8033), .ZN(n9190) );
  NAND2_X1 U10503 ( .A1(n9190), .A2(n9189), .ZN(n9195) );
  NOR2_X1 U10504 ( .A1(n9227), .A2(n9685), .ZN(n9193) );
  NOR2_X1 U10505 ( .A1(n9191), .A2(n9683), .ZN(n9192) );
  INV_X1 U10506 ( .A(n9214), .ZN(n9197) );
  AOI211_X1 U10507 ( .C1(n9388), .C2(n9197), .A(n9753), .B(n9196), .ZN(n9387)
         );
  NAND2_X1 U10508 ( .A1(n9387), .A2(n9340), .ZN(n9201) );
  INV_X1 U10509 ( .A(n9198), .ZN(n9199) );
  AOI22_X1 U10510 ( .A1(n9199), .A2(n9357), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4381), .ZN(n9200) );
  OAI211_X1 U10511 ( .C1(n9202), .C2(n9694), .A(n9201), .B(n9200), .ZN(n9203)
         );
  AOI21_X1 U10512 ( .B1(n9386), .B2(n9692), .A(n9203), .ZN(n9204) );
  OAI21_X1 U10513 ( .B1(n9205), .B2(n9370), .A(n9204), .ZN(P1_U3263) );
  XOR2_X1 U10514 ( .A(n9208), .B(n9206), .Z(n9394) );
  AOI22_X1 U10515 ( .A1(n9392), .A2(n9309), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4381), .ZN(n9219) );
  OAI211_X1 U10516 ( .C1(n9209), .C2(n9208), .A(n9207), .B(n9189), .ZN(n9212)
         );
  NAND2_X1 U10517 ( .A1(n9210), .A2(n9664), .ZN(n9211) );
  OAI211_X1 U10518 ( .C1(n9213), .C2(n9685), .A(n9212), .B(n9211), .ZN(n9390)
         );
  AOI211_X1 U10519 ( .C1(n9392), .C2(n9228), .A(n9753), .B(n9214), .ZN(n9391)
         );
  INV_X1 U10520 ( .A(n9391), .ZN(n9216) );
  OAI22_X1 U10521 ( .A1(n9216), .A2(n9670), .B1(n9693), .B2(n9215), .ZN(n9217)
         );
  OAI21_X1 U10522 ( .B1(n9390), .B2(n9217), .A(n9692), .ZN(n9218) );
  OAI211_X1 U10523 ( .C1(n9394), .C2(n9370), .A(n9219), .B(n9218), .ZN(
        P1_U3264) );
  XNOR2_X1 U10524 ( .A(n9220), .B(n9223), .ZN(n9399) );
  NAND2_X1 U10525 ( .A1(n9222), .A2(n9221), .ZN(n9224) );
  XNOR2_X1 U10526 ( .A(n9224), .B(n9223), .ZN(n9225) );
  OAI222_X1 U10527 ( .A1(n9683), .A2(n9227), .B1(n9685), .B2(n9226), .C1(n9672), .C2(n9225), .ZN(n9395) );
  AOI211_X1 U10528 ( .C1(n9397), .C2(n9236), .A(n9753), .B(n4609), .ZN(n9396)
         );
  NAND2_X1 U10529 ( .A1(n9396), .A2(n9340), .ZN(n9231) );
  AOI22_X1 U10530 ( .A1(n9229), .A2(n9357), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4381), .ZN(n9230) );
  OAI211_X1 U10531 ( .C1(n9232), .C2(n9694), .A(n9231), .B(n9230), .ZN(n9233)
         );
  AOI21_X1 U10532 ( .B1(n9395), .B2(n9692), .A(n9233), .ZN(n9234) );
  OAI21_X1 U10533 ( .B1(n9399), .B2(n9370), .A(n9234), .ZN(P1_U3265) );
  XOR2_X1 U10534 ( .A(n9243), .B(n9235), .Z(n9404) );
  INV_X1 U10535 ( .A(n9252), .ZN(n9237) );
  AOI21_X1 U10536 ( .B1(n9400), .B2(n9237), .A(n4610), .ZN(n9401) );
  INV_X1 U10537 ( .A(n9238), .ZN(n9239) );
  AOI22_X1 U10538 ( .A1(n9239), .A2(n9357), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4381), .ZN(n9240) );
  OAI21_X1 U10539 ( .B1(n9241), .B2(n9694), .A(n9240), .ZN(n9249) );
  NAND2_X1 U10540 ( .A1(n9258), .A2(n9242), .ZN(n9244) );
  XNOR2_X1 U10541 ( .A(n9244), .B(n9243), .ZN(n9247) );
  AOI222_X1 U10542 ( .A1(n9189), .A2(n9247), .B1(n9246), .B2(n9664), .C1(n9245), .C2(n9363), .ZN(n9403) );
  NOR2_X1 U10543 ( .A1(n9403), .A2(n4381), .ZN(n9248) );
  AOI211_X1 U10544 ( .C1(n9401), .C2(n9679), .A(n9249), .B(n9248), .ZN(n9250)
         );
  OAI21_X1 U10545 ( .B1(n9404), .B2(n9370), .A(n9250), .ZN(P1_U3266) );
  XOR2_X1 U10546 ( .A(n9251), .B(n9260), .Z(n9409) );
  INV_X1 U10547 ( .A(n9274), .ZN(n9253) );
  AOI211_X1 U10548 ( .C1(n9406), .C2(n9253), .A(n9753), .B(n9252), .ZN(n9405)
         );
  INV_X1 U10549 ( .A(n9254), .ZN(n9255) );
  AOI22_X1 U10550 ( .A1(n9255), .A2(n9357), .B1(n4381), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9256) );
  OAI21_X1 U10551 ( .B1(n9257), .B2(n9694), .A(n9256), .ZN(n9265) );
  OAI21_X1 U10552 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9263) );
  AOI222_X1 U10553 ( .A1(n9189), .A2(n9263), .B1(n9262), .B2(n9664), .C1(n9261), .C2(n9363), .ZN(n9408) );
  NOR2_X1 U10554 ( .A1(n9408), .A2(n4381), .ZN(n9264) );
  AOI211_X1 U10555 ( .C1(n9405), .C2(n9340), .A(n9265), .B(n9264), .ZN(n9266)
         );
  OAI21_X1 U10556 ( .B1(n9409), .B2(n9370), .A(n9266), .ZN(P1_U3267) );
  XNOR2_X1 U10557 ( .A(n9268), .B(n9267), .ZN(n9414) );
  XNOR2_X1 U10558 ( .A(n9270), .B(n9269), .ZN(n9271) );
  OAI222_X1 U10559 ( .A1(n9683), .A2(n9273), .B1(n9685), .B2(n9272), .C1(n9672), .C2(n9271), .ZN(n9410) );
  AOI211_X1 U10560 ( .C1(n9412), .C2(n9283), .A(n9753), .B(n9274), .ZN(n9411)
         );
  NAND2_X1 U10561 ( .A1(n9411), .A2(n9340), .ZN(n9278) );
  INV_X1 U10562 ( .A(n9275), .ZN(n9276) );
  AOI22_X1 U10563 ( .A1(n4381), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9276), .B2(
        n9357), .ZN(n9277) );
  OAI211_X1 U10564 ( .C1(n9279), .C2(n9694), .A(n9278), .B(n9277), .ZN(n9280)
         );
  AOI21_X1 U10565 ( .B1(n9410), .B2(n9692), .A(n9280), .ZN(n9281) );
  OAI21_X1 U10566 ( .B1(n9414), .B2(n9370), .A(n9281), .ZN(P1_U3268) );
  XOR2_X1 U10567 ( .A(n9290), .B(n9282), .Z(n9419) );
  INV_X1 U10568 ( .A(n9283), .ZN(n9284) );
  AOI211_X1 U10569 ( .C1(n9417), .C2(n9302), .A(n9753), .B(n9284), .ZN(n9416)
         );
  NOR2_X1 U10570 ( .A1(n9285), .A2(n9694), .ZN(n9289) );
  OAI22_X1 U10571 ( .A1(n9692), .A2(n9287), .B1(n9286), .B2(n9693), .ZN(n9288)
         );
  AOI211_X1 U10572 ( .C1(n9416), .C2(n9340), .A(n9289), .B(n9288), .ZN(n9296)
         );
  XNOR2_X1 U10573 ( .A(n9291), .B(n9290), .ZN(n9292) );
  OAI222_X1 U10574 ( .A1(n9683), .A2(n9294), .B1(n9685), .B2(n9293), .C1(n9292), .C2(n9672), .ZN(n9415) );
  NAND2_X1 U10575 ( .A1(n9415), .A2(n9692), .ZN(n9295) );
  OAI211_X1 U10576 ( .C1(n9419), .C2(n9370), .A(n9296), .B(n9295), .ZN(
        P1_U3269) );
  OAI21_X1 U10577 ( .B1(n9307), .B2(n9298), .A(n9297), .ZN(n9301) );
  AOI222_X1 U10578 ( .A1(n9189), .A2(n9301), .B1(n9300), .B2(n9664), .C1(n9299), .C2(n9363), .ZN(n9424) );
  INV_X1 U10579 ( .A(n9314), .ZN(n9303) );
  AOI211_X1 U10580 ( .C1(n9422), .C2(n9303), .A(n9753), .B(n4601), .ZN(n9421)
         );
  AOI22_X1 U10581 ( .A1(n9421), .A2(n9305), .B1(n9357), .B2(n9304), .ZN(n9306)
         );
  AND2_X1 U10582 ( .A1(n9424), .A2(n9306), .ZN(n9312) );
  NAND2_X1 U10583 ( .A1(n9308), .A2(n9307), .ZN(n9420) );
  NAND3_X1 U10584 ( .A1(n4794), .A2(n7395), .A3(n9420), .ZN(n9311) );
  AOI22_X1 U10585 ( .A1(n9422), .A2(n9309), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n4381), .ZN(n9310) );
  OAI211_X1 U10586 ( .C1(n4381), .C2(n9312), .A(n9311), .B(n9310), .ZN(
        P1_U3270) );
  XNOR2_X1 U10587 ( .A(n9313), .B(n9320), .ZN(n9431) );
  INV_X1 U10588 ( .A(n9338), .ZN(n9315) );
  AOI21_X1 U10589 ( .B1(n9427), .B2(n9315), .A(n9314), .ZN(n9428) );
  INV_X1 U10590 ( .A(n9316), .ZN(n9317) );
  AOI22_X1 U10591 ( .A1(n4381), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9317), .B2(
        n9357), .ZN(n9318) );
  OAI21_X1 U10592 ( .B1(n9319), .B2(n9694), .A(n9318), .ZN(n9326) );
  XNOR2_X1 U10593 ( .A(n9321), .B(n9320), .ZN(n9324) );
  AOI222_X1 U10594 ( .A1(n9189), .A2(n9324), .B1(n9323), .B2(n9664), .C1(n9322), .C2(n9363), .ZN(n9430) );
  NOR2_X1 U10595 ( .A1(n9430), .A2(n4381), .ZN(n9325) );
  AOI211_X1 U10596 ( .C1(n9428), .C2(n9679), .A(n9326), .B(n9325), .ZN(n9327)
         );
  OAI21_X1 U10597 ( .B1(n9370), .B2(n9431), .A(n9327), .ZN(P1_U3271) );
  XNOR2_X1 U10598 ( .A(n9328), .B(n9329), .ZN(n9436) );
  NOR2_X1 U10599 ( .A1(n4720), .A2(n4719), .ZN(n9333) );
  AOI21_X1 U10600 ( .B1(n9333), .B2(n9332), .A(n9331), .ZN(n9334) );
  OAI222_X1 U10601 ( .A1(n9683), .A2(n9336), .B1(n9685), .B2(n9335), .C1(n9672), .C2(n9334), .ZN(n9432) );
  INV_X1 U10602 ( .A(n9337), .ZN(n9339) );
  AOI211_X1 U10603 ( .C1(n9434), .C2(n9339), .A(n9753), .B(n9338), .ZN(n9433)
         );
  NAND2_X1 U10604 ( .A1(n9433), .A2(n9340), .ZN(n9344) );
  INV_X1 U10605 ( .A(n9341), .ZN(n9342) );
  AOI22_X1 U10606 ( .A1(n4381), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9342), .B2(
        n9357), .ZN(n9343) );
  OAI211_X1 U10607 ( .C1(n9345), .C2(n9694), .A(n9344), .B(n9343), .ZN(n9346)
         );
  AOI21_X1 U10608 ( .B1(n9432), .B2(n9692), .A(n9346), .ZN(n9347) );
  OAI21_X1 U10609 ( .B1(n9436), .B2(n9370), .A(n9347), .ZN(P1_U3272) );
  OR2_X1 U10610 ( .A1(n7912), .A2(n9348), .ZN(n9350) );
  NAND2_X1 U10611 ( .A1(n9350), .A2(n9349), .ZN(n9352) );
  XNOR2_X1 U10612 ( .A(n9352), .B(n9351), .ZN(n9446) );
  INV_X1 U10613 ( .A(n9353), .ZN(n9354) );
  AOI21_X1 U10614 ( .B1(n9442), .B2(n9355), .A(n9354), .ZN(n9443) );
  INV_X1 U10615 ( .A(n9356), .ZN(n9358) );
  AOI22_X1 U10616 ( .A1(n4381), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9358), .B2(
        n9357), .ZN(n9359) );
  OAI21_X1 U10617 ( .B1(n9360), .B2(n9694), .A(n9359), .ZN(n9368) );
  XNOR2_X1 U10618 ( .A(n9362), .B(n9361), .ZN(n9366) );
  AOI222_X1 U10619 ( .A1(n9189), .A2(n9366), .B1(n9365), .B2(n9664), .C1(n9364), .C2(n9363), .ZN(n9445) );
  NOR2_X1 U10620 ( .A1(n9445), .A2(n4381), .ZN(n9367) );
  AOI211_X1 U10621 ( .C1(n9443), .C2(n9679), .A(n9368), .B(n9367), .ZN(n9369)
         );
  OAI21_X1 U10622 ( .B1(n9370), .B2(n9446), .A(n9369), .ZN(P1_U3274) );
  AOI21_X1 U10623 ( .B1(n9371), .B2(n9727), .A(n9557), .ZN(n9372) );
  OAI21_X1 U10624 ( .B1(n9373), .B2(n9753), .A(n9372), .ZN(n9456) );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9456), .S(n9772), .Z(
        P1_U3554) );
  INV_X1 U10626 ( .A(n9374), .ZN(n9375) );
  NAND2_X1 U10627 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  NAND2_X1 U10628 ( .A1(n9378), .A2(n9755), .ZN(n9384) );
  NAND2_X1 U10629 ( .A1(n9384), .A2(n9383), .ZN(n9457) );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9457), .S(n9772), .Z(
        P1_U3552) );
  NAND2_X1 U10631 ( .A1(n9385), .A2(n9755), .ZN(n9389) );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9458), .S(n9772), .Z(
        P1_U3551) );
  AOI211_X1 U10633 ( .C1(n9727), .C2(n9392), .A(n9391), .B(n9390), .ZN(n9393)
         );
  OAI21_X1 U10634 ( .B1(n9394), .B2(n9740), .A(n9393), .ZN(n9459) );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9459), .S(n9772), .Z(
        P1_U3550) );
  AOI211_X1 U10636 ( .C1(n9727), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9398)
         );
  OAI21_X1 U10637 ( .B1(n9399), .B2(n9740), .A(n9398), .ZN(n9460) );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9460), .S(n9772), .Z(
        P1_U3549) );
  AOI22_X1 U10639 ( .A1(n9401), .A2(n9728), .B1(n9727), .B2(n9400), .ZN(n9402)
         );
  OAI211_X1 U10640 ( .C1(n9404), .C2(n9740), .A(n9403), .B(n9402), .ZN(n9461)
         );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9461), .S(n9772), .Z(
        P1_U3548) );
  AOI21_X1 U10642 ( .B1(n9727), .B2(n9406), .A(n9405), .ZN(n9407) );
  OAI211_X1 U10643 ( .C1(n9409), .C2(n9740), .A(n9408), .B(n9407), .ZN(n9462)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9462), .S(n9772), .Z(
        P1_U3547) );
  AOI211_X1 U10645 ( .C1(n9727), .C2(n9412), .A(n9411), .B(n9410), .ZN(n9413)
         );
  OAI21_X1 U10646 ( .B1(n9414), .B2(n9740), .A(n9413), .ZN(n9463) );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9463), .S(n9772), .Z(
        P1_U3546) );
  AOI211_X1 U10648 ( .C1(n9727), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9418)
         );
  OAI21_X1 U10649 ( .B1(n9419), .B2(n9740), .A(n9418), .ZN(n9464) );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9464), .S(n9772), .Z(
        P1_U3545) );
  NAND2_X1 U10651 ( .A1(n9420), .A2(n9755), .ZN(n9425) );
  AOI21_X1 U10652 ( .B1(n9727), .B2(n9422), .A(n9421), .ZN(n9423) );
  OAI211_X1 U10653 ( .C1(n9426), .C2(n9425), .A(n9424), .B(n9423), .ZN(n9465)
         );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9465), .S(n9772), .Z(
        P1_U3544) );
  AOI22_X1 U10655 ( .A1(n9428), .A2(n9728), .B1(n9727), .B2(n9427), .ZN(n9429)
         );
  OAI211_X1 U10656 ( .C1(n9431), .C2(n9740), .A(n9430), .B(n9429), .ZN(n9466)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9466), .S(n9772), .Z(
        P1_U3543) );
  AOI211_X1 U10658 ( .C1(n9727), .C2(n9434), .A(n9433), .B(n9432), .ZN(n9435)
         );
  OAI21_X1 U10659 ( .B1(n9740), .B2(n9436), .A(n9435), .ZN(n9467) );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9467), .S(n9772), .Z(
        P1_U3542) );
  AOI22_X1 U10661 ( .A1(n9438), .A2(n9728), .B1(n9727), .B2(n9437), .ZN(n9439)
         );
  OAI211_X1 U10662 ( .C1(n9441), .C2(n9740), .A(n9440), .B(n9439), .ZN(n9468)
         );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9468), .S(n9772), .Z(
        P1_U3541) );
  AOI22_X1 U10664 ( .A1(n9443), .A2(n9728), .B1(n9727), .B2(n9442), .ZN(n9444)
         );
  OAI211_X1 U10665 ( .C1(n9446), .C2(n9740), .A(n9445), .B(n9444), .ZN(n9469)
         );
  MUX2_X1 U10666 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9469), .S(n9772), .Z(
        P1_U3540) );
  AOI211_X1 U10667 ( .C1(n9727), .C2(n7905), .A(n9448), .B(n9447), .ZN(n9449)
         );
  OAI21_X1 U10668 ( .B1(n9740), .B2(n9450), .A(n9449), .ZN(n9470) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9470), .S(n9772), .Z(
        P1_U3539) );
  AOI211_X1 U10670 ( .C1(n9727), .C2(n9453), .A(n9452), .B(n9451), .ZN(n9454)
         );
  OAI21_X1 U10671 ( .B1(n9455), .B2(n9740), .A(n9454), .ZN(n9471) );
  MUX2_X1 U10672 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9471), .S(n9772), .Z(
        P1_U3538) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9456), .S(n9759), .Z(
        P1_U3522) );
  MUX2_X1 U10674 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9457), .S(n9759), .Z(
        P1_U3520) );
  MUX2_X1 U10675 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9459), .S(n9759), .Z(
        P1_U3518) );
  MUX2_X1 U10676 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9460), .S(n9759), .Z(
        P1_U3517) );
  MUX2_X1 U10677 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9461), .S(n9759), .Z(
        P1_U3516) );
  MUX2_X1 U10678 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9462), .S(n9759), .Z(
        P1_U3515) );
  MUX2_X1 U10679 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9463), .S(n9759), .Z(
        P1_U3514) );
  MUX2_X1 U10680 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9464), .S(n9759), .Z(
        P1_U3513) );
  MUX2_X1 U10681 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9465), .S(n9759), .Z(
        P1_U3512) );
  MUX2_X1 U10682 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9466), .S(n9759), .Z(
        P1_U3511) );
  MUX2_X1 U10683 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9467), .S(n9759), .Z(
        P1_U3510) );
  MUX2_X1 U10684 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9468), .S(n9759), .Z(
        P1_U3508) );
  MUX2_X1 U10685 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9469), .S(n9759), .Z(
        P1_U3505) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9470), .S(n9759), .Z(
        P1_U3502) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9471), .S(n9759), .Z(
        P1_U3499) );
  NOR4_X1 U10688 ( .A1(n9472), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n4595), .ZN(n9473) );
  AOI21_X1 U10689 ( .B1(n9474), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9473), .ZN(
        n9475) );
  OAI21_X1 U10690 ( .B1(n9476), .B2(n9479), .A(n9475), .ZN(P1_U3322) );
  OAI222_X1 U10691 ( .A1(n7945), .A2(n10227), .B1(n9479), .B2(n9478), .C1(
        P1_U3084), .C2(n9477), .ZN(P1_U3323) );
  MUX2_X1 U10692 ( .A(n9480), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10693 ( .A1(n9775), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9491) );
  OR2_X1 U10694 ( .A1(n9777), .A2(n9481), .ZN(n9485) );
  OAI211_X1 U10695 ( .C1(n9483), .C2(n9482), .A(n9773), .B(n4645), .ZN(n9484)
         );
  AND2_X1 U10696 ( .A1(n9485), .A2(n9484), .ZN(n9490) );
  OAI211_X1 U10697 ( .C1(n9488), .C2(n9487), .A(n9774), .B(n9486), .ZN(n9489)
         );
  NAND3_X1 U10698 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(P2_U3247) );
  OAI21_X1 U10699 ( .B1(n9493), .B2(n9742), .A(n9492), .ZN(n9494) );
  AOI211_X1 U10700 ( .C1(n9496), .C2(n9755), .A(n9495), .B(n9494), .ZN(n9498)
         );
  INV_X1 U10701 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9497) );
  AOI22_X1 U10702 ( .A1(n9759), .A2(n9498), .B1(n9497), .B2(n9757), .ZN(
        P1_U3484) );
  AOI22_X1 U10703 ( .A1(n9772), .A2(n9498), .B1(n6878), .B2(n9770), .ZN(
        P1_U3533) );
  NAND2_X1 U10704 ( .A1(n9500), .A2(n9499), .ZN(n9502) );
  OAI211_X1 U10705 ( .C1(n9504), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9505)
         );
  INV_X1 U10706 ( .A(n9505), .ZN(n9515) );
  NOR2_X1 U10707 ( .A1(n9506), .A2(n9742), .ZN(n9574) );
  NAND2_X1 U10708 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  AOI21_X1 U10709 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9512) );
  AOI21_X1 U10710 ( .B1(n9513), .B2(n9574), .A(n9512), .ZN(n9514) );
  OAI211_X1 U10711 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9514), .ZN(
        P1_U3222) );
  INV_X1 U10712 ( .A(n9518), .ZN(n9520) );
  OAI21_X1 U10713 ( .B1(n9520), .B2(n9542), .A(n9519), .ZN(n9543) );
  INV_X1 U10714 ( .A(n9543), .ZN(n9522) );
  AOI22_X1 U10715 ( .A1(n9522), .A2(n9521), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n9808), .ZN(n9540) );
  OAI21_X1 U10716 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9546) );
  INV_X1 U10717 ( .A(n9526), .ZN(n9527) );
  NOR2_X1 U10718 ( .A1(n9542), .A2(n9527), .ZN(n9536) );
  XNOR2_X1 U10719 ( .A(n9528), .B(n9529), .ZN(n9530) );
  OAI222_X1 U10720 ( .A1(n9535), .A2(n9534), .B1(n9533), .B2(n9532), .C1(n9531), .C2(n9530), .ZN(n9544) );
  AOI211_X1 U10721 ( .C1(n9537), .C2(n9546), .A(n9536), .B(n9544), .ZN(n9538)
         );
  OR2_X1 U10722 ( .A1(n9538), .A2(n9808), .ZN(n9539) );
  OAI211_X1 U10723 ( .C1(n9541), .C2(n9793), .A(n9540), .B(n9539), .ZN(
        P2_U3281) );
  OAI22_X1 U10724 ( .A1(n9543), .A2(n9900), .B1(n9542), .B2(n9899), .ZN(n9545)
         );
  AOI211_X1 U10725 ( .C1(n9904), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9553)
         );
  AOI22_X1 U10726 ( .A1(n9924), .A2(n9553), .B1(n10145), .B2(n9922), .ZN(
        P2_U3535) );
  OAI21_X1 U10727 ( .B1(n9548), .B2(n9899), .A(n9547), .ZN(n9550) );
  AOI211_X1 U10728 ( .C1(n9551), .C2(n9904), .A(n9550), .B(n9549), .ZN(n9554)
         );
  AOI22_X1 U10729 ( .A1(n9924), .A2(n9554), .B1(n9552), .B2(n9922), .ZN(
        P2_U3534) );
  INV_X1 U10730 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U10731 ( .A1(n9908), .A2(n9553), .B1(n9983), .B2(n9906), .ZN(
        P2_U3496) );
  INV_X1 U10732 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U10733 ( .A1(n9908), .A2(n9554), .B1(n10187), .B2(n9906), .ZN(
        P2_U3493) );
  NOR2_X1 U10734 ( .A1(n9555), .A2(n9753), .ZN(n9556) );
  AOI211_X1 U10735 ( .C1(n9727), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9581)
         );
  INV_X1 U10736 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10737 ( .A1(n9772), .A2(n9581), .B1(n9559), .B2(n9770), .ZN(
        P1_U3553) );
  OAI21_X1 U10738 ( .B1(n9561), .B2(n9742), .A(n9560), .ZN(n9562) );
  AOI211_X1 U10739 ( .C1(n9564), .C2(n9755), .A(n9563), .B(n9562), .ZN(n9583)
         );
  AOI22_X1 U10740 ( .A1(n9772), .A2(n9583), .B1(n7491), .B2(n9770), .ZN(
        P1_U3537) );
  INV_X1 U10741 ( .A(n9565), .ZN(n9566) );
  OAI21_X1 U10742 ( .B1(n9567), .B2(n9753), .A(n9566), .ZN(n9568) );
  AOI211_X1 U10743 ( .C1(n9570), .C2(n9755), .A(n9569), .B(n9568), .ZN(n9584)
         );
  AOI22_X1 U10744 ( .A1(n9772), .A2(n9584), .B1(n7179), .B2(n9770), .ZN(
        P1_U3536) );
  NOR2_X1 U10745 ( .A1(n9571), .A2(n9740), .ZN(n9575) );
  NOR4_X1 U10746 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n9585)
         );
  AOI22_X1 U10747 ( .A1(n9772), .A2(n9585), .B1(n6985), .B2(n9770), .ZN(
        P1_U3535) );
  OAI22_X1 U10748 ( .A1(n9577), .A2(n9753), .B1(n9576), .B2(n9742), .ZN(n9578)
         );
  AOI211_X1 U10749 ( .C1(n9580), .C2(n9755), .A(n9579), .B(n9578), .ZN(n9586)
         );
  AOI22_X1 U10750 ( .A1(n9772), .A2(n9586), .B1(n5317), .B2(n9770), .ZN(
        P1_U3534) );
  INV_X1 U10751 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U10752 ( .A1(n9759), .A2(n9581), .B1(n10176), .B2(n9757), .ZN(
        P1_U3521) );
  INV_X1 U10753 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9582) );
  AOI22_X1 U10754 ( .A1(n9759), .A2(n9583), .B1(n9582), .B2(n9757), .ZN(
        P1_U3496) );
  INV_X1 U10755 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U10756 ( .A1(n9759), .A2(n9584), .B1(n10075), .B2(n9757), .ZN(
        P1_U3493) );
  INV_X1 U10757 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U10758 ( .A1(n9759), .A2(n9585), .B1(n10194), .B2(n9757), .ZN(
        P1_U3490) );
  INV_X1 U10759 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U10760 ( .A1(n9759), .A2(n9586), .B1(n10069), .B2(n9757), .ZN(
        P1_U3487) );
  XNOR2_X1 U10761 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10762 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U10764 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6708), .S(n9587), .Z(n9590)
         );
  NAND3_X1 U10765 ( .A1(n9590), .A2(n9589), .A3(n9588), .ZN(n9591) );
  AND3_X1 U10766 ( .A1(n9593), .A2(n9592), .A3(n9591), .ZN(n9602) );
  INV_X1 U10767 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9600) );
  OAI211_X1 U10768 ( .C1(n9596), .C2(n9595), .A(n9653), .B(n9594), .ZN(n9599)
         );
  NAND2_X1 U10769 ( .A1(n9654), .A2(n9597), .ZN(n9598) );
  OAI211_X1 U10770 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9600), .A(n9599), .B(
        n9598), .ZN(n9601) );
  NOR2_X1 U10771 ( .A1(n9602), .A2(n9601), .ZN(n9610) );
  MUX2_X1 U10772 ( .A(n9605), .B(n9604), .S(n9603), .Z(n9607) );
  NAND2_X1 U10773 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  OAI211_X1 U10774 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9609), .A(n9608), .B(
        P1_U4006), .ZN(n9627) );
  OAI211_X1 U10775 ( .C1(n9611), .C2(n9629), .A(n9610), .B(n9627), .ZN(
        P1_U3243) );
  INV_X1 U10776 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U10777 ( .A1(n9613), .A2(n9612), .ZN(n9614) );
  NOR2_X1 U10778 ( .A1(n9615), .A2(n9614), .ZN(n9625) );
  AND2_X1 U10779 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  OAI21_X1 U10780 ( .B1(n9619), .B2(n9618), .A(n9653), .ZN(n9624) );
  INV_X1 U10781 ( .A(n9620), .ZN(n9622) );
  AOI21_X1 U10782 ( .B1(n9654), .B2(n9622), .A(n9621), .ZN(n9623) );
  OAI211_X1 U10783 ( .C1(n9625), .C2(n9647), .A(n9624), .B(n9623), .ZN(n9626)
         );
  INV_X1 U10784 ( .A(n9626), .ZN(n9628) );
  OAI211_X1 U10785 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(
        P1_U3245) );
  OAI21_X1 U10786 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9639) );
  AOI211_X1 U10787 ( .C1(n9636), .C2(n9635), .A(n9647), .B(n9634), .ZN(n9637)
         );
  AOI211_X1 U10788 ( .C1(n9653), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9642)
         );
  AOI22_X1 U10789 ( .A1(n9656), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9640), .B2(
        n9654), .ZN(n9641) );
  NAND2_X1 U10790 ( .A1(n9642), .A2(n9641), .ZN(P1_U3250) );
  OAI21_X1 U10791 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9652) );
  AOI211_X1 U10792 ( .C1(n9649), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9650)
         );
  AOI211_X1 U10793 ( .C1(n9653), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9658)
         );
  AOI22_X1 U10794 ( .A1(n9656), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9655), .B2(
        n9654), .ZN(n9657) );
  NAND2_X1 U10795 ( .A1(n9658), .A2(n9657), .ZN(P1_U3251) );
  XNOR2_X1 U10796 ( .A(n9660), .B(n9659), .ZN(n9725) );
  AOI21_X1 U10797 ( .B1(n9661), .B2(n9668), .A(n9753), .ZN(n9663) );
  NAND2_X1 U10798 ( .A1(n9663), .A2(n9662), .ZN(n9721) );
  NAND2_X1 U10799 ( .A1(n9665), .A2(n9664), .ZN(n9720) );
  OAI21_X1 U10800 ( .B1(n9693), .B2(n9666), .A(n9720), .ZN(n9667) );
  AOI21_X1 U10801 ( .B1(n5008), .B2(n9668), .A(n9667), .ZN(n9669) );
  OAI21_X1 U10802 ( .B1(n9721), .B2(n9670), .A(n9669), .ZN(n9674) );
  XNOR2_X1 U10803 ( .A(n9671), .B(n7208), .ZN(n9673) );
  OAI22_X1 U10804 ( .A1(n9673), .A2(n9672), .B1(n9684), .B2(n9685), .ZN(n9723)
         );
  AOI211_X1 U10805 ( .C1(n9675), .C2(n9725), .A(n9674), .B(n9723), .ZN(n9676)
         );
  AOI22_X1 U10806 ( .A1(n4381), .A2(n5166), .B1(n9676), .B2(n9692), .ZN(
        P1_U3286) );
  OAI21_X1 U10807 ( .B1(n9678), .B2(n9709), .A(n9677), .ZN(n9710) );
  INV_X1 U10808 ( .A(n9710), .ZN(n9680) );
  NAND2_X1 U10809 ( .A1(n9680), .A2(n9679), .ZN(n9698) );
  XNOR2_X1 U10810 ( .A(n9681), .B(n4566), .ZN(n9691) );
  XNOR2_X1 U10811 ( .A(n9682), .B(n4566), .ZN(n9688) );
  OAI22_X1 U10812 ( .A1(n9686), .A2(n9685), .B1(n9684), .B2(n9683), .ZN(n9687)
         );
  AOI21_X1 U10813 ( .B1(n9688), .B2(n9189), .A(n9687), .ZN(n9689) );
  OAI21_X1 U10814 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9711) );
  MUX2_X1 U10815 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9711), .S(n9692), .Z(n9696)
         );
  OAI22_X1 U10816 ( .A1(n9694), .A2(n9709), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9693), .ZN(n9695) );
  NOR2_X1 U10817 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  NAND2_X1 U10818 ( .A1(n9698), .A2(n9697), .ZN(P1_U3288) );
  AND2_X1 U10819 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9700), .ZN(P1_U3292) );
  AND2_X1 U10820 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9700), .ZN(P1_U3293) );
  AND2_X1 U10821 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9700), .ZN(P1_U3294) );
  AND2_X1 U10822 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9700), .ZN(P1_U3295) );
  AND2_X1 U10823 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9700), .ZN(P1_U3296) );
  AND2_X1 U10824 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9700), .ZN(P1_U3297) );
  AND2_X1 U10825 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9700), .ZN(P1_U3298) );
  INV_X1 U10826 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9993) );
  NOR2_X1 U10827 ( .A1(n9699), .A2(n9993), .ZN(P1_U3299) );
  AND2_X1 U10828 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9700), .ZN(P1_U3300) );
  AND2_X1 U10829 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9700), .ZN(P1_U3301) );
  AND2_X1 U10830 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9700), .ZN(P1_U3302) );
  INV_X1 U10831 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9979) );
  NOR2_X1 U10832 ( .A1(n9699), .A2(n9979), .ZN(P1_U3303) );
  INV_X1 U10833 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10020) );
  NOR2_X1 U10834 ( .A1(n9699), .A2(n10020), .ZN(P1_U3304) );
  AND2_X1 U10835 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9700), .ZN(P1_U3305) );
  AND2_X1 U10836 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9700), .ZN(P1_U3306) );
  AND2_X1 U10837 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9700), .ZN(P1_U3307) );
  AND2_X1 U10838 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9700), .ZN(P1_U3308) );
  AND2_X1 U10839 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9700), .ZN(P1_U3309) );
  INV_X1 U10840 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U10841 ( .A1(n9699), .A2(n9954), .ZN(P1_U3310) );
  INV_X1 U10842 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U10843 ( .A1(n9699), .A2(n9956), .ZN(P1_U3311) );
  AND2_X1 U10844 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9700), .ZN(P1_U3312) );
  AND2_X1 U10845 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9700), .ZN(P1_U3313) );
  AND2_X1 U10846 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9700), .ZN(P1_U3314) );
  AND2_X1 U10847 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9700), .ZN(P1_U3315) );
  INV_X1 U10848 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U10849 ( .A1(n9699), .A2(n10123), .ZN(P1_U3316) );
  INV_X1 U10850 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U10851 ( .A1(n9699), .A2(n10067), .ZN(P1_U3317) );
  AND2_X1 U10852 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9700), .ZN(P1_U3318) );
  INV_X1 U10853 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U10854 ( .A1(n9699), .A2(n10184), .ZN(P1_U3319) );
  AND2_X1 U10855 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9700), .ZN(P1_U3320) );
  AND2_X1 U10856 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9700), .ZN(P1_U3321) );
  NAND2_X1 U10857 ( .A1(n9702), .A2(n9701), .ZN(n9704) );
  AOI211_X1 U10858 ( .C1(n9705), .C2(n9755), .A(n9704), .B(n9703), .ZN(n9761)
         );
  INV_X1 U10859 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9706) );
  AOI22_X1 U10860 ( .A1(n9759), .A2(n9761), .B1(n9706), .B2(n9757), .ZN(
        P1_U3457) );
  INV_X1 U10861 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U10862 ( .A1(n9759), .A2(n9708), .B1(n9707), .B2(n9757), .ZN(
        P1_U3460) );
  OAI22_X1 U10863 ( .A1(n9710), .A2(n9753), .B1(n9709), .B2(n9742), .ZN(n9712)
         );
  NOR2_X1 U10864 ( .A1(n9712), .A2(n9711), .ZN(n9763) );
  INV_X1 U10865 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U10866 ( .A1(n9759), .A2(n9763), .B1(n9713), .B2(n9757), .ZN(
        P1_U3463) );
  OAI22_X1 U10867 ( .A1(n9715), .A2(n9753), .B1(n9714), .B2(n9742), .ZN(n9716)
         );
  INV_X1 U10868 ( .A(n9716), .ZN(n9717) );
  AND2_X1 U10869 ( .A1(n9718), .A2(n9717), .ZN(n9764) );
  INV_X1 U10870 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10871 ( .A1(n9759), .A2(n9764), .B1(n9719), .B2(n9757), .ZN(
        P1_U3466) );
  OAI211_X1 U10872 ( .C1(n9722), .C2(n9742), .A(n9721), .B(n9720), .ZN(n9724)
         );
  AOI211_X1 U10873 ( .C1(n9755), .C2(n9725), .A(n9724), .B(n9723), .ZN(n9765)
         );
  INV_X1 U10874 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U10875 ( .A1(n9759), .A2(n9765), .B1(n10195), .B2(n9757), .ZN(
        P1_U3469) );
  AOI22_X1 U10876 ( .A1(n9729), .A2(n9728), .B1(n9727), .B2(n9726), .ZN(n9730)
         );
  OAI211_X1 U10877 ( .C1(n9740), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9733)
         );
  INV_X1 U10878 ( .A(n9733), .ZN(n9766) );
  INV_X1 U10879 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9734) );
  AOI22_X1 U10880 ( .A1(n9759), .A2(n9766), .B1(n9734), .B2(n9757), .ZN(
        P1_U3472) );
  OAI21_X1 U10881 ( .B1(n9736), .B2(n9742), .A(n9735), .ZN(n9738) );
  AOI211_X1 U10882 ( .C1(n9755), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9767)
         );
  INV_X1 U10883 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U10884 ( .A1(n9759), .A2(n9767), .B1(n10217), .B2(n9757), .ZN(
        P1_U3475) );
  NOR2_X1 U10885 ( .A1(n9741), .A2(n9740), .ZN(n9748) );
  OAI22_X1 U10886 ( .A1(n9744), .A2(n9753), .B1(n9743), .B2(n9742), .ZN(n9746)
         );
  AOI211_X1 U10887 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9769)
         );
  INV_X1 U10888 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U10889 ( .A1(n9759), .A2(n9769), .B1(n10085), .B2(n9757), .ZN(
        P1_U3478) );
  INV_X1 U10890 ( .A(n9749), .ZN(n9750) );
  OAI211_X1 U10891 ( .C1(n9753), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9754)
         );
  AOI21_X1 U10892 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9771) );
  INV_X1 U10893 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U10894 ( .A1(n9759), .A2(n9771), .B1(n9758), .B2(n9757), .ZN(
        P1_U3481) );
  INV_X1 U10895 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9760) );
  AOI22_X1 U10896 ( .A1(n9772), .A2(n9761), .B1(n9760), .B2(n9770), .ZN(
        P1_U3524) );
  INV_X1 U10897 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9762) );
  AOI22_X1 U10898 ( .A1(n9772), .A2(n9763), .B1(n9762), .B2(n9770), .ZN(
        P1_U3526) );
  AOI22_X1 U10899 ( .A1(n9772), .A2(n9764), .B1(n6701), .B2(n9770), .ZN(
        P1_U3527) );
  AOI22_X1 U10900 ( .A1(n9772), .A2(n9765), .B1(n6702), .B2(n9770), .ZN(
        P1_U3528) );
  AOI22_X1 U10901 ( .A1(n9772), .A2(n9766), .B1(n10012), .B2(n9770), .ZN(
        P1_U3529) );
  AOI22_X1 U10902 ( .A1(n9772), .A2(n9767), .B1(n6745), .B2(n9770), .ZN(
        P1_U3530) );
  INV_X1 U10903 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10904 ( .A1(n9772), .A2(n9769), .B1(n9768), .B2(n9770), .ZN(
        P1_U3531) );
  AOI22_X1 U10905 ( .A1(n9772), .A2(n9771), .B1(n5272), .B2(n9770), .ZN(
        P1_U3532) );
  AOI22_X1 U10906 ( .A1(n9774), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9773), .ZN(n9783) );
  AOI22_X1 U10907 ( .A1(n9775), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9782) );
  NOR2_X1 U10908 ( .A1(n9776), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9780) );
  OAI21_X1 U10909 ( .B1(n9778), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9777), .ZN(
        n9779) );
  OAI21_X1 U10910 ( .B1(n9780), .B2(n9779), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9781) );
  OAI211_X1 U10911 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9783), .A(n9782), .B(
        n9781), .ZN(P2_U3245) );
  XOR2_X1 U10912 ( .A(n9803), .B(n9784), .Z(n9789) );
  AOI222_X1 U10913 ( .A1(n9790), .A2(n9789), .B1(n9788), .B2(n9787), .C1(n4402), .C2(n9785), .ZN(n9862) );
  OAI22_X1 U10914 ( .A1(n9793), .A2(n9792), .B1(n6796), .B2(n9791), .ZN(n9794)
         );
  INV_X1 U10915 ( .A(n9794), .ZN(n9807) );
  NAND2_X1 U10916 ( .A1(n9795), .A2(n9799), .ZN(n9796) );
  NAND2_X1 U10917 ( .A1(n9796), .A2(n9883), .ZN(n9798) );
  OR2_X1 U10918 ( .A1(n9798), .A2(n9797), .ZN(n9801) );
  NAND2_X1 U10919 ( .A1(n9799), .A2(n9882), .ZN(n9800) );
  NAND2_X1 U10920 ( .A1(n9801), .A2(n9800), .ZN(n9864) );
  XNOR2_X1 U10921 ( .A(n9802), .B(n9803), .ZN(n9865) );
  AOI22_X1 U10922 ( .A1(n9805), .A2(n9864), .B1(n9804), .B2(n9865), .ZN(n9806)
         );
  OAI211_X1 U10923 ( .C1(n9808), .C2(n9862), .A(n9807), .B(n9806), .ZN(
        P2_U3292) );
  NOR2_X1 U10924 ( .A1(n9835), .A2(n10039), .ZN(P2_U3297) );
  INV_X1 U10925 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U10926 ( .A1(n9835), .A2(n9811), .ZN(P2_U3298) );
  INV_X1 U10927 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U10928 ( .A1(n9835), .A2(n9812), .ZN(P2_U3299) );
  NOR2_X1 U10929 ( .A1(n9835), .A2(n10138), .ZN(P2_U3300) );
  INV_X1 U10930 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10931 ( .A1(n9820), .A2(n9813), .ZN(P2_U3301) );
  INV_X1 U10932 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U10933 ( .A1(n9820), .A2(n9814), .ZN(P2_U3302) );
  INV_X1 U10934 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U10935 ( .A1(n9820), .A2(n9815), .ZN(P2_U3303) );
  INV_X1 U10936 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U10937 ( .A1(n9820), .A2(n9816), .ZN(P2_U3304) );
  INV_X1 U10938 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U10939 ( .A1(n9820), .A2(n10030), .ZN(P2_U3305) );
  INV_X1 U10940 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U10941 ( .A1(n9820), .A2(n10047), .ZN(P2_U3306) );
  INV_X1 U10942 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U10943 ( .A1(n9820), .A2(n10183), .ZN(P2_U3307) );
  INV_X1 U10944 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U10945 ( .A1(n9820), .A2(n9817), .ZN(P2_U3308) );
  INV_X1 U10946 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U10947 ( .A1(n9820), .A2(n9818), .ZN(P2_U3309) );
  INV_X1 U10948 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U10949 ( .A1(n9820), .A2(n9819), .ZN(P2_U3310) );
  INV_X1 U10950 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U10951 ( .A1(n9835), .A2(n9821), .ZN(P2_U3311) );
  INV_X1 U10952 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U10953 ( .A1(n9835), .A2(n9822), .ZN(P2_U3312) );
  INV_X1 U10954 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10139) );
  NOR2_X1 U10955 ( .A1(n9835), .A2(n10139), .ZN(P2_U3313) );
  INV_X1 U10956 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U10957 ( .A1(n9835), .A2(n9823), .ZN(P2_U3314) );
  INV_X1 U10958 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U10959 ( .A1(n9835), .A2(n9824), .ZN(P2_U3315) );
  INV_X1 U10960 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U10961 ( .A1(n9835), .A2(n9825), .ZN(P2_U3316) );
  INV_X1 U10962 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U10963 ( .A1(n9835), .A2(n9826), .ZN(P2_U3317) );
  INV_X1 U10964 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U10965 ( .A1(n9835), .A2(n9827), .ZN(P2_U3318) );
  NOR2_X1 U10966 ( .A1(n9835), .A2(n10144), .ZN(P2_U3319) );
  NOR2_X1 U10967 ( .A1(n9835), .A2(n9968), .ZN(P2_U3320) );
  INV_X1 U10968 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9991) );
  NOR2_X1 U10969 ( .A1(n9835), .A2(n9991), .ZN(P2_U3321) );
  INV_X1 U10970 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U10971 ( .A1(n9835), .A2(n9828), .ZN(P2_U3322) );
  INV_X1 U10972 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U10973 ( .A1(n9835), .A2(n9829), .ZN(P2_U3323) );
  INV_X1 U10974 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9980) );
  NOR2_X1 U10975 ( .A1(n9835), .A2(n9980), .ZN(P2_U3324) );
  INV_X1 U10976 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U10977 ( .A1(n9835), .A2(n10057), .ZN(P2_U3325) );
  INV_X1 U10978 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U10979 ( .A1(n9835), .A2(n9830), .ZN(P2_U3326) );
  OAI22_X1 U10980 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9835), .B1(n9831), .B2(
        n9833), .ZN(n9832) );
  INV_X1 U10981 ( .A(n9832), .ZN(P2_U3437) );
  OAI22_X1 U10982 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9835), .B1(n9834), .B2(
        n9833), .ZN(n9836) );
  INV_X1 U10983 ( .A(n9836), .ZN(P2_U3438) );
  AOI22_X1 U10984 ( .A1(n9838), .A2(n9904), .B1(n6399), .B2(n9837), .ZN(n9839)
         );
  AND2_X1 U10985 ( .A1(n9840), .A2(n9839), .ZN(n9909) );
  INV_X1 U10986 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U10987 ( .A1(n9908), .A2(n9909), .B1(n10197), .B2(n9906), .ZN(
        P2_U3451) );
  NOR3_X1 U10988 ( .A1(n9842), .A2(n9841), .A3(n9900), .ZN(n9843) );
  AOI21_X1 U10989 ( .B1(n9882), .B2(n9844), .A(n9843), .ZN(n9845) );
  OAI211_X1 U10990 ( .C1(n9871), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9848)
         );
  INV_X1 U10991 ( .A(n9848), .ZN(n9910) );
  INV_X1 U10992 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U10993 ( .A1(n9908), .A2(n9910), .B1(n10203), .B2(n9906), .ZN(
        P2_U3454) );
  OAI211_X1 U10994 ( .C1(n9851), .C2(n9899), .A(n9850), .B(n9849), .ZN(n9852)
         );
  AOI21_X1 U10995 ( .B1(n9904), .B2(n9853), .A(n9852), .ZN(n9912) );
  INV_X1 U10996 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10997 ( .A1(n9908), .A2(n9912), .B1(n9854), .B2(n9906), .ZN(
        P2_U3457) );
  AOI22_X1 U10998 ( .A1(n9856), .A2(n9883), .B1(n9882), .B2(n9855), .ZN(n9857)
         );
  OAI211_X1 U10999 ( .C1(n9859), .C2(n9890), .A(n9858), .B(n9857), .ZN(n9860)
         );
  INV_X1 U11000 ( .A(n9860), .ZN(n9914) );
  INV_X1 U11001 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U11002 ( .A1(n9908), .A2(n9914), .B1(n9861), .B2(n9906), .ZN(
        P2_U3460) );
  INV_X1 U11003 ( .A(n9862), .ZN(n9863) );
  AOI211_X1 U11004 ( .C1(n9904), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9916)
         );
  INV_X1 U11005 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9866) );
  AOI22_X1 U11006 ( .A1(n9908), .A2(n9916), .B1(n9866), .B2(n9906), .ZN(
        P2_U3463) );
  AOI211_X1 U11007 ( .C1(n9882), .C2(n4821), .A(n9868), .B(n9867), .ZN(n9869)
         );
  OAI21_X1 U11008 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9872) );
  INV_X1 U11009 ( .A(n9872), .ZN(n9918) );
  INV_X1 U11010 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9873) );
  AOI22_X1 U11011 ( .A1(n9908), .A2(n9918), .B1(n9873), .B2(n9906), .ZN(
        P2_U3466) );
  AND2_X1 U11012 ( .A1(n9874), .A2(n9904), .ZN(n9880) );
  NAND2_X1 U11013 ( .A1(n9875), .A2(n9883), .ZN(n9876) );
  OAI21_X1 U11014 ( .B1(n9877), .B2(n9899), .A(n9876), .ZN(n9878) );
  NOR3_X1 U11015 ( .A1(n9880), .A2(n9879), .A3(n9878), .ZN(n9919) );
  INV_X1 U11016 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11017 ( .A1(n9908), .A2(n9919), .B1(n9959), .B2(n9906), .ZN(
        P2_U3469) );
  AOI22_X1 U11018 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9881), .ZN(n9885)
         );
  OAI21_X1 U11019 ( .B1(n9886), .B2(n9890), .A(n9885), .ZN(n9887) );
  NOR2_X1 U11020 ( .A1(n9888), .A2(n9887), .ZN(n9920) );
  INV_X1 U11021 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U11022 ( .A1(n9908), .A2(n9920), .B1(n9889), .B2(n9906), .ZN(
        P2_U3475) );
  INV_X1 U11023 ( .A(n9890), .ZN(n9897) );
  INV_X1 U11024 ( .A(n9891), .ZN(n9896) );
  OAI22_X1 U11025 ( .A1(n9893), .A2(n9900), .B1(n9892), .B2(n9899), .ZN(n9895)
         );
  AOI211_X1 U11026 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9921)
         );
  INV_X1 U11027 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U11028 ( .A1(n9908), .A2(n9921), .B1(n9898), .B2(n9906), .ZN(
        P2_U3481) );
  OAI22_X1 U11029 ( .A1(n9901), .A2(n9900), .B1(n4806), .B2(n9899), .ZN(n9903)
         );
  AOI211_X1 U11030 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9923)
         );
  INV_X1 U11031 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U11032 ( .A1(n9908), .A2(n9923), .B1(n9907), .B2(n9906), .ZN(
        P2_U3487) );
  INV_X1 U11033 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U11034 ( .A1(n9924), .A2(n9909), .B1(n10186), .B2(n9922), .ZN(
        P2_U3520) );
  AOI22_X1 U11035 ( .A1(n9924), .A2(n9910), .B1(n6769), .B2(n9922), .ZN(
        P2_U3521) );
  INV_X1 U11036 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U11037 ( .A1(n9924), .A2(n9912), .B1(n9911), .B2(n9922), .ZN(
        P2_U3522) );
  INV_X1 U11038 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U11039 ( .A1(n9924), .A2(n9914), .B1(n9913), .B2(n9922), .ZN(
        P2_U3523) );
  INV_X1 U11040 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U11041 ( .A1(n9924), .A2(n9916), .B1(n9915), .B2(n9922), .ZN(
        P2_U3524) );
  INV_X1 U11042 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U11043 ( .A1(n9924), .A2(n9918), .B1(n9917), .B2(n9922), .ZN(
        P2_U3525) );
  AOI22_X1 U11044 ( .A1(n9924), .A2(n9919), .B1(n6774), .B2(n9922), .ZN(
        P2_U3526) );
  AOI22_X1 U11045 ( .A1(n9924), .A2(n9920), .B1(n6777), .B2(n9922), .ZN(
        P2_U3528) );
  AOI22_X1 U11046 ( .A1(n9924), .A2(n9921), .B1(n7126), .B2(n9922), .ZN(
        P2_U3530) );
  AOI22_X1 U11047 ( .A1(n9924), .A2(n9923), .B1(n7512), .B2(n9922), .ZN(
        P2_U3532) );
  INV_X1 U11048 ( .A(n9925), .ZN(n9926) );
  NAND2_X1 U11049 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  XNOR2_X1 U11050 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9928), .ZN(ADD_1071_U5) );
  XOR2_X1 U11051 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11052 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(ADD_1071_U56) );
  OAI21_X1 U11053 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(ADD_1071_U57) );
  OAI21_X1 U11054 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(ADD_1071_U58) );
  AOI21_X1 U11055 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(ADD_1071_U59) );
  OAI21_X1 U11056 ( .B1(n9943), .B2(n9942), .A(n9941), .ZN(ADD_1071_U60) );
  OAI21_X1 U11057 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(ADD_1071_U61) );
  AOI21_X1 U11058 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(ADD_1071_U62) );
  AOI21_X1 U11059 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(ADD_1071_U63) );
  AOI22_X1 U11060 ( .A1(n10216), .A2(keyinput93), .B1(n9954), .B2(keyinput111), 
        .ZN(n9953) );
  OAI221_X1 U11061 ( .B1(n10216), .B2(keyinput93), .C1(n9954), .C2(keyinput111), .A(n9953), .ZN(n9965) );
  AOI22_X1 U11062 ( .A1(n9956), .A2(keyinput80), .B1(keyinput67), .B2(n10217), 
        .ZN(n9955) );
  OAI221_X1 U11063 ( .B1(n9956), .B2(keyinput80), .C1(n10217), .C2(keyinput67), 
        .A(n9955), .ZN(n9964) );
  AOI22_X1 U11064 ( .A1(n9959), .A2(keyinput34), .B1(n9958), .B2(keyinput70), 
        .ZN(n9957) );
  OAI221_X1 U11065 ( .B1(n9959), .B2(keyinput34), .C1(n9958), .C2(keyinput70), 
        .A(n9957), .ZN(n9963) );
  XOR2_X1 U11066 ( .A(n5024), .B(keyinput102), .Z(n9961) );
  XNOR2_X1 U11067 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput54), .ZN(n9960) );
  NAND2_X1 U11068 ( .A1(n9961), .A2(n9960), .ZN(n9962) );
  NOR4_X1 U11069 ( .A1(n9965), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(n10005)
         );
  INV_X1 U11070 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U11071 ( .A1(n10215), .A2(keyinput75), .B1(n5059), .B2(keyinput124), 
        .ZN(n9966) );
  OAI221_X1 U11072 ( .B1(n10215), .B2(keyinput75), .C1(n5059), .C2(keyinput124), .A(n9966), .ZN(n9977) );
  AOI22_X1 U11073 ( .A1(n9968), .A2(keyinput49), .B1(n10214), .B2(keyinput29), 
        .ZN(n9967) );
  OAI221_X1 U11074 ( .B1(n9968), .B2(keyinput49), .C1(n10214), .C2(keyinput29), 
        .A(n9967), .ZN(n9976) );
  AOI22_X1 U11075 ( .A1(n9971), .A2(keyinput103), .B1(n9970), .B2(keyinput26), 
        .ZN(n9969) );
  OAI221_X1 U11076 ( .B1(n9971), .B2(keyinput103), .C1(n9970), .C2(keyinput26), 
        .A(n9969), .ZN(n9975) );
  INV_X1 U11077 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11078 ( .A1(n10220), .A2(keyinput23), .B1(n9973), .B2(keyinput84), 
        .ZN(n9972) );
  OAI221_X1 U11079 ( .B1(n10220), .B2(keyinput23), .C1(n9973), .C2(keyinput84), 
        .A(n9972), .ZN(n9974) );
  NOR4_X1 U11080 ( .A1(n9977), .A2(n9976), .A3(n9975), .A4(n9974), .ZN(n10004)
         );
  AOI22_X1 U11081 ( .A1(n9980), .A2(keyinput113), .B1(n9979), .B2(keyinput76), 
        .ZN(n9978) );
  OAI221_X1 U11082 ( .B1(n9980), .B2(keyinput113), .C1(n9979), .C2(keyinput76), 
        .A(n9978), .ZN(n9989) );
  AOI22_X1 U11083 ( .A1(n6788), .A2(keyinput56), .B1(n10219), .B2(keyinput28), 
        .ZN(n9981) );
  OAI221_X1 U11084 ( .B1(n6788), .B2(keyinput56), .C1(n10219), .C2(keyinput28), 
        .A(n9981), .ZN(n9988) );
  AOI22_X1 U11085 ( .A1(n10218), .A2(keyinput95), .B1(keyinput97), .B2(n9983), 
        .ZN(n9982) );
  OAI221_X1 U11086 ( .B1(n10218), .B2(keyinput95), .C1(n9983), .C2(keyinput97), 
        .A(n9982), .ZN(n9987) );
  INV_X1 U11087 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9985) );
  INV_X1 U11088 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11089 ( .A1(n9985), .A2(keyinput39), .B1(keyinput96), .B2(n10266), 
        .ZN(n9984) );
  OAI221_X1 U11090 ( .B1(n9985), .B2(keyinput39), .C1(n10266), .C2(keyinput96), 
        .A(n9984), .ZN(n9986) );
  NOR4_X1 U11091 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n10003)
         );
  AOI22_X1 U11092 ( .A1(n10205), .A2(keyinput107), .B1(keyinput110), .B2(n9991), .ZN(n9990) );
  OAI221_X1 U11093 ( .B1(n10205), .B2(keyinput107), .C1(n9991), .C2(
        keyinput110), .A(n9990), .ZN(n10001) );
  INV_X1 U11094 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11095 ( .A1(n9994), .A2(keyinput35), .B1(n9993), .B2(keyinput30), 
        .ZN(n9992) );
  OAI221_X1 U11096 ( .B1(n9994), .B2(keyinput35), .C1(n9993), .C2(keyinput30), 
        .A(n9992), .ZN(n10000) );
  XNOR2_X1 U11097 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput25), .ZN(n9998) );
  XNOR2_X1 U11098 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput115), .ZN(n9997) );
  XNOR2_X1 U11099 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput83), .ZN(n9996) );
  XNOR2_X1 U11100 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput123), .ZN(n9995) );
  NAND4_X1 U11101 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n9999)
         );
  NOR3_X1 U11102 ( .A1(n10001), .A2(n10000), .A3(n9999), .ZN(n10002) );
  NAND4_X1 U11103 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n10164) );
  INV_X1 U11104 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U11105 ( .A1(n10168), .A2(keyinput81), .B1(n10007), .B2(keyinput121), .ZN(n10006) );
  OAI221_X1 U11106 ( .B1(n10168), .B2(keyinput81), .C1(n10007), .C2(
        keyinput121), .A(n10006), .ZN(n10016) );
  AOI22_X1 U11107 ( .A1(n10251), .A2(keyinput48), .B1(keyinput12), .B2(n6754), 
        .ZN(n10008) );
  OAI221_X1 U11108 ( .B1(n10251), .B2(keyinput48), .C1(n6754), .C2(keyinput12), 
        .A(n10008), .ZN(n10015) );
  AOI22_X1 U11109 ( .A1(n10206), .A2(keyinput58), .B1(keyinput11), .B2(n7926), 
        .ZN(n10009) );
  OAI221_X1 U11110 ( .B1(n10206), .B2(keyinput58), .C1(n7926), .C2(keyinput11), 
        .A(n10009), .ZN(n10014) );
  AOI22_X1 U11111 ( .A1(n10012), .A2(keyinput6), .B1(n10011), .B2(keyinput8), 
        .ZN(n10010) );
  OAI221_X1 U11112 ( .B1(n10012), .B2(keyinput6), .C1(n10011), .C2(keyinput8), 
        .A(n10010), .ZN(n10013) );
  NOR4_X1 U11113 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10055) );
  AOI22_X1 U11114 ( .A1(n6335), .A2(keyinput4), .B1(n6709), .B2(keyinput0), 
        .ZN(n10017) );
  OAI221_X1 U11115 ( .B1(n6335), .B2(keyinput4), .C1(n6709), .C2(keyinput0), 
        .A(n10017), .ZN(n10026) );
  INV_X1 U11116 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U11117 ( .A1(n10203), .A2(keyinput122), .B1(keyinput106), .B2(
        n10173), .ZN(n10018) );
  OAI221_X1 U11118 ( .B1(n10203), .B2(keyinput122), .C1(n10173), .C2(
        keyinput106), .A(n10018), .ZN(n10025) );
  AOI22_X1 U11119 ( .A1(n10204), .A2(keyinput78), .B1(n10020), .B2(keyinput38), 
        .ZN(n10019) );
  OAI221_X1 U11120 ( .B1(n10204), .B2(keyinput78), .C1(n10020), .C2(keyinput38), .A(n10019), .ZN(n10024) );
  AOI22_X1 U11121 ( .A1(n10022), .A2(keyinput50), .B1(keyinput22), .B2(n10176), 
        .ZN(n10021) );
  OAI221_X1 U11122 ( .B1(n10022), .B2(keyinput50), .C1(n10176), .C2(keyinput22), .A(n10021), .ZN(n10023) );
  NOR4_X1 U11123 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10054) );
  AOI22_X1 U11124 ( .A1(n5317), .A2(keyinput105), .B1(keyinput1), .B2(n6956), 
        .ZN(n10027) );
  OAI221_X1 U11125 ( .B1(n5317), .B2(keyinput105), .C1(n6956), .C2(keyinput1), 
        .A(n10027), .ZN(n10037) );
  AOI22_X1 U11126 ( .A1(n5091), .A2(keyinput104), .B1(keyinput61), .B2(n8270), 
        .ZN(n10028) );
  OAI221_X1 U11127 ( .B1(n5091), .B2(keyinput104), .C1(n8270), .C2(keyinput61), 
        .A(n10028), .ZN(n10036) );
  AOI22_X1 U11128 ( .A1(n10031), .A2(keyinput89), .B1(keyinput51), .B2(n10030), 
        .ZN(n10029) );
  OAI221_X1 U11129 ( .B1(n10031), .B2(keyinput89), .C1(n10030), .C2(keyinput51), .A(n10029), .ZN(n10035) );
  XNOR2_X1 U11130 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput44), .ZN(n10033)
         );
  XNOR2_X1 U11131 ( .A(P1_REG3_REG_3__SCAN_IN), .B(keyinput2), .ZN(n10032) );
  NAND2_X1 U11132 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  NOR4_X1 U11133 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10053) );
  AOI22_X1 U11134 ( .A1(n5781), .A2(keyinput21), .B1(n10039), .B2(keyinput116), 
        .ZN(n10038) );
  OAI221_X1 U11135 ( .B1(n5781), .B2(keyinput21), .C1(n10039), .C2(keyinput116), .A(n10038), .ZN(n10051) );
  INV_X1 U11136 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10042) );
  INV_X1 U11137 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11138 ( .A1(n10042), .A2(keyinput9), .B1(keyinput32), .B2(n10041), 
        .ZN(n10040) );
  OAI221_X1 U11139 ( .B1(n10042), .B2(keyinput9), .C1(n10041), .C2(keyinput32), 
        .A(n10040), .ZN(n10050) );
  INV_X1 U11140 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11141 ( .A1(n10234), .A2(keyinput118), .B1(keyinput14), .B2(n10044), .ZN(n10043) );
  OAI221_X1 U11142 ( .B1(n10234), .B2(keyinput118), .C1(n10044), .C2(
        keyinput14), .A(n10043), .ZN(n10049) );
  INV_X1 U11143 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11144 ( .A1(n10047), .A2(keyinput24), .B1(keyinput33), .B2(n10046), 
        .ZN(n10045) );
  OAI221_X1 U11145 ( .B1(n10047), .B2(keyinput24), .C1(n10046), .C2(keyinput33), .A(n10045), .ZN(n10048) );
  NOR4_X1 U11146 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10052) );
  NAND4_X1 U11147 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10163) );
  AOI22_X1 U11148 ( .A1(n7673), .A2(keyinput87), .B1(keyinput27), .B2(n10057), 
        .ZN(n10056) );
  OAI221_X1 U11149 ( .B1(n7673), .B2(keyinput87), .C1(n10057), .C2(keyinput27), 
        .A(n10056), .ZN(n10065) );
  AOI22_X1 U11150 ( .A1(n10225), .A2(keyinput72), .B1(n5070), .B2(keyinput101), 
        .ZN(n10058) );
  OAI221_X1 U11151 ( .B1(n10225), .B2(keyinput72), .C1(n5070), .C2(keyinput101), .A(n10058), .ZN(n10064) );
  XNOR2_X1 U11152 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput90), .ZN(n10062)
         );
  XNOR2_X1 U11153 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput68), .ZN(n10061) );
  XNOR2_X1 U11154 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput88), .ZN(n10060) );
  XNOR2_X1 U11155 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput126), .ZN(n10059) );
  NAND4_X1 U11156 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10063) );
  NOR3_X1 U11157 ( .A1(n10065), .A2(n10064), .A3(n10063), .ZN(n10107) );
  AOI22_X1 U11158 ( .A1(n10067), .A2(keyinput98), .B1(keyinput100), .B2(n10226), .ZN(n10066) );
  OAI221_X1 U11159 ( .B1(n10067), .B2(keyinput98), .C1(n10226), .C2(
        keyinput100), .A(n10066), .ZN(n10080) );
  AOI22_X1 U11160 ( .A1(n10070), .A2(keyinput125), .B1(keyinput46), .B2(n10069), .ZN(n10068) );
  OAI221_X1 U11161 ( .B1(n10070), .B2(keyinput125), .C1(n10069), .C2(
        keyinput46), .A(n10068), .ZN(n10079) );
  INV_X1 U11162 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10073) );
  INV_X1 U11163 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U11164 ( .A1(n10073), .A2(keyinput62), .B1(keyinput64), .B2(n10072), 
        .ZN(n10071) );
  OAI221_X1 U11165 ( .B1(n10073), .B2(keyinput62), .C1(n10072), .C2(keyinput64), .A(n10071), .ZN(n10078) );
  AOI22_X1 U11166 ( .A1(n10076), .A2(keyinput82), .B1(keyinput109), .B2(n10075), .ZN(n10074) );
  OAI221_X1 U11167 ( .B1(n10076), .B2(keyinput82), .C1(n10075), .C2(
        keyinput109), .A(n10074), .ZN(n10077) );
  NOR4_X1 U11168 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10106) );
  AOI22_X1 U11169 ( .A1(n10083), .A2(keyinput15), .B1(n10082), .B2(keyinput71), 
        .ZN(n10081) );
  OAI221_X1 U11170 ( .B1(n10083), .B2(keyinput15), .C1(n10082), .C2(keyinput71), .A(n10081), .ZN(n10093) );
  AOI22_X1 U11171 ( .A1(n10228), .A2(keyinput85), .B1(keyinput120), .B2(n10085), .ZN(n10084) );
  OAI221_X1 U11172 ( .B1(n10228), .B2(keyinput85), .C1(n10085), .C2(
        keyinput120), .A(n10084), .ZN(n10092) );
  INV_X1 U11173 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U11174 ( .A1(n10165), .A2(keyinput60), .B1(n4988), .B2(keyinput42), 
        .ZN(n10086) );
  OAI221_X1 U11175 ( .B1(n10165), .B2(keyinput60), .C1(n4988), .C2(keyinput42), 
        .A(n10086), .ZN(n10091) );
  INV_X1 U11176 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11177 ( .A1(n10089), .A2(keyinput45), .B1(n10088), .B2(keyinput55), 
        .ZN(n10087) );
  OAI221_X1 U11178 ( .B1(n10089), .B2(keyinput45), .C1(n10088), .C2(keyinput55), .A(n10087), .ZN(n10090) );
  NOR4_X1 U11179 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n10105) );
  AOI22_X1 U11180 ( .A1(n10227), .A2(keyinput41), .B1(n10095), .B2(keyinput43), 
        .ZN(n10094) );
  OAI221_X1 U11181 ( .B1(n10227), .B2(keyinput41), .C1(n10095), .C2(keyinput43), .A(n10094), .ZN(n10103) );
  INV_X1 U11182 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U11183 ( .A1(n10177), .A2(keyinput3), .B1(keyinput74), .B2(n10195), 
        .ZN(n10096) );
  OAI221_X1 U11184 ( .B1(n10177), .B2(keyinput3), .C1(n10195), .C2(keyinput74), 
        .A(n10096), .ZN(n10102) );
  AOI22_X1 U11185 ( .A1(n5691), .A2(keyinput127), .B1(keyinput77), .B2(n6796), 
        .ZN(n10097) );
  OAI221_X1 U11186 ( .B1(n5691), .B2(keyinput127), .C1(n6796), .C2(keyinput77), 
        .A(n10097), .ZN(n10101) );
  AOI22_X1 U11187 ( .A1(n10099), .A2(keyinput19), .B1(keyinput18), .B2(n10194), 
        .ZN(n10098) );
  OAI221_X1 U11188 ( .B1(n10099), .B2(keyinput19), .C1(n10194), .C2(keyinput18), .A(n10098), .ZN(n10100) );
  NOR4_X1 U11189 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10104) );
  NAND4_X1 U11190 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n10162) );
  INV_X1 U11191 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11192 ( .A1(n10193), .A2(keyinput16), .B1(keyinput40), .B2(n7539), 
        .ZN(n10108) );
  OAI221_X1 U11193 ( .B1(n10193), .B2(keyinput16), .C1(n7539), .C2(keyinput40), 
        .A(n10108), .ZN(n10117) );
  AOI22_X1 U11194 ( .A1(n10110), .A2(keyinput63), .B1(n6702), .B2(keyinput47), 
        .ZN(n10109) );
  OAI221_X1 U11195 ( .B1(n10110), .B2(keyinput63), .C1(n6702), .C2(keyinput47), 
        .A(n10109), .ZN(n10116) );
  AOI22_X1 U11196 ( .A1(n6769), .A2(keyinput108), .B1(n10112), .B2(keyinput69), 
        .ZN(n10111) );
  OAI221_X1 U11197 ( .B1(n6769), .B2(keyinput108), .C1(n10112), .C2(keyinput69), .A(n10111), .ZN(n10115) );
  AOI22_X1 U11198 ( .A1(n10198), .A2(keyinput86), .B1(n6062), .B2(keyinput117), 
        .ZN(n10113) );
  OAI221_X1 U11199 ( .B1(n10198), .B2(keyinput86), .C1(n6062), .C2(keyinput117), .A(n10113), .ZN(n10114) );
  NOR4_X1 U11200 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10160) );
  AOI22_X1 U11201 ( .A1(n10196), .A2(keyinput53), .B1(keyinput37), .B2(n10197), 
        .ZN(n10118) );
  OAI221_X1 U11202 ( .B1(n10196), .B2(keyinput53), .C1(n10197), .C2(keyinput37), .A(n10118), .ZN(n10130) );
  AOI22_X1 U11203 ( .A1(n10121), .A2(keyinput79), .B1(n10120), .B2(keyinput5), 
        .ZN(n10119) );
  OAI221_X1 U11204 ( .B1(n10121), .B2(keyinput79), .C1(n10120), .C2(keyinput5), 
        .A(n10119), .ZN(n10129) );
  AOI22_X1 U11205 ( .A1(n10124), .A2(keyinput73), .B1(n10123), .B2(keyinput13), 
        .ZN(n10122) );
  OAI221_X1 U11206 ( .B1(n10124), .B2(keyinput73), .C1(n10123), .C2(keyinput13), .A(n10122), .ZN(n10128) );
  AOI22_X1 U11207 ( .A1(n10186), .A2(keyinput112), .B1(n10126), .B2(
        keyinput119), .ZN(n10125) );
  OAI221_X1 U11208 ( .B1(n10186), .B2(keyinput112), .C1(n10126), .C2(
        keyinput119), .A(n10125), .ZN(n10127) );
  NOR4_X1 U11209 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10159) );
  AOI22_X1 U11210 ( .A1(n10183), .A2(keyinput92), .B1(n10185), .B2(keyinput59), 
        .ZN(n10131) );
  OAI221_X1 U11211 ( .B1(n10183), .B2(keyinput92), .C1(n10185), .C2(keyinput59), .A(n10131), .ZN(n10134) );
  XNOR2_X1 U11212 ( .A(n10184), .B(keyinput17), .ZN(n10133) );
  XNOR2_X1 U11213 ( .A(n5019), .B(keyinput94), .ZN(n10132) );
  OR3_X1 U11214 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n10142) );
  AOI22_X1 U11215 ( .A1(n10136), .A2(keyinput10), .B1(keyinput52), .B2(n10172), 
        .ZN(n10135) );
  OAI221_X1 U11216 ( .B1(n10136), .B2(keyinput10), .C1(n10172), .C2(keyinput52), .A(n10135), .ZN(n10141) );
  AOI22_X1 U11217 ( .A1(n10139), .A2(keyinput31), .B1(n10138), .B2(keyinput36), 
        .ZN(n10137) );
  OAI221_X1 U11218 ( .B1(n10139), .B2(keyinput31), .C1(n10138), .C2(keyinput36), .A(n10137), .ZN(n10140) );
  NOR3_X1 U11219 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(n10158) );
  AOI22_X1 U11220 ( .A1(n10145), .A2(keyinput20), .B1(n10144), .B2(keyinput65), 
        .ZN(n10143) );
  OAI221_X1 U11221 ( .B1(n10145), .B2(keyinput20), .C1(n10144), .C2(keyinput65), .A(n10143), .ZN(n10156) );
  INV_X1 U11222 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U11223 ( .A1(n10188), .A2(keyinput99), .B1(keyinput114), .B2(n10147), .ZN(n10146) );
  OAI221_X1 U11224 ( .B1(n10188), .B2(keyinput99), .C1(n10147), .C2(
        keyinput114), .A(n10146), .ZN(n10155) );
  AOI22_X1 U11225 ( .A1(n10187), .A2(keyinput91), .B1(n10149), .B2(keyinput7), 
        .ZN(n10148) );
  OAI221_X1 U11226 ( .B1(n10187), .B2(keyinput91), .C1(n10149), .C2(keyinput7), 
        .A(n10148), .ZN(n10154) );
  AOI22_X1 U11227 ( .A1(n10152), .A2(keyinput66), .B1(keyinput57), .B2(n10151), 
        .ZN(n10150) );
  OAI221_X1 U11228 ( .B1(n10152), .B2(keyinput66), .C1(n10151), .C2(keyinput57), .A(n10150), .ZN(n10153) );
  NOR4_X1 U11229 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n10157) );
  NAND4_X1 U11230 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10161) );
  NOR4_X1 U11231 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10249) );
  NAND4_X1 U11232 ( .A1(n10167), .A2(n10166), .A3(P2_ADDR_REG_8__SCAN_IN), 
        .A4(n10165), .ZN(n10171) );
  NOR4_X1 U11233 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .A3(P1_ADDR_REG_7__SCAN_IN), .A4(n10168), .ZN(n10169) );
  NAND3_X1 U11234 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .A3(n10169), .ZN(n10170) );
  NOR4_X1 U11235 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), 
        .A3(n10171), .A4(n10170), .ZN(n10182) );
  NAND2_X1 U11236 ( .A1(n10173), .A2(n10172), .ZN(n10174) );
  NOR4_X1 U11237 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        n10175), .A4(n10174), .ZN(n10181) );
  NOR4_X1 U11238 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P2_DATAO_REG_24__SCAN_IN), 
        .A3(P2_REG0_REG_6__SCAN_IN), .A4(n10176), .ZN(n10178) );
  NAND3_X1 U11239 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(n10178), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n10179) );
  NOR3_X1 U11240 ( .A1(n10179), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_21__SCAN_IN), .ZN(n10180) );
  NAND3_X1 U11241 ( .A1(n10182), .A2(n10181), .A3(n10180), .ZN(n10247) );
  NOR4_X1 U11242 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n10185), .A3(n10184), 
        .A4(n10183), .ZN(n10192) );
  NOR4_X1 U11243 ( .A1(P1_D_REG_7__SCAN_IN), .A2(SI_10_), .A3(
        P1_DATAO_REG_0__SCAN_IN), .A4(n10186), .ZN(n10191) );
  NOR4_X1 U11244 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG2_REG_8__SCAN_IN), 
        .A3(P1_DATAO_REG_31__SCAN_IN), .A4(n10187), .ZN(n10190) );
  NOR4_X1 U11245 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(P1_REG1_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_15__SCAN_IN), .A4(n10188), .ZN(n10189) );
  NAND4_X1 U11246 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10246) );
  NOR4_X1 U11247 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG2_REG_10__SCAN_IN), 
        .A3(n10194), .A4(n10193), .ZN(n10202) );
  NOR4_X1 U11248 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(n10195), .A4(n6796), .ZN(n10201) );
  NOR4_X1 U11249 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(P2_DATAO_REG_31__SCAN_IN), 
        .A3(n10197), .A4(n10196), .ZN(n10200) );
  NOR4_X1 U11250 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n6702), .A3(n6769), .A4(
        n10198), .ZN(n10199) );
  NAND4_X1 U11251 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10245) );
  NAND4_X1 U11252 ( .A1(n10204), .A2(n6709), .A3(n6335), .A4(n10203), .ZN(
        n10213) );
  NAND4_X1 U11253 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P2_REG0_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_30__SCAN_IN), .A4(n10205), .ZN(n10212) );
  NAND4_X1 U11254 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P1_REG1_REG_6__SCAN_IN), 
        .A3(n10206), .A4(n7926), .ZN(n10211) );
  NAND4_X1 U11255 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(
        P2_IR_REG_3__SCAN_IN), .ZN(n10210) );
  NOR4_X1 U11256 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10243) );
  NAND4_X1 U11257 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P2_RD_REG_SCAN_IN), 
        .A3(P2_REG1_REG_29__SCAN_IN), .A4(n10214), .ZN(n10224) );
  NAND4_X1 U11258 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10217), .A3(n10216), .A4(
        n10215), .ZN(n10223) );
  NAND4_X1 U11259 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(n10219), .A3(n10218), 
        .A4(n6788), .ZN(n10222) );
  NAND4_X1 U11260 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), 
        .A3(P2_D_REG_4__SCAN_IN), .A4(n10220), .ZN(n10221) );
  NOR4_X1 U11261 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(
        n10242) );
  NAND4_X1 U11262 ( .A1(SI_21_), .A2(P1_REG0_REG_13__SCAN_IN), .A3(
        P2_REG1_REG_20__SCAN_IN), .A4(P2_REG1_REG_31__SCAN_IN), .ZN(n10232) );
  NAND4_X1 U11263 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P1_REG0_REG_11__SCAN_IN), 
        .A3(n10226), .A4(n10225), .ZN(n10231) );
  NAND4_X1 U11264 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(SI_15_), .A3(
        P2_REG1_REG_18__SCAN_IN), .A4(n10227), .ZN(n10230) );
  NAND4_X1 U11265 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(P2_REG2_REG_7__SCAN_IN), 
        .A3(n10228), .A4(n4988), .ZN(n10229) );
  NOR4_X1 U11266 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10241) );
  NAND4_X1 U11267 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_9__SCAN_IN), .A4(n10233), .ZN(n10239) );
  NAND4_X1 U11268 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), 
        .A3(n5317), .A4(n8270), .ZN(n10238) );
  NAND4_X1 U11269 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(P1_REG3_REG_1__SCAN_IN), 
        .A3(n10235), .A4(n10234), .ZN(n10237) );
  NAND4_X1 U11270 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG0_REG_18__SCAN_IN), .A4(n5781), .ZN(n10236) );
  NOR4_X1 U11271 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  NAND4_X1 U11272 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10244) );
  NOR4_X1 U11273 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  XNOR2_X1 U11274 ( .A(n10249), .B(n10248), .ZN(n10253) );
  MUX2_X1 U11275 ( .A(n10251), .B(n10250), .S(P1_U4006), .Z(n10252) );
  XOR2_X1 U11276 ( .A(n10253), .B(n10252), .Z(P1_U3585) );
  XOR2_X1 U11277 ( .A(n10254), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11278 ( .A(n10255), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11279 ( .A1(n10257), .A2(n10256), .ZN(n10258) );
  XOR2_X1 U11280 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10258), .Z(ADD_1071_U51) );
  OAI21_X1 U11281 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(n10262) );
  XNOR2_X1 U11282 ( .A(n10262), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11283 ( .B1(n10265), .B2(n10264), .A(n10263), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11284 ( .A(n10267), .B(n10266), .ZN(ADD_1071_U48) );
  XOR2_X1 U11285 ( .A(n10269), .B(n10268), .Z(ADD_1071_U54) );
  XOR2_X1 U11286 ( .A(n10271), .B(n10270), .Z(ADD_1071_U53) );
  XNOR2_X1 U11287 ( .A(n10273), .B(n10272), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4892 ( .A(n6421), .Z(n6538) );
  CLKBUF_X1 U4895 ( .A(n5821), .Z(n6658) );
  CLKBUF_X1 U4897 ( .A(n6658), .Z(n4406) );
  CLKBUF_X1 U4915 ( .A(n5815), .Z(n5974) );
  CLKBUF_X1 U4917 ( .A(n5747), .Z(n4378) );
  CLKBUF_X1 U4923 ( .A(n9786), .Z(n4402) );
endmodule

