

module b21_C_AntiSAT_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031;

  NAND2_X1 U4814 ( .A1(n8904), .A2(n4323), .ZN(n8854) );
  INV_X2 U4815 ( .A(n5468), .ZN(n6175) );
  AND3_X1 U4816 ( .A1(n4954), .A2(n4953), .A3(n4952), .ZN(n6594) );
  INV_X1 U4817 ( .A(n6129), .ZN(n8350) );
  NAND2_X2 U4818 ( .A1(n5600), .A2(n6209), .ZN(n6058) );
  BUF_X1 U4819 ( .A(n5518), .Z(n4312) );
  AND2_X4 U4820 ( .A1(n9053), .A2(n9057), .ZN(n4964) );
  OR2_X1 U4822 ( .A1(n6735), .A2(n6749), .ZN(n6747) );
  INV_X1 U4823 ( .A(n4947), .ZN(n5291) );
  INV_X1 U4824 ( .A(n4926), .ZN(n6244) );
  NAND2_X1 U4825 ( .A1(n4630), .A2(n4628), .ZN(n9335) );
  INV_X1 U4826 ( .A(n7132), .ZN(n9818) );
  INV_X1 U4827 ( .A(n8382), .ZN(n6174) );
  OAI22_X1 U4828 ( .A1(n8812), .A2(n4558), .B1(n8697), .B2(n8968), .ZN(n8800)
         );
  AND2_X1 U4829 ( .A1(n7448), .A2(n7497), .ZN(n7505) );
  NAND2_X1 U4830 ( .A1(n4312), .A2(n8379), .ZN(n5526) );
  INV_X1 U4831 ( .A(n8379), .ZN(n5290) );
  INV_X1 U4832 ( .A(n6756), .ZN(n6760) );
  NAND2_X1 U4833 ( .A1(n5407), .A2(n5406), .ZN(n8629) );
  NAND2_X1 U4834 ( .A1(n5271), .A2(n5270), .ZN(n9000) );
  NAND2_X1 U4835 ( .A1(n4667), .A2(n4664), .ZN(n8812) );
  OAI21_X1 U4836 ( .B1(n8946), .B2(n9963), .A(n4678), .ZN(n4677) );
  NAND2_X2 U4838 ( .A1(n6154), .A2(n6311), .ZN(n8002) );
  OAI21_X1 U4839 ( .B1(n9105), .B2(n4609), .A(n4337), .ZN(n6134) );
  OR3_X1 U4840 ( .A1(n7518), .A2(n7321), .A3(n7467), .ZN(n6209) );
  AND2_X1 U4841 ( .A1(n4709), .A2(n4389), .ZN(n6196) );
  XNOR2_X1 U4842 ( .A(n5491), .B(n7927), .ZN(n5519) );
  INV_X1 U4843 ( .A(n8296), .ZN(n9283) );
  NOR2_X2 U4844 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4927) );
  OAI222_X1 U4845 ( .A1(n9060), .A2(n6232), .B1(n9058), .B2(n6231), .C1(
        P2_U3152), .C2(n6405), .ZN(P2_U3352) );
  OAI222_X1 U4846 ( .A1(n9609), .A2(n6230), .B1(n9613), .B2(n6231), .C1(
        P1_U3084), .C2(n6450), .ZN(P1_U3347) );
  OR2_X2 U4847 ( .A1(n5717), .A2(n6231), .ZN(n5704) );
  XNOR2_X1 U4849 ( .A(n4874), .B(n4899), .ZN(n5530) );
  AOI22_X1 U4850 ( .A1(n6593), .A2(n6592), .B1(n4961), .B2(n4960), .ZN(n6608)
         );
  XNOR2_X2 U4851 ( .A(n5116), .B(n4856), .ZN(n6269) );
  AOI21_X2 U4852 ( .B1(n5283), .B2(n4391), .A(n4769), .ZN(n5344) );
  OAI21_X2 U4853 ( .B1(n5268), .B2(n5267), .A(n5266), .ZN(n5283) );
  NAND2_X2 U4854 ( .A1(n6359), .A2(n5530), .ZN(n4926) );
  AOI21_X2 U4855 ( .B1(n9335), .B2(n8152), .A(n7735), .ZN(n9299) );
  OAI22_X2 U4856 ( .A1(n8611), .A2(n8610), .B1(n5067), .B2(n5066), .ZN(n6868)
         );
  NOR2_X2 U4857 ( .A1(n6813), .A2(n8382), .ZN(n6814) );
  NAND2_X2 U4858 ( .A1(n8191), .A2(n6725), .ZN(n6735) );
  NAND2_X2 U4859 ( .A1(n8350), .A2(n9283), .ZN(n6727) );
  NAND2_X1 U4860 ( .A1(n4992), .A2(n4991), .ZN(n5006) );
  XNOR2_X1 U4862 ( .A(n5605), .B(n5604), .ZN(n6129) );
  NAND2_X2 U4863 ( .A1(n5519), .A2(n8409), .ZN(n5516) );
  NAND2_X2 U4864 ( .A1(n4480), .A2(n5641), .ZN(n6756) );
  INV_X1 U4865 ( .A(n9892), .ZN(n6283) );
  AND2_X2 U4866 ( .A1(n8366), .A2(n5592), .ZN(n5644) );
  XNOR2_X1 U4869 ( .A(n4611), .B(n5583), .ZN(n6154) );
  NAND2_X1 U4870 ( .A1(n8001), .A2(P1_U3084), .ZN(n9609) );
  OAI21_X1 U4871 ( .B1(n8582), .B2(n4751), .A(n6245), .ZN(n4750) );
  AOI21_X1 U4872 ( .B1(n4674), .B2(n9983), .A(n4673), .ZN(n4672) );
  OR2_X1 U4873 ( .A1(n4565), .A2(n8959), .ZN(n9034) );
  NAND2_X1 U4874 ( .A1(n4842), .A2(n4841), .ZN(n8354) );
  NAND2_X1 U4875 ( .A1(n4371), .A2(n8572), .ZN(n4838) );
  AOI211_X1 U4876 ( .C1(n9897), .C2(n9627), .A(n9626), .B(n9625), .ZN(n9630)
         );
  NAND2_X1 U4877 ( .A1(n9407), .A2(n9408), .ZN(n9406) );
  AND3_X1 U4878 ( .A1(n4552), .A2(n8543), .A3(n4553), .ZN(n8803) );
  OAI21_X1 U4879 ( .B1(n8887), .B2(n8029), .A(n8028), .ZN(n8853) );
  XNOR2_X1 U4880 ( .A(n7995), .B(n7994), .ZN(n8004) );
  OAI21_X1 U4881 ( .B1(n7608), .B2(n4407), .A(n4405), .ZN(n8024) );
  AOI21_X1 U4882 ( .B1(n7576), .B2(n8503), .A(n7575), .ZN(n7606) );
  NAND2_X1 U4883 ( .A1(n5394), .A2(n5393), .ZN(n8968) );
  OR2_X1 U4884 ( .A1(n7433), .A2(n8498), .ZN(n7504) );
  OAI21_X1 U4885 ( .B1(n5392), .B2(n4766), .A(n4764), .ZN(n6087) );
  INV_X1 U4886 ( .A(n8507), .ZN(n4311) );
  OR2_X1 U4887 ( .A1(n7328), .A2(n7282), .ZN(n7284) );
  NAND2_X1 U4888 ( .A1(n5258), .A2(n5257), .ZN(n9007) );
  NAND2_X1 U4889 ( .A1(n7002), .A2(n4357), .ZN(n7019) );
  NAND2_X1 U4890 ( .A1(n6847), .A2(n8463), .ZN(n7002) );
  AND2_X1 U4891 ( .A1(n4522), .A2(n6860), .ZN(n7116) );
  INV_X2 U4892 ( .A(n8933), .ZN(n8931) );
  NAND2_X2 U4893 ( .A1(n6813), .A2(n8844), .ZN(n8933) );
  NAND2_X1 U4894 ( .A1(n5099), .A2(n5098), .ZN(n9941) );
  NOR2_X1 U4895 ( .A1(n9983), .A2(n6183), .ZN(n4673) );
  NAND2_X1 U4896 ( .A1(n6850), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U4897 ( .A1(n5030), .A2(n5029), .ZN(n6975) );
  INV_X1 U4898 ( .A(n7102), .ZN(n6825) );
  INV_X4 U4899 ( .A(n6744), .ZN(n6024) );
  AND2_X1 U4900 ( .A1(n4994), .A2(n4993), .ZN(n7102) );
  AND3_X1 U4901 ( .A1(n4982), .A2(n4981), .A3(n4980), .ZN(n9905) );
  NAND2_X1 U4902 ( .A1(n4894), .A2(n6285), .ZN(n4898) );
  NAND2_X2 U4903 ( .A1(n6726), .A2(n6209), .ZN(n6055) );
  CLKBUF_X1 U4904 ( .A(n6130), .Z(n8292) );
  NAND2_X1 U4905 ( .A1(n8588), .A2(n5290), .ZN(n6285) );
  OR2_X2 U4906 ( .A1(n6130), .A2(n8340), .ZN(n6726) );
  NAND2_X1 U4907 ( .A1(n6277), .A2(n6528), .ZN(n8440) );
  AND2_X1 U4908 ( .A1(n5516), .A2(n8409), .ZN(n4894) );
  NAND2_X1 U4909 ( .A1(n5603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5605) );
  AND2_X1 U4910 ( .A1(n4725), .A2(n4728), .ZN(n6528) );
  XNOR2_X1 U4911 ( .A(n4890), .B(n4889), .ZN(n8409) );
  AND3_X1 U4912 ( .A1(n4931), .A2(n4930), .A3(n4929), .ZN(n6532) );
  AND2_X2 U4913 ( .A1(n5594), .A2(n5592), .ZN(n6067) );
  NAND2_X1 U4914 ( .A1(n4893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4896) );
  OAI21_X1 U4915 ( .B1(n4888), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U4916 ( .A1(n5568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U4917 ( .A1(n9604), .A2(n5588), .ZN(n9611) );
  XNOR2_X1 U4918 ( .A(n4901), .B(n4900), .ZN(n9053) );
  XNOR2_X1 U4919 ( .A(n4903), .B(n4559), .ZN(n9057) );
  XNOR2_X1 U4920 ( .A(n5584), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5594) );
  MUX2_X1 U4921 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5587), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5588) );
  NAND2_X1 U4922 ( .A1(n4902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4903) );
  XNOR2_X1 U4923 ( .A(n4610), .B(n5559), .ZN(n6311) );
  OR2_X1 U4924 ( .A1(n5585), .A2(n5557), .ZN(n5584) );
  OR2_X1 U4925 ( .A1(n5558), .A2(n4811), .ZN(n5586) );
  AND2_X1 U4926 ( .A1(n4822), .A2(n5618), .ZN(n5560) );
  AND3_X1 U4927 ( .A1(n4732), .A2(n4733), .A3(n4883), .ZN(n5236) );
  OR2_X2 U4928 ( .A1(n4870), .A2(n4978), .ZN(n4332) );
  NAND2_X2 U4929 ( .A1(n4412), .A2(n4411), .ZN(n4919) );
  AND4_X1 U4930 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n4847)
         );
  AND3_X1 U4931 ( .A1(n5567), .A2(n5908), .A3(n5604), .ZN(n5556) );
  NAND3_X1 U4932 ( .A1(n4877), .A2(n4413), .A3(n4414), .ZN(n4412) );
  NOR2_X1 U4933 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4533) );
  INV_X1 U4934 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4889) );
  INV_X4 U4935 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X2 U4936 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4568) );
  INV_X1 U4937 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5702) );
  INV_X1 U4938 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4413) );
  INV_X1 U4939 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5119) );
  NOR2_X1 U4940 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4865) );
  INV_X1 U4941 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U4942 ( .A1(n5594), .A2(n9611), .ZN(n8010) );
  XNOR2_X1 U4943 ( .A(n4729), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5518) );
  AND2_X4 U4944 ( .A1(n9053), .A2(n4905), .ZN(n4955) );
  AND2_X4 U4945 ( .A1(n4904), .A2(n9057), .ZN(n4995) );
  AOI22_X2 U4946 ( .A1(n6697), .A2(n6696), .B1(n5040), .B2(n5039), .ZN(n8611)
         );
  NAND2_X1 U4947 ( .A1(n4926), .A2(n8377), .ZN(n4317) );
  XNOR2_X2 U4948 ( .A(n4876), .B(n4875), .ZN(n6359) );
  INV_X1 U4949 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5231) );
  INV_X1 U4950 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5230) );
  OR2_X1 U4951 ( .A1(n8990), .A2(n8025), .ZN(n8528) );
  NAND2_X1 U4952 ( .A1(n4657), .A2(n8384), .ZN(n4656) );
  INV_X1 U4953 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4452) );
  AND2_X1 U4954 ( .A1(n5579), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U4955 ( .A1(n5283), .A2(n5282), .ZN(n4773) );
  INV_X1 U4956 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5548) );
  NOR2_X1 U4957 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5550) );
  NOR2_X1 U4958 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5549) );
  NAND2_X1 U4959 ( .A1(n5105), .A2(n5106), .ZN(n4692) );
  INV_X1 U4960 ( .A(n4956), .ZN(n6180) );
  OR2_X1 U4961 ( .A1(n8965), .A2(n8696), .ZN(n8030) );
  NAND2_X1 U4962 ( .A1(n8552), .A2(n8555), .ZN(n8788) );
  NAND2_X1 U4963 ( .A1(n8002), .A2(n8377), .ZN(n5717) );
  AOI21_X1 U4964 ( .B1(n4802), .B2(n4801), .A(n4366), .ZN(n4800) );
  INV_X1 U4965 ( .A(n4806), .ZN(n4801) );
  NAND2_X1 U4966 ( .A1(n8491), .A2(n4339), .ZN(n4505) );
  AOI21_X1 U4967 ( .B1(n8517), .B2(n8533), .A(n8516), .ZN(n8521) );
  AOI21_X1 U4968 ( .B1(n4473), .B2(n8134), .A(n8138), .ZN(n4472) );
  NAND2_X1 U4969 ( .A1(n9941), .A2(n7111), .ZN(n8417) );
  INV_X1 U4970 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4823) );
  NOR2_X1 U4971 ( .A1(n4758), .A2(n4755), .ZN(n4754) );
  INV_X1 U4972 ( .A(n5091), .ZN(n4755) );
  INV_X1 U4973 ( .A(n4759), .ZN(n4758) );
  INV_X1 U4974 ( .A(n4661), .ZN(n4407) );
  NAND2_X1 U4975 ( .A1(n4316), .A2(n8433), .ZN(n6811) );
  OR2_X1 U4976 ( .A1(n8586), .A2(n6352), .ZN(n6804) );
  NOR2_X1 U4977 ( .A1(n5499), .A2(n7546), .ZN(n5510) );
  AND2_X1 U4978 ( .A1(n7465), .A2(n5495), .ZN(n5499) );
  INV_X1 U4979 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4899) );
  INV_X1 U4980 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4885) );
  NOR2_X1 U4981 ( .A1(n4978), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4732) );
  OR2_X1 U4982 ( .A1(n5061), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5097) );
  OR3_X1 U4983 ( .A1(n7226), .A2(n7126), .A3(n7228), .ZN(n4851) );
  AND2_X1 U4984 ( .A1(n4594), .A2(n7563), .ZN(n4593) );
  INV_X1 U4985 ( .A(n6055), .ZN(n4606) );
  INV_X1 U4986 ( .A(n9611), .ZN(n5592) );
  NOR2_X1 U4987 ( .A1(n9323), .A2(n4818), .ZN(n4817) );
  INV_X1 U4988 ( .A(n7716), .ZN(n4818) );
  OR2_X1 U4989 ( .A1(n9513), .A2(n7717), .ZN(n8286) );
  AND2_X1 U4990 ( .A1(n8286), .A2(n8183), .ZN(n9323) );
  NOR2_X1 U4991 ( .A1(n7715), .A2(n4629), .ZN(n4628) );
  INV_X1 U4992 ( .A(n8253), .ZN(n4629) );
  INV_X1 U4993 ( .A(n7703), .ZN(n4776) );
  NOR2_X1 U4994 ( .A1(n9193), .A2(n9570), .ZN(n4495) );
  NAND2_X1 U4995 ( .A1(n4763), .A2(n5413), .ZN(n5461) );
  NAND2_X1 U4996 ( .A1(n5392), .A2(n4767), .ZN(n4763) );
  NAND2_X1 U4997 ( .A1(n5347), .A2(n5346), .ZN(n5369) );
  OR2_X1 U4998 ( .A1(n5344), .A2(n5343), .ZN(n5347) );
  AND2_X1 U4999 ( .A1(n5253), .A2(n5235), .ZN(n5251) );
  XNOR2_X1 U5000 ( .A(n4910), .B(n4731), .ZN(n6345) );
  INV_X1 U5001 ( .A(n4911), .ZN(n4731) );
  OR2_X1 U5002 ( .A1(n5354), .A2(n8671), .ZN(n5377) );
  INV_X1 U5003 ( .A(n6867), .ZN(n4689) );
  AND3_X1 U5004 ( .A1(n5322), .A2(n5321), .A3(n5320), .ZN(n8025) );
  NOR2_X1 U5005 ( .A1(n6486), .A2(n6485), .ZN(n6484) );
  AND2_X1 U5006 ( .A1(n8788), .A2(n4403), .ZN(n4402) );
  OR2_X1 U5007 ( .A1(n8802), .A2(n4404), .ZN(n4403) );
  INV_X1 U5008 ( .A(n8030), .ZN(n4404) );
  AOI21_X1 U5009 ( .B1(n7949), .B2(n4543), .A(n4542), .ZN(n4541) );
  INV_X1 U5010 ( .A(n8524), .ZN(n4542) );
  NAND2_X1 U5011 ( .A1(n7114), .A2(n8394), .ZN(n7213) );
  INV_X2 U5012 ( .A(n4939), .ZN(n8370) );
  INV_X1 U5013 ( .A(n8915), .ZN(n8861) );
  NAND2_X1 U5014 ( .A1(n4653), .A2(n4655), .ZN(n4651) );
  AND2_X1 U5015 ( .A1(n8459), .A2(n8452), .ZN(n6833) );
  OR2_X1 U5016 ( .A1(n8359), .A2(n6180), .ZN(n5540) );
  NAND2_X1 U5017 ( .A1(n8362), .A2(n8559), .ZN(n8363) );
  AND2_X1 U5018 ( .A1(n6350), .A2(n9885), .ZN(n9879) );
  AND2_X1 U5019 ( .A1(n5925), .A2(n5944), .ZN(n4604) );
  NAND2_X1 U5020 ( .A1(n9741), .A2(n9740), .ZN(n9739) );
  NAND2_X1 U5021 ( .A1(n4821), .A2(n7717), .ZN(n4820) );
  NOR2_X1 U5022 ( .A1(n7710), .A2(n4807), .ZN(n4806) );
  INV_X1 U5023 ( .A(n7707), .ZN(n4807) );
  OR2_X1 U5024 ( .A1(n9399), .A2(n7706), .ZN(n7708) );
  NAND2_X1 U5025 ( .A1(n7653), .A2(n4638), .ZN(n7627) );
  AND2_X1 U5026 ( .A1(n8110), .A2(n8103), .ZN(n4638) );
  AOI21_X1 U5027 ( .B1(n4789), .B2(n8315), .A(n4386), .ZN(n4788) );
  OR2_X1 U5028 ( .A1(n9616), .A2(n7378), .ZN(n8204) );
  INV_X1 U5029 ( .A(n8006), .ZN(n5928) );
  INV_X1 U5030 ( .A(n8002), .ZN(n5927) );
  OAI21_X1 U5031 ( .B1(n7068), .B2(n4795), .A(n4793), .ZN(n7250) );
  INV_X1 U5032 ( .A(n4794), .ZN(n4793) );
  OAI21_X1 U5033 ( .B1(n4335), .B2(n4795), .A(n8311), .ZN(n4794) );
  INV_X1 U5034 ( .A(n7070), .ZN(n4795) );
  NAND2_X1 U5035 ( .A1(n7068), .A2(n4335), .ZN(n7149) );
  NAND2_X1 U5036 ( .A1(n6724), .A2(n8341), .ZN(n9488) );
  NAND2_X1 U5037 ( .A1(n7725), .A2(n7724), .ZN(n9499) );
  OAI21_X1 U5038 ( .B1(n5558), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4611) );
  XNOR2_X1 U5039 ( .A(n5025), .B(SI_6_), .ZN(n5023) );
  OR3_X1 U5040 ( .A1(n7324), .A2(n7465), .A3(n7546), .ZN(n6350) );
  AND2_X1 U5041 ( .A1(n8221), .A2(n8171), .ZN(n4464) );
  AND2_X1 U5042 ( .A1(n4507), .A2(n8504), .ZN(n4506) );
  OR2_X1 U5043 ( .A1(n8397), .A2(n4508), .ZN(n4507) );
  AOI21_X1 U5044 ( .B1(n4327), .B2(n8114), .A(n4462), .ZN(n4461) );
  OAI211_X1 U5045 ( .C1(n8102), .C2(n8101), .A(n4459), .B(n4458), .ZN(n4457)
         );
  INV_X1 U5046 ( .A(n8113), .ZN(n4462) );
  NAND2_X1 U5047 ( .A1(n4513), .A2(n8556), .ZN(n8540) );
  OAI21_X1 U5048 ( .B1(n8521), .B2(n8518), .A(n4514), .ZN(n4513) );
  NOR2_X1 U5049 ( .A1(n8820), .A2(n8520), .ZN(n4514) );
  INV_X1 U5050 ( .A(n5326), .ZN(n4715) );
  AND2_X1 U5051 ( .A1(n8137), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U5052 ( .A1(n4472), .A2(n4470), .ZN(n4469) );
  INV_X1 U5053 ( .A(n4472), .ZN(n4471) );
  INV_X1 U5054 ( .A(n8142), .ZN(n4467) );
  AOI21_X1 U5055 ( .B1(n8553), .B2(n8552), .A(n8551), .ZN(n4499) );
  NAND2_X1 U5056 ( .A1(n4558), .A2(n8541), .ZN(n4557) );
  NAND2_X1 U5057 ( .A1(n4387), .A2(n5413), .ZN(n4766) );
  NOR2_X1 U5058 ( .A1(n5409), .A2(n4768), .ZN(n4767) );
  INV_X1 U5059 ( .A(n5391), .ZN(n4768) );
  AND2_X1 U5060 ( .A1(n5329), .A2(n5328), .ZN(n5331) );
  INV_X1 U5061 ( .A(n4856), .ZN(n4757) );
  NOR2_X1 U5062 ( .A1(n5130), .A2(n4760), .ZN(n4759) );
  INV_X1 U5063 ( .A(n5117), .ZN(n4760) );
  NAND2_X1 U5064 ( .A1(n5090), .A2(n4855), .ZN(n5092) );
  INV_X1 U5065 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4414) );
  AOI21_X1 U5066 ( .B1(n4713), .B2(n4716), .A(n4343), .ZN(n4712) );
  AND2_X1 U5067 ( .A1(n5480), .A2(n5479), .ZN(n6179) );
  INV_X1 U5068 ( .A(n5126), .ZN(n4691) );
  INV_X1 U5069 ( .A(n7136), .ZN(n4685) );
  INV_X1 U5070 ( .A(n4333), .ZN(n4683) );
  OR2_X1 U5071 ( .A1(n8949), .A2(n8776), .ZN(n8562) );
  NAND2_X1 U5072 ( .A1(n8043), .A2(n8033), .ZN(n4518) );
  OR2_X1 U5073 ( .A1(n8980), .A2(n8837), .ZN(n8834) );
  NOR2_X1 U5074 ( .A1(n8996), .A2(n8990), .ZN(n4520) );
  OR2_X1 U5075 ( .A1(n9020), .A2(n7600), .ZN(n8494) );
  NOR2_X1 U5076 ( .A1(n7028), .A2(n8615), .ZN(n4524) );
  OR2_X1 U5077 ( .A1(n7028), .A2(n7008), .ZN(n8419) );
  INV_X1 U5078 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4873) );
  NOR2_X1 U5079 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4528) );
  INV_X1 U5080 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5081 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4530) );
  NOR2_X1 U5082 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4531) );
  NOR2_X1 U5083 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n4532) );
  INV_X1 U5084 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5176) );
  INV_X1 U5085 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5205) );
  AND2_X1 U5086 ( .A1(n4732), .A2(n4733), .ZN(n5166) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4867) );
  NOR2_X1 U5088 ( .A1(n4590), .A2(n4587), .ZN(n4586) );
  INV_X1 U5089 ( .A(n5830), .ZN(n4587) );
  NAND2_X1 U5090 ( .A1(n4448), .A2(n4446), .ZN(n8172) );
  NAND2_X1 U5091 ( .A1(n8153), .A2(n4449), .ZN(n4448) );
  AND2_X1 U5092 ( .A1(n8159), .A2(n4447), .ZN(n4446) );
  AND2_X1 U5093 ( .A1(n8151), .A2(n8152), .ZN(n4449) );
  OR2_X1 U5094 ( .A1(n9499), .A2(n9505), .ZN(n4488) );
  INV_X1 U5095 ( .A(n8099), .ZN(n4618) );
  AND2_X1 U5096 ( .A1(n4616), .A2(n8094), .ZN(n4615) );
  NAND2_X1 U5097 ( .A1(n8099), .A2(n4617), .ZN(n4616) );
  OR2_X1 U5098 ( .A1(n7275), .A2(n7078), .ZN(n4492) );
  INV_X1 U5099 ( .A(n8197), .ZN(n4624) );
  INV_X1 U5100 ( .A(n7057), .ZN(n4456) );
  NOR2_X1 U5101 ( .A1(n6890), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5102 ( .A1(n6735), .A2(n6737), .ZN(n6736) );
  OR2_X1 U5103 ( .A1(n5717), .A2(n6218), .ZN(n5640) );
  OR2_X1 U5104 ( .A1(n8006), .A2(n6216), .ZN(n5641) );
  NAND2_X1 U5105 ( .A1(n4367), .A2(n8002), .ZN(n4476) );
  INV_X1 U5106 ( .A(n8292), .ZN(n8332) );
  NAND2_X1 U5107 ( .A1(n7719), .A2(n7718), .ZN(n7987) );
  NOR2_X1 U5108 ( .A1(n5566), .A2(n5565), .ZN(n5606) );
  NAND2_X1 U5109 ( .A1(n4850), .A2(n5564), .ZN(n5565) );
  AOI21_X1 U5110 ( .B1(n5200), .B2(n4739), .A(n4735), .ZN(n4734) );
  NAND2_X1 U5111 ( .A1(n4736), .A2(n5253), .ZN(n4735) );
  NAND2_X1 U5112 ( .A1(n4739), .A2(n4741), .ZN(n4736) );
  NAND2_X1 U5113 ( .A1(n5560), .A2(n5561), .ZN(n5566) );
  AND2_X1 U5114 ( .A1(n5867), .A2(n5865), .ZN(n5561) );
  AND2_X1 U5115 ( .A1(n5551), .A2(n4351), .ZN(n4822) );
  OAI21_X1 U5116 ( .B1(n5160), .B2(n5159), .A(n5158), .ZN(n5174) );
  OAI21_X1 U5117 ( .B1(n5069), .B2(n5068), .A(n5070), .ZN(n5090) );
  OAI21_X1 U5118 ( .B1(n8377), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4512), .ZN(
        n5025) );
  NAND2_X1 U5119 ( .A1(n8377), .A2(n6230), .ZN(n4512) );
  OAI21_X1 U5120 ( .B1(n8377), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4946), .ZN(
        n4971) );
  NAND2_X1 U5121 ( .A1(n8377), .A2(n6217), .ZN(n4946) );
  OAI211_X1 U5122 ( .C1(n4919), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n4879), .B(
        SI_0_), .ZN(n4922) );
  NAND2_X1 U5123 ( .A1(n4919), .A2(n4878), .ZN(n4879) );
  AND2_X1 U5124 ( .A1(n5022), .A2(n4701), .ZN(n4693) );
  OR2_X1 U5125 ( .A1(n5152), .A2(n7090), .ZN(n5182) );
  INV_X1 U5126 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5181) );
  OR2_X1 U5127 ( .A1(n5377), .A2(n5376), .ZN(n5397) );
  INV_X1 U5128 ( .A(n4706), .ZN(n4705) );
  OAI21_X1 U5129 ( .B1(n4708), .B2(n4707), .A(n8678), .ZN(n4706) );
  INV_X1 U5130 ( .A(n5262), .ZN(n4707) );
  NAND2_X1 U5131 ( .A1(n8377), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4727) );
  NAND2_X1 U5132 ( .A1(n4917), .A2(n6283), .ZN(n4918) );
  NAND2_X1 U5133 ( .A1(n5468), .A2(n9892), .ZN(n4730) );
  NOR2_X1 U5134 ( .A1(n5216), .A2(n7595), .ZN(n4723) );
  INV_X1 U5135 ( .A(n4719), .ZN(n4718) );
  OAI21_X1 U5136 ( .B1(n4724), .B2(n4722), .A(n4720), .ZN(n4719) );
  OR2_X1 U5137 ( .A1(n5182), .A2(n5181), .ZN(n5221) );
  NAND2_X1 U5138 ( .A1(n5335), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U5139 ( .A1(n5078), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5110) );
  XNOR2_X1 U5140 ( .A(n8925), .B(n4932), .ZN(n4910) );
  NOR2_X1 U5141 ( .A1(n4985), .A2(n6562), .ZN(n4701) );
  NOR2_X1 U5142 ( .A1(n6647), .A2(n4698), .ZN(n4697) );
  INV_X1 U5143 ( .A(n4700), .ZN(n4698) );
  OR2_X1 U5144 ( .A1(n6808), .A2(n5512), .ZN(n5529) );
  AND2_X1 U5145 ( .A1(n5215), .A2(n5192), .ZN(n4724) );
  OR2_X1 U5146 ( .A1(n6484), .A2(n4382), .ZN(n4418) );
  AND2_X1 U5147 ( .A1(n4418), .A2(n4417), .ZN(n6395) );
  INV_X1 U5148 ( .A(n6396), .ZN(n4417) );
  OR2_X1 U5149 ( .A1(n6510), .A2(n4392), .ZN(n4430) );
  AND2_X1 U5150 ( .A1(n4430), .A2(n4429), .ZN(n6622) );
  INV_X1 U5151 ( .A(n6513), .ZN(n4429) );
  NOR2_X1 U5152 ( .A1(n6791), .A2(n6790), .ZN(n7039) );
  NOR2_X1 U5153 ( .A1(n7039), .A2(n4442), .ZN(n7041) );
  AND2_X1 U5154 ( .A1(n7047), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4442) );
  NOR2_X1 U5155 ( .A1(n7972), .A2(n7973), .ZN(n8715) );
  NAND2_X1 U5156 ( .A1(n8715), .A2(n8714), .ZN(n8713) );
  AND2_X1 U5157 ( .A1(n5471), .A2(n5444), .ZN(n8793) );
  INV_X1 U5158 ( .A(n4665), .ZN(n4664) );
  OAI21_X1 U5159 ( .B1(n8833), .B2(n4666), .A(n4853), .ZN(n4665) );
  NOR2_X1 U5160 ( .A1(n8833), .A2(n4669), .ZN(n4668) );
  INV_X1 U5161 ( .A(n4671), .ZN(n4669) );
  OR2_X1 U5162 ( .A1(n8853), .A2(n8048), .ZN(n4670) );
  OR2_X1 U5163 ( .A1(n8980), .A2(n8882), .ZN(n4671) );
  INV_X1 U5164 ( .A(n8528), .ZN(n8045) );
  AND2_X1 U5165 ( .A1(n8522), .A2(n8526), .ZN(n7952) );
  INV_X1 U5166 ( .A(n4406), .ZN(n4405) );
  OAI21_X1 U5167 ( .B1(n4407), .B2(n7577), .A(n4660), .ZN(n4406) );
  AOI21_X1 U5168 ( .B1(n8507), .B2(n4661), .A(n4324), .ZN(n4660) );
  OR2_X1 U5169 ( .A1(n9007), .A2(n8686), .ZN(n8910) );
  AND2_X1 U5170 ( .A1(n8511), .A2(n8524), .ZN(n8914) );
  AND4_X1 U5171 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n7948)
         );
  NAND2_X1 U5172 ( .A1(n4663), .A2(n4311), .ZN(n7941) );
  NAND2_X1 U5173 ( .A1(n4537), .A2(n4539), .ZN(n4534) );
  AND2_X1 U5174 ( .A1(n8395), .A2(n7212), .ZN(n4415) );
  NAND2_X1 U5175 ( .A1(n7116), .A2(n9949), .ZN(n7215) );
  NAND2_X1 U5176 ( .A1(n7019), .A2(n4360), .ZN(n7113) );
  AND4_X1 U5177 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n6854)
         );
  INV_X1 U5178 ( .A(n6581), .ZN(n4659) );
  OR2_X1 U5179 ( .A1(n8449), .A2(n4827), .ZN(n4824) );
  NAND2_X1 U5180 ( .A1(n8424), .A2(n6830), .ZN(n6955) );
  NAND2_X1 U5181 ( .A1(n6956), .A2(n6955), .ZN(n6954) );
  OR2_X1 U5182 ( .A1(n9030), .A2(n8433), .ZN(n6809) );
  AND2_X1 U5183 ( .A1(n5140), .A2(n5139), .ZN(n9956) );
  INV_X1 U5184 ( .A(n6528), .ZN(n8925) );
  AND2_X1 U5185 ( .A1(n8579), .A2(n5526), .ZN(n9897) );
  AND2_X1 U5186 ( .A1(n8579), .A2(n4316), .ZN(n9898) );
  AND2_X1 U5187 ( .A1(n4845), .A2(n4873), .ZN(n4844) );
  AND2_X1 U5188 ( .A1(n4899), .A2(n4875), .ZN(n4845) );
  NAND2_X1 U5189 ( .A1(n5492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5514) );
  INV_X1 U5190 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5513) );
  INV_X1 U5191 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4884) );
  NOR2_X1 U5192 ( .A1(n4571), .A2(n6009), .ZN(n4570) );
  NOR2_X1 U5193 ( .A1(n5634), .A2(n5633), .ZN(n5659) );
  NAND2_X1 U5194 ( .A1(n6061), .A2(n4608), .ZN(n4607) );
  INV_X1 U5195 ( .A(n9106), .ZN(n4608) );
  NAND2_X1 U5196 ( .A1(n7181), .A2(n4598), .ZN(n5727) );
  NAND2_X1 U5197 ( .A1(n9123), .A2(n6029), .ZN(n9105) );
  NAND2_X1 U5198 ( .A1(n4578), .A2(n9182), .ZN(n9644) );
  NAND2_X1 U5199 ( .A1(n5881), .A2(n9185), .ZN(n4579) );
  NAND2_X1 U5200 ( .A1(n4577), .A2(n4576), .ZN(n9123) );
  INV_X1 U5201 ( .A(n9125), .ZN(n4576) );
  NAND2_X1 U5202 ( .A1(n6703), .A2(n5677), .ZN(n6200) );
  NAND2_X1 U5203 ( .A1(n5651), .A2(n5650), .ZN(n6557) );
  AND2_X1 U5204 ( .A1(n6750), .A2(n6101), .ZN(n4605) );
  NAND2_X1 U5205 ( .A1(n5829), .A2(n7456), .ZN(n4594) );
  NOR2_X1 U5206 ( .A1(n9134), .A2(n4602), .ZN(n4601) );
  INV_X1 U5207 ( .A(n5947), .ZN(n4602) );
  OR2_X1 U5208 ( .A1(n5882), .A2(n5881), .ZN(n9183) );
  AND2_X1 U5209 ( .A1(n6040), .A2(n6039), .ZN(n9176) );
  OR2_X1 U5210 ( .A1(n9697), .A2(n9696), .ZN(n4643) );
  NAND2_X1 U5211 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5212 ( .A1(n9694), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4642) );
  AND2_X1 U5213 ( .A1(n4641), .A2(n4640), .ZN(n6329) );
  INV_X1 U5214 ( .A(n6330), .ZN(n4640) );
  NOR2_X1 U5215 ( .A1(n9726), .A2(n4639), .ZN(n9741) );
  NOR2_X1 U5216 ( .A1(n6450), .A2(n6449), .ZN(n4639) );
  INV_X1 U5217 ( .A(n4488), .ZN(n4487) );
  NOR2_X1 U5218 ( .A1(n9317), .A2(n4488), .ZN(n9289) );
  INV_X1 U5219 ( .A(n4817), .ZN(n4813) );
  OR2_X1 U5220 ( .A1(n9317), .A2(n9505), .ZN(n9305) );
  INV_X1 U5221 ( .A(n9323), .ZN(n9315) );
  INV_X1 U5222 ( .A(n4628), .ZN(n4627) );
  AOI21_X1 U5223 ( .B1(n4628), .B2(n4626), .A(n8181), .ZN(n4625) );
  OR2_X1 U5224 ( .A1(n9523), .A2(n9176), .ZN(n8253) );
  AND2_X1 U5225 ( .A1(n9334), .A2(n9344), .ZN(n9329) );
  AND2_X1 U5226 ( .A1(n9358), .A2(n9348), .ZN(n9344) );
  NAND2_X1 U5227 ( .A1(n4798), .A2(n4796), .ZN(n9343) );
  AND2_X1 U5228 ( .A1(n4797), .A2(n7712), .ZN(n4796) );
  NOR2_X1 U5229 ( .A1(n9373), .A2(n9528), .ZN(n9358) );
  INV_X1 U5230 ( .A(n7709), .ZN(n4804) );
  AND2_X1 U5231 ( .A1(n8142), .A2(n9349), .ZN(n9365) );
  OR2_X1 U5232 ( .A1(n9386), .A2(n9532), .ZN(n9373) );
  NAND2_X1 U5233 ( .A1(n4777), .A2(n7705), .ZN(n9399) );
  OAI21_X1 U5234 ( .B1(n7702), .B2(n4776), .A(n4774), .ZN(n4777) );
  AND2_X1 U5235 ( .A1(n7693), .A2(n9454), .ZN(n9428) );
  NAND2_X1 U5236 ( .A1(n7702), .A2(n7701), .ZN(n9429) );
  OR2_X1 U5237 ( .A1(n9471), .A2(n9560), .ZN(n9457) );
  INV_X1 U5238 ( .A(n7631), .ZN(n7671) );
  AND4_X1 U5239 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n9631)
         );
  INV_X1 U5240 ( .A(n7527), .ZN(n4791) );
  NOR2_X1 U5241 ( .A1(n7155), .A2(n7078), .ZN(n7258) );
  NAND2_X1 U5242 ( .A1(n8067), .A2(n8263), .ZN(n8311) );
  INV_X1 U5243 ( .A(n6899), .ZN(n4784) );
  NAND2_X1 U5244 ( .A1(n4780), .A2(n6900), .ZN(n4779) );
  AND4_X1 U5245 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n7184)
         );
  OR2_X1 U5246 ( .A1(n4314), .A2(n6449), .ZN(n5698) );
  AND2_X1 U5247 ( .A1(n7147), .A2(n8269), .ZN(n8306) );
  NAND2_X1 U5248 ( .A1(n4479), .A2(n9811), .ZN(n6939) );
  INV_X1 U5249 ( .A(n6918), .ZN(n4479) );
  OR2_X1 U5250 ( .A1(n8061), .A2(n8347), .ZN(n7744) );
  AND2_X1 U5251 ( .A1(n6729), .A2(n8347), .ZN(n9483) );
  INV_X1 U5252 ( .A(n7744), .ZN(n9485) );
  NAND2_X1 U5253 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  INV_X1 U5254 ( .A(n9334), .ZN(n9517) );
  NAND2_X1 U5255 ( .A1(n5972), .A2(n5971), .ZN(n9543) );
  NAND2_X1 U5256 ( .A1(n5786), .A2(n5785), .ZN(n9582) );
  OR2_X1 U5257 ( .A1(n8168), .A2(n8340), .ZN(n9805) );
  OR2_X1 U5258 ( .A1(n6111), .A2(n7518), .ZN(n9602) );
  NAND2_X1 U5259 ( .A1(n4810), .A2(n4809), .ZN(n4808) );
  INV_X1 U5260 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4809) );
  INV_X1 U5261 ( .A(n4811), .ZN(n4810) );
  NAND2_X1 U5262 ( .A1(n6089), .A2(n6088), .ZN(n7719) );
  NAND2_X1 U5263 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  INV_X1 U5264 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5577) );
  XNOR2_X1 U5265 ( .A(n5439), .B(n5438), .ZN(n7516) );
  INV_X1 U5266 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5581) );
  INV_X1 U5267 ( .A(n5686), .ZN(n4451) );
  INV_X1 U5268 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U5269 ( .A1(n5392), .A2(n5391), .ZN(n5410) );
  OAI21_X1 U5270 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5390) );
  AND2_X1 U5271 ( .A1(n5391), .A2(n5373), .ZN(n5389) );
  OR2_X1 U5272 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  XNOR2_X1 U5273 ( .A(n5574), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8340) );
  XNOR2_X1 U5274 ( .A(n5314), .B(n5313), .ZN(n6926) );
  NAND2_X1 U5275 ( .A1(n4773), .A2(n4771), .ZN(n5332) );
  INV_X1 U5276 ( .A(n4737), .ZN(n5252) );
  AOI21_X1 U5277 ( .B1(n5200), .B2(n4738), .A(n4741), .ZN(n4737) );
  INV_X1 U5278 ( .A(n4742), .ZN(n4738) );
  NOR2_X1 U5279 ( .A1(n5737), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5766) );
  OAI21_X1 U5280 ( .B1(n7539), .B2(n7540), .A(n5172), .ZN(n7493) );
  NAND2_X1 U5281 ( .A1(n5169), .A2(n5171), .ZN(n5172) );
  OAI22_X1 U5282 ( .A1(n6472), .A2(n6473), .B1(n4938), .B2(n4937), .ZN(n6593)
         );
  NAND2_X1 U5283 ( .A1(n5327), .A2(n5326), .ZN(n8621) );
  NAND2_X1 U5284 ( .A1(n6608), .A2(n6607), .ZN(n6606) );
  NAND2_X1 U5285 ( .A1(n4690), .A2(n4692), .ZN(n4688) );
  NAND2_X1 U5286 ( .A1(n6945), .A2(n5088), .ZN(n4690) );
  NAND2_X1 U5287 ( .A1(n4687), .A2(n4333), .ZN(n4686) );
  OR2_X1 U5288 ( .A1(n5004), .A2(n5003), .ZN(n4700) );
  NAND2_X1 U5289 ( .A1(n6606), .A2(n4701), .ZN(n4699) );
  INV_X1 U5290 ( .A(n8633), .ZN(n8680) );
  AND2_X1 U5291 ( .A1(n9879), .A2(n5527), .ZN(n8586) );
  AND2_X1 U5292 ( .A1(n6246), .A2(n5541), .ZN(n8915) );
  OAI21_X1 U5293 ( .B1(n8577), .B2(n8578), .A(n4752), .ZN(n4751) );
  NAND2_X1 U5294 ( .A1(n8584), .A2(n8583), .ZN(n4752) );
  INV_X1 U5295 ( .A(n5519), .ZN(n8588) );
  INV_X1 U5296 ( .A(n8037), .ZN(n8692) );
  OR2_X1 U5297 ( .A1(n5521), .A2(n6180), .ZN(n5478) );
  INV_X1 U5298 ( .A(n8837), .ZN(n8882) );
  INV_X1 U5299 ( .A(n8025), .ZN(n8881) );
  INV_X1 U5300 ( .A(n7210), .ZN(n8704) );
  INV_X1 U5301 ( .A(n6854), .ZN(n8708) );
  NAND2_X1 U5302 ( .A1(n4956), .A2(n6599), .ZN(n4831) );
  NAND2_X1 U5303 ( .A1(n4955), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5304 ( .A1(n4955), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4906) );
  NOR2_X1 U5305 ( .A1(n6363), .A2(n6362), .ZN(n6510) );
  NAND2_X1 U5306 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  OR2_X1 U5307 ( .A1(n7979), .A2(n7977), .ZN(n4435) );
  OR2_X1 U5308 ( .A1(n7978), .A2(n9871), .ZN(n4434) );
  AOI21_X1 U5309 ( .B1(n7980), .B2(n4440), .A(n8379), .ZN(n4439) );
  INV_X1 U5310 ( .A(n4441), .ZN(n4440) );
  OAI21_X1 U5311 ( .B1(n7981), .B2(n9871), .A(n9869), .ZN(n4441) );
  OAI21_X1 U5312 ( .B1(n8745), .B2(n4413), .A(n7982), .ZN(n4437) );
  NAND2_X1 U5313 ( .A1(n8950), .A2(n6814), .ZN(n4410) );
  NAND2_X1 U5314 ( .A1(n8363), .A2(n4359), .ZN(n8948) );
  NAND2_X1 U5315 ( .A1(n8799), .A2(n8030), .ZN(n8784) );
  NAND2_X1 U5316 ( .A1(n4563), .A2(n4561), .ZN(n8959) );
  AOI21_X1 U5317 ( .B1(n8694), .B2(n8917), .A(n4562), .ZN(n4561) );
  OAI21_X1 U5318 ( .B1(n8786), .B2(n4564), .A(n8920), .ZN(n4563) );
  NOR2_X1 U5319 ( .A1(n8822), .A2(n8861), .ZN(n4562) );
  OR2_X1 U5320 ( .A1(n6231), .A2(n4939), .ZN(n4416) );
  INV_X1 U5321 ( .A(n6814), .ZN(n8850) );
  NAND2_X1 U5322 ( .A1(n8933), .A2(n6824), .ZN(n8924) );
  NAND2_X1 U5323 ( .A1(n9963), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4678) );
  XNOR2_X1 U5324 ( .A(n8038), .B(n8565), .ZN(n8947) );
  INV_X1 U5325 ( .A(n7078), .ZN(n9830) );
  OR2_X1 U5326 ( .A1(n9307), .A2(n6147), .ZN(n6100) );
  NAND2_X1 U5327 ( .A1(n5854), .A2(n5853), .ZN(n9570) );
  INV_X1 U5328 ( .A(n6134), .ZN(n9065) );
  OR2_X1 U5329 ( .A1(n6653), .A2(n6654), .ZN(n4582) );
  INV_X1 U5330 ( .A(n4581), .ZN(n6655) );
  NAND2_X1 U5331 ( .A1(n5815), .A2(n5814), .ZN(n9574) );
  INV_X1 U5332 ( .A(n9446), .ZN(n9635) );
  AND4_X1 U5333 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n7378)
         );
  NAND2_X1 U5334 ( .A1(n5963), .A2(n5962), .ZN(n9537) );
  NAND2_X1 U5335 ( .A1(n6054), .A2(n6053), .ZN(n9352) );
  OR2_X1 U5336 ( .A1(n9331), .A2(n6147), .ZN(n6054) );
  INV_X1 U5337 ( .A(n9162), .ZN(n9447) );
  NAND2_X1 U5338 ( .A1(n9757), .A2(n9758), .ZN(n6451) );
  AND2_X1 U5339 ( .A1(n8003), .A2(n8002), .ZN(n9495) );
  NAND2_X1 U5340 ( .A1(n4816), .A2(n4814), .ZN(n9297) );
  NAND2_X1 U5341 ( .A1(n4816), .A2(n4820), .ZN(n9295) );
  NAND2_X1 U5342 ( .A1(n8418), .A2(n4500), .ZN(n8472) );
  AOI21_X1 U5343 ( .B1(n4502), .B2(n8570), .A(n4501), .ZN(n4500) );
  NAND2_X1 U5344 ( .A1(n8417), .A2(n8423), .ZN(n4502) );
  NOR2_X1 U5345 ( .A1(n8419), .A2(n8570), .ZN(n4501) );
  INV_X1 U5346 ( .A(n8502), .ZN(n4508) );
  AND2_X1 U5347 ( .A1(n4510), .A2(n8502), .ZN(n4509) );
  INV_X1 U5348 ( .A(n8497), .ZN(n4510) );
  NOR2_X1 U5349 ( .A1(n4463), .A2(n4460), .ZN(n4459) );
  OR2_X1 U5350 ( .A1(n4464), .A2(n4374), .ZN(n4460) );
  INV_X1 U5351 ( .A(n8114), .ZN(n4463) );
  NOR2_X1 U5352 ( .A1(n4347), .A2(n4474), .ZN(n4473) );
  AND2_X1 U5353 ( .A1(n8133), .A2(n4475), .ZN(n4474) );
  INV_X1 U5354 ( .A(n8119), .ZN(n8118) );
  INV_X1 U5355 ( .A(n4473), .ZN(n4470) );
  AND2_X1 U5356 ( .A1(n5366), .A2(n4714), .ZN(n4713) );
  NAND2_X1 U5357 ( .A1(n4715), .A2(n8622), .ZN(n4714) );
  INV_X1 U5358 ( .A(n8622), .ZN(n4716) );
  AND2_X1 U5359 ( .A1(n9298), .A2(n8158), .ZN(n4447) );
  AOI21_X1 U5360 ( .B1(n4468), .B2(n4471), .A(n4467), .ZN(n4466) );
  OR2_X1 U5361 ( .A1(n9435), .A2(n9428), .ZN(n7697) );
  AOI21_X1 U5362 ( .B1(n4742), .B2(n5227), .A(n4740), .ZN(n4739) );
  INV_X1 U5363 ( .A(n5251), .ZN(n4740) );
  INV_X1 U5364 ( .A(SI_16_), .ZN(n5232) );
  NAND2_X1 U5365 ( .A1(n4746), .A2(n5023), .ZN(n4511) );
  INV_X1 U5366 ( .A(n5008), .ZN(n4746) );
  NAND2_X1 U5367 ( .A1(n5216), .A2(n4721), .ZN(n4720) );
  INV_X1 U5368 ( .A(n5192), .ZN(n4721) );
  INV_X1 U5369 ( .A(n7595), .ZN(n4722) );
  AND2_X1 U5370 ( .A1(n9627), .A2(n4395), .ZN(n4840) );
  NAND2_X1 U5371 ( .A1(n8941), .A2(n8755), .ZN(n8571) );
  AOI21_X1 U5372 ( .B1(n4498), .B2(n4497), .A(n4496), .ZN(n8574) );
  AND2_X1 U5373 ( .A1(n8565), .A2(n8564), .ZN(n4497) );
  XNOR2_X1 U5374 ( .A(n6394), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U5375 ( .A1(n7417), .A2(n4420), .ZN(n7970) );
  NAND2_X1 U5376 ( .A1(n7196), .A2(n4421), .ZN(n4420) );
  AND2_X1 U5377 ( .A1(n8942), .A2(n8037), .ZN(n8051) );
  AND2_X1 U5378 ( .A1(n8043), .A2(n8692), .ZN(n8368) );
  AND2_X1 U5379 ( .A1(n8562), .A2(n8563), .ZN(n8405) );
  NOR2_X1 U5380 ( .A1(n4557), .A2(n4836), .ZN(n4556) );
  NAND2_X1 U5381 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  INV_X1 U5382 ( .A(n8537), .ZN(n4554) );
  INV_X1 U5383 ( .A(n4557), .ZN(n4555) );
  NAND2_X1 U5384 ( .A1(n8048), .A2(n4671), .ZN(n4666) );
  NOR2_X1 U5385 ( .A1(n4544), .A2(n4550), .ZN(n4543) );
  INV_X1 U5386 ( .A(n4547), .ZN(n4544) );
  INV_X1 U5387 ( .A(n7940), .ZN(n4662) );
  NAND2_X1 U5388 ( .A1(n4550), .A2(n4548), .ZN(n4547) );
  INV_X1 U5389 ( .A(n4837), .ZN(n4548) );
  AND2_X1 U5390 ( .A1(n4352), .A2(n7582), .ZN(n4837) );
  AND2_X1 U5391 ( .A1(n4352), .A2(n8505), .ZN(n8504) );
  INV_X1 U5392 ( .A(n4538), .ZN(n4537) );
  OAI21_X1 U5393 ( .B1(n4540), .B2(n4539), .A(n8489), .ZN(n4538) );
  INV_X1 U5394 ( .A(n8484), .ZN(n4539) );
  AND2_X1 U5395 ( .A1(n8478), .A2(n4348), .ZN(n4540) );
  AND2_X1 U5396 ( .A1(n4658), .A2(n4325), .ZN(n4653) );
  OR2_X1 U5397 ( .A1(n8711), .A2(n9905), .ZN(n8424) );
  NAND2_X1 U5398 ( .A1(n4829), .A2(n4828), .ZN(n8428) );
  INV_X1 U5399 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4892) );
  OR2_X1 U5400 ( .A1(n7179), .A2(n7178), .ZN(n4598) );
  INV_X1 U5401 ( .A(n9640), .ZN(n4580) );
  INV_X1 U5402 ( .A(n9078), .ZN(n4575) );
  AND2_X1 U5403 ( .A1(n8172), .A2(n4444), .ZN(n8165) );
  NOR2_X1 U5404 ( .A1(n8164), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U5405 ( .A1(n8289), .A2(n8160), .ZN(n4445) );
  NOR2_X1 U5406 ( .A1(n7169), .A2(n4644), .ZN(n9213) );
  AND2_X1 U5407 ( .A1(n7170), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4644) );
  OR2_X1 U5408 ( .A1(n9505), .A2(n9071), .ZN(n8179) );
  INV_X1 U5409 ( .A(n7734), .ZN(n4626) );
  AND2_X1 U5410 ( .A1(n4800), .A2(n4345), .ZN(n4799) );
  NAND2_X1 U5411 ( .A1(n4326), .A2(n9419), .ZN(n4482) );
  OAI21_X1 U5412 ( .B1(n7701), .B2(n4776), .A(n7704), .ZN(n4775) );
  NOR2_X1 U5413 ( .A1(n4489), .A2(n7155), .ZN(n7286) );
  OR2_X1 U5414 ( .A1(n4490), .A2(n9616), .ZN(n4489) );
  NAND2_X1 U5415 ( .A1(n4491), .A2(n9842), .ZN(n4490) );
  INV_X1 U5416 ( .A(n4492), .ZN(n4491) );
  AND2_X1 U5417 ( .A1(n7060), .A2(n7058), .ZN(n8276) );
  NAND2_X1 U5418 ( .A1(n9207), .A2(n9823), .ZN(n8271) );
  NOR2_X1 U5419 ( .A1(n4784), .A2(n4783), .ZN(n4782) );
  OR2_X1 U5420 ( .A1(n5709), .A2(n5697), .ZN(n5699) );
  NAND2_X1 U5421 ( .A1(n6717), .A2(n6760), .ZN(n8191) );
  NAND2_X1 U5422 ( .A1(n4819), .A2(n9483), .ZN(n7746) );
  NAND2_X1 U5423 ( .A1(n7653), .A2(n8103), .ZN(n7663) );
  INV_X1 U5424 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5583) );
  INV_X1 U5425 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5426 ( .B1(n4766), .B2(n4767), .A(n5460), .ZN(n4765) );
  OR2_X1 U5427 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  AND2_X1 U5428 ( .A1(n6088), .A2(n5465), .ZN(n6086) );
  NAND2_X1 U5429 ( .A1(n5570), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5572) );
  INV_X1 U5430 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5569) );
  INV_X1 U5431 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5571) );
  OAI21_X1 U5432 ( .B1(n4771), .B2(n4770), .A(n5330), .ZN(n4769) );
  INV_X1 U5433 ( .A(n5331), .ZN(n4770) );
  NOR2_X1 U5434 ( .A1(n5308), .A2(n4772), .ZN(n4771) );
  INV_X1 U5435 ( .A(n5285), .ZN(n4772) );
  INV_X1 U5436 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U5437 ( .A1(n4743), .A2(n5199), .ZN(n4742) );
  INV_X1 U5438 ( .A(n5228), .ZN(n4743) );
  INV_X1 U5439 ( .A(n5227), .ZN(n4741) );
  AND2_X1 U5440 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  AOI21_X1 U5441 ( .B1(n4757), .B2(n4759), .A(n4368), .ZN(n4756) );
  NAND2_X1 U5442 ( .A1(n5053), .A2(n5052), .ZN(n5069) );
  NAND3_X1 U5443 ( .A1(n4762), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4411) );
  INV_X1 U5444 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4762) );
  OR2_X1 U5445 ( .A1(n5272), .A2(n8681), .ZN(n5298) );
  NAND2_X1 U5446 ( .A1(n5296), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5318) );
  INV_X1 U5447 ( .A(n5298), .ZN(n5296) );
  OR2_X1 U5448 ( .A1(n5318), .A2(n5317), .ZN(n5337) );
  AOI21_X1 U5449 ( .B1(n4684), .B2(n4683), .A(n4369), .ZN(n4682) );
  NAND2_X1 U5450 ( .A1(n5218), .A2(n5217), .ZN(n5245) );
  INV_X1 U5451 ( .A(n5221), .ZN(n5218) );
  AND2_X1 U5452 ( .A1(n5524), .A2(n5523), .ZN(n6341) );
  NOR2_X1 U5453 ( .A1(n8641), .A2(n5242), .ZN(n4708) );
  NAND2_X1 U5454 ( .A1(n8382), .A2(n8381), .ZN(n8583) );
  INV_X1 U5455 ( .A(n6285), .ZN(n8580) );
  INV_X1 U5456 ( .A(n5516), .ZN(n8579) );
  NAND2_X1 U5457 ( .A1(n4964), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4907) );
  AND2_X1 U5458 ( .A1(n4428), .A2(n4427), .ZN(n6385) );
  NOR2_X1 U5459 ( .A1(n9876), .A2(n9966), .ZN(n4427) );
  INV_X1 U5460 ( .A(n4428), .ZN(n4425) );
  AOI21_X1 U5461 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6367), .A(n6385), .ZN(
        n6504) );
  AOI21_X1 U5462 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6507), .A(n6502), .ZN(
        n6462) );
  NOR2_X1 U5463 ( .A1(n6417), .A2(n4419), .ZN(n6486) );
  AND2_X1 U5464 ( .A1(n6356), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4419) );
  AOI21_X1 U5465 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6377), .A(n6395), .ZN(
        n6408) );
  NOR2_X1 U5466 ( .A1(n6787), .A2(n4443), .ZN(n6791) );
  AND2_X1 U5467 ( .A1(n6788), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5468 ( .A1(n7041), .A2(n7040), .ZN(n7086) );
  NAND2_X1 U5469 ( .A1(n7089), .A2(n7088), .ZN(n7197) );
  NAND2_X1 U5470 ( .A1(n7197), .A2(n4422), .ZN(n7199) );
  NAND2_X1 U5471 ( .A1(n7092), .A2(n7778), .ZN(n4422) );
  NAND2_X1 U5472 ( .A1(n7199), .A2(n7200), .ZN(n7417) );
  NAND2_X1 U5473 ( .A1(n8713), .A2(n7974), .ZN(n8734) );
  NOR2_X1 U5474 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  AOI21_X1 U5475 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8732), .A(n8733), .ZN(
        n8743) );
  NOR2_X1 U5476 ( .A1(n9627), .A2(n4518), .ZN(n4517) );
  INV_X1 U5477 ( .A(n8368), .ZN(n8567) );
  INV_X1 U5478 ( .A(n4518), .ZN(n4516) );
  OR2_X1 U5479 ( .A1(n8954), .A2(n8694), .ZN(n8032) );
  AOI21_X1 U5480 ( .B1(n4319), .B2(n8788), .A(n4372), .ZN(n4841) );
  INV_X1 U5481 ( .A(n8405), .ZN(n8559) );
  NAND2_X1 U5482 ( .A1(n8783), .A2(n8031), .ZN(n8768) );
  NAND2_X1 U5483 ( .A1(n8039), .A2(n8775), .ZN(n8031) );
  AND2_X1 U5484 ( .A1(n8787), .A2(n8788), .ZN(n4564) );
  NAND2_X1 U5485 ( .A1(n8800), .A2(n8802), .ZN(n8799) );
  NAND2_X1 U5486 ( .A1(n4552), .A2(n4553), .ZN(n8819) );
  AND2_X1 U5487 ( .A1(n5428), .A2(n5427), .ZN(n8822) );
  AND2_X1 U5488 ( .A1(n5361), .A2(n5360), .ZN(n8837) );
  AND2_X1 U5489 ( .A1(n8832), .A2(n8537), .ZN(n8835) );
  AND3_X1 U5490 ( .A1(n5341), .A2(n5340), .A3(n5339), .ZN(n8862) );
  NAND2_X1 U5491 ( .A1(n8904), .A2(n4320), .ZN(n8872) );
  OAI21_X1 U5492 ( .B1(n8024), .B2(n8023), .A(n8022), .ZN(n8887) );
  NAND2_X1 U5493 ( .A1(n8904), .A2(n7947), .ZN(n8892) );
  INV_X1 U5494 ( .A(n7952), .ZN(n8401) );
  NAND2_X1 U5495 ( .A1(n7583), .A2(n4837), .ZN(n4551) );
  NAND2_X1 U5496 ( .A1(n4551), .A2(n4550), .ZN(n8911) );
  NAND2_X1 U5497 ( .A1(n7608), .A2(n7577), .ZN(n7579) );
  INV_X1 U5498 ( .A(n8504), .ZN(n7605) );
  NAND2_X1 U5499 ( .A1(n7429), .A2(n4358), .ZN(n7444) );
  INV_X1 U5500 ( .A(n8489), .ZN(n8396) );
  AND2_X1 U5501 ( .A1(n8487), .A2(n8480), .ZN(n8489) );
  OAI21_X1 U5502 ( .B1(n7208), .B2(n4539), .A(n4537), .ZN(n7441) );
  NAND2_X1 U5503 ( .A1(n4536), .A2(n8484), .ZN(n7442) );
  NAND2_X1 U5504 ( .A1(n7208), .A2(n4540), .ZN(n4536) );
  AND4_X1 U5505 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n7430)
         );
  NOR2_X1 U5506 ( .A1(n9941), .A2(n4523), .ZN(n4522) );
  INV_X1 U5507 ( .A(n4524), .ZN(n4523) );
  AND4_X1 U5508 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n7210)
         );
  NAND2_X1 U5509 ( .A1(n6860), .A2(n4524), .ZN(n7029) );
  NAND2_X1 U5510 ( .A1(n6860), .A2(n9927), .ZN(n7027) );
  AND2_X1 U5511 ( .A1(n8419), .A2(n8423), .ZN(n8390) );
  AND4_X1 U5512 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n7111)
         );
  AND4_X1 U5513 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n7008)
         );
  NAND2_X1 U5514 ( .A1(n4515), .A2(n9913), .ZN(n6971) );
  NOR2_X1 U5515 ( .A1(n6537), .A2(n4828), .ZN(n6958) );
  NAND2_X1 U5516 ( .A1(n6958), .A2(n9905), .ZN(n6957) );
  NAND2_X1 U5517 ( .A1(n8428), .A2(n8448), .ZN(n6540) );
  INV_X1 U5518 ( .A(n6542), .ZN(n8383) );
  NAND2_X1 U5519 ( .A1(n6280), .A2(n8379), .ZN(n7609) );
  NAND2_X1 U5520 ( .A1(n5180), .A2(n5179), .ZN(n9020) );
  INV_X1 U5521 ( .A(n9897), .ZN(n9955) );
  INV_X1 U5522 ( .A(n9898), .ZN(n9957) );
  INV_X1 U5523 ( .A(n6429), .ZN(n6805) );
  AND2_X1 U5524 ( .A1(n6808), .A2(n6275), .ZN(n6430) );
  INV_X1 U5525 ( .A(n5510), .ZN(n9878) );
  NOR2_X1 U5526 ( .A1(n4529), .A2(n4525), .ZN(n4871) );
  XNOR2_X1 U5527 ( .A(n5514), .B(n5513), .ZN(n6242) );
  NAND2_X1 U5528 ( .A1(n4891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5269) );
  AND3_X1 U5529 ( .A1(n4882), .A2(n5205), .A3(n5176), .ZN(n4883) );
  AND2_X1 U5530 ( .A1(n5062), .A2(n5097), .ZN(n6511) );
  AND2_X1 U5531 ( .A1(n4927), .A2(n4865), .ZN(n4975) );
  NAND2_X1 U5532 ( .A1(n4599), .A2(n4597), .ZN(n4596) );
  NOR2_X1 U5533 ( .A1(n5721), .A2(n4859), .ZN(n5726) );
  INV_X1 U5534 ( .A(n9352), .ZN(n9068) );
  INV_X1 U5535 ( .A(n4589), .ZN(n4588) );
  OAI21_X1 U5536 ( .B1(n4593), .B2(n4590), .A(n5862), .ZN(n4589) );
  NAND2_X1 U5537 ( .A1(n5873), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U5538 ( .A1(n4569), .A2(n4573), .ZN(n4577) );
  NAND2_X1 U5539 ( .A1(n6008), .A2(n4575), .ZN(n4573) );
  NAND3_X1 U5540 ( .A1(n9147), .A2(n6007), .A3(n4574), .ZN(n4569) );
  OR2_X1 U5541 ( .A1(n6008), .A2(n4575), .ZN(n4574) );
  AOI21_X1 U5542 ( .B1(n7295), .B2(n5747), .A(n5746), .ZN(n7400) );
  INV_X1 U5543 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5751) );
  OR2_X1 U5544 ( .A1(n5952), .A2(n9135), .ZN(n5973) );
  INV_X1 U5545 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U5546 ( .A1(n5914), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5932) );
  INV_X1 U5547 ( .A(n5916), .ZN(n5914) );
  OR2_X1 U5548 ( .A1(n5894), .A2(n5893), .ZN(n5916) );
  INV_X1 U5549 ( .A(n9632), .ZN(n9160) );
  NAND2_X1 U5550 ( .A1(n4600), .A2(n6198), .ZN(n7225) );
  OR2_X1 U5551 ( .A1(n6200), .A2(n6197), .ZN(n4600) );
  OR2_X1 U5552 ( .A1(n8061), .A2(n6139), .ZN(n6741) );
  INV_X1 U5553 ( .A(n5644), .ZN(n7742) );
  INV_X1 U5554 ( .A(n6067), .ZN(n6147) );
  AND4_X1 U5555 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n7665)
         );
  INV_X1 U5556 ( .A(n5709), .ZN(n7738) );
  NOR2_X1 U5557 ( .A1(n9764), .A2(n4646), .ZN(n6454) );
  AND2_X1 U5558 ( .A1(n9769), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4646) );
  NOR2_X1 U5559 ( .A1(n6454), .A2(n6453), .ZN(n6678) );
  NOR2_X1 U5560 ( .A1(n6678), .A2(n4645), .ZN(n9781) );
  AND2_X1 U5561 ( .A1(n6679), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4645) );
  NAND2_X1 U5562 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  NOR2_X1 U5563 ( .A1(n6773), .A2(n4396), .ZN(n6777) );
  NOR2_X1 U5564 ( .A1(n6777), .A2(n6776), .ZN(n7169) );
  XNOR2_X1 U5565 ( .A(n9213), .B(n9212), .ZN(n7172) );
  NOR2_X1 U5566 ( .A1(n9265), .A2(n4650), .ZN(n9268) );
  AND2_X1 U5567 ( .A1(n9266), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5568 ( .A1(n9268), .A2(n9267), .ZN(n9274) );
  XNOR2_X1 U5569 ( .A(n4648), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9282) );
  OR2_X1 U5570 ( .A1(n9274), .A2(n4649), .ZN(n4648) );
  AND2_X1 U5571 ( .A1(n9276), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4649) );
  INV_X1 U5572 ( .A(SI_21_), .ZN(n7919) );
  NAND2_X1 U5573 ( .A1(n9329), .A2(n4821), .ZN(n9317) );
  AND2_X1 U5574 ( .A1(n8254), .A2(n9322), .ZN(n9336) );
  AND2_X1 U5575 ( .A1(n8253), .A2(n8249), .ZN(n9350) );
  INV_X1 U5576 ( .A(n9350), .ZN(n9342) );
  NAND2_X1 U5577 ( .A1(n9379), .A2(n8245), .ZN(n9364) );
  INV_X1 U5578 ( .A(n9371), .ZN(n7733) );
  AOI21_X1 U5579 ( .B1(n9406), .B2(n7732), .A(n8242), .ZN(n4863) );
  NAND2_X1 U5580 ( .A1(n4863), .A2(n7733), .ZN(n9379) );
  NAND2_X1 U5581 ( .A1(n7730), .A2(n8298), .ZN(n9407) );
  AND2_X1 U5582 ( .A1(n8239), .A2(n9390), .ZN(n9408) );
  NOR2_X1 U5583 ( .A1(n9457), .A2(n9552), .ZN(n9432) );
  NAND2_X1 U5584 ( .A1(n8126), .A2(n8122), .ZN(n9452) );
  INV_X1 U5585 ( .A(n4495), .ZN(n4493) );
  NAND2_X1 U5586 ( .A1(n9638), .A2(n4495), .ZN(n4494) );
  NAND2_X1 U5587 ( .A1(n7626), .A2(n8322), .ZN(n9480) );
  AND2_X1 U5588 ( .A1(n5871), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U5589 ( .A1(n4786), .A2(n4785), .ZN(n7662) );
  AOI21_X1 U5590 ( .B1(n4329), .B2(n4790), .A(n4384), .ZN(n4785) );
  NOR2_X1 U5591 ( .A1(n7649), .A2(n9570), .ZN(n7631) );
  AND2_X1 U5592 ( .A1(n4614), .A2(n8315), .ZN(n4613) );
  NAND2_X1 U5593 ( .A1(n4615), .A2(n4618), .ZN(n4614) );
  NOR2_X1 U5594 ( .A1(n7481), .A2(n9574), .ZN(n7529) );
  OAI21_X1 U5595 ( .B1(n7308), .B2(n4618), .A(n4615), .ZN(n7519) );
  INV_X1 U5596 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5788) );
  NOR2_X1 U5597 ( .A1(n5789), .A2(n5788), .ZN(n5816) );
  AOI21_X1 U5598 ( .B1(n7306), .B2(n7307), .A(n7279), .ZN(n7471) );
  OR2_X1 U5599 ( .A1(n5770), .A2(n6443), .ZN(n5789) );
  NOR2_X1 U5600 ( .A1(n7155), .A2(n4492), .ZN(n7335) );
  NAND2_X1 U5601 ( .A1(n7061), .A2(n7060), .ZN(n8197) );
  INV_X1 U5602 ( .A(n8311), .ZN(n8075) );
  OR2_X1 U5603 ( .A1(n7153), .A2(n7157), .ZN(n7155) );
  AND2_X1 U5604 ( .A1(n8073), .A2(n8271), .ZN(n8305) );
  AND4_X1 U5605 ( .A1(n5617), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(n7298)
         );
  OAI211_X1 U5606 ( .C1(n7063), .C2(n7059), .A(n4453), .B(n8306), .ZN(n7148)
         );
  INV_X1 U5607 ( .A(n4455), .ZN(n4454) );
  NOR2_X1 U5608 ( .A1(n6939), .A2(n6993), .ZN(n6938) );
  NAND2_X1 U5609 ( .A1(n7063), .A2(n7057), .ZN(n6931) );
  NAND2_X1 U5610 ( .A1(n6929), .A2(n8304), .ZN(n6928) );
  NAND2_X1 U5611 ( .A1(n6911), .A2(n6899), .ZN(n6929) );
  AND4_X1 U5612 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n6913)
         );
  AND4_X1 U5613 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(n6912)
         );
  NAND2_X1 U5614 ( .A1(n6736), .A2(n6719), .ZN(n6720) );
  AND4_X1 U5615 ( .A1(n4376), .A2(n4480), .A3(n5641), .A4(n5631), .ZN(n4478)
         );
  NAND2_X1 U5616 ( .A1(n8193), .A2(n8195), .ZN(n8303) );
  AND4_X1 U5617 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n6930)
         );
  NAND2_X1 U5618 ( .A1(n6031), .A2(n6030), .ZN(n9523) );
  NAND2_X1 U5619 ( .A1(n5892), .A2(n5891), .ZN(n9565) );
  NAND2_X1 U5620 ( .A1(n6137), .A2(n6131), .ZN(n9615) );
  AND2_X1 U5621 ( .A1(n6723), .A2(n8295), .ZN(n9655) );
  INV_X1 U5622 ( .A(n9615), .ZN(n9841) );
  AND3_X1 U5623 ( .A1(n4340), .A2(n5631), .A3(n4476), .ZN(n6896) );
  XNOR2_X1 U5624 ( .A(n6127), .B(n4632), .ZN(n6210) );
  XNOR2_X1 U5625 ( .A(n8004), .B(SI_30_), .ZN(n8371) );
  NAND2_X1 U5626 ( .A1(n5583), .A2(n5559), .ZN(n4811) );
  NAND4_X1 U5627 ( .A1(n4321), .A2(n4847), .A3(n5551), .A4(n4450), .ZN(n5558)
         );
  NOR2_X1 U5628 ( .A1(n4361), .A2(n5686), .ZN(n4450) );
  XNOR2_X1 U5629 ( .A(n7723), .B(n7722), .ZN(n9056) );
  XNOR2_X1 U5630 ( .A(n6087), .B(n6086), .ZN(n7547) );
  INV_X1 U5631 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U5632 ( .A1(n5572), .A2(n5571), .ZN(n5603) );
  XNOR2_X1 U5633 ( .A(n5608), .B(P1_IR_REG_19__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U5634 ( .A1(n4773), .A2(n5285), .ZN(n5309) );
  INV_X1 U5635 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U5636 ( .A(n5268), .B(n5263), .ZN(n6666) );
  INV_X1 U5637 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5867) );
  INV_X1 U5638 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5865) );
  INV_X1 U5639 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5552) );
  AND2_X1 U5640 ( .A1(n5618), .A2(n5551), .ZN(n5812) );
  NAND2_X1 U5641 ( .A1(n4761), .A2(n5117), .ZN(n5131) );
  NAND2_X1 U5642 ( .A1(n5116), .A2(n4856), .ZN(n4761) );
  NAND2_X1 U5643 ( .A1(n4974), .A2(n4973), .ZN(n4989) );
  NOR2_X2 U5644 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5630) );
  NOR2_X1 U5645 ( .A1(n10015), .A2(n7357), .ZN(n7358) );
  NAND2_X1 U5646 ( .A1(n4696), .A2(n5022), .ZN(n4695) );
  INV_X1 U5647 ( .A(n4697), .ZN(n4696) );
  AND4_X1 U5648 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n6970)
         );
  AND4_X1 U5649 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n7023)
         );
  NAND2_X1 U5650 ( .A1(n6164), .A2(n5484), .ZN(n4710) );
  NOR2_X1 U5651 ( .A1(n5485), .A2(n5483), .ZN(n5484) );
  AND4_X1 U5652 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n8499)
         );
  NOR2_X1 U5653 ( .A1(n6866), .A2(n5089), .ZN(n6946) );
  AOI21_X1 U5654 ( .B1(n4705), .B2(n4707), .A(n4354), .ZN(n4703) );
  NAND2_X1 U5655 ( .A1(n6173), .A2(n6172), .ZN(n8949) );
  NAND2_X1 U5656 ( .A1(n4926), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5657 ( .A1(n4349), .A2(n4727), .ZN(n4726) );
  INV_X1 U5658 ( .A(n9956), .ZN(n7270) );
  AND4_X1 U5659 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n8646)
         );
  NAND2_X1 U5660 ( .A1(n7678), .A2(n5243), .ZN(n8642) );
  NOR2_X1 U5661 ( .A1(n6868), .A2(n6867), .ZN(n6866) );
  NAND2_X1 U5662 ( .A1(n5316), .A2(n5315), .ZN(n8990) );
  NAND2_X1 U5663 ( .A1(n5168), .A2(n5167), .ZN(n9025) );
  NAND2_X1 U5664 ( .A1(n8621), .A2(n8622), .ZN(n8666) );
  NAND2_X1 U5665 ( .A1(n6343), .A2(n4334), .ZN(n6472) );
  AND2_X1 U5666 ( .A1(n8634), .A2(n8917), .ZN(n8682) );
  AND2_X1 U5667 ( .A1(n8634), .A2(n8915), .ZN(n8623) );
  AND4_X1 U5668 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n8686)
         );
  NAND2_X1 U5669 ( .A1(n4704), .A2(n5262), .ZN(n8679) );
  NAND2_X1 U5670 ( .A1(n7678), .A2(n4708), .ZN(n4704) );
  AND4_X1 U5671 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n7600)
         );
  NAND2_X1 U5672 ( .A1(n7491), .A2(n4724), .ZN(n7594) );
  NAND2_X1 U5673 ( .A1(n4717), .A2(n5216), .ZN(n7593) );
  NAND2_X1 U5674 ( .A1(n7491), .A2(n5192), .ZN(n4717) );
  NAND2_X1 U5675 ( .A1(n5210), .A2(n5209), .ZN(n9015) );
  AOI21_X1 U5676 ( .B1(n5383), .B2(n4956), .A(n5382), .ZN(n8864) );
  INV_X1 U5677 ( .A(n8862), .ZN(n8897) );
  INV_X1 U5678 ( .A(n8661), .ZN(n8918) );
  INV_X1 U5679 ( .A(n8499), .ZN(n8700) );
  INV_X1 U5680 ( .A(n7430), .ZN(n8702) );
  INV_X1 U5681 ( .A(P2_U3966), .ZN(n8712) );
  INV_X1 U5682 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4878) );
  NOR2_X1 U5683 ( .A1(n7977), .A2(n4423), .ZN(n6387) );
  NAND2_X1 U5684 ( .A1(n4426), .A2(n4424), .ZN(n4423) );
  NAND2_X1 U5685 ( .A1(n4425), .A2(n6386), .ZN(n4424) );
  INV_X1 U5686 ( .A(n6385), .ZN(n4426) );
  INV_X1 U5687 ( .A(n4418), .ZN(n6397) );
  NOR2_X1 U5688 ( .A1(n6406), .A2(n4431), .ZN(n6363) );
  AND2_X1 U5689 ( .A1(n6365), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4431) );
  INV_X1 U5690 ( .A(n4430), .ZN(n6514) );
  AOI21_X1 U5691 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n6626), .A(n6622), .ZN(
        n6625) );
  OAI21_X1 U5692 ( .B1(n9048), .B2(n8377), .A(n4747), .ZN(n8941) );
  NOR2_X1 U5693 ( .A1(n6244), .A2(n4748), .ZN(n4747) );
  AND2_X1 U5694 ( .A1(n8377), .A2(n4749), .ZN(n4748) );
  INV_X1 U5695 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n4749) );
  XNOR2_X1 U5696 ( .A(n8760), .B(n8941), .ZN(n8938) );
  NAND2_X1 U5697 ( .A1(n4843), .A2(n4319), .ZN(n8778) );
  NAND2_X1 U5698 ( .A1(n5419), .A2(n5418), .ZN(n8965) );
  NAND2_X1 U5699 ( .A1(n4670), .A2(n4668), .ZN(n8831) );
  NAND2_X1 U5700 ( .A1(n4670), .A2(n4671), .ZN(n8829) );
  NAND2_X1 U5701 ( .A1(n5375), .A2(n5374), .ZN(n8848) );
  CLKBUF_X1 U5702 ( .A(n8044), .Z(n7951) );
  NAND2_X1 U5703 ( .A1(n7941), .A2(n7940), .ZN(n8902) );
  NAND2_X1 U5704 ( .A1(n5239), .A2(n5238), .ZN(n9010) );
  AND2_X1 U5705 ( .A1(n7213), .A2(n7212), .ZN(n7214) );
  NAND2_X1 U5706 ( .A1(n7019), .A2(n7004), .ZN(n7005) );
  NAND2_X1 U5707 ( .A1(n4654), .A2(n4655), .ZN(n6845) );
  OR2_X1 U5708 ( .A1(n6956), .A2(n4658), .ZN(n4654) );
  NAND2_X1 U5709 ( .A1(n4826), .A2(n8426), .ZN(n6832) );
  NAND2_X1 U5710 ( .A1(n6831), .A2(n8449), .ZN(n4826) );
  NAND2_X1 U5711 ( .A1(n6954), .A2(n6581), .ZN(n6829) );
  NAND2_X1 U5712 ( .A1(n9879), .A2(n6810), .ZN(n8844) );
  INV_X1 U5713 ( .A(n6809), .ZN(n6810) );
  NAND2_X1 U5714 ( .A1(n6981), .A2(n4331), .ZN(n6982) );
  INV_X1 U5715 ( .A(n8844), .ZN(n8929) );
  INV_X1 U5716 ( .A(n8908), .ZN(n8926) );
  INV_X1 U5717 ( .A(n8946), .ZN(n4674) );
  AND2_X2 U5718 ( .A1(n6430), .A2(n6429), .ZN(n9983) );
  OAI21_X1 U5719 ( .B1(n8962), .B2(n9890), .A(n4566), .ZN(n4565) );
  NOR2_X1 U5720 ( .A1(n8960), .A2(n4567), .ZN(n4566) );
  AND2_X1 U5721 ( .A1(n8961), .A2(n9897), .ZN(n4567) );
  AND2_X1 U5722 ( .A1(n6242), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9885) );
  INV_X1 U5723 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U5724 ( .A1(n4560), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4901) );
  INV_X1 U5725 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U5726 ( .A1(n5498), .A2(n5497), .ZN(n7546) );
  INV_X1 U5727 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U5728 ( .A1(n5493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5729 ( .A1(n5514), .A2(n5513), .ZN(n5493) );
  INV_X1 U5730 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7244) );
  INV_X1 U5731 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8021) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7854) );
  AOI21_X1 U5733 ( .B1(n4896), .B2(n4895), .A(n9049), .ZN(n4729) );
  INV_X1 U5734 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6800) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7863) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6552) );
  INV_X1 U5737 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6499) );
  INV_X1 U5738 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6270) );
  INV_X1 U5739 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4950) );
  NOR2_X1 U5740 ( .A1(n6209), .A2(n7246), .ZN(n6259) );
  AND4_X1 U5741 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n7251)
         );
  INV_X1 U5742 ( .A(n4572), .ZN(n9076) );
  NAND2_X1 U5743 ( .A1(n5997), .A2(n5996), .ZN(n9532) );
  NAND2_X1 U5744 ( .A1(n6688), .A2(n5660), .ZN(n6704) );
  AND2_X1 U5745 ( .A1(n5926), .A2(n5925), .ZN(n9088) );
  INV_X1 U5746 ( .A(n6061), .ZN(n4609) );
  AND2_X1 U5747 ( .A1(n6047), .A2(n6034), .ZN(n9346) );
  NAND2_X1 U5748 ( .A1(n9183), .A2(n9185), .ZN(n9639) );
  AND4_X1 U5749 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n9119)
         );
  INV_X1 U5750 ( .A(n4577), .ZN(n9126) );
  NAND2_X1 U5751 ( .A1(n6011), .A2(n6010), .ZN(n9528) );
  AND4_X1 U5752 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n7236)
         );
  NAND2_X1 U5753 ( .A1(n4603), .A2(n5947), .ZN(n9133) );
  NOR2_X1 U5754 ( .A1(n4592), .A2(n4591), .ZN(n7562) );
  INV_X1 U5755 ( .A(n4594), .ZN(n4591) );
  INV_X1 U5756 ( .A(n4595), .ZN(n4592) );
  INV_X1 U5757 ( .A(n6896), .ZN(n6876) );
  NAND2_X1 U5758 ( .A1(n9115), .A2(n5907), .ZN(n9159) );
  NAND2_X1 U5759 ( .A1(n5913), .A2(n5912), .ZN(n9560) );
  INV_X1 U5760 ( .A(n9650), .ZN(n9164) );
  NAND2_X1 U5761 ( .A1(n9168), .A2(n6061), .ZN(n9172) );
  AND2_X1 U5762 ( .A1(n9646), .A2(n9615), .ZN(n9192) );
  INV_X1 U5763 ( .A(n9176), .ZN(n9366) );
  INV_X1 U5764 ( .A(n9119), .ZN(n9486) );
  INV_X1 U5765 ( .A(n7378), .ZN(n9203) );
  INV_X1 U5766 ( .A(n7251), .ZN(n9205) );
  INV_X1 U5767 ( .A(n6913), .ZN(n9211) );
  INV_X1 U5768 ( .A(n6718), .ZN(n6717) );
  NAND4_X1 U5769 ( .A1(n5648), .A2(n5647), .A3(n5646), .A4(n5645), .ZN(n6750)
         );
  OR2_X1 U5770 ( .A1(n4314), .A2(n5643), .ZN(n5648) );
  NAND2_X1 U5771 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4647) );
  XNOR2_X1 U5772 ( .A(n9682), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9687) );
  INV_X1 U5773 ( .A(n4643), .ZN(n9695) );
  INV_X1 U5774 ( .A(n4641), .ZN(n6331) );
  NOR2_X1 U5775 ( .A1(n6329), .A2(n4338), .ZN(n9713) );
  NAND2_X1 U5776 ( .A1(n9739), .A2(n4381), .ZN(n9757) );
  INV_X1 U5777 ( .A(n9786), .ZN(n9750) );
  INV_X1 U5778 ( .A(n9787), .ZN(n9763) );
  XNOR2_X1 U5779 ( .A(n9495), .B(n4342), .ZN(n9497) );
  NOR2_X1 U5780 ( .A1(n9290), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U5781 ( .A1(n4487), .A2(n4821), .ZN(n4486) );
  NOR2_X1 U5782 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  AOI21_X1 U5783 ( .B1(n9500), .B2(n9441), .A(n7753), .ZN(n7754) );
  AOI21_X1 U5784 ( .B1(n4814), .B2(n4813), .A(n4388), .ZN(n4812) );
  NAND2_X1 U5785 ( .A1(n9327), .A2(n7716), .ZN(n9316) );
  AND2_X1 U5786 ( .A1(n4637), .A2(n4636), .ZN(n9515) );
  AOI21_X1 U5787 ( .B1(n4819), .B2(n9485), .A(n4385), .ZN(n4636) );
  NAND2_X1 U5788 ( .A1(n9325), .A2(n9488), .ZN(n4637) );
  AND2_X1 U5789 ( .A1(n6045), .A2(n6044), .ZN(n9334) );
  INV_X1 U5790 ( .A(n9523), .ZN(n9348) );
  OAI21_X1 U5791 ( .B1(n7708), .B2(n4803), .A(n4800), .ZN(n9357) );
  NAND2_X1 U5792 ( .A1(n4805), .A2(n7709), .ZN(n9372) );
  NAND2_X1 U5793 ( .A1(n7708), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5794 ( .A1(n7708), .A2(n7707), .ZN(n9385) );
  NAND2_X1 U5795 ( .A1(n9429), .A2(n7703), .ZN(n9414) );
  INV_X1 U5796 ( .A(n9565), .ZN(n9478) );
  NAND2_X1 U5797 ( .A1(n5870), .A2(n5869), .ZN(n9193) );
  NAND2_X1 U5798 ( .A1(n4787), .A2(n4788), .ZN(n7648) );
  OR2_X1 U5799 ( .A1(n7526), .A2(n4790), .ZN(n4787) );
  NAND2_X1 U5800 ( .A1(n5834), .A2(n5833), .ZN(n7622) );
  NAND2_X1 U5801 ( .A1(n4792), .A2(n7527), .ZN(n7624) );
  NAND2_X1 U5802 ( .A1(n7526), .A2(n7525), .ZN(n4792) );
  NAND2_X1 U5803 ( .A1(n9313), .A2(n6746), .ZN(n9494) );
  NAND2_X1 U5804 ( .A1(n7308), .A2(n8204), .ZN(n7474) );
  NAND2_X1 U5805 ( .A1(n5622), .A2(n5621), .ZN(n7078) );
  AND2_X1 U5806 ( .A1(n5620), .A2(n4848), .ZN(n5621) );
  NAND2_X1 U5807 ( .A1(n7149), .A2(n7070), .ZN(n7071) );
  AOI21_X1 U5808 ( .B1(n8304), .B2(n4784), .A(n4783), .ZN(n4778) );
  INV_X1 U5809 ( .A(n9494), .ZN(n9456) );
  OR2_X1 U5810 ( .A1(n9805), .A2(n6743), .ZN(n7669) );
  NAND2_X1 U5811 ( .A1(n9313), .A2(n6758), .ZN(n9477) );
  INV_X1 U5812 ( .A(n9477), .ZN(n8017) );
  OR2_X1 U5813 ( .A1(n9504), .A2(n9661), .ZN(n9511) );
  INV_X2 U5814 ( .A(n9849), .ZN(n9850) );
  AND2_X1 U5815 ( .A1(n9804), .A2(n9602), .ZN(n9801) );
  INV_X1 U5816 ( .A(n5594), .ZN(n8366) );
  XNOR2_X1 U5817 ( .A(n7719), .B(n7718), .ZN(n7557) );
  XNOR2_X1 U5818 ( .A(n5578), .B(n5577), .ZN(n7518) );
  NAND2_X1 U5819 ( .A1(n5576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U5820 ( .A(n5582), .B(n5581), .ZN(n7467) );
  INV_X1 U5821 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7320) );
  XNOR2_X1 U5822 ( .A(n5580), .B(n5579), .ZN(n7321) );
  INV_X1 U5823 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7248) );
  AND2_X1 U5824 ( .A1(n8377), .A2(P1_U3084), .ZN(n7556) );
  INV_X1 U5825 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6927) );
  INV_X1 U5826 ( .A(n8340), .ZN(n8295) );
  INV_X1 U5827 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6802) );
  INV_X1 U5828 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6527) );
  INV_X1 U5829 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6271) );
  INV_X1 U5830 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7868) );
  AND2_X1 U5831 ( .A1(n5740), .A2(n5739), .ZN(n9756) );
  XNOR2_X1 U5832 ( .A(n5024), .B(n5023), .ZN(n6231) );
  NAND2_X1 U5833 ( .A1(n4745), .A2(n5008), .ZN(n5024) );
  NOR2_X1 U5834 ( .A1(n7368), .A2(n10021), .ZN(n10011) );
  AOI21_X1 U5835 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10009), .ZN(n10008) );
  NOR2_X1 U5836 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  AOI21_X1 U5837 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10006), .ZN(n10005) );
  OAI21_X1 U5838 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10003), .ZN(n10001) );
  NAND2_X1 U5839 ( .A1(n6606), .A2(n4986), .ZN(n6563) );
  NAND2_X1 U5840 ( .A1(n4686), .A2(n4688), .ZN(n7137) );
  NAND2_X1 U5841 ( .A1(n4699), .A2(n4700), .ZN(n6646) );
  OAI21_X1 U5842 ( .B1(n8039), .B2(n7687), .A(n6168), .ZN(n6169) );
  NAND2_X1 U5843 ( .A1(n4750), .A2(n8589), .ZN(P2_U3244) );
  INV_X1 U5844 ( .A(n4437), .ZN(n4436) );
  INV_X1 U5845 ( .A(n4439), .ZN(n4438) );
  NAND2_X1 U5846 ( .A1(n4433), .A2(n8379), .ZN(n4432) );
  AOI21_X1 U5847 ( .B1(n8948), .B2(n8928), .A(n4408), .ZN(n8365) );
  NAND2_X1 U5848 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  INV_X1 U5849 ( .A(n8364), .ZN(n4409) );
  NAND2_X1 U5850 ( .A1(n9965), .A2(n9962), .ZN(n4679) );
  INV_X1 U5851 ( .A(n4677), .ZN(n4676) );
  INV_X1 U5852 ( .A(n4582), .ZN(n6659) );
  OAI21_X1 U5853 ( .B1(n9515), .B2(n9489), .A(n4633), .ZN(P1_U3264) );
  AOI21_X1 U5854 ( .B1(n9512), .B2(n9492), .A(n4634), .ZN(n4633) );
  OAI21_X1 U5855 ( .B1(n9516), .B2(n9494), .A(n4635), .ZN(n4634) );
  INV_X1 U5856 ( .A(n9326), .ZN(n4635) );
  OR2_X1 U5857 ( .A1(n8941), .A2(n8755), .ZN(n8572) );
  INV_X1 U5858 ( .A(n4790), .ZN(n4789) );
  OR2_X1 U5859 ( .A1(n7623), .A2(n4791), .ZN(n4790) );
  INV_X1 U5860 ( .A(n4995), .ZN(n5381) );
  AND2_X1 U5861 ( .A1(n8555), .A2(n8554), .ZN(n4319) );
  INV_X1 U5862 ( .A(n8304), .ZN(n4780) );
  AND2_X1 U5863 ( .A1(n4520), .A2(n8877), .ZN(n4320) );
  INV_X1 U5864 ( .A(n8820), .ZN(n4558) );
  INV_X1 U5865 ( .A(n4803), .ZN(n4802) );
  OR2_X1 U5866 ( .A1(n7711), .A2(n4804), .ZN(n4803) );
  AND3_X1 U5867 ( .A1(n4631), .A2(n4351), .A3(n4452), .ZN(n4321) );
  NAND2_X1 U5868 ( .A1(n4416), .A2(n5010), .ZN(n6841) );
  INV_X1 U5869 ( .A(n6841), .ZN(n9913) );
  INV_X1 U5870 ( .A(n6594), .ZN(n4828) );
  OR2_X1 U5871 ( .A1(n4857), .A2(n4395), .ZN(n4322) );
  AND2_X1 U5872 ( .A1(n4320), .A2(n4519), .ZN(n4323) );
  AND2_X1 U5873 ( .A1(n9000), .A2(n8698), .ZN(n4324) );
  OR2_X1 U5874 ( .A1(n9913), .A2(n6970), .ZN(n4325) );
  AND2_X1 U5875 ( .A1(n9405), .A2(n4483), .ZN(n4326) );
  NAND2_X1 U5876 ( .A1(n8108), .A2(n8109), .ZN(n4327) );
  AND2_X1 U5877 ( .A1(n5726), .A2(n6198), .ZN(n4328) );
  AND2_X1 U5878 ( .A1(n4788), .A2(n4383), .ZN(n4329) );
  INV_X1 U5879 ( .A(n7525), .ZN(n8315) );
  NAND2_X1 U5880 ( .A1(n6064), .A2(n6063), .ZN(n9513) );
  INV_X1 U5881 ( .A(n9513), .ZN(n4821) );
  NAND2_X1 U5882 ( .A1(n5478), .A2(n5477), .ZN(n8694) );
  AND2_X1 U5883 ( .A1(n6100), .A2(n6099), .ZN(n9071) );
  INV_X1 U5884 ( .A(n9071), .ZN(n4819) );
  NAND2_X1 U5885 ( .A1(n4584), .A2(n4583), .ZN(n4581) );
  NAND2_X1 U5886 ( .A1(n6961), .A2(n8384), .ZN(n6831) );
  OR2_X1 U5887 ( .A1(n7649), .A2(n4493), .ZN(n4330) );
  OR2_X1 U5888 ( .A1(n6980), .A2(n6542), .ZN(n4331) );
  NOR2_X1 U5889 ( .A1(n5558), .A2(n4808), .ZN(n5585) );
  NAND4_X1 U5890 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n6277)
         );
  NAND2_X1 U5891 ( .A1(n4926), .A2(n8001), .ZN(n4939) );
  NAND2_X1 U5892 ( .A1(n8878), .A2(n4835), .ZN(n8832) );
  XNOR2_X1 U5893 ( .A(n4881), .B(n4880), .ZN(n6394) );
  NAND2_X1 U5894 ( .A1(n5949), .A2(n5948), .ZN(n9548) );
  AND2_X1 U5895 ( .A1(n4689), .A2(n4692), .ZN(n4333) );
  OR2_X1 U5896 ( .A1(n4910), .A2(n4911), .ZN(n4334) );
  NAND4_X1 U5897 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n6531)
         );
  AND2_X1 U5898 ( .A1(n7069), .A2(n7067), .ZN(n4335) );
  NOR2_X1 U5899 ( .A1(n7942), .A2(n4662), .ZN(n4661) );
  NOR2_X1 U5900 ( .A1(n5987), .A2(n9098), .ZN(n4336) );
  AND2_X1 U5901 ( .A1(n4607), .A2(n6085), .ZN(n4337) );
  INV_X1 U5902 ( .A(n7108), .ZN(n8391) );
  AND2_X1 U5903 ( .A1(n6320), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4338) );
  AND2_X1 U5904 ( .A1(n8498), .A2(n8570), .ZN(n4339) );
  OR2_X1 U5905 ( .A1(n8002), .A2(n6213), .ZN(n4340) );
  NOR2_X1 U5906 ( .A1(n8985), .A2(n8897), .ZN(n4341) );
  NAND2_X1 U5907 ( .A1(n9329), .A2(n4485), .ZN(n4342) );
  AND2_X1 U5908 ( .A1(n8667), .A2(n8668), .ZN(n4343) );
  INV_X1 U5909 ( .A(n8860), .ZN(n8048) );
  AND2_X1 U5910 ( .A1(n5005), .A2(n5023), .ZN(n4344) );
  INV_X1 U5911 ( .A(n8298), .ZN(n4475) );
  OR2_X1 U5912 ( .A1(n9528), .A2(n9380), .ZN(n4345) );
  AND2_X1 U5913 ( .A1(n8202), .A2(n8171), .ZN(n4346) );
  AND2_X1 U5914 ( .A1(n8201), .A2(n8168), .ZN(n4347) );
  NAND2_X1 U5915 ( .A1(n8878), .A2(n8532), .ZN(n8858) );
  NAND2_X1 U5916 ( .A1(n9956), .A2(n8703), .ZN(n4348) );
  OR2_X1 U5917 ( .A1(n6218), .A2(n8377), .ZN(n4349) );
  AND3_X1 U5918 ( .A1(n6827), .A2(n4656), .A3(n4325), .ZN(n4350) );
  AND2_X1 U5919 ( .A1(n5552), .A2(n4823), .ZN(n4351) );
  OR2_X1 U5920 ( .A1(n9010), .A2(n8646), .ZN(n4352) );
  INV_X1 U5921 ( .A(n4658), .ZN(n4657) );
  OR2_X1 U5922 ( .A1(n6828), .A2(n4659), .ZN(n4658) );
  NAND3_X1 U5923 ( .A1(n4832), .A2(n4831), .A3(n4830), .ZN(n6534) );
  INV_X1 U5924 ( .A(n6534), .ZN(n4829) );
  NAND2_X1 U5925 ( .A1(n5293), .A2(n5292), .ZN(n8996) );
  OR2_X1 U5926 ( .A1(n8369), .A2(n8368), .ZN(n4353) );
  AND2_X1 U5927 ( .A1(n5280), .A2(n5279), .ZN(n4354) );
  AND2_X1 U5928 ( .A1(n4630), .A2(n8253), .ZN(n4355) );
  INV_X1 U5929 ( .A(n4550), .ZN(n4549) );
  NOR2_X1 U5930 ( .A1(n4311), .A2(n7584), .ZN(n4550) );
  NAND2_X1 U5931 ( .A1(n8373), .A2(n8372), .ZN(n9627) );
  NAND2_X1 U5932 ( .A1(n8571), .A2(n8569), .ZN(n4356) );
  AND2_X1 U5933 ( .A1(n7003), .A2(n7001), .ZN(n4357) );
  AND2_X1 U5934 ( .A1(n8396), .A2(n7428), .ZN(n4358) );
  OR2_X1 U5935 ( .A1(n8362), .A2(n8559), .ZN(n4359) );
  INV_X1 U5936 ( .A(n9290), .ZN(n9652) );
  NAND2_X1 U5937 ( .A1(n8008), .A2(n8007), .ZN(n9290) );
  AND2_X1 U5938 ( .A1(n7108), .A2(n7004), .ZN(n4360) );
  NAND2_X1 U5939 ( .A1(n5581), .A2(n5577), .ZN(n4361) );
  NAND2_X1 U5940 ( .A1(n4843), .A2(n8555), .ZN(n4362) );
  INV_X1 U5941 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5942 ( .A1(n5334), .A2(n5333), .ZN(n8985) );
  AND2_X1 U5943 ( .A1(n7561), .A2(n7564), .ZN(n4363) );
  NAND2_X1 U5944 ( .A1(n5433), .A2(n5432), .ZN(n4364) );
  AND2_X1 U5945 ( .A1(n8910), .A2(n8413), .ZN(n8507) );
  NAND2_X1 U5946 ( .A1(n8036), .A2(n8035), .ZN(n8942) );
  OR2_X1 U5947 ( .A1(n6126), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4365) );
  INV_X1 U5948 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5949 ( .A1(n8048), .A2(n8532), .ZN(n4836) );
  NOR2_X1 U5950 ( .A1(n9532), .A2(n9394), .ZN(n4366) );
  NOR2_X1 U5951 ( .A1(n6220), .A2(n8001), .ZN(n4367) );
  AND2_X1 U5952 ( .A1(n8179), .A2(n8184), .ZN(n9298) );
  AND2_X1 U5953 ( .A1(n5129), .A2(SI_11_), .ZN(n4368) );
  INV_X1 U5954 ( .A(n8039), .ZN(n8961) );
  AND2_X1 U5955 ( .A1(n5441), .A2(n5440), .ZN(n8039) );
  AND2_X1 U5956 ( .A1(n5125), .A2(n4691), .ZN(n4369) );
  OR2_X1 U5957 ( .A1(n9941), .A2(n7111), .ZN(n8418) );
  NAND2_X1 U5958 ( .A1(n5026), .A2(SI_6_), .ZN(n4370) );
  OR2_X1 U5959 ( .A1(n4356), .A2(n4840), .ZN(n4371) );
  NOR2_X1 U5960 ( .A1(n8954), .A2(n8789), .ZN(n4372) );
  INV_X1 U5961 ( .A(n7275), .ZN(n9835) );
  OR2_X1 U5962 ( .A1(n8002), .A2(n6215), .ZN(n4373) );
  BUF_X8 U5963 ( .A(n4919), .Z(n8377) );
  INV_X1 U5964 ( .A(n4919), .ZN(n8001) );
  INV_X1 U5965 ( .A(n7510), .ZN(n8498) );
  AND2_X1 U5966 ( .A1(n4346), .A2(n8095), .ZN(n4374) );
  INV_X1 U5967 ( .A(n8426), .ZN(n4827) );
  OR2_X1 U5968 ( .A1(n8710), .A2(n7102), .ZN(n8426) );
  AND2_X1 U5969 ( .A1(n4370), .A2(n4511), .ZN(n4375) );
  INV_X1 U5970 ( .A(n5725), .ZN(n4599) );
  NAND2_X1 U5971 ( .A1(n4851), .A2(n5724), .ZN(n5725) );
  AND2_X1 U5972 ( .A1(n4340), .A2(n4476), .ZN(n4376) );
  INV_X1 U5973 ( .A(n4815), .ZN(n4814) );
  NAND2_X1 U5974 ( .A1(n7736), .A2(n4820), .ZN(n4815) );
  AND2_X1 U5975 ( .A1(n4685), .A2(n4688), .ZN(n4684) );
  NAND2_X1 U5976 ( .A1(n4580), .A2(n4579), .ZN(n4377) );
  INV_X1 U5977 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4875) );
  OR2_X1 U5978 ( .A1(n9288), .A2(n9287), .ZN(P1_U3260) );
  NAND2_X1 U5979 ( .A1(n5930), .A2(n5929), .ZN(n9552) );
  INV_X1 U5980 ( .A(n9552), .ZN(n4483) );
  INV_X1 U5981 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4895) );
  INV_X1 U5982 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5983 ( .A1(n6129), .A2(n8296), .ZN(n8168) );
  NOR3_X1 U5984 ( .A1(n9457), .A2(n9548), .A3(n9552), .ZN(n9400) );
  NAND2_X1 U5985 ( .A1(n4833), .A2(n4834), .ZN(n4379) );
  AND2_X1 U5986 ( .A1(n7949), .A2(n4547), .ZN(n4546) );
  INV_X1 U5987 ( .A(n4964), .ZN(n5015) );
  NAND2_X1 U5988 ( .A1(n7250), .A2(n7249), .ZN(n7274) );
  NOR2_X1 U5989 ( .A1(n9204), .A2(n7337), .ZN(n4380) );
  NAND2_X1 U5990 ( .A1(n7504), .A2(n7503), .ZN(n7576) );
  NAND2_X1 U5991 ( .A1(n7583), .A2(n7582), .ZN(n7604) );
  OR2_X1 U5992 ( .A1(n9738), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4381) );
  AND2_X1 U5993 ( .A1(n6489), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4382) );
  INV_X1 U5994 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4897) );
  OAI21_X1 U5995 ( .B1(n7583), .B2(n4549), .A(n4546), .ZN(n8912) );
  NAND2_X1 U5996 ( .A1(n4595), .A2(n4593), .ZN(n7561) );
  OR2_X1 U5997 ( .A1(n9570), .A2(n9199), .ZN(n4383) );
  AND2_X1 U5998 ( .A1(n9570), .A2(n9199), .ZN(n4384) );
  NAND2_X1 U5999 ( .A1(n4834), .A2(n4871), .ZN(n5488) );
  NAND2_X1 U6000 ( .A1(n5812), .A2(n5552), .ZN(n5831) );
  NAND2_X1 U6001 ( .A1(n4545), .A2(n4541), .ZN(n7950) );
  NAND2_X1 U6002 ( .A1(n9644), .A2(n5887), .ZN(n9114) );
  NOR3_X1 U6003 ( .A1(n9457), .A2(n9537), .A3(n4482), .ZN(n4484) );
  NAND2_X1 U6004 ( .A1(n8904), .A2(n4520), .ZN(n4521) );
  INV_X1 U6005 ( .A(n7717), .ZN(n9337) );
  AND2_X1 U6006 ( .A1(n6073), .A2(n6072), .ZN(n7717) );
  AND2_X1 U6007 ( .A1(n9352), .A2(n9483), .ZN(n4385) );
  NAND2_X1 U6008 ( .A1(n5467), .A2(n5466), .ZN(n8954) );
  INV_X1 U6009 ( .A(n4481), .ZN(n9401) );
  NOR2_X1 U6010 ( .A1(n9457), .A2(n4482), .ZN(n4481) );
  INV_X1 U6011 ( .A(n6900), .ZN(n4783) );
  NAND2_X1 U6012 ( .A1(n6091), .A2(n6090), .ZN(n9505) );
  NOR2_X1 U6013 ( .A1(n7622), .A2(n9200), .ZN(n4386) );
  NOR2_X1 U6014 ( .A1(n5455), .A2(n5459), .ZN(n4387) );
  AND2_X1 U6015 ( .A1(n9505), .A2(n4819), .ZN(n4388) );
  INV_X1 U6016 ( .A(n8204), .ZN(n4617) );
  OR2_X1 U6017 ( .A1(n5487), .A2(n5486), .ZN(n4389) );
  AND2_X1 U6018 ( .A1(n8001), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4390) );
  AND2_X1 U6019 ( .A1(n5282), .A2(n5331), .ZN(n4391) );
  AND2_X1 U6020 ( .A1(n6511), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4392) );
  AND2_X1 U6021 ( .A1(n7429), .A2(n7428), .ZN(n4393) );
  AND2_X1 U6022 ( .A1(n4551), .A2(n8505), .ZN(n4394) );
  NOR2_X1 U6023 ( .A1(n8755), .A2(n8409), .ZN(n4395) );
  AND2_X2 U6024 ( .A1(n6430), .A2(n6805), .ZN(n9965) );
  AND2_X1 U6025 ( .A1(n6774), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4396) );
  INV_X1 U6026 ( .A(n8266), .ZN(n4621) );
  NOR2_X1 U6027 ( .A1(n7278), .A2(n7277), .ZN(n7306) );
  NAND2_X1 U6028 ( .A1(n5353), .A2(n5352), .ZN(n8980) );
  INV_X1 U6029 ( .A(n8980), .ZN(n4519) );
  INV_X1 U6030 ( .A(n7564), .ZN(n4590) );
  NOR2_X1 U6031 ( .A1(n7649), .A2(n4494), .ZN(n7749) );
  NAND2_X1 U6032 ( .A1(n7213), .A2(n4415), .ZN(n7429) );
  NAND2_X1 U6033 ( .A1(n7002), .A2(n7001), .ZN(n7018) );
  OR2_X1 U6034 ( .A1(n4490), .A2(n7155), .ZN(n4397) );
  INV_X1 U6035 ( .A(n6197), .ZN(n4597) );
  AND2_X1 U6036 ( .A1(n6582), .A2(n8428), .ZN(n6961) );
  INV_X1 U6037 ( .A(n4477), .ZN(n8264) );
  NAND2_X1 U6038 ( .A1(n4622), .A2(n8193), .ZN(n4477) );
  INV_X1 U6039 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4526) );
  AND2_X1 U6040 ( .A1(n7068), .A2(n7067), .ZN(n4398) );
  AND2_X1 U6041 ( .A1(n4619), .A2(n4623), .ZN(n4399) );
  AND2_X1 U6042 ( .A1(n4582), .A2(n4581), .ZN(n4400) );
  INV_X1 U6043 ( .A(n6657), .ZN(n4583) );
  NAND2_X1 U6044 ( .A1(n6246), .A2(n4310), .ZN(n8863) );
  INV_X1 U6045 ( .A(n8863), .ZN(n8917) );
  OR3_X1 U6046 ( .A1(n6554), .A2(n9615), .A3(n6729), .ZN(n9642) );
  INV_X1 U6047 ( .A(n9642), .ZN(n9173) );
  INV_X1 U6048 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4632) );
  OR2_X1 U6049 ( .A1(n6957), .A2(n6825), .ZN(n6836) );
  INV_X1 U6050 ( .A(n6836), .ZN(n4515) );
  AND2_X1 U6051 ( .A1(n4699), .A2(n4697), .ZN(n4401) );
  AND2_X1 U6052 ( .A1(n6541), .A2(n8440), .ZN(n6980) );
  INV_X1 U6053 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n4421) );
  INV_X2 U6054 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X2 U6055 ( .B1(n8800), .B2(n4404), .A(n4402), .ZN(n8783) );
  NAND3_X1 U6056 ( .A1(n4438), .A2(n4436), .A3(n4432), .ZN(P2_U3264) );
  NAND4_X1 U6057 ( .A1(n4321), .A2(n4847), .A3(n5551), .A4(n4451), .ZN(n5575)
         );
  NOR2_X2 U6058 ( .A1(n5686), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5618) );
  NOR2_X1 U6059 ( .A1(n8304), .A2(n4456), .ZN(n4455) );
  NAND2_X1 U6060 ( .A1(n6933), .A2(n8267), .ZN(n6892) );
  NAND2_X1 U6061 ( .A1(n7063), .A2(n4455), .ZN(n6933) );
  NAND2_X1 U6062 ( .A1(n4454), .A2(n8267), .ZN(n4453) );
  NAND2_X1 U6063 ( .A1(n8097), .A2(n8168), .ZN(n4458) );
  NAND2_X1 U6064 ( .A1(n4457), .A2(n4461), .ZN(n8119) );
  NAND2_X1 U6065 ( .A1(n8132), .A2(n4468), .ZN(n4465) );
  NAND2_X1 U6066 ( .A1(n4465), .A2(n4466), .ZN(n8141) );
  NAND2_X2 U6067 ( .A1(n8002), .A2(n8001), .ZN(n8006) );
  NAND2_X1 U6068 ( .A1(n8002), .A2(n4390), .ZN(n5631) );
  AND2_X1 U6069 ( .A1(n5640), .A2(n4373), .ZN(n4480) );
  NAND2_X1 U6070 ( .A1(n4478), .A2(n6721), .ZN(n6918) );
  INV_X1 U6071 ( .A(n4484), .ZN(n9386) );
  NAND3_X1 U6072 ( .A1(n8568), .A2(n8569), .A3(n4857), .ZN(n4496) );
  OAI21_X1 U6073 ( .B1(n4499), .B2(n8561), .A(n8560), .ZN(n4498) );
  NAND2_X1 U6074 ( .A1(n4503), .A2(n4506), .ZN(n8508) );
  NAND3_X1 U6075 ( .A1(n4505), .A2(n4509), .A3(n4504), .ZN(n4503) );
  NAND3_X1 U6076 ( .A1(n8492), .A2(n8556), .A3(n8498), .ZN(n4504) );
  AND2_X1 U6077 ( .A1(n8770), .A2(n4516), .ZN(n8761) );
  NAND2_X1 U6078 ( .A1(n8770), .A2(n8033), .ZN(n8356) );
  NAND2_X1 U6079 ( .A1(n8770), .A2(n4517), .ZN(n8760) );
  INV_X1 U6080 ( .A(n4521), .ZN(n8891) );
  NAND4_X1 U6081 ( .A1(n4528), .A2(n4889), .A3(n4527), .A4(n4526), .ZN(n4525)
         );
  NAND4_X1 U6082 ( .A1(n4533), .A2(n4532), .A3(n4531), .A4(n4530), .ZN(n4529)
         );
  NAND2_X1 U6083 ( .A1(n4537), .A2(n7208), .ZN(n4535) );
  NAND3_X1 U6084 ( .A1(n4535), .A2(n8480), .A3(n4534), .ZN(n7511) );
  NAND2_X1 U6085 ( .A1(n7208), .A2(n8478), .ZN(n7436) );
  NAND2_X1 U6086 ( .A1(n4546), .A2(n7583), .ZN(n4545) );
  NAND2_X1 U6087 ( .A1(n8878), .A2(n4556), .ZN(n4552) );
  NAND3_X1 U6088 ( .A1(n4833), .A2(n4834), .A3(n4844), .ZN(n4902) );
  NAND4_X1 U6089 ( .A1(n4833), .A2(n4834), .A3(n4844), .A4(n4559), .ZN(n4560)
         );
  NAND3_X2 U6090 ( .A1(n5630), .A2(n4568), .A3(n5547), .ZN(n5686) );
  NAND2_X1 U6091 ( .A1(n4568), .A2(n5630), .ZN(n5684) );
  NAND2_X1 U6092 ( .A1(n4570), .A2(n9147), .ZN(n9075) );
  INV_X1 U6093 ( .A(n6007), .ZN(n4571) );
  AOI21_X1 U6094 ( .B1(n9147), .B2(n6007), .A(n6008), .ZN(n4572) );
  AOI21_X1 U6095 ( .B1(n5882), .B2(n9185), .A(n4377), .ZN(n4578) );
  NAND3_X1 U6096 ( .A1(n4581), .A2(n4582), .A3(n6689), .ZN(n6688) );
  NAND2_X1 U6097 ( .A1(n6653), .A2(n6654), .ZN(n4584) );
  NAND2_X1 U6098 ( .A1(n7455), .A2(n5830), .ZN(n4595) );
  NAND2_X1 U6099 ( .A1(n4585), .A2(n4588), .ZN(n7637) );
  NAND2_X1 U6100 ( .A1(n7455), .A2(n4586), .ZN(n4585) );
  OAI22_X1 U6101 ( .A1(n6200), .A2(n4596), .B1(n5725), .B2(n4328), .ZN(n7181)
         );
  NAND2_X2 U6102 ( .A1(n4603), .A2(n4601), .ZN(n9143) );
  NAND2_X2 U6103 ( .A1(n5926), .A2(n4604), .ZN(n4603) );
  INV_X2 U6104 ( .A(n6101), .ZN(n6057) );
  NOR2_X1 U6105 ( .A1(n5656), .A2(n4605), .ZN(n6558) );
  AND2_X4 U6106 ( .A1(n4606), .A2(n5610), .ZN(n6101) );
  NAND2_X1 U6107 ( .A1(n9105), .A2(n9106), .ZN(n9168) );
  NAND2_X1 U6108 ( .A1(n5558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U6109 ( .A1(n7308), .A2(n4615), .ZN(n4612) );
  NAND2_X1 U6110 ( .A1(n4612), .A2(n4613), .ZN(n7522) );
  NAND2_X1 U6111 ( .A1(n8189), .A2(n6891), .ZN(n4622) );
  NAND3_X1 U6112 ( .A1(n4619), .A2(n4623), .A3(n8067), .ZN(n7280) );
  NAND3_X1 U6113 ( .A1(n7063), .A2(n8075), .A3(n8276), .ZN(n4619) );
  NAND2_X2 U6114 ( .A1(n4622), .A2(n4620), .ZN(n7063) );
  NAND2_X1 U6115 ( .A1(n4624), .A2(n8075), .ZN(n4623) );
  OAI21_X1 U6116 ( .B1(n9363), .B2(n4627), .A(n4625), .ZN(n9324) );
  NAND2_X1 U6117 ( .A1(n9363), .A2(n7734), .ZN(n4630) );
  NAND3_X1 U6118 ( .A1(n4822), .A2(n5618), .A3(n4847), .ZN(n6126) );
  NAND2_X1 U6119 ( .A1(n7627), .A2(n8222), .ZN(n7626) );
  NAND2_X1 U6120 ( .A1(n7286), .A2(n7413), .ZN(n7481) );
  XNOR2_X1 U6121 ( .A(n5642), .B(n6024), .ZN(n6654) );
  OAI211_X2 U6122 ( .C1(n8002), .C2(n6450), .A(n5705), .B(n5704), .ZN(n7157)
         );
  NAND2_X1 U6123 ( .A1(n5657), .A2(n6556), .ZN(n6653) );
  NAND2_X1 U6124 ( .A1(n5573), .A2(n5603), .ZN(n6130) );
  NAND2_X1 U6125 ( .A1(n6557), .A2(n6558), .ZN(n6556) );
  INV_X2 U6126 ( .A(n7157), .ZN(n9823) );
  XNOR2_X2 U6127 ( .A(n4647), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U6128 ( .A1(n6956), .A2(n4350), .ZN(n4652) );
  NAND3_X1 U6129 ( .A1(n4652), .A2(n6844), .A3(n4651), .ZN(n6966) );
  AND2_X1 U6130 ( .A1(n6827), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U6131 ( .A1(n7444), .A2(n7431), .ZN(n7433) );
  INV_X1 U6132 ( .A(n7579), .ZN(n4663) );
  NAND2_X1 U6133 ( .A1(n8853), .A2(n4668), .ZN(n4667) );
  OAI21_X1 U6134 ( .B1(n8947), .B2(n4675), .A(n4672), .ZN(P2_U3549) );
  OAI21_X1 U6135 ( .B1(n8947), .B2(n4679), .A(n4676), .ZN(P2_U3517) );
  NAND2_X1 U6136 ( .A1(n9983), .A2(n9962), .ZN(n4675) );
  NAND2_X1 U6137 ( .A1(n4680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4874) );
  NAND4_X1 U6138 ( .A1(n4833), .A2(n4834), .A3(n4875), .A4(n4873), .ZN(n4680)
         );
  NAND3_X1 U6139 ( .A1(n4833), .A2(n4834), .A3(n4873), .ZN(n5498) );
  INV_X1 U6140 ( .A(n6868), .ZN(n4687) );
  NAND2_X1 U6141 ( .A1(n4681), .A2(n4682), .ZN(n5150) );
  NAND2_X1 U6142 ( .A1(n4684), .A2(n6868), .ZN(n4681) );
  NAND2_X1 U6143 ( .A1(n4693), .A2(n6606), .ZN(n4694) );
  NAND2_X1 U6144 ( .A1(n4694), .A2(n4695), .ZN(n6697) );
  NAND2_X1 U6145 ( .A1(n7678), .A2(n4705), .ZN(n4702) );
  NAND2_X1 U6146 ( .A1(n4702), .A2(n4703), .ZN(n8602) );
  NAND3_X1 U6147 ( .A1(n5433), .A2(n5432), .A3(n5453), .ZN(n6164) );
  NAND3_X1 U6148 ( .A1(n5433), .A2(n5432), .A3(n4862), .ZN(n4709) );
  NAND3_X1 U6149 ( .A1(n6196), .A2(n8612), .A3(n4710), .ZN(n5546) );
  NAND2_X1 U6150 ( .A1(n4711), .A2(n4712), .ZN(n5384) );
  NAND2_X1 U6151 ( .A1(n5327), .A2(n4713), .ZN(n4711) );
  OAI21_X2 U6152 ( .B1(n7491), .B2(n4723), .A(n4718), .ZN(n7679) );
  NAND2_X1 U6153 ( .A1(n4926), .A2(n8377), .ZN(n4947) );
  NAND3_X1 U6154 ( .A1(n6359), .A2(n4310), .A3(n6367), .ZN(n4728) );
  NAND2_X1 U6155 ( .A1(n6345), .A2(n6344), .ZN(n6343) );
  NAND2_X1 U6156 ( .A1(n4918), .A2(n4730), .ZN(n6344) );
  INV_X1 U6157 ( .A(n4870), .ZN(n4733) );
  INV_X1 U6158 ( .A(n4734), .ZN(n5268) );
  NAND2_X1 U6159 ( .A1(n5200), .A2(n5199), .ZN(n5229) );
  NAND2_X1 U6160 ( .A1(n5006), .A2(n4344), .ZN(n4744) );
  NAND2_X1 U6161 ( .A1(n4744), .A2(n4375), .ZN(n5050) );
  NAND2_X1 U6162 ( .A1(n5006), .A2(n5005), .ZN(n4745) );
  XNOR2_X2 U6163 ( .A(n8000), .B(n7999), .ZN(n9048) );
  NAND2_X1 U6164 ( .A1(n5092), .A2(n4754), .ZN(n4753) );
  NAND2_X1 U6165 ( .A1(n5092), .A2(n5091), .ZN(n5116) );
  NAND2_X1 U6166 ( .A1(n4753), .A2(n4756), .ZN(n5160) );
  INV_X1 U6167 ( .A(n4775), .ZN(n4774) );
  OAI21_X1 U6168 ( .B1(n6911), .B2(n4780), .A(n4778), .ZN(n6903) );
  NAND2_X1 U6169 ( .A1(n4781), .A2(n4779), .ZN(n6902) );
  NAND2_X1 U6170 ( .A1(n6911), .A2(n4782), .ZN(n4781) );
  NAND2_X1 U6171 ( .A1(n7526), .A2(n4329), .ZN(n4786) );
  NAND2_X1 U6172 ( .A1(n7708), .A2(n4799), .ZN(n4798) );
  NAND3_X1 U6173 ( .A1(n4800), .A2(n4803), .A3(n4345), .ZN(n4797) );
  OAI21_X1 U6174 ( .B1(n9327), .B2(n4815), .A(n4812), .ZN(n7726) );
  NAND2_X1 U6175 ( .A1(n9327), .A2(n4817), .ZN(n4816) );
  NAND3_X1 U6176 ( .A1(n4825), .A2(n6833), .A3(n4824), .ZN(n6967) );
  NAND3_X1 U6177 ( .A1(n8426), .A2(n6961), .A3(n8384), .ZN(n4825) );
  NAND2_X1 U6178 ( .A1(n6534), .A2(n6594), .ZN(n8448) );
  AND2_X1 U6179 ( .A1(n4958), .A2(n4957), .ZN(n4832) );
  AND2_X1 U6180 ( .A1(n4871), .A2(n4872), .ZN(n4833) );
  INV_X2 U6181 ( .A(n4332), .ZN(n4834) );
  NAND2_X2 U6182 ( .A1(n8879), .A2(n8880), .ZN(n8878) );
  OAI21_X1 U6183 ( .B1(n4353), .B2(n4839), .A(n4838), .ZN(n8380) );
  NAND2_X1 U6184 ( .A1(n8572), .A2(n4322), .ZN(n4839) );
  NAND2_X1 U6185 ( .A1(n8787), .A2(n4319), .ZN(n4842) );
  OR2_X1 U6186 ( .A1(n8787), .A2(n8788), .ZN(n4843) );
  INV_X1 U6187 ( .A(n4843), .ZN(n8786) );
  NAND3_X1 U6188 ( .A1(n4927), .A2(n4865), .A3(n4866), .ZN(n4978) );
  XNOR2_X1 U6189 ( .A(n7737), .B(n8329), .ZN(n7748) );
  NAND2_X1 U6190 ( .A1(n4364), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U6191 ( .A1(n5882), .A2(n5881), .ZN(n9182) );
  NAND2_X1 U6192 ( .A1(n6718), .A2(n6756), .ZN(n6725) );
  XNOR2_X1 U6193 ( .A(n7726), .B(n8329), .ZN(n9503) );
  NAND2_X1 U6194 ( .A1(n4956), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4908) );
  AOI21_X2 U6195 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8945) );
  NOR2_X2 U6196 ( .A1(n8178), .A2(n8177), .ZN(n8345) );
  AND2_X1 U6197 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  INV_X1 U6198 ( .A(n8688), .ZN(n7687) );
  AND2_X1 U6199 ( .A1(n5524), .A2(n5520), .ZN(n8688) );
  AND3_X1 U6200 ( .A1(n4895), .A2(n4892), .A3(n4897), .ZN(n4846) );
  AND2_X2 U6201 ( .A1(n6259), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND2_X2 U6202 ( .A1(n6755), .A2(n7669), .ZN(n9489) );
  INV_X1 U6203 ( .A(n9489), .ZN(n9313) );
  OR2_X1 U6204 ( .A1(n8002), .A2(n6445), .ZN(n4848) );
  INV_X1 U6205 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4882) );
  AND2_X1 U6206 ( .A1(n6132), .A2(n9173), .ZN(n4849) );
  AND2_X1 U6207 ( .A1(n5908), .A2(n5888), .ZN(n4850) );
  NOR2_X1 U6208 ( .A1(n5810), .A2(n7404), .ZN(n4852) );
  OR2_X1 U6209 ( .A1(n8974), .A2(n8864), .ZN(n4853) );
  AND2_X1 U6210 ( .A1(n5545), .A2(n5544), .ZN(n4854) );
  AND2_X1 U6211 ( .A1(n5091), .A2(n5074), .ZN(n4855) );
  AND2_X1 U6212 ( .A1(n5117), .A2(n5096), .ZN(n4856) );
  AND2_X1 U6213 ( .A1(n5540), .A2(n5539), .ZN(n8776) );
  INV_X1 U6214 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5567) );
  OR2_X1 U6215 ( .A1(n9627), .A2(n8378), .ZN(n4857) );
  NAND2_X1 U6216 ( .A1(n7337), .A2(n9204), .ZN(n4858) );
  AND2_X1 U6217 ( .A1(n7226), .A2(n7126), .ZN(n4859) );
  INV_X1 U6218 ( .A(n8949), .ZN(n8033) );
  AND3_X1 U6219 ( .A1(n6189), .A2(n6190), .A3(n8612), .ZN(n4860) );
  AND3_X1 U6220 ( .A1(n6136), .A2(n9173), .A3(n6135), .ZN(n4861) );
  INV_X1 U6221 ( .A(n8889), .ZN(n8046) );
  INV_X1 U6222 ( .A(n8305), .ZN(n7069) );
  INV_X1 U6223 ( .A(n9336), .ZN(n7715) );
  NOR2_X1 U6224 ( .A1(n6163), .A2(n5487), .ZN(n4862) );
  NOR2_X1 U6225 ( .A1(n5994), .A2(n9144), .ZN(n4864) );
  OAI21_X1 U6226 ( .B1(n8667), .B2(n8668), .A(n8665), .ZN(n5365) );
  INV_X1 U6227 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5564) );
  INV_X1 U6228 ( .A(n5365), .ZN(n5366) );
  INV_X1 U6229 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5611) );
  INV_X1 U6230 ( .A(n5337), .ZN(n5335) );
  INV_X1 U6231 ( .A(n5142), .ZN(n5141) );
  NOR2_X1 U6232 ( .A1(n8052), .A2(n8051), .ZN(n8369) );
  OAI21_X1 U6233 ( .B1(n7109), .B2(n7108), .A(n8418), .ZN(n7207) );
  INV_X1 U6234 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4872) );
  INV_X1 U6235 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4866) );
  INV_X1 U6236 ( .A(n5674), .ZN(n5675) );
  INV_X1 U6237 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7167) );
  OR2_X1 U6238 ( .A1(n6065), .A2(n9067), .ZN(n6093) );
  INV_X1 U6239 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5254) );
  AND4_X1 U6240 ( .A1(n5550), .A2(n5549), .A3(n5702), .A4(n5548), .ZN(n5551)
         );
  OR2_X1 U6241 ( .A1(n5736), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5737) );
  INV_X1 U6242 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5041) );
  OR2_X1 U6243 ( .A1(n5443), .A2(n5442), .ZN(n5471) );
  NAND2_X1 U6244 ( .A1(n5141), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5152) );
  AND2_X1 U6245 ( .A1(n9879), .A2(n5515), .ZN(n6352) );
  INV_X1 U6246 ( .A(n8409), .ZN(n8433) );
  OR2_X1 U6247 ( .A1(n8996), .A2(n8918), .ZN(n8022) );
  INV_X1 U6248 ( .A(n8390), .ZN(n7003) );
  INV_X1 U6249 ( .A(n8848), .ZN(n8974) );
  OAI21_X1 U6250 ( .B1(n7511), .B2(n7510), .A(n8494), .ZN(n7581) );
  OR2_X1 U6251 ( .A1(n6557), .A2(n6024), .ZN(n5657) );
  NAND2_X1 U6252 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  OR2_X1 U6253 ( .A1(n5973), .A2(n5964), .ZN(n5999) );
  NOR2_X1 U6254 ( .A1(n5855), .A2(n7167), .ZN(n5871) );
  NAND2_X1 U6255 ( .A1(n4313), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5639) );
  INV_X1 U6256 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6443) );
  INV_X1 U6257 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7927) );
  AND2_X1 U6258 ( .A1(n6093), .A2(n6066), .ZN(n9320) );
  OR2_X1 U6259 ( .A1(n7691), .A2(n7690), .ZN(n9450) );
  INV_X1 U6260 ( .A(n7286), .ZN(n7313) );
  OR2_X1 U6261 ( .A1(n9602), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6125) );
  INV_X1 U6262 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6263 ( .A1(n8954), .A2(n8688), .ZN(n5545) );
  OR2_X1 U6264 ( .A1(n5042), .A2(n5041), .ZN(n5080) );
  INV_X1 U6265 ( .A(n8682), .ZN(n8672) );
  OR2_X1 U6266 ( .A1(n5110), .A2(n5109), .ZN(n5142) );
  INV_X1 U6267 ( .A(n8623), .ZN(n8685) );
  OR2_X1 U6268 ( .A1(n6352), .A2(n6351), .ZN(n6361) );
  INV_X1 U6269 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7090) );
  INV_X1 U6270 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8681) );
  AND2_X1 U6271 ( .A1(n8588), .A2(n8433), .ZN(n6246) );
  NOR2_X2 U6272 ( .A1(n7449), .A2(n9025), .ZN(n7448) );
  OR2_X1 U6273 ( .A1(n6808), .A2(n6807), .ZN(n6813) );
  AND2_X1 U6274 ( .A1(n5510), .A2(n9883), .ZN(n5511) );
  AND2_X1 U6275 ( .A1(n6285), .A2(n8381), .ZN(n8859) );
  OAI21_X1 U6276 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n9878), .A(n9887), .ZN(n6808)
         );
  INV_X1 U6277 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U6278 ( .A1(n4363), .A2(n5863), .ZN(n7638) );
  NAND2_X1 U6279 ( .A1(n6704), .A2(n6705), .ZN(n6703) );
  AOI21_X1 U6280 ( .B1(n7400), .B2(n5811), .A(n4852), .ZN(n7455) );
  OR2_X1 U6281 ( .A1(n6033), .A2(n6032), .ZN(n6047) );
  AND3_X1 U6282 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5707) );
  OR2_X1 U6283 ( .A1(n5752), .A2(n5751), .ZN(n5770) );
  OR2_X1 U6284 ( .A1(n5836), .A2(n5835), .ZN(n5855) );
  NAND2_X1 U6285 ( .A1(n8350), .A2(n8332), .ZN(n8061) );
  INV_X1 U6286 ( .A(n9778), .ZN(n9264) );
  OR2_X1 U6287 ( .A1(n6620), .A2(n8295), .ZN(n6137) );
  INV_X1 U6288 ( .A(n7754), .ZN(n7755) );
  OAI21_X1 U6289 ( .B1(n9343), .B2(n9350), .A(n7713), .ZN(n7714) );
  INV_X1 U6290 ( .A(n6154), .ZN(n8347) );
  AND2_X1 U6291 ( .A1(n8080), .A2(n8218), .ZN(n8308) );
  NAND2_X1 U6292 ( .A1(n6902), .A2(n6901), .ZN(n7068) );
  OR2_X1 U6293 ( .A1(n9602), .A2(n6639), .ZN(n6640) );
  AND2_X1 U6294 ( .A1(n5194), .A2(n5165), .ZN(n5173) );
  NOR2_X1 U6295 ( .A1(n5529), .A2(n5528), .ZN(n8634) );
  NOR2_X1 U6296 ( .A1(n5529), .A2(n5517), .ZN(n8612) );
  AND2_X1 U6297 ( .A1(n6186), .A2(n6185), .ZN(n8037) );
  AND3_X1 U6298 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n8661) );
  NAND2_X1 U6299 ( .A1(n6361), .A2(n6360), .ZN(n7977) );
  INV_X1 U6300 ( .A(n9871), .ZN(n9867) );
  INV_X1 U6301 ( .A(n7977), .ZN(n9868) );
  AND2_X1 U6302 ( .A1(n8529), .A2(n8532), .ZN(n8880) );
  INV_X1 U6303 ( .A(n8859), .ZN(n8920) );
  NOR2_X1 U6304 ( .A1(n9884), .A2(n5511), .ZN(n6429) );
  AND2_X1 U6305 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  AND2_X1 U6306 ( .A1(n7609), .A2(n9030), .ZN(n9890) );
  INV_X1 U6307 ( .A(n9890), .ZN(n9962) );
  NAND2_X1 U6308 ( .A1(n6155), .A2(n6154), .ZN(n9636) );
  AND3_X1 U6309 ( .A1(n8014), .A2(n8013), .A3(n8012), .ZN(n8062) );
  AND4_X1 U6310 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n9162)
         );
  AND4_X1 U6311 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n7570)
         );
  AND2_X1 U6312 ( .A1(n6313), .A2(n6304), .ZN(n9787) );
  AND2_X1 U6313 ( .A1(n6313), .A2(n6312), .ZN(n9778) );
  AND2_X1 U6314 ( .A1(n6313), .A2(n6260), .ZN(n9786) );
  AND2_X1 U6315 ( .A1(n9443), .A2(n8300), .ZN(n9481) );
  AND2_X1 U6316 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  OR2_X1 U6317 ( .A1(n7274), .A2(n8308), .ZN(n7326) );
  AND2_X1 U6318 ( .A1(n9492), .A2(n9655), .ZN(n9441) );
  INV_X1 U6319 ( .A(n9655), .ZN(n9843) );
  AND2_X1 U6320 ( .A1(n9498), .A2(n9805), .ZN(n9661) );
  OR2_X1 U6321 ( .A1(n6617), .A2(n6616), .ZN(n6642) );
  AND2_X1 U6322 ( .A1(n6210), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6128) );
  INV_X1 U6323 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7867) );
  INV_X1 U6324 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7918) );
  OAI21_X1 U6325 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9988), .ZN(n10018) );
  INV_X1 U6326 ( .A(n9885), .ZN(n9888) );
  NAND2_X1 U6327 ( .A1(n5525), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8633) );
  INV_X1 U6328 ( .A(n6169), .ZN(n6170) );
  INV_X1 U6329 ( .A(n8612), .ZN(n8690) );
  INV_X1 U6330 ( .A(n8822), .ZN(n8696) );
  INV_X1 U6331 ( .A(n7948), .ZN(n8698) );
  NAND2_X1 U6332 ( .A1(n6380), .A2(n4310), .ZN(n9869) );
  NAND2_X1 U6333 ( .A1(n6380), .A2(n6379), .ZN(n9871) );
  AND2_X1 U6334 ( .A1(n6248), .A2(n6247), .ZN(n8745) );
  NAND2_X1 U6335 ( .A1(n8933), .A2(n6819), .ZN(n8908) );
  INV_X1 U6336 ( .A(n9983), .ZN(n9980) );
  INV_X1 U6337 ( .A(n9965), .ZN(n9963) );
  NAND2_X1 U6338 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  XNOR2_X1 U6339 ( .A(n5494), .B(n4526), .ZN(n7324) );
  INV_X1 U6340 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U6341 ( .A1(n4861), .A2(n6159), .ZN(n6160) );
  INV_X1 U6342 ( .A(n9543), .ZN(n9405) );
  AND2_X1 U6343 ( .A1(n6145), .A2(n6144), .ZN(n9650) );
  INV_X1 U6344 ( .A(n7622), .ZN(n9673) );
  INV_X1 U6345 ( .A(n9192), .ZN(n9181) );
  INV_X1 U6346 ( .A(n8062), .ZN(n9196) );
  OR2_X1 U6347 ( .A1(n5956), .A2(n5955), .ZN(n9437) );
  INV_X1 U6348 ( .A(n7665), .ZN(n9484) );
  INV_X1 U6349 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9725) );
  OR2_X1 U6350 ( .A1(P1_U3083), .A2(n6259), .ZN(n9792) );
  INV_X1 U6351 ( .A(n9313), .ZN(n9465) );
  OR2_X1 U6352 ( .A1(n6642), .A2(n6618), .ZN(n9864) );
  AND2_X1 U6353 ( .A1(n9669), .A2(n9668), .ZN(n9679) );
  OR2_X1 U6354 ( .A1(n6642), .A2(n6740), .ZN(n9849) );
  INV_X1 U6355 ( .A(n9801), .ZN(n9798) );
  AND2_X1 U6356 ( .A1(n6209), .A2(n6128), .ZN(n9804) );
  INV_X1 U6357 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7517) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7242) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6615) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6274) );
  NOR2_X1 U6361 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  OAI21_X1 U6362 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10000), .ZN(n9998) );
  NOR2_X1 U6363 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4869) );
  NOR2_X1 U6364 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4868) );
  NAND4_X1 U6365 ( .A1(n4869), .A2(n4868), .A3(n4867), .A4(n5119), .ZN(n4870)
         );
  NAND2_X1 U6366 ( .A1(n5498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4876) );
  XNOR2_X1 U6367 ( .A(n4922), .B(SI_1_), .ZN(n4921) );
  MUX2_X1 U6368 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4919), .Z(n4920) );
  XNOR2_X1 U6369 ( .A(n4921), .B(n4920), .ZN(n6218) );
  INV_X1 U6370 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6219) );
  INV_X1 U6371 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U6372 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4880) );
  NAND2_X1 U6373 ( .A1(n5236), .A2(n4884), .ZN(n5255) );
  INV_X1 U6374 ( .A(n5255), .ZN(n4886) );
  NAND2_X1 U6375 ( .A1(n4886), .A2(n4885), .ZN(n4891) );
  INV_X1 U6376 ( .A(n4891), .ZN(n4887) );
  NAND2_X1 U6377 ( .A1(n4887), .A2(n4846), .ZN(n4888) );
  NAND2_X1 U6378 ( .A1(n4888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U6379 ( .A1(n5269), .A2(n4892), .ZN(n4893) );
  XNOR2_X2 U6380 ( .A(n4896), .B(n4895), .ZN(n8379) );
  NAND2_X2 U6381 ( .A1(n4898), .A2(n6811), .ZN(n4932) );
  INV_X1 U6382 ( .A(n9053), .ZN(n4904) );
  NAND2_X1 U6383 ( .A1(n4995), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4909) );
  INV_X1 U6384 ( .A(n9057), .ZN(n4905) );
  AND2_X2 U6385 ( .A1(n4904), .A2(n4905), .ZN(n4956) );
  OR2_X4 U6386 ( .A1(n5526), .A2(n5516), .ZN(n8382) );
  AND2_X1 U6387 ( .A1(n6277), .A2(n8382), .ZN(n4911) );
  NAND2_X1 U6388 ( .A1(n4995), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U6389 ( .A1(n4955), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6390 ( .A1(n4956), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U6391 ( .A1(n4964), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4912) );
  NAND4_X1 U6392 ( .A1(n4915), .A2(n4914), .A3(n4913), .A4(n4912), .ZN(n6281)
         );
  NAND2_X1 U6393 ( .A1(n6281), .A2(n8382), .ZN(n4917) );
  INV_X1 U6394 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U6395 ( .A1(n8001), .A2(SI_0_), .ZN(n4916) );
  XNOR2_X1 U6396 ( .A(n4916), .B(n6479), .ZN(n9061) );
  MUX2_X1 U6397 ( .A(n9876), .B(n9061), .S(n4926), .Z(n9892) );
  BUF_X4 U6398 ( .A(n4932), .Z(n5468) );
  INV_X1 U6399 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6221) );
  INV_X1 U6400 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6214) );
  MUX2_X1 U6401 ( .A(n6221), .B(n6214), .S(n4919), .Z(n4942) );
  XNOR2_X1 U6402 ( .A(n4942), .B(SI_2_), .ZN(n4940) );
  NAND2_X1 U6403 ( .A1(n4921), .A2(n4920), .ZN(n4925) );
  INV_X1 U6404 ( .A(n4922), .ZN(n4923) );
  NAND2_X1 U6405 ( .A1(n4923), .A2(SI_1_), .ZN(n4924) );
  NAND2_X1 U6406 ( .A1(n4925), .A2(n4924), .ZN(n4941) );
  XNOR2_X1 U6407 ( .A(n4940), .B(n4941), .ZN(n6220) );
  OR2_X1 U6408 ( .A1(n4939), .A2(n6220), .ZN(n4931) );
  OR2_X1 U6409 ( .A1(n4317), .A2(n6221), .ZN(n4930) );
  OR2_X1 U6410 ( .A1(n4927), .A2(n9049), .ZN(n4928) );
  INV_X1 U6411 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4948) );
  XNOR2_X1 U6412 ( .A(n4928), .B(n4948), .ZN(n6371) );
  OR2_X1 U6413 ( .A1(n4926), .A2(n6371), .ZN(n4929) );
  XNOR2_X1 U6414 ( .A(n6532), .B(n4932), .ZN(n4938) );
  NAND2_X1 U6415 ( .A1(n4995), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4936) );
  NAND2_X1 U6416 ( .A1(n4955), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6417 ( .A1(n4956), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U6418 ( .A1(n4964), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4933) );
  INV_X1 U6419 ( .A(n6531), .ZN(n6596) );
  NAND2_X1 U6420 ( .A1(n6531), .A2(n8382), .ZN(n4937) );
  XNOR2_X1 U6421 ( .A(n4938), .B(n4937), .ZN(n6473) );
  NAND2_X1 U6422 ( .A1(n4941), .A2(n4940), .ZN(n4945) );
  INV_X1 U6423 ( .A(n4942), .ZN(n4943) );
  NAND2_X1 U6424 ( .A1(n4943), .A2(SI_2_), .ZN(n4944) );
  NAND2_X1 U6425 ( .A1(n4945), .A2(n4944), .ZN(n4970) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6223) );
  INV_X1 U6427 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U6428 ( .A(n4971), .B(SI_3_), .ZN(n4969) );
  XNOR2_X1 U6429 ( .A(n4970), .B(n4969), .ZN(n6222) );
  OR2_X1 U6430 ( .A1(n4939), .A2(n6222), .ZN(n4954) );
  OR2_X1 U6431 ( .A1(n4947), .A2(n6223), .ZN(n4953) );
  AND2_X1 U6432 ( .A1(n4927), .A2(n4948), .ZN(n4949) );
  OR2_X1 U6433 ( .A1(n4949), .A2(n9049), .ZN(n4951) );
  XNOR2_X1 U6434 ( .A(n4951), .B(n4950), .ZN(n6471) );
  OR2_X1 U6435 ( .A1(n4926), .A2(n6471), .ZN(n4952) );
  XNOR2_X1 U6436 ( .A(n5468), .B(n6594), .ZN(n4959) );
  NAND2_X1 U6437 ( .A1(n4995), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4958) );
  INV_X1 U6438 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U6439 ( .A1(n4964), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4957) );
  AND2_X1 U6440 ( .A1(n6534), .A2(n8382), .ZN(n4961) );
  XNOR2_X1 U6441 ( .A(n4959), .B(n4961), .ZN(n6592) );
  INV_X1 U6442 ( .A(n4959), .ZN(n4960) );
  INV_X1 U6443 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n4962) );
  OR2_X1 U6444 ( .A1(n5381), .A2(n4962), .ZN(n4968) );
  NAND2_X1 U6445 ( .A1(n4955), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6446 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n4997) );
  OAI21_X1 U6447 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n4997), .ZN(n6959) );
  INV_X1 U6448 ( .A(n6959), .ZN(n4963) );
  NAND2_X1 U6449 ( .A1(n4956), .A2(n4963), .ZN(n4966) );
  NAND2_X1 U6450 ( .A1(n4964), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4965) );
  NAND4_X1 U6451 ( .A1(n4968), .A2(n4967), .A3(n4966), .A4(n4965), .ZN(n8711)
         );
  INV_X1 U6452 ( .A(n8711), .ZN(n6595) );
  NOR2_X1 U6453 ( .A1(n6595), .A2(n6174), .ZN(n4984) );
  NAND2_X1 U6454 ( .A1(n4970), .A2(n4969), .ZN(n4974) );
  INV_X1 U6455 ( .A(n4971), .ZN(n4972) );
  NAND2_X1 U6456 ( .A1(n4972), .A2(SI_3_), .ZN(n4973) );
  MUX2_X1 U6457 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8377), .Z(n4990) );
  INV_X1 U6458 ( .A(SI_4_), .ZN(n7771) );
  XNOR2_X1 U6459 ( .A(n4990), .B(n7771), .ZN(n4988) );
  XNOR2_X1 U6460 ( .A(n4989), .B(n4988), .ZN(n6225) );
  OR2_X1 U6461 ( .A1(n4939), .A2(n6225), .ZN(n4982) );
  INV_X1 U6462 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6224) );
  OR2_X1 U6463 ( .A1(n4947), .A2(n6224), .ZN(n4981) );
  NOR2_X1 U6464 ( .A1(n4975), .A2(n9049), .ZN(n4976) );
  MUX2_X1 U6465 ( .A(n9049), .B(n4976), .S(P2_IR_REG_4__SCAN_IN), .Z(n4977) );
  INV_X1 U6466 ( .A(n4977), .ZN(n4979) );
  NAND2_X1 U6467 ( .A1(n4979), .A2(n4978), .ZN(n6428) );
  OR2_X1 U6468 ( .A1(n4926), .A2(n6428), .ZN(n4980) );
  XOR2_X1 U6469 ( .A(n5468), .B(n9905), .Z(n4983) );
  NOR2_X1 U6470 ( .A1(n4983), .A2(n4984), .ZN(n4985) );
  AOI21_X1 U6471 ( .B1(n4984), .B2(n4983), .A(n4985), .ZN(n6607) );
  INV_X1 U6472 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6473 ( .A1(n4978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4987) );
  XNOR2_X1 U6474 ( .A(n4987), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6489) );
  AOI22_X1 U6475 ( .A1(n5291), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6244), .B2(
        n6489), .ZN(n4994) );
  NAND2_X1 U6476 ( .A1(n4989), .A2(n4988), .ZN(n4992) );
  NAND2_X1 U6477 ( .A1(n4990), .A2(SI_4_), .ZN(n4991) );
  MUX2_X1 U6478 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8377), .Z(n5007) );
  INV_X1 U6479 ( .A(SI_5_), .ZN(n7760) );
  XNOR2_X1 U6480 ( .A(n5007), .B(n7760), .ZN(n5005) );
  XNOR2_X1 U6481 ( .A(n5006), .B(n5005), .ZN(n6228) );
  OR2_X1 U6482 ( .A1(n6228), .A2(n4939), .ZN(n4993) );
  XNOR2_X1 U6483 ( .A(n5468), .B(n7102), .ZN(n5004) );
  NAND2_X1 U6484 ( .A1(n4995), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6485 ( .A1(n4955), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5001) );
  INV_X1 U6486 ( .A(n4997), .ZN(n4996) );
  NAND2_X1 U6487 ( .A1(n4996), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5013) );
  INV_X1 U6488 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U6489 ( .A1(n4997), .A2(n6568), .ZN(n4998) );
  AND2_X1 U6490 ( .A1(n5013), .A2(n4998), .ZN(n7099) );
  NAND2_X1 U6491 ( .A1(n4956), .A2(n7099), .ZN(n5000) );
  NAND2_X1 U6492 ( .A1(n4964), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4999) );
  NAND4_X1 U6493 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n8710)
         );
  NAND2_X1 U6494 ( .A1(n8710), .A2(n8382), .ZN(n5003) );
  XNOR2_X1 U6495 ( .A(n5004), .B(n5003), .ZN(n6562) );
  NAND2_X1 U6496 ( .A1(n5007), .A2(SI_5_), .ZN(n5008) );
  INV_X1 U6497 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6232) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6230) );
  OR2_X1 U6499 ( .A1(n4978), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6500 ( .A1(n5027), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5009) );
  XNOR2_X1 U6501 ( .A(n5009), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6377) );
  AOI22_X1 U6502 ( .A1(n5291), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6244), .B2(
        n6377), .ZN(n5010) );
  XNOR2_X1 U6503 ( .A(n6175), .B(n6841), .ZN(n5021) );
  NAND2_X1 U6504 ( .A1(n4995), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6505 ( .A1(n4955), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5018) );
  INV_X1 U6506 ( .A(n5013), .ZN(n5011) );
  NAND2_X1 U6507 ( .A1(n5011), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5032) );
  INV_X1 U6508 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6509 ( .A1(n5013), .A2(n5012), .ZN(n5014) );
  AND2_X1 U6510 ( .A1(n5032), .A2(n5014), .ZN(n6838) );
  NAND2_X1 U6511 ( .A1(n4956), .A2(n6838), .ZN(n5017) );
  NAND2_X1 U6512 ( .A1(n4964), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5016) );
  OR2_X1 U6513 ( .A1(n6970), .A2(n6174), .ZN(n5020) );
  NAND2_X1 U6514 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  OAI21_X1 U6515 ( .B1(n5021), .B2(n5020), .A(n5022), .ZN(n6647) );
  INV_X1 U6516 ( .A(n5025), .ZN(n5026) );
  MUX2_X1 U6517 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8377), .Z(n5051) );
  XNOR2_X1 U6518 ( .A(n5051), .B(SI_7_), .ZN(n5048) );
  XNOR2_X1 U6519 ( .A(n5050), .B(n5048), .ZN(n6233) );
  NAND2_X1 U6520 ( .A1(n6233), .A2(n8370), .ZN(n5030) );
  NOR2_X1 U6521 ( .A1(n5027), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5059) );
  OR2_X1 U6522 ( .A1(n5059), .A2(n9049), .ZN(n5028) );
  XNOR2_X1 U6523 ( .A(n5028), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U6524 ( .A1(n5291), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6244), .B2(
        n6365), .ZN(n5029) );
  XNOR2_X1 U6525 ( .A(n6975), .B(n6175), .ZN(n5038) );
  NAND2_X1 U6526 ( .A1(n4995), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6527 ( .A1(n4955), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5036) );
  INV_X1 U6528 ( .A(n5032), .ZN(n5031) );
  NAND2_X1 U6529 ( .A1(n5031), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5042) );
  INV_X1 U6530 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U6531 ( .A1(n5032), .A2(n6698), .ZN(n5033) );
  AND2_X1 U6532 ( .A1(n5042), .A2(n5033), .ZN(n6972) );
  NAND2_X1 U6533 ( .A1(n4956), .A2(n6972), .ZN(n5035) );
  NAND2_X1 U6534 ( .A1(n4964), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5034) );
  NOR2_X1 U6535 ( .A1(n6854), .A2(n6174), .ZN(n5040) );
  XNOR2_X1 U6536 ( .A(n5038), .B(n5040), .ZN(n6696) );
  INV_X1 U6537 ( .A(n5038), .ZN(n5039) );
  NAND2_X1 U6538 ( .A1(n4964), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6539 ( .A1(n4995), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6540 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  AND2_X1 U6541 ( .A1(n5080), .A2(n5043), .ZN(n8616) );
  NAND2_X1 U6542 ( .A1(n4956), .A2(n8616), .ZN(n5045) );
  NAND2_X1 U6543 ( .A1(n4955), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5044) );
  INV_X1 U6544 ( .A(n7023), .ZN(n8707) );
  NAND2_X1 U6545 ( .A1(n8707), .A2(n8382), .ZN(n5066) );
  INV_X1 U6546 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6547 ( .A1(n5050), .A2(n5049), .ZN(n5053) );
  NAND2_X1 U6548 ( .A1(n5051), .A2(SI_7_), .ZN(n5052) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6241) );
  MUX2_X1 U6550 ( .A(n6241), .B(n7868), .S(n8377), .Z(n5055) );
  INV_X1 U6551 ( .A(SI_8_), .ZN(n5054) );
  NAND2_X1 U6552 ( .A1(n5055), .A2(n5054), .ZN(n5070) );
  INV_X1 U6553 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6554 ( .A1(n5056), .A2(SI_8_), .ZN(n5057) );
  NAND2_X1 U6555 ( .A1(n5070), .A2(n5057), .ZN(n5068) );
  XNOR2_X1 U6556 ( .A(n5069), .B(n5068), .ZN(n6238) );
  NAND2_X1 U6557 ( .A1(n6238), .A2(n8370), .ZN(n5064) );
  INV_X1 U6558 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6559 ( .A1(n5059), .A2(n5058), .ZN(n5061) );
  NAND2_X1 U6560 ( .A1(n5061), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5060) );
  MUX2_X1 U6561 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5060), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5062) );
  AOI22_X1 U6562 ( .A1(n5291), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6244), .B2(
        n6511), .ZN(n5063) );
  NAND2_X1 U6563 ( .A1(n5064), .A2(n5063), .ZN(n8615) );
  XNOR2_X1 U6564 ( .A(n8615), .B(n5468), .ZN(n5065) );
  XOR2_X1 U6565 ( .A(n5066), .B(n5065), .Z(n8610) );
  INV_X1 U6566 ( .A(n5065), .ZN(n5067) );
  INV_X1 U6567 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6256) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6250) );
  MUX2_X1 U6569 ( .A(n6256), .B(n6250), .S(n8377), .Z(n5072) );
  INV_X1 U6570 ( .A(SI_9_), .ZN(n5071) );
  NAND2_X1 U6571 ( .A1(n5072), .A2(n5071), .ZN(n5091) );
  INV_X1 U6572 ( .A(n5072), .ZN(n5073) );
  NAND2_X1 U6573 ( .A1(n5073), .A2(SI_9_), .ZN(n5074) );
  XNOR2_X1 U6574 ( .A(n5090), .B(n4855), .ZN(n6249) );
  NAND2_X1 U6575 ( .A1(n6249), .A2(n8370), .ZN(n5077) );
  NAND2_X1 U6576 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5075) );
  XNOR2_X1 U6577 ( .A(n5075), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U6578 ( .A1(n5291), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6244), .B2(
        n6626), .ZN(n5076) );
  NAND2_X1 U6579 ( .A1(n5077), .A2(n5076), .ZN(n7028) );
  XNOR2_X1 U6580 ( .A(n7028), .B(n6175), .ZN(n5087) );
  NAND2_X1 U6581 ( .A1(n4995), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6582 ( .A1(n4955), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5084) );
  INV_X1 U6583 ( .A(n5080), .ZN(n5078) );
  INV_X1 U6584 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6585 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  AND2_X1 U6586 ( .A1(n5110), .A2(n5081), .ZN(n7031) );
  NAND2_X1 U6587 ( .A1(n4956), .A2(n7031), .ZN(n5083) );
  NAND2_X1 U6588 ( .A1(n4964), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5082) );
  OR2_X1 U6589 ( .A1(n7008), .A2(n6174), .ZN(n5086) );
  NAND2_X1 U6590 ( .A1(n5087), .A2(n5086), .ZN(n5088) );
  OAI21_X1 U6591 ( .B1(n5087), .B2(n5086), .A(n5088), .ZN(n6867) );
  INV_X1 U6592 ( .A(n5088), .ZN(n5089) );
  MUX2_X1 U6593 ( .A(n6270), .B(n6274), .S(n8377), .Z(n5094) );
  INV_X1 U6594 ( .A(SI_10_), .ZN(n5093) );
  NAND2_X1 U6595 ( .A1(n5094), .A2(n5093), .ZN(n5117) );
  INV_X1 U6596 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6597 ( .A1(n5095), .A2(SI_10_), .ZN(n5096) );
  NAND2_X1 U6598 ( .A1(n6269), .A2(n8370), .ZN(n5099) );
  OAI21_X1 U6599 ( .B1(n5097), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U6600 ( .A(n5120), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U6601 ( .A1(n5291), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6244), .B2(
        n6788), .ZN(n5098) );
  XNOR2_X1 U6602 ( .A(n9941), .B(n5468), .ZN(n5105) );
  NAND2_X1 U6603 ( .A1(n4995), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6604 ( .A1(n4964), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U6605 ( .A(n5110), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U6606 ( .A1(n4956), .A2(n6947), .ZN(n5101) );
  NAND2_X1 U6607 ( .A1(n4955), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5100) );
  INV_X1 U6608 ( .A(n7111), .ZN(n8705) );
  NAND2_X1 U6609 ( .A1(n8705), .A2(n8382), .ZN(n5104) );
  XNOR2_X1 U6610 ( .A(n5105), .B(n5104), .ZN(n6945) );
  INV_X1 U6611 ( .A(n5104), .ZN(n5106) );
  NAND2_X1 U6612 ( .A1(n4995), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6613 ( .A1(n4955), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5114) );
  INV_X1 U6614 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5108) );
  INV_X1 U6615 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5107) );
  OAI21_X1 U6616 ( .B1(n5110), .B2(n5108), .A(n5107), .ZN(n5111) );
  NAND2_X1 U6617 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5109) );
  AND2_X1 U6618 ( .A1(n5111), .A2(n5142), .ZN(n7142) );
  NAND2_X1 U6619 ( .A1(n4956), .A2(n7142), .ZN(n5113) );
  NAND2_X1 U6620 ( .A1(n4964), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6621 ( .A1(n8704), .A2(n8382), .ZN(n5126) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5118) );
  MUX2_X1 U6623 ( .A(n5118), .B(n6271), .S(n8377), .Z(n5128) );
  XNOR2_X1 U6624 ( .A(n5128), .B(SI_11_), .ZN(n5127) );
  XNOR2_X1 U6625 ( .A(n5131), .B(n5127), .ZN(n6257) );
  NAND2_X1 U6626 ( .A1(n6257), .A2(n8370), .ZN(n5124) );
  NAND2_X1 U6627 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  NAND2_X1 U6628 ( .A1(n5121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6629 ( .A(n5122), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7047) );
  AOI22_X1 U6630 ( .A1(n5291), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6244), .B2(
        n7047), .ZN(n5123) );
  NAND2_X1 U6631 ( .A1(n5124), .A2(n5123), .ZN(n7211) );
  XNOR2_X1 U6632 ( .A(n7211), .B(n5468), .ZN(n5125) );
  XOR2_X1 U6633 ( .A(n5126), .B(n5125), .Z(n7136) );
  INV_X1 U6634 ( .A(n5127), .ZN(n5130) );
  INV_X1 U6635 ( .A(n5128), .ZN(n5129) );
  INV_X1 U6636 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5133) );
  INV_X1 U6637 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5132) );
  MUX2_X1 U6638 ( .A(n5133), .B(n5132), .S(n8377), .Z(n5135) );
  INV_X1 U6639 ( .A(SI_12_), .ZN(n5134) );
  NAND2_X1 U6640 ( .A1(n5135), .A2(n5134), .ZN(n5158) );
  INV_X1 U6641 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6642 ( .A1(n5136), .A2(SI_12_), .ZN(n5137) );
  NAND2_X1 U6643 ( .A1(n5158), .A2(n5137), .ZN(n5159) );
  XNOR2_X1 U6644 ( .A(n5160), .B(n5159), .ZN(n6300) );
  NAND2_X1 U6645 ( .A1(n6300), .A2(n8370), .ZN(n5140) );
  NAND2_X1 U6646 ( .A1(n4332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  XNOR2_X1 U6647 ( .A(n5138), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U6648 ( .A1(n5291), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6244), .B2(
        n7087), .ZN(n5139) );
  XNOR2_X1 U6649 ( .A(n9956), .B(n5468), .ZN(n5148) );
  XNOR2_X1 U6650 ( .A(n5150), .B(n5148), .ZN(n7264) );
  NAND2_X1 U6651 ( .A1(n4995), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6652 ( .A1(n4964), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5146) );
  INV_X1 U6653 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U6654 ( .A1(n5142), .A2(n7784), .ZN(n5143) );
  AND2_X1 U6655 ( .A1(n5152), .A2(n5143), .ZN(n7217) );
  NAND2_X1 U6656 ( .A1(n4956), .A2(n7217), .ZN(n5145) );
  NAND2_X1 U6657 ( .A1(n4955), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5144) );
  NAND4_X1 U6658 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n8703)
         );
  INV_X1 U6659 ( .A(n8703), .ZN(n7443) );
  NOR2_X1 U6660 ( .A1(n7443), .A2(n6174), .ZN(n7265) );
  INV_X1 U6661 ( .A(n5148), .ZN(n5149) );
  AOI21_X1 U6662 ( .B1(n7264), .B2(n7265), .A(n5151), .ZN(n7539) );
  NAND2_X1 U6663 ( .A1(n4995), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6664 ( .A1(n4964), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6665 ( .A1(n5152), .A2(n7090), .ZN(n5153) );
  AND2_X1 U6666 ( .A1(n5182), .A2(n5153), .ZN(n7534) );
  NAND2_X1 U6667 ( .A1(n4956), .A2(n7534), .ZN(n5155) );
  NAND2_X1 U6668 ( .A1(n4955), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6669 ( .A1(n8702), .A2(n8382), .ZN(n5170) );
  INV_X1 U6670 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U6671 ( .A(n6499), .B(n5161), .S(n8377), .Z(n5163) );
  INV_X1 U6672 ( .A(SI_13_), .ZN(n5162) );
  NAND2_X1 U6673 ( .A1(n5163), .A2(n5162), .ZN(n5194) );
  INV_X1 U6674 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6675 ( .A1(n5164), .A2(SI_13_), .ZN(n5165) );
  XNOR2_X1 U6676 ( .A(n5174), .B(n5173), .ZN(n6480) );
  NAND2_X1 U6677 ( .A1(n6480), .A2(n8370), .ZN(n5168) );
  OR2_X1 U6678 ( .A1(n5166), .A2(n9049), .ZN(n5177) );
  XNOR2_X1 U6679 ( .A(n5177), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7198) );
  AOI22_X1 U6680 ( .A1(n5291), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6244), .B2(
        n7198), .ZN(n5167) );
  XNOR2_X1 U6681 ( .A(n9025), .B(n5468), .ZN(n5169) );
  XOR2_X1 U6682 ( .A(n5170), .B(n5169), .Z(n7540) );
  INV_X1 U6683 ( .A(n5170), .ZN(n5171) );
  INV_X1 U6684 ( .A(n7493), .ZN(n5191) );
  NAND2_X1 U6685 ( .A1(n5174), .A2(n5173), .ZN(n5196) );
  NAND2_X1 U6686 ( .A1(n5196), .A2(n5194), .ZN(n5175) );
  MUX2_X1 U6687 ( .A(n6552), .B(n6527), .S(n8377), .Z(n5197) );
  XNOR2_X1 U6688 ( .A(n5197), .B(SI_14_), .ZN(n5193) );
  XNOR2_X1 U6689 ( .A(n5175), .B(n5193), .ZN(n6526) );
  NAND2_X1 U6690 ( .A1(n6526), .A2(n8370), .ZN(n5180) );
  NAND2_X1 U6691 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6692 ( .A1(n5178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6693 ( .A(n5206), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U6694 ( .A1(n5291), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6244), .B2(
        n7418), .ZN(n5179) );
  XNOR2_X1 U6695 ( .A(n9020), .B(n6175), .ZN(n5189) );
  NAND2_X1 U6696 ( .A1(n4995), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6697 ( .A1(n4964), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6698 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  AND2_X1 U6699 ( .A1(n5221), .A2(n5183), .ZN(n7500) );
  NAND2_X1 U6700 ( .A1(n4956), .A2(n7500), .ZN(n5185) );
  NAND2_X1 U6701 ( .A1(n4955), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6702 ( .A1(n7600), .A2(n6174), .ZN(n5188) );
  NAND2_X1 U6703 ( .A1(n5189), .A2(n5188), .ZN(n5192) );
  OAI21_X1 U6704 ( .B1(n5189), .B2(n5188), .A(n5192), .ZN(n7494) );
  INV_X1 U6705 ( .A(n7494), .ZN(n5190) );
  NAND2_X2 U6706 ( .A1(n5191), .A2(n5190), .ZN(n7491) );
  NAND2_X1 U6707 ( .A1(n5196), .A2(n5195), .ZN(n5200) );
  INV_X1 U6708 ( .A(n5197), .ZN(n5198) );
  NAND2_X1 U6709 ( .A1(n5198), .A2(SI_14_), .ZN(n5199) );
  MUX2_X1 U6710 ( .A(n6613), .B(n6615), .S(n8377), .Z(n5202) );
  INV_X1 U6711 ( .A(SI_15_), .ZN(n5201) );
  NAND2_X1 U6712 ( .A1(n5202), .A2(n5201), .ZN(n5227) );
  INV_X1 U6713 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6714 ( .A1(n5203), .A2(SI_15_), .ZN(n5204) );
  NAND2_X1 U6715 ( .A1(n5227), .A2(n5204), .ZN(n5228) );
  XNOR2_X1 U6716 ( .A(n5229), .B(n5228), .ZN(n6612) );
  NAND2_X1 U6717 ( .A1(n6612), .A2(n8370), .ZN(n5210) );
  NAND2_X1 U6718 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  NAND2_X1 U6719 ( .A1(n5207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6720 ( .A(n5208), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7960) );
  AOI22_X1 U6721 ( .A1(n5291), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6244), .B2(
        n7960), .ZN(n5209) );
  XNOR2_X1 U6722 ( .A(n9015), .B(n5468), .ZN(n5215) );
  NAND2_X1 U6723 ( .A1(n4964), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6724 ( .A1(n4995), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6725 ( .A(n5221), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U6726 ( .A1(n4956), .A2(n7597), .ZN(n5212) );
  NAND2_X1 U6727 ( .A1(n4955), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6728 ( .A1(n8700), .A2(n8382), .ZN(n7595) );
  INV_X1 U6729 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6730 ( .A1(n4964), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6731 ( .A1(n4995), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5225) );
  AND2_X1 U6732 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5217) );
  INV_X1 U6733 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5220) );
  INV_X1 U6734 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5219) );
  OAI21_X1 U6735 ( .B1(n5221), .B2(n5220), .A(n5219), .ZN(n5222) );
  AND2_X1 U6736 ( .A1(n5245), .A2(n5222), .ZN(n7684) );
  NAND2_X1 U6737 ( .A1(n4956), .A2(n7684), .ZN(n5224) );
  NAND2_X1 U6738 ( .A1(n4955), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5223) );
  NOR2_X1 U6739 ( .A1(n8646), .A2(n6174), .ZN(n5241) );
  MUX2_X1 U6740 ( .A(n5231), .B(n5230), .S(n8377), .Z(n5233) );
  NAND2_X1 U6741 ( .A1(n5233), .A2(n5232), .ZN(n5253) );
  INV_X1 U6742 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6743 ( .A1(n5234), .A2(SI_16_), .ZN(n5235) );
  XNOR2_X1 U6744 ( .A(n5252), .B(n5251), .ZN(n6575) );
  NAND2_X1 U6745 ( .A1(n6575), .A2(n8370), .ZN(n5239) );
  OR2_X1 U6746 ( .A1(n5236), .A2(n9049), .ZN(n5237) );
  XNOR2_X1 U6747 ( .A(n5237), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8720) );
  AOI22_X1 U6748 ( .A1(n5291), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6244), .B2(
        n8720), .ZN(n5238) );
  XNOR2_X1 U6749 ( .A(n9010), .B(n5468), .ZN(n5240) );
  NOR2_X1 U6750 ( .A1(n5240), .A2(n5241), .ZN(n5242) );
  AOI21_X1 U6751 ( .B1(n5241), .B2(n5240), .A(n5242), .ZN(n7680) );
  NAND2_X1 U6752 ( .A1(n7679), .A2(n7680), .ZN(n7678) );
  INV_X1 U6753 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6754 ( .A1(n4995), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6755 ( .A1(n4955), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5249) );
  INV_X1 U6756 ( .A(n5245), .ZN(n5244) );
  NAND2_X1 U6757 ( .A1(n5244), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5272) );
  INV_X1 U6758 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U6759 ( .A1(n5245), .A2(n8730), .ZN(n5246) );
  AND2_X1 U6760 ( .A1(n5272), .A2(n5246), .ZN(n8643) );
  NAND2_X1 U6761 ( .A1(n4956), .A2(n8643), .ZN(n5248) );
  NAND2_X1 U6762 ( .A1(n4964), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5247) );
  INV_X1 U6763 ( .A(n8686), .ZN(n8916) );
  NAND2_X1 U6764 ( .A1(n8916), .A2(n8382), .ZN(n5259) );
  MUX2_X1 U6765 ( .A(n7863), .B(n5254), .S(n8377), .Z(n5264) );
  XNOR2_X1 U6766 ( .A(n5264), .B(SI_17_), .ZN(n5263) );
  NAND2_X1 U6767 ( .A1(n6666), .A2(n8370), .ZN(n5258) );
  NAND2_X1 U6768 ( .A1(n5255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5256) );
  XNOR2_X1 U6769 ( .A(n5256), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8732) );
  AOI22_X1 U6770 ( .A1(n5291), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6244), .B2(
        n8732), .ZN(n5257) );
  XNOR2_X1 U6771 ( .A(n9007), .B(n5468), .ZN(n5261) );
  XOR2_X1 U6772 ( .A(n5259), .B(n5261), .Z(n8641) );
  INV_X1 U6773 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6774 ( .A1(n5261), .A2(n5260), .ZN(n5262) );
  INV_X1 U6775 ( .A(n5263), .ZN(n5267) );
  INV_X1 U6776 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6777 ( .A1(n5265), .A2(SI_17_), .ZN(n5266) );
  MUX2_X1 U6778 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8377), .Z(n5284) );
  XNOR2_X1 U6779 ( .A(n5284), .B(SI_18_), .ZN(n5281) );
  XNOR2_X1 U6780 ( .A(n5283), .B(n5281), .ZN(n6713) );
  NAND2_X1 U6781 ( .A1(n6713), .A2(n8370), .ZN(n5271) );
  XNOR2_X1 U6782 ( .A(n5269), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8749) );
  AOI22_X1 U6783 ( .A1(n5291), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6244), .B2(
        n8749), .ZN(n5270) );
  XNOR2_X1 U6784 ( .A(n9000), .B(n5468), .ZN(n5280) );
  NAND2_X1 U6785 ( .A1(n4964), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6786 ( .A1(n4995), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6787 ( .A1(n5272), .A2(n8681), .ZN(n5273) );
  AND2_X1 U6788 ( .A1(n5298), .A2(n5273), .ZN(n8906) );
  NAND2_X1 U6789 ( .A1(n4956), .A2(n8906), .ZN(n5275) );
  NAND2_X1 U6790 ( .A1(n4955), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6791 ( .A1(n8698), .A2(n8382), .ZN(n5278) );
  XNOR2_X1 U6792 ( .A(n5280), .B(n5278), .ZN(n8678) );
  INV_X1 U6793 ( .A(n5278), .ZN(n5279) );
  INV_X1 U6794 ( .A(n5281), .ZN(n5282) );
  NAND2_X1 U6795 ( .A1(n5284), .A2(SI_18_), .ZN(n5285) );
  MUX2_X1 U6796 ( .A(n6800), .B(n6802), .S(n8377), .Z(n5287) );
  INV_X1 U6797 ( .A(SI_19_), .ZN(n5286) );
  NAND2_X1 U6798 ( .A1(n5287), .A2(n5286), .ZN(n5329) );
  INV_X1 U6799 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6800 ( .A1(n5288), .A2(SI_19_), .ZN(n5289) );
  NAND2_X1 U6801 ( .A1(n5329), .A2(n5289), .ZN(n5308) );
  XNOR2_X1 U6802 ( .A(n5309), .B(n5308), .ZN(n6799) );
  NAND2_X1 U6803 ( .A1(n6799), .A2(n8370), .ZN(n5293) );
  AOI22_X1 U6804 ( .A1(n5291), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5290), .B2(
        n6244), .ZN(n5292) );
  XNOR2_X1 U6805 ( .A(n8996), .B(n6175), .ZN(n5303) );
  NAND2_X1 U6806 ( .A1(n4995), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6807 ( .A1(n4964), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5294) );
  AND2_X1 U6808 ( .A1(n5295), .A2(n5294), .ZN(n5302) );
  INV_X1 U6809 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6810 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6811 ( .A1(n5318), .A2(n5299), .ZN(n8606) );
  OR2_X1 U6812 ( .A1(n8606), .A2(n6180), .ZN(n5301) );
  NAND2_X1 U6813 ( .A1(n4955), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6814 ( .A1(n8918), .A2(n8382), .ZN(n5304) );
  NAND2_X1 U6815 ( .A1(n5303), .A2(n5304), .ZN(n8601) );
  NAND2_X1 U6816 ( .A1(n8602), .A2(n8601), .ZN(n5307) );
  INV_X1 U6817 ( .A(n5303), .ZN(n5306) );
  INV_X1 U6818 ( .A(n5304), .ZN(n5305) );
  NAND2_X1 U6819 ( .A1(n5306), .A2(n5305), .ZN(n8600) );
  NAND2_X1 U6820 ( .A1(n5307), .A2(n8600), .ZN(n8658) );
  NAND2_X1 U6821 ( .A1(n5332), .A2(n5329), .ZN(n5314) );
  MUX2_X1 U6822 ( .A(n7854), .B(n6927), .S(n8377), .Z(n5311) );
  INV_X1 U6823 ( .A(SI_20_), .ZN(n5310) );
  NAND2_X1 U6824 ( .A1(n5311), .A2(n5310), .ZN(n5328) );
  INV_X1 U6825 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6826 ( .A1(n5312), .A2(SI_20_), .ZN(n5330) );
  AND2_X1 U6827 ( .A1(n5328), .A2(n5330), .ZN(n5313) );
  NAND2_X1 U6828 ( .A1(n6926), .A2(n8370), .ZN(n5316) );
  OR2_X1 U6829 ( .A1(n4947), .A2(n7854), .ZN(n5315) );
  XNOR2_X1 U6830 ( .A(n8990), .B(n5468), .ZN(n5325) );
  INV_X1 U6831 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6832 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  AND2_X1 U6833 ( .A1(n5337), .A2(n5319), .ZN(n8893) );
  NAND2_X1 U6834 ( .A1(n8893), .A2(n4956), .ZN(n5322) );
  AOI22_X1 U6835 ( .A1(n4995), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n4964), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6836 ( .A1(n4955), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6837 ( .A1(n8881), .A2(n8382), .ZN(n5323) );
  XNOR2_X1 U6838 ( .A(n5325), .B(n5323), .ZN(n8657) );
  NAND2_X1 U6839 ( .A1(n8658), .A2(n8657), .ZN(n5327) );
  INV_X1 U6840 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U6841 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  MUX2_X1 U6842 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8377), .Z(n5345) );
  XNOR2_X1 U6843 ( .A(n5345), .B(n7919), .ZN(n5342) );
  XNOR2_X1 U6844 ( .A(n5344), .B(n5342), .ZN(n7037) );
  NAND2_X1 U6845 ( .A1(n7037), .A2(n8370), .ZN(n5334) );
  INV_X1 U6846 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7038) );
  OR2_X1 U6847 ( .A1(n4947), .A2(n7038), .ZN(n5333) );
  XNOR2_X1 U6848 ( .A(n8985), .B(n5468), .ZN(n5364) );
  INV_X1 U6849 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6850 ( .A1(n5337), .A2(n5336), .ZN(n5338) );
  NAND2_X1 U6851 ( .A1(n5354), .A2(n5338), .ZN(n8874) );
  OR2_X1 U6852 ( .A1(n8874), .A2(n6180), .ZN(n5341) );
  AOI22_X1 U6853 ( .A1(n4955), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n4995), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6854 ( .A1(n4964), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6855 ( .A1(n8897), .A2(n8382), .ZN(n5362) );
  XNOR2_X1 U6856 ( .A(n5364), .B(n5362), .ZN(n8622) );
  INV_X1 U6857 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6858 ( .A1(n5345), .A2(SI_21_), .ZN(n5346) );
  MUX2_X1 U6859 ( .A(n8021), .B(n7242), .S(n8377), .Z(n5349) );
  INV_X1 U6860 ( .A(SI_22_), .ZN(n5348) );
  NAND2_X1 U6861 ( .A1(n5349), .A2(n5348), .ZN(n5367) );
  INV_X1 U6862 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6863 ( .A1(n5350), .A2(SI_22_), .ZN(n5351) );
  NAND2_X1 U6864 ( .A1(n5367), .A2(n5351), .ZN(n5368) );
  XNOR2_X1 U6865 ( .A(n5369), .B(n5368), .ZN(n7241) );
  NAND2_X1 U6866 ( .A1(n7241), .A2(n8370), .ZN(n5353) );
  OR2_X1 U6867 ( .A1(n4947), .A2(n8021), .ZN(n5352) );
  XNOR2_X1 U6868 ( .A(n8980), .B(n6175), .ZN(n8667) );
  INV_X1 U6869 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U6870 ( .A1(n5354), .A2(n8671), .ZN(n5355) );
  AND2_X1 U6871 ( .A1(n5377), .A2(n5355), .ZN(n8856) );
  NAND2_X1 U6872 ( .A1(n8856), .A2(n4956), .ZN(n5361) );
  INV_X1 U6873 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7871) );
  INV_X1 U6874 ( .A(n4955), .ZN(n5358) );
  NAND2_X1 U6875 ( .A1(n4995), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6876 ( .A1(n4964), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5356) );
  OAI211_X1 U6877 ( .C1(n7871), .C2(n5358), .A(n5357), .B(n5356), .ZN(n5359)
         );
  INV_X1 U6878 ( .A(n5359), .ZN(n5360) );
  OR2_X1 U6879 ( .A1(n8837), .A2(n6174), .ZN(n8668) );
  INV_X1 U6880 ( .A(n5362), .ZN(n5363) );
  NAND2_X1 U6881 ( .A1(n5364), .A2(n5363), .ZN(n8665) );
  MUX2_X1 U6882 ( .A(n7244), .B(n7248), .S(n8377), .Z(n5371) );
  INV_X1 U6883 ( .A(SI_23_), .ZN(n5370) );
  NAND2_X1 U6884 ( .A1(n5371), .A2(n5370), .ZN(n5391) );
  INV_X1 U6885 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6886 ( .A1(n5372), .A2(SI_23_), .ZN(n5373) );
  XNOR2_X1 U6887 ( .A(n5390), .B(n5389), .ZN(n7245) );
  NAND2_X1 U6888 ( .A1(n7245), .A2(n8370), .ZN(n5375) );
  OR2_X1 U6889 ( .A1(n4947), .A2(n7244), .ZN(n5374) );
  XNOR2_X1 U6890 ( .A(n8974), .B(n5468), .ZN(n5385) );
  NAND2_X1 U6891 ( .A1(n5384), .A2(n5385), .ZN(n8591) );
  INV_X1 U6892 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6893 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6894 ( .A1(n5397), .A2(n5378), .ZN(n8845) );
  INV_X1 U6895 ( .A(n8845), .ZN(n5383) );
  INV_X1 U6896 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U6897 ( .A1(n4964), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6898 ( .A1(n4955), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5379) );
  OAI211_X1 U6899 ( .C1(n5381), .C2(n8846), .A(n5380), .B(n5379), .ZN(n5382)
         );
  NOR2_X1 U6900 ( .A1(n8864), .A2(n6174), .ZN(n8594) );
  NAND2_X1 U6901 ( .A1(n8591), .A2(n8594), .ZN(n5388) );
  INV_X1 U6902 ( .A(n5384), .ZN(n5387) );
  INV_X1 U6903 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6904 ( .A1(n5387), .A2(n5386), .ZN(n8592) );
  NAND2_X1 U6905 ( .A1(n5388), .A2(n8592), .ZN(n5403) );
  NAND2_X1 U6906 ( .A1(n5390), .A2(n5389), .ZN(n5392) );
  MUX2_X1 U6907 ( .A(n7322), .B(n7320), .S(n8377), .Z(n5411) );
  XNOR2_X1 U6908 ( .A(n5411), .B(SI_24_), .ZN(n5408) );
  XNOR2_X1 U6909 ( .A(n5410), .B(n5408), .ZN(n7319) );
  NAND2_X1 U6910 ( .A1(n7319), .A2(n8370), .ZN(n5394) );
  OR2_X1 U6911 ( .A1(n4317), .A2(n7322), .ZN(n5393) );
  XNOR2_X1 U6912 ( .A(n8968), .B(n6175), .ZN(n5404) );
  XNOR2_X1 U6913 ( .A(n5403), .B(n5404), .ZN(n8650) );
  INV_X1 U6914 ( .A(n5397), .ZN(n5395) );
  NAND2_X1 U6915 ( .A1(n5395), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5421) );
  INV_X1 U6916 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6917 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  AND2_X1 U6918 ( .A1(n5421), .A2(n5398), .ZN(n8816) );
  INV_X1 U6919 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6920 ( .A1(n4995), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6921 ( .A1(n4955), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5399) );
  OAI211_X1 U6922 ( .C1(n5401), .C2(n5015), .A(n5400), .B(n5399), .ZN(n5402)
         );
  AOI21_X1 U6923 ( .B1(n8816), .B2(n4956), .A(n5402), .ZN(n8838) );
  NOR2_X1 U6924 ( .A1(n8838), .A2(n6174), .ZN(n8651) );
  NAND2_X1 U6925 ( .A1(n8650), .A2(n8651), .ZN(n5407) );
  INV_X1 U6926 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6927 ( .A1(n5403), .A2(n5405), .ZN(n5406) );
  INV_X1 U6928 ( .A(n5408), .ZN(n5409) );
  INV_X1 U6929 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6930 ( .A1(n5412), .A2(SI_24_), .ZN(n5413) );
  INV_X1 U6931 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7466) );
  INV_X1 U6932 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7469) );
  MUX2_X1 U6933 ( .A(n7466), .B(n7469), .S(n8377), .Z(n5415) );
  INV_X1 U6934 ( .A(SI_25_), .ZN(n5414) );
  NAND2_X1 U6935 ( .A1(n5415), .A2(n5414), .ZN(n5457) );
  INV_X1 U6936 ( .A(n5415), .ZN(n5416) );
  NAND2_X1 U6937 ( .A1(n5416), .A2(SI_25_), .ZN(n5417) );
  NAND2_X1 U6938 ( .A1(n5457), .A2(n5417), .ZN(n5455) );
  XNOR2_X1 U6939 ( .A(n5461), .B(n5455), .ZN(n7464) );
  NAND2_X1 U6940 ( .A1(n7464), .A2(n8370), .ZN(n5419) );
  OR2_X1 U6941 ( .A1(n4947), .A2(n7466), .ZN(n5418) );
  XNOR2_X1 U6942 ( .A(n8965), .B(n5468), .ZN(n8631) );
  NAND2_X1 U6943 ( .A1(n8629), .A2(n8631), .ZN(n5429) );
  INV_X1 U6944 ( .A(n5421), .ZN(n5420) );
  NAND2_X1 U6945 ( .A1(n5420), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5443) );
  INV_X1 U6946 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U6947 ( .A1(n5421), .A2(n8635), .ZN(n5422) );
  NAND2_X1 U6948 ( .A1(n5443), .A2(n5422), .ZN(n8807) );
  OR2_X1 U6949 ( .A1(n8807), .A2(n6180), .ZN(n5428) );
  INV_X1 U6950 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6951 ( .A1(n4955), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6952 ( .A1(n4995), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5423) );
  OAI211_X1 U6953 ( .C1(n5015), .C2(n5425), .A(n5424), .B(n5423), .ZN(n5426)
         );
  INV_X1 U6954 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6955 ( .A1(n8696), .A2(n8382), .ZN(n8630) );
  NAND2_X1 U6956 ( .A1(n5429), .A2(n8630), .ZN(n5433) );
  INV_X1 U6957 ( .A(n8629), .ZN(n5431) );
  INV_X1 U6958 ( .A(n8631), .ZN(n5430) );
  NAND2_X1 U6959 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  OR2_X1 U6960 ( .A1(n5461), .A2(n5455), .ZN(n5434) );
  NAND2_X1 U6961 ( .A1(n5434), .A2(n5457), .ZN(n5439) );
  MUX2_X1 U6962 ( .A(n7762), .B(n7517), .S(n8377), .Z(n5436) );
  INV_X1 U6963 ( .A(SI_26_), .ZN(n5435) );
  NAND2_X1 U6964 ( .A1(n5436), .A2(n5435), .ZN(n5456) );
  INV_X1 U6965 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6966 ( .A1(n5437), .A2(SI_26_), .ZN(n5454) );
  AND2_X1 U6967 ( .A1(n5456), .A2(n5454), .ZN(n5438) );
  NAND2_X1 U6968 ( .A1(n7516), .A2(n8370), .ZN(n5441) );
  OR2_X1 U6969 ( .A1(n4947), .A2(n7762), .ZN(n5440) );
  XNOR2_X1 U6970 ( .A(n8039), .B(n6175), .ZN(n5452) );
  INV_X1 U6971 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6972 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  NAND2_X1 U6973 ( .A1(n8793), .A2(n4956), .ZN(n5450) );
  INV_X1 U6974 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6975 ( .A1(n4964), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6976 ( .A1(n4995), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5445) );
  OAI211_X1 U6977 ( .C1(n5447), .C2(n5358), .A(n5446), .B(n5445), .ZN(n5448)
         );
  INV_X1 U6978 ( .A(n5448), .ZN(n5449) );
  NAND2_X1 U6979 ( .A1(n5450), .A2(n5449), .ZN(n8695) );
  AND2_X1 U6980 ( .A1(n8695), .A2(n8382), .ZN(n5451) );
  NAND2_X1 U6981 ( .A1(n5452), .A2(n5451), .ZN(n5486) );
  OAI21_X1 U6982 ( .B1(n5452), .B2(n5451), .A(n5486), .ZN(n6163) );
  INV_X1 U6983 ( .A(n6163), .ZN(n5453) );
  INV_X1 U6984 ( .A(n5454), .ZN(n5459) );
  AND2_X1 U6985 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  INV_X1 U6986 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7551) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6062) );
  MUX2_X1 U6988 ( .A(n7551), .B(n6062), .S(n8377), .Z(n5463) );
  INV_X1 U6989 ( .A(SI_27_), .ZN(n5462) );
  NAND2_X1 U6990 ( .A1(n5463), .A2(n5462), .ZN(n6088) );
  INV_X1 U6991 ( .A(n5463), .ZN(n5464) );
  NAND2_X1 U6992 ( .A1(n5464), .A2(SI_27_), .ZN(n5465) );
  NAND2_X1 U6993 ( .A1(n7547), .A2(n8370), .ZN(n5467) );
  OR2_X1 U6994 ( .A1(n4317), .A2(n7551), .ZN(n5466) );
  XNOR2_X1 U6995 ( .A(n8954), .B(n5468), .ZN(n5480) );
  INV_X1 U6996 ( .A(n5480), .ZN(n5482) );
  INV_X1 U6997 ( .A(n5471), .ZN(n5469) );
  NAND2_X1 U6998 ( .A1(n5469), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5533) );
  INV_X1 U6999 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7000 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U7001 ( .A1(n5533), .A2(n5472), .ZN(n5521) );
  INV_X1 U7002 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7003 ( .A1(n4964), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7004 ( .A1(n4995), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5473) );
  OAI211_X1 U7005 ( .C1(n5475), .C2(n5358), .A(n5474), .B(n5473), .ZN(n5476)
         );
  INV_X1 U7006 ( .A(n5476), .ZN(n5477) );
  AND2_X1 U7007 ( .A1(n8694), .A2(n8382), .ZN(n5479) );
  INV_X1 U7008 ( .A(n5479), .ZN(n5481) );
  AOI21_X1 U7009 ( .B1(n5482), .B2(n5481), .A(n6179), .ZN(n5485) );
  INV_X1 U7010 ( .A(n5486), .ZN(n5483) );
  INV_X1 U7011 ( .A(n5485), .ZN(n5487) );
  NAND2_X1 U7012 ( .A1(n5488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5489) );
  MUX2_X1 U7013 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5489), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5490) );
  NAND2_X1 U7014 ( .A1(n5490), .A2(n4379), .ZN(n7465) );
  NAND2_X1 U7015 ( .A1(n5491), .A2(n7927), .ZN(n5492) );
  XNOR2_X1 U7016 ( .A(n7324), .B(P2_B_REG_SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7017 ( .A1(n4379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5496) );
  MUX2_X1 U7018 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5496), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5497) );
  NAND2_X1 U7019 ( .A1(n7465), .A2(n7546), .ZN(n9887) );
  NOR4_X1 U7020 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5508) );
  OR4_X1 U7021 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5505) );
  NOR4_X1 U7022 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5503) );
  NOR4_X1 U7023 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5502) );
  NOR4_X1 U7024 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5501) );
  NOR4_X1 U7025 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5500) );
  NAND4_X1 U7026 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .ZN(n5504)
         );
  NOR4_X1 U7027 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5505), .A4(n5504), .ZN(n5507) );
  NOR4_X1 U7028 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5506) );
  NAND3_X1 U7029 ( .A1(n5508), .A2(n5507), .A3(n5506), .ZN(n5509) );
  NAND2_X1 U7030 ( .A1(n5509), .A2(n5510), .ZN(n6806) );
  AND2_X1 U7031 ( .A1(n7324), .A2(n7546), .ZN(n9884) );
  INV_X1 U7032 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U7033 ( .A1(n6806), .A2(n6429), .ZN(n5512) );
  INV_X1 U7034 ( .A(n6246), .ZN(n5515) );
  NAND2_X1 U7035 ( .A1(n6352), .A2(n9955), .ZN(n5517) );
  INV_X1 U7036 ( .A(n8954), .ZN(n8773) );
  NAND3_X1 U7037 ( .A1(n4316), .A2(n5290), .A3(n5519), .ZN(n9030) );
  NAND2_X1 U7038 ( .A1(n5529), .A2(n6809), .ZN(n5524) );
  AND2_X1 U7039 ( .A1(n9879), .A2(n9897), .ZN(n5520) );
  INV_X1 U7040 ( .A(n5521), .ZN(n8771) );
  NAND2_X1 U7041 ( .A1(n5526), .A2(n6246), .ZN(n5522) );
  AND2_X1 U7042 ( .A1(n6350), .A2(n5522), .ZN(n5523) );
  NAND2_X1 U7043 ( .A1(n6341), .A2(n6242), .ZN(n5525) );
  INV_X1 U7044 ( .A(n8695), .ZN(n8775) );
  INV_X1 U7045 ( .A(n5526), .ZN(n5527) );
  INV_X1 U7046 ( .A(n8586), .ZN(n5528) );
  INV_X1 U7047 ( .A(n4310), .ZN(n5541) );
  INV_X1 U7048 ( .A(n5533), .ZN(n5531) );
  NAND2_X1 U7049 ( .A1(n5531), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8040) );
  INV_X1 U7050 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7051 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7052 ( .A1(n8040), .A2(n5534), .ZN(n8359) );
  INV_X1 U7053 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7054 ( .A1(n4964), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7055 ( .A1(n4995), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U7056 ( .C1(n5537), .C2(n5358), .A(n5536), .B(n5535), .ZN(n5538)
         );
  INV_X1 U7057 ( .A(n5538), .ZN(n5539) );
  INV_X1 U7058 ( .A(n8776), .ZN(n8693) );
  AOI22_X1 U7059 ( .A1(n8693), .A2(n8682), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n5542) );
  OAI21_X1 U7060 ( .B1(n8775), .B2(n8685), .A(n5542), .ZN(n5543) );
  AOI21_X1 U7061 ( .B1(n8771), .B2(n8680), .A(n5543), .ZN(n5544) );
  NAND2_X1 U7062 ( .A1(n5546), .A2(n4854), .ZN(P2_U3216) );
  NOR2_X1 U7063 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5555) );
  NOR2_X1 U7064 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5554) );
  NOR2_X1 U7065 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5553) );
  INV_X1 U7066 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5557) );
  INV_X2 U7067 ( .A(n5717), .ZN(n8005) );
  NAND2_X1 U7068 ( .A1(n6575), .A2(n8005), .ZN(n5563) );
  INV_X1 U7069 ( .A(n5560), .ZN(n5851) );
  NAND2_X1 U7070 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7071 ( .A(n5889), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9249) );
  AOI22_X1 U7072 ( .A1(n5928), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5927), .B2(
        n9249), .ZN(n5562) );
  NAND2_X1 U7073 ( .A1(n5563), .A2(n5562), .ZN(n7689) );
  NAND2_X1 U7074 ( .A1(n5606), .A2(n5567), .ZN(n5568) );
  NAND2_X1 U7075 ( .A1(n5574), .A2(n5569), .ZN(n5570) );
  NAND2_X1 U7076 ( .A1(n5575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7077 ( .A1(n5582), .A2(n5581), .ZN(n5576) );
  NAND2_X1 U7078 ( .A1(n4365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5580) );
  INV_X2 U7079 ( .A(n6055), .ZN(n6106) );
  NAND2_X1 U7080 ( .A1(n7689), .A2(n6106), .ZN(n5602) );
  INV_X1 U7081 ( .A(n5585), .ZN(n9604) );
  NAND2_X1 U7082 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7083 ( .A1(n5707), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5696) );
  NOR2_X1 U7084 ( .A1(n5696), .A2(n5611), .ZN(n5730) );
  NAND2_X1 U7085 ( .A1(n5730), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7086 ( .A1(n5816), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5836) );
  INV_X1 U7087 ( .A(n5873), .ZN(n5590) );
  INV_X1 U7088 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7089 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7090 ( .A1(n5894), .A2(n5591), .ZN(n9649) );
  INV_X1 U7091 ( .A(n9649), .ZN(n7632) );
  NAND2_X1 U7092 ( .A1(n6067), .A2(n7632), .ZN(n5599) );
  NAND2_X1 U7093 ( .A1(n5644), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5598) );
  NAND2_X2 U7094 ( .A1(n8366), .A2(n9611), .ZN(n5709) );
  INV_X1 U7095 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5593) );
  OR2_X1 U7096 ( .A1(n5709), .A2(n5593), .ZN(n5597) );
  INV_X1 U7097 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5595) );
  OR2_X1 U7098 ( .A1(n4315), .A2(n5595), .ZN(n5596) );
  INV_X1 U7099 ( .A(n6726), .ZN(n5600) );
  BUF_X4 U7100 ( .A(n5652), .Z(n6105) );
  NAND2_X1 U7101 ( .A1(n9484), .A2(n6105), .ZN(n5601) );
  NAND2_X1 U7102 ( .A1(n5602), .A2(n5601), .ZN(n5609) );
  INV_X1 U7103 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7104 ( .A1(n5607), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5608) );
  NAND2_X4 U7105 ( .A1(n6727), .A2(n6726), .ZN(n6744) );
  XNOR2_X1 U7106 ( .A(n5609), .B(n6744), .ZN(n5883) );
  INV_X1 U7107 ( .A(n7689), .ZN(n9638) );
  NAND2_X1 U7108 ( .A1(n6129), .A2(n8295), .ZN(n5610) );
  OAI22_X1 U7109 ( .A1(n9638), .A2(n6058), .B1(n7665), .B2(n6057), .ZN(n5884)
         );
  XNOR2_X1 U7110 ( .A(n5883), .B(n5884), .ZN(n9640) );
  NAND2_X1 U7111 ( .A1(n5644), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5617) );
  AND2_X1 U7112 ( .A1(n5696), .A2(n5611), .ZN(n5612) );
  NOR2_X1 U7113 ( .A1(n5730), .A2(n5612), .ZN(n7072) );
  NAND2_X1 U7114 ( .A1(n6067), .A2(n7072), .ZN(n5616) );
  INV_X1 U7115 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5613) );
  OR2_X1 U7116 ( .A1(n5709), .A2(n5613), .ZN(n5615) );
  INV_X1 U7117 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7073) );
  OR2_X1 U7118 ( .A1(n4315), .A2(n7073), .ZN(n5614) );
  NAND2_X1 U7119 ( .A1(n6233), .A2(n8005), .ZN(n5622) );
  INV_X1 U7120 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6236) );
  OR2_X1 U7121 ( .A1(n8006), .A2(n6236), .ZN(n5620) );
  NAND2_X1 U7122 ( .A1(n5618), .A2(n5702), .ZN(n5736) );
  NAND2_X1 U7123 ( .A1(n5736), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5619) );
  XNOR2_X1 U7124 ( .A(n5619), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9738) );
  INV_X1 U7125 ( .A(n9738), .ZN(n6445) );
  OAI22_X1 U7126 ( .A1(n7298), .A2(n6058), .B1(n9830), .B2(n6055), .ZN(n5623)
         );
  XNOR2_X1 U7127 ( .A(n5623), .B(n6744), .ZN(n7179) );
  INV_X1 U7128 ( .A(n7179), .ZN(n5729) );
  OAI22_X1 U7129 ( .A1(n7298), .A2(n6057), .B1(n9830), .B2(n6058), .ZN(n7178)
         );
  INV_X1 U7130 ( .A(n7178), .ZN(n5728) );
  NAND2_X1 U7131 ( .A1(n5644), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7132 ( .A1(n6067), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5628) );
  INV_X1 U7133 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5624) );
  OR2_X1 U7134 ( .A1(n5709), .A2(n5624), .ZN(n5627) );
  INV_X1 U7135 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5625) );
  OR2_X1 U7136 ( .A1(n4315), .A2(n5625), .ZN(n5626) );
  OR2_X1 U7137 ( .A1(n5630), .A2(n5557), .ZN(n5667) );
  XNOR2_X1 U7138 ( .A(n5667), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9694) );
  INV_X1 U7139 ( .A(n9694), .ZN(n6213) );
  OAI22_X1 U7140 ( .A1(n6913), .A2(n6058), .B1(n6896), .B2(n6055), .ZN(n5632)
         );
  XNOR2_X1 U7141 ( .A(n5632), .B(n6744), .ZN(n5634) );
  OAI22_X1 U7142 ( .A1(n6913), .A2(n6057), .B1(n6896), .B2(n6058), .ZN(n5633)
         );
  AOI21_X1 U7143 ( .B1(n5634), .B2(n5633), .A(n5659), .ZN(n6689) );
  NAND2_X1 U7144 ( .A1(n6067), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5638) );
  INV_X1 U7145 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5635) );
  OR2_X1 U7146 ( .A1(n5709), .A2(n5635), .ZN(n5637) );
  NAND2_X1 U7147 ( .A1(n5644), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5636) );
  AND4_X2 U7148 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(n6718)
         );
  INV_X1 U7149 ( .A(n9682), .ZN(n6215) );
  INV_X1 U7150 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6216) );
  OAI22_X1 U7151 ( .A1(n6718), .A2(n6058), .B1(n6760), .B2(n6055), .ZN(n5642)
         );
  INV_X1 U7152 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7153 ( .A1(n6067), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5647) );
  INV_X1 U7154 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6645) );
  OR2_X1 U7155 ( .A1(n5709), .A2(n6645), .ZN(n5646) );
  NAND2_X1 U7156 ( .A1(n5644), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5645) );
  INV_X1 U7157 ( .A(n6058), .ZN(n5652) );
  NAND2_X1 U7158 ( .A1(n6750), .A2(n5652), .ZN(n5651) );
  NAND2_X1 U7159 ( .A1(n8377), .A2(SI_0_), .ZN(n5649) );
  XNOR2_X1 U7160 ( .A(n5649), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9614) );
  MUX2_X1 U7161 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9614), .S(n8002), .Z(n6764) );
  INV_X1 U7162 ( .A(n6209), .ZN(n5653) );
  AOI22_X1 U7163 ( .A1(n6764), .A2(n6106), .B1(n5653), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7164 ( .A1(n6764), .A2(n5652), .ZN(n5655) );
  NAND2_X1 U7165 ( .A1(n5653), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7166 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  AND2_X1 U7167 ( .A1(n6756), .A2(n5652), .ZN(n5658) );
  AOI21_X1 U7168 ( .B1(n6717), .B2(n6101), .A(n5658), .ZN(n6657) );
  INV_X1 U7169 ( .A(n5659), .ZN(n5660) );
  INV_X1 U7170 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U7171 ( .A1(n6067), .A2(n6920), .ZN(n5666) );
  NAND2_X1 U7172 ( .A1(n5644), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5665) );
  INV_X1 U7173 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5661) );
  OR2_X1 U7174 ( .A1(n5709), .A2(n5661), .ZN(n5664) );
  INV_X1 U7175 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5662) );
  OR2_X1 U7176 ( .A1(n4314), .A2(n5662), .ZN(n5663) );
  INV_X1 U7177 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U7178 ( .A1(n5667), .A2(n7914), .ZN(n5668) );
  NAND2_X1 U7179 ( .A1(n5668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U7180 ( .A(n5669), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6320) );
  INV_X1 U7181 ( .A(n6320), .ZN(n6335) );
  OR2_X1 U7182 ( .A1(n5717), .A2(n6222), .ZN(n5671) );
  OR2_X1 U7183 ( .A1(n8006), .A2(n6217), .ZN(n5670) );
  OAI211_X1 U7184 ( .C1(n8002), .C2(n6335), .A(n5671), .B(n5670), .ZN(n6921)
         );
  INV_X1 U7185 ( .A(n6921), .ZN(n9811) );
  OAI22_X1 U7186 ( .A1(n6930), .A2(n6057), .B1(n9811), .B2(n6058), .ZN(n5674)
         );
  OAI22_X1 U7187 ( .A1(n6930), .A2(n6058), .B1(n9811), .B2(n6055), .ZN(n5672)
         );
  XNOR2_X1 U7188 ( .A(n5672), .B(n6744), .ZN(n5673) );
  XOR2_X1 U7189 ( .A(n5674), .B(n5673), .Z(n6705) );
  INV_X1 U7190 ( .A(n5673), .ZN(n5676) );
  NAND2_X1 U7191 ( .A1(n5644), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5683) );
  INV_X1 U7192 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U7193 ( .A(n5678), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7194 ( .A1(n6067), .A2(n6202), .ZN(n5682) );
  INV_X1 U7195 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5679) );
  OR2_X1 U7196 ( .A1(n5709), .A2(n5679), .ZN(n5681) );
  INV_X1 U7197 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6937) );
  OR2_X1 U7198 ( .A1(n4314), .A2(n6937), .ZN(n5680) );
  NAND2_X1 U7199 ( .A1(n5684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5685) );
  MUX2_X1 U7200 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5685), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5687) );
  NAND2_X1 U7201 ( .A1(n5687), .A2(n5686), .ZN(n6316) );
  INV_X1 U7202 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7203 ( .A1(n8006), .A2(n6226), .ZN(n5689) );
  OR2_X1 U7204 ( .A1(n5717), .A2(n6225), .ZN(n5688) );
  OAI211_X1 U7205 ( .C1(n8002), .C2(n6316), .A(n5689), .B(n5688), .ZN(n6993)
         );
  INV_X1 U7206 ( .A(n6993), .ZN(n6941) );
  OAI22_X1 U7207 ( .A1(n6912), .A2(n6058), .B1(n6941), .B2(n6055), .ZN(n5690)
         );
  XNOR2_X1 U7208 ( .A(n5690), .B(n6024), .ZN(n5692) );
  INV_X1 U7209 ( .A(n6912), .ZN(n9209) );
  AND2_X1 U7210 ( .A1(n6993), .A2(n6105), .ZN(n5691) );
  AOI21_X1 U7211 ( .B1(n9209), .B2(n6101), .A(n5691), .ZN(n5693) );
  AND2_X1 U7212 ( .A1(n5692), .A2(n5693), .ZN(n6197) );
  INV_X1 U7213 ( .A(n5692), .ZN(n5695) );
  INV_X1 U7214 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7215 ( .A1(n5695), .A2(n5694), .ZN(n6198) );
  NAND2_X1 U7216 ( .A1(n5644), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5701) );
  OAI21_X1 U7217 ( .B1(n5707), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5696), .ZN(
        n7232) );
  INV_X1 U7218 ( .A(n7232), .ZN(n7156) );
  NAND2_X1 U7219 ( .A1(n6067), .A2(n7156), .ZN(n5700) );
  INV_X1 U7220 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5697) );
  INV_X1 U7221 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6449) );
  OR2_X1 U7222 ( .A1(n5618), .A2(n5557), .ZN(n5703) );
  XNOR2_X1 U7223 ( .A(n5703), .B(n5702), .ZN(n6450) );
  OR2_X1 U7224 ( .A1(n8006), .A2(n6230), .ZN(n5705) );
  OAI22_X1 U7225 ( .A1(n7184), .A2(n6058), .B1(n9823), .B2(n6055), .ZN(n5706)
         );
  XNOR2_X1 U7226 ( .A(n5706), .B(n6024), .ZN(n7227) );
  INV_X1 U7227 ( .A(n7184), .ZN(n9207) );
  AOI22_X1 U7228 ( .A1(n9207), .A2(n6101), .B1(n6105), .B2(n7157), .ZN(n5722)
         );
  NOR2_X1 U7229 ( .A1(n7227), .A2(n5722), .ZN(n5721) );
  NAND2_X1 U7230 ( .A1(n5644), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5715) );
  AOI21_X1 U7231 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5708) );
  NOR2_X1 U7232 ( .A1(n5708), .A2(n5707), .ZN(n7125) );
  NAND2_X1 U7233 ( .A1(n6067), .A2(n7125), .ZN(n5714) );
  INV_X1 U7234 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5710) );
  OR2_X1 U7235 ( .A1(n5709), .A2(n5710), .ZN(n5713) );
  INV_X1 U7236 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5711) );
  OR2_X1 U7237 ( .A1(n4314), .A2(n5711), .ZN(n5712) );
  NAND2_X1 U7238 ( .A1(n5686), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5716) );
  XNOR2_X1 U7239 ( .A(n5716), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6446) );
  INV_X1 U7240 ( .A(n6446), .ZN(n6315) );
  OR2_X1 U7241 ( .A1(n5717), .A2(n6228), .ZN(n5719) );
  INV_X1 U7242 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6229) );
  OR2_X1 U7243 ( .A1(n8006), .A2(n6229), .ZN(n5718) );
  OAI211_X1 U7244 ( .C1(n8002), .C2(n6315), .A(n5719), .B(n5718), .ZN(n7132)
         );
  OAI22_X1 U7245 ( .A1(n7236), .A2(n6058), .B1(n9818), .B2(n6055), .ZN(n5720)
         );
  XNOR2_X1 U7246 ( .A(n5720), .B(n6744), .ZN(n7226) );
  OAI22_X1 U7247 ( .A1(n7236), .A2(n6057), .B1(n9818), .B2(n6058), .ZN(n7126)
         );
  INV_X1 U7248 ( .A(n5722), .ZN(n7228) );
  OAI21_X1 U7249 ( .B1(n7226), .B2(n7126), .A(n7228), .ZN(n5723) );
  NAND2_X1 U7250 ( .A1(n5723), .A2(n7227), .ZN(n5724) );
  OAI21_X1 U7251 ( .B1(n5729), .B2(n5728), .A(n5727), .ZN(n7295) );
  NAND2_X1 U7252 ( .A1(n5644), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5735) );
  OR2_X1 U7253 ( .A1(n5730), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5731) );
  AND2_X1 U7254 ( .A1(n5752), .A2(n5731), .ZN(n7256) );
  NAND2_X1 U7255 ( .A1(n6067), .A2(n7256), .ZN(n5734) );
  OR2_X1 U7256 ( .A1(n5709), .A2(n9840), .ZN(n5733) );
  INV_X1 U7257 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7257) );
  OR2_X1 U7258 ( .A1(n4314), .A2(n7257), .ZN(n5732) );
  NAND2_X1 U7259 ( .A1(n6238), .A2(n8005), .ZN(n5742) );
  INV_X1 U7260 ( .A(n5766), .ZN(n5740) );
  NAND2_X1 U7261 ( .A1(n5737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5738) );
  MUX2_X1 U7262 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5738), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5739) );
  AOI22_X1 U7263 ( .A1(n5928), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5927), .B2(
        n9756), .ZN(n5741) );
  NAND2_X1 U7264 ( .A1(n5742), .A2(n5741), .ZN(n7275) );
  NAND2_X1 U7265 ( .A1(n7275), .A2(n6106), .ZN(n5743) );
  OAI21_X1 U7266 ( .B1(n7251), .B2(n6058), .A(n5743), .ZN(n5744) );
  XNOR2_X1 U7267 ( .A(n5744), .B(n6024), .ZN(n7293) );
  AND2_X1 U7268 ( .A1(n7275), .A2(n6105), .ZN(n5745) );
  AOI21_X1 U7269 ( .B1(n9205), .B2(n6101), .A(n5745), .ZN(n7292) );
  NAND2_X1 U7270 ( .A1(n7293), .A2(n7292), .ZN(n5747) );
  NOR2_X1 U7271 ( .A1(n7293), .A2(n7292), .ZN(n5746) );
  NAND2_X1 U7272 ( .A1(n6249), .A2(n8005), .ZN(n5750) );
  OR2_X1 U7273 ( .A1(n5766), .A2(n5557), .ZN(n5748) );
  XNOR2_X1 U7274 ( .A(n5748), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U7275 ( .A1(n5928), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5927), .B2(
        n9769), .ZN(n5749) );
  NAND2_X1 U7276 ( .A1(n5750), .A2(n5749), .ZN(n7337) );
  NAND2_X1 U7277 ( .A1(n7337), .A2(n6106), .ZN(n5760) );
  NAND2_X1 U7278 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  AND2_X1 U7279 ( .A1(n5770), .A2(n5753), .ZN(n7380) );
  NAND2_X1 U7280 ( .A1(n6067), .A2(n7380), .ZN(n5758) );
  INV_X1 U7281 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7282 ( .A1(n5709), .A2(n5754), .ZN(n5757) );
  NAND2_X1 U7283 ( .A1(n4313), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7284 ( .A1(n5644), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5755) );
  NAND4_X1 U7285 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n9204)
         );
  NAND2_X1 U7286 ( .A1(n9204), .A2(n6105), .ZN(n5759) );
  NAND2_X1 U7287 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  XNOR2_X1 U7288 ( .A(n5761), .B(n6024), .ZN(n5763) );
  AOI22_X1 U7289 ( .A1(n7337), .A2(n6105), .B1(n6101), .B2(n9204), .ZN(n5762)
         );
  NAND2_X1 U7290 ( .A1(n5763), .A2(n5762), .ZN(n7383) );
  OAI21_X1 U7291 ( .B1(n5763), .B2(n5762), .A(n7383), .ZN(n5764) );
  INV_X1 U7292 ( .A(n5764), .ZN(n7375) );
  NAND2_X1 U7293 ( .A1(n6269), .A2(n8005), .ZN(n5769) );
  INV_X1 U7294 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7295 ( .A1(n5766), .A2(n5765), .ZN(n5783) );
  NAND2_X1 U7296 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U7297 ( .A(n5767), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U7298 ( .A1(n5928), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5927), .B2(
        n6679), .ZN(n5768) );
  NAND2_X2 U7299 ( .A1(n5769), .A2(n5768), .ZN(n9616) );
  NAND2_X1 U7300 ( .A1(n9616), .A2(n6106), .ZN(n5779) );
  NAND2_X1 U7301 ( .A1(n5644), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7302 ( .A1(n5770), .A2(n6443), .ZN(n5771) );
  AND2_X1 U7303 ( .A1(n5789), .A2(n5771), .ZN(n7389) );
  NAND2_X1 U7304 ( .A1(n6067), .A2(n7389), .ZN(n5776) );
  INV_X1 U7305 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5772) );
  OR2_X1 U7306 ( .A1(n5709), .A2(n5772), .ZN(n5775) );
  INV_X1 U7307 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5773) );
  OR2_X1 U7308 ( .A1(n4315), .A2(n5773), .ZN(n5774) );
  NAND2_X1 U7309 ( .A1(n9203), .A2(n6105), .ZN(n5778) );
  NAND2_X1 U7310 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  XNOR2_X1 U7311 ( .A(n5780), .B(n6744), .ZN(n5801) );
  NAND2_X1 U7312 ( .A1(n9616), .A2(n6105), .ZN(n5782) );
  NAND2_X1 U7313 ( .A1(n9203), .A2(n6101), .ZN(n5781) );
  NAND2_X1 U7314 ( .A1(n5782), .A2(n5781), .ZN(n5802) );
  NAND2_X1 U7315 ( .A1(n5801), .A2(n5802), .ZN(n7386) );
  AND2_X1 U7316 ( .A1(n7375), .A2(n7386), .ZN(n7399) );
  NAND2_X1 U7317 ( .A1(n6257), .A2(n8005), .ZN(n5786) );
  OAI21_X1 U7318 ( .B1(n5783), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U7319 ( .A(n5784), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U7320 ( .A1(n5928), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5927), .B2(
        n9777), .ZN(n5785) );
  NAND2_X1 U7321 ( .A1(n9582), .A2(n6106), .ZN(n5796) );
  NAND2_X1 U7322 ( .A1(n5644), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5794) );
  INV_X1 U7323 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5787) );
  OR2_X1 U7324 ( .A1(n4315), .A2(n5787), .ZN(n5793) );
  NAND2_X1 U7325 ( .A1(n7738), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5792) );
  AND2_X1 U7326 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  NOR2_X1 U7327 ( .A1(n5816), .A2(n5790), .ZN(n7410) );
  NAND2_X1 U7328 ( .A1(n6067), .A2(n7410), .ZN(n5791) );
  NAND4_X1 U7329 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n9202)
         );
  NAND2_X1 U7330 ( .A1(n9202), .A2(n6105), .ZN(n5795) );
  NAND2_X1 U7331 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  XNOR2_X1 U7332 ( .A(n5797), .B(n6744), .ZN(n5807) );
  AND2_X1 U7333 ( .A1(n9202), .A2(n6101), .ZN(n5798) );
  AOI21_X1 U7334 ( .B1(n9582), .B2(n6105), .A(n5798), .ZN(n5808) );
  INV_X1 U7335 ( .A(n5808), .ZN(n5799) );
  NAND2_X1 U7336 ( .A1(n5807), .A2(n5799), .ZN(n5800) );
  AND2_X1 U7337 ( .A1(n7399), .A2(n5800), .ZN(n5811) );
  INV_X1 U7338 ( .A(n5800), .ZN(n5810) );
  INV_X1 U7339 ( .A(n7386), .ZN(n5806) );
  INV_X1 U7340 ( .A(n5801), .ZN(n5804) );
  INV_X1 U7341 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7342 ( .A1(n5804), .A2(n5803), .ZN(n7385) );
  AND2_X1 U7343 ( .A1(n7383), .A2(n7385), .ZN(n5805) );
  OR2_X1 U7344 ( .A1(n5806), .A2(n5805), .ZN(n7401) );
  XOR2_X1 U7345 ( .A(n5808), .B(n5807), .Z(n7402) );
  INV_X1 U7346 ( .A(n7402), .ZN(n5809) );
  AND2_X1 U7347 ( .A1(n7401), .A2(n5809), .ZN(n7404) );
  NAND2_X1 U7348 ( .A1(n6300), .A2(n8005), .ZN(n5815) );
  OR2_X1 U7349 ( .A1(n5812), .A2(n5557), .ZN(n5813) );
  XNOR2_X1 U7350 ( .A(n5813), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7351 ( .A1(n5928), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5927), .B2(
        n6774), .ZN(n5814) );
  NAND2_X1 U7352 ( .A1(n9574), .A2(n6106), .ZN(n5825) );
  NAND2_X1 U7353 ( .A1(n5644), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7354 ( .A1(n5816), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5817) );
  AND2_X1 U7355 ( .A1(n5817), .A2(n5836), .ZN(n7484) );
  NAND2_X1 U7356 ( .A1(n6067), .A2(n7484), .ZN(n5822) );
  INV_X1 U7357 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5818) );
  OR2_X1 U7358 ( .A1(n5709), .A2(n5818), .ZN(n5821) );
  INV_X1 U7359 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5819) );
  OR2_X1 U7360 ( .A1(n4314), .A2(n5819), .ZN(n5820) );
  INV_X1 U7361 ( .A(n7570), .ZN(n9201) );
  NAND2_X1 U7362 ( .A1(n9201), .A2(n6105), .ZN(n5824) );
  NAND2_X1 U7363 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  XNOR2_X1 U7364 ( .A(n5826), .B(n6024), .ZN(n7457) );
  NOR2_X1 U7365 ( .A1(n7570), .A2(n6057), .ZN(n5827) );
  AOI21_X1 U7366 ( .B1(n9574), .B2(n6105), .A(n5827), .ZN(n5828) );
  NAND2_X1 U7367 ( .A1(n7457), .A2(n5828), .ZN(n5830) );
  INV_X1 U7368 ( .A(n7457), .ZN(n5829) );
  INV_X1 U7369 ( .A(n5828), .ZN(n7456) );
  NAND2_X1 U7370 ( .A1(n6480), .A2(n8005), .ZN(n5834) );
  NAND2_X1 U7371 ( .A1(n5831), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5832) );
  XNOR2_X1 U7372 ( .A(n5832), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7170) );
  AOI22_X1 U7373 ( .A1(n5928), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5927), .B2(
        n7170), .ZN(n5833) );
  NAND2_X1 U7374 ( .A1(n7622), .A2(n6106), .ZN(n5843) );
  NAND2_X1 U7375 ( .A1(n5644), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5841) );
  INV_X1 U7376 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6775) );
  OR2_X1 U7377 ( .A1(n4315), .A2(n6775), .ZN(n5840) );
  NAND2_X1 U7378 ( .A1(n7738), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7379 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  AND2_X1 U7380 ( .A1(n5855), .A2(n5837), .ZN(n7572) );
  NAND2_X1 U7381 ( .A1(n6067), .A2(n7572), .ZN(n5838) );
  NAND4_X1 U7382 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n9200)
         );
  NAND2_X1 U7383 ( .A1(n9200), .A2(n6105), .ZN(n5842) );
  NAND2_X1 U7384 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  XNOR2_X1 U7385 ( .A(n5844), .B(n6744), .ZN(n5847) );
  NAND2_X1 U7386 ( .A1(n7622), .A2(n6105), .ZN(n5846) );
  NAND2_X1 U7387 ( .A1(n9200), .A2(n6101), .ZN(n5845) );
  NAND2_X1 U7388 ( .A1(n5846), .A2(n5845), .ZN(n5848) );
  NAND2_X1 U7389 ( .A1(n5847), .A2(n5848), .ZN(n7563) );
  INV_X1 U7390 ( .A(n5847), .ZN(n5850) );
  INV_X1 U7391 ( .A(n5848), .ZN(n5849) );
  NAND2_X1 U7392 ( .A1(n5850), .A2(n5849), .ZN(n7564) );
  NAND2_X1 U7393 ( .A1(n6526), .A2(n8005), .ZN(n5854) );
  NAND2_X1 U7394 ( .A1(n5851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7395 ( .A(n5852), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9219) );
  AOI22_X1 U7396 ( .A1(n5928), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5927), .B2(
        n9219), .ZN(n5853) );
  NAND2_X1 U7397 ( .A1(n7738), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7398 ( .A1(n5644), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5859) );
  AND2_X1 U7399 ( .A1(n5855), .A2(n7167), .ZN(n5856) );
  NOR2_X1 U7400 ( .A1(n5871), .A2(n5856), .ZN(n7650) );
  NAND2_X1 U7401 ( .A1(n6067), .A2(n7650), .ZN(n5858) );
  NAND2_X1 U7402 ( .A1(n4313), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5857) );
  NAND4_X1 U7403 ( .A1(n5860), .A2(n5859), .A3(n5858), .A4(n5857), .ZN(n9199)
         );
  AOI22_X1 U7404 ( .A1(n9570), .A2(n6106), .B1(n6105), .B2(n9199), .ZN(n5861)
         );
  XNOR2_X1 U7405 ( .A(n5861), .B(n6744), .ZN(n5862) );
  INV_X1 U7406 ( .A(n9570), .ZN(n7652) );
  INV_X1 U7407 ( .A(n9199), .ZN(n9186) );
  OAI22_X1 U7408 ( .A1(n7652), .A2(n6058), .B1(n9186), .B2(n6057), .ZN(n7640)
         );
  NAND2_X1 U7409 ( .A1(n7637), .A2(n7640), .ZN(n5864) );
  INV_X1 U7410 ( .A(n5862), .ZN(n5863) );
  NAND2_X1 U7411 ( .A1(n5864), .A2(n7638), .ZN(n5882) );
  NAND2_X1 U7412 ( .A1(n6612), .A2(n8005), .ZN(n5870) );
  AND2_X1 U7413 ( .A1(n5560), .A2(n5865), .ZN(n5866) );
  OR2_X1 U7414 ( .A1(n5866), .A2(n5557), .ZN(n5868) );
  XNOR2_X1 U7415 ( .A(n5868), .B(n5867), .ZN(n9234) );
  INV_X1 U7416 ( .A(n9234), .ZN(n9223) );
  AOI22_X1 U7417 ( .A1(n5928), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5927), .B2(
        n9223), .ZN(n5869) );
  NAND2_X1 U7418 ( .A1(n5644), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5879) );
  NOR2_X1 U7419 ( .A1(n5871), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7420 ( .A1(n5873), .A2(n5872), .ZN(n9190) );
  INV_X1 U7421 ( .A(n9190), .ZN(n5874) );
  NAND2_X1 U7422 ( .A1(n6067), .A2(n5874), .ZN(n5878) );
  INV_X1 U7423 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5875) );
  OR2_X1 U7424 ( .A1(n5709), .A2(n5875), .ZN(n5877) );
  INV_X1 U7425 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7670) );
  OR2_X1 U7426 ( .A1(n4314), .A2(n7670), .ZN(n5876) );
  INV_X1 U7427 ( .A(n9631), .ZN(n9198) );
  AOI22_X1 U7428 ( .A1(n9193), .A2(n6106), .B1(n6105), .B2(n9198), .ZN(n5880)
         );
  XOR2_X1 U7429 ( .A(n6744), .B(n5880), .Z(n5881) );
  INV_X1 U7430 ( .A(n9193), .ZN(n9663) );
  OAI22_X1 U7431 ( .A1(n9663), .A2(n6058), .B1(n9631), .B2(n6057), .ZN(n9185)
         );
  INV_X1 U7432 ( .A(n5883), .ZN(n5886) );
  INV_X1 U7433 ( .A(n5884), .ZN(n5885) );
  NAND2_X1 U7434 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7435 ( .A1(n6666), .A2(n8005), .ZN(n5892) );
  NAND2_X1 U7436 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U7437 ( .A1(n5890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7438 ( .A(n5909), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9266) );
  AOI22_X1 U7439 ( .A1(n5928), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5927), .B2(
        n9266), .ZN(n5891) );
  NAND2_X1 U7440 ( .A1(n5644), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7441 ( .A1(n7738), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5898) );
  INV_X1 U7442 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7443 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  AND2_X1 U7444 ( .A1(n5916), .A2(n5895), .ZN(n9475) );
  NAND2_X1 U7445 ( .A1(n6067), .A2(n9475), .ZN(n5897) );
  NAND2_X1 U7446 ( .A1(n4313), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5896) );
  NAND4_X1 U7447 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n9446)
         );
  OAI22_X1 U7448 ( .A1(n9478), .A2(n6058), .B1(n9635), .B2(n6057), .ZN(n5904)
         );
  NAND2_X1 U7449 ( .A1(n9565), .A2(n6106), .ZN(n5901) );
  NAND2_X1 U7450 ( .A1(n9446), .A2(n6105), .ZN(n5900) );
  NAND2_X1 U7451 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  XNOR2_X1 U7452 ( .A(n5902), .B(n6744), .ZN(n5903) );
  XOR2_X1 U7453 ( .A(n5904), .B(n5903), .Z(n9116) );
  NAND2_X1 U7454 ( .A1(n9114), .A2(n9116), .ZN(n9115) );
  INV_X1 U7455 ( .A(n5903), .ZN(n5906) );
  INV_X1 U7456 ( .A(n5904), .ZN(n5905) );
  NAND2_X1 U7457 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7458 ( .A1(n6713), .A2(n8005), .ZN(n5913) );
  NAND2_X1 U7459 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  NAND2_X1 U7460 ( .A1(n5910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U7461 ( .A(n5911), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9276) );
  AOI22_X1 U7462 ( .A1(n5928), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5927), .B2(
        n9276), .ZN(n5912) );
  INV_X1 U7463 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7464 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  AND2_X1 U7465 ( .A1(n5932), .A2(n5917), .ZN(n9459) );
  NAND2_X1 U7466 ( .A1(n6067), .A2(n9459), .ZN(n5923) );
  NAND2_X1 U7467 ( .A1(n5644), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5922) );
  INV_X1 U7468 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7469 ( .A1(n5709), .A2(n5918), .ZN(n5921) );
  INV_X1 U7470 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5919) );
  OR2_X1 U7471 ( .A1(n4314), .A2(n5919), .ZN(n5920) );
  AOI22_X1 U7472 ( .A1(n9560), .A2(n6106), .B1(n6105), .B2(n9486), .ZN(n5924)
         );
  XNOR2_X1 U7473 ( .A(n5924), .B(n6744), .ZN(n9157) );
  AOI22_X1 U7474 ( .A1(n9560), .A2(n6105), .B1(n6101), .B2(n9486), .ZN(n9156)
         );
  OAI21_X1 U7475 ( .B1(n9159), .B2(n9157), .A(n9156), .ZN(n5926) );
  NAND2_X1 U7476 ( .A1(n9159), .A2(n9157), .ZN(n5925) );
  NAND2_X1 U7477 ( .A1(n6799), .A2(n8005), .ZN(n5930) );
  AOI22_X1 U7478 ( .A1(n5928), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8296), .B2(
        n5927), .ZN(n5929) );
  NAND2_X1 U7479 ( .A1(n9552), .A2(n6106), .ZN(n5941) );
  NAND2_X1 U7480 ( .A1(n5644), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5939) );
  INV_X1 U7481 ( .A(n5932), .ZN(n5931) );
  NAND2_X1 U7482 ( .A1(n5931), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5952) );
  INV_X1 U7483 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U7484 ( .A1(n5932), .A2(n7913), .ZN(n5933) );
  AND2_X1 U7485 ( .A1(n5952), .A2(n5933), .ZN(n9433) );
  NAND2_X1 U7486 ( .A1(n6067), .A2(n9433), .ZN(n5938) );
  INV_X1 U7487 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5934) );
  OR2_X1 U7488 ( .A1(n5709), .A2(n5934), .ZN(n5937) );
  INV_X1 U7489 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7490 ( .A1(n4314), .A2(n5935), .ZN(n5936) );
  NAND2_X1 U7491 ( .A1(n9447), .A2(n6105), .ZN(n5940) );
  NAND2_X1 U7492 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  XNOR2_X1 U7493 ( .A(n5942), .B(n6024), .ZN(n9086) );
  NOR2_X1 U7494 ( .A1(n9162), .A2(n6057), .ZN(n5943) );
  AOI21_X1 U7495 ( .B1(n9552), .B2(n6105), .A(n5943), .ZN(n5945) );
  NAND2_X1 U7496 ( .A1(n9086), .A2(n5945), .ZN(n5944) );
  INV_X1 U7497 ( .A(n9086), .ZN(n5946) );
  INV_X1 U7498 ( .A(n5945), .ZN(n9085) );
  NAND2_X1 U7499 ( .A1(n5946), .A2(n9085), .ZN(n5947) );
  NAND2_X1 U7500 ( .A1(n6926), .A2(n8005), .ZN(n5949) );
  OR2_X1 U7501 ( .A1(n8006), .A2(n6927), .ZN(n5948) );
  NAND2_X1 U7502 ( .A1(n9548), .A2(n6106), .ZN(n5958) );
  INV_X1 U7503 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7504 ( .A1(n7738), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5950) );
  OAI21_X1 U7505 ( .B1(n5951), .B2(n7742), .A(n5950), .ZN(n5956) );
  INV_X1 U7506 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U7507 ( .A1(n5952), .A2(n9135), .ZN(n5953) );
  NAND2_X1 U7508 ( .A1(n5973), .A2(n5953), .ZN(n9416) );
  NAND2_X1 U7509 ( .A1(n4313), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U7510 ( .B1(n9416), .B2(n6147), .A(n5954), .ZN(n5955) );
  NAND2_X1 U7511 ( .A1(n9437), .A2(n6105), .ZN(n5957) );
  NAND2_X1 U7512 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7513 ( .A(n5959), .B(n6024), .ZN(n5961) );
  AOI22_X1 U7514 ( .A1(n9548), .A2(n6105), .B1(n6101), .B2(n9437), .ZN(n5960)
         );
  NAND2_X1 U7515 ( .A1(n5961), .A2(n5960), .ZN(n9095) );
  OAI21_X1 U7516 ( .B1(n5961), .B2(n5960), .A(n9095), .ZN(n9134) );
  NAND2_X1 U7517 ( .A1(n7241), .A2(n8005), .ZN(n5963) );
  OR2_X1 U7518 ( .A1(n8006), .A2(n7242), .ZN(n5962) );
  INV_X1 U7519 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7520 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5964) );
  INV_X1 U7521 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5966) );
  INV_X1 U7522 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U7523 ( .B1(n5973), .B2(n5966), .A(n5965), .ZN(n5967) );
  AND2_X1 U7524 ( .A1(n5999), .A2(n5967), .ZN(n9387) );
  NAND2_X1 U7525 ( .A1(n9387), .A2(n6067), .ZN(n5969) );
  AOI22_X1 U7526 ( .A1(n5644), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n7738), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5968) );
  OAI211_X1 U7527 ( .C1(n4315), .C2(n5970), .A(n5969), .B(n5968), .ZN(n9409)
         );
  AOI22_X1 U7528 ( .A1(n9537), .A2(n6105), .B1(n6101), .B2(n9409), .ZN(n5993)
         );
  NAND2_X1 U7529 ( .A1(n7037), .A2(n8005), .ZN(n5972) );
  INV_X1 U7530 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7145) );
  OR2_X1 U7531 ( .A1(n8006), .A2(n7145), .ZN(n5971) );
  NAND2_X1 U7532 ( .A1(n9543), .A2(n6106), .ZN(n5980) );
  INV_X1 U7533 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7534 ( .A(n5973), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U7535 ( .A1(n9403), .A2(n6067), .ZN(n5977) );
  NAND2_X1 U7536 ( .A1(n7738), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7537 ( .A1(n4313), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5974) );
  AND2_X1 U7538 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  OAI211_X1 U7539 ( .C1(n7742), .C2(n5978), .A(n5977), .B(n5976), .ZN(n9422)
         );
  NAND2_X1 U7540 ( .A1(n9422), .A2(n6105), .ZN(n5979) );
  NAND2_X1 U7541 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  XNOR2_X1 U7542 ( .A(n5981), .B(n6744), .ZN(n5985) );
  INV_X1 U7543 ( .A(n5985), .ZN(n5983) );
  INV_X1 U7544 ( .A(n9422), .ZN(n9136) );
  OAI22_X1 U7545 ( .A1(n9405), .A2(n6058), .B1(n9136), .B2(n6057), .ZN(n5986)
         );
  INV_X1 U7546 ( .A(n5986), .ZN(n5982) );
  NAND2_X1 U7547 ( .A1(n5983), .A2(n5982), .ZN(n5989) );
  INV_X1 U7548 ( .A(n5989), .ZN(n5991) );
  NOR2_X1 U7549 ( .A1(n5993), .A2(n5991), .ZN(n5984) );
  AND2_X1 U7550 ( .A1(n9095), .A2(n5984), .ZN(n5988) );
  INV_X1 U7551 ( .A(n5984), .ZN(n5987) );
  XOR2_X1 U7552 ( .A(n5986), .B(n5985), .Z(n9098) );
  AOI21_X2 U7553 ( .B1(n9143), .B2(n5988), .A(n4336), .ZN(n9147) );
  AND2_X1 U7554 ( .A1(n9095), .A2(n5989), .ZN(n9142) );
  AOI22_X1 U7555 ( .A1(n9537), .A2(n6106), .B1(n6105), .B2(n9409), .ZN(n5990)
         );
  XOR2_X1 U7556 ( .A(n6744), .B(n5990), .Z(n9149) );
  AND2_X1 U7557 ( .A1(n9142), .A2(n9149), .ZN(n5995) );
  INV_X1 U7558 ( .A(n9149), .ZN(n5994) );
  OR2_X1 U7559 ( .A1(n5991), .A2(n9098), .ZN(n5992) );
  AND2_X1 U7560 ( .A1(n5993), .A2(n5992), .ZN(n9144) );
  AOI21_X2 U7561 ( .B1(n9143), .B2(n5995), .A(n4864), .ZN(n6007) );
  NAND2_X1 U7562 ( .A1(n7245), .A2(n8005), .ZN(n5997) );
  OR2_X1 U7563 ( .A1(n8006), .A2(n7248), .ZN(n5996) );
  NAND2_X1 U7564 ( .A1(n9532), .A2(n6106), .ZN(n6005) );
  INV_X1 U7565 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6003) );
  INV_X1 U7566 ( .A(n5999), .ZN(n5998) );
  NAND2_X1 U7567 ( .A1(n5998), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6014) );
  INV_X1 U7568 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U7569 ( .A1(n5999), .A2(n9079), .ZN(n6000) );
  NAND2_X1 U7570 ( .A1(n6014), .A2(n6000), .ZN(n9375) );
  OR2_X1 U7571 ( .A1(n9375), .A2(n6147), .ZN(n6002) );
  AOI22_X1 U7572 ( .A1(n4313), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n7738), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n6001) );
  OAI211_X1 U7573 ( .C1(n7742), .C2(n6003), .A(n6002), .B(n6001), .ZN(n9394)
         );
  NAND2_X1 U7574 ( .A1(n9394), .A2(n6105), .ZN(n6004) );
  NAND2_X1 U7575 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  XNOR2_X1 U7576 ( .A(n6006), .B(n6024), .ZN(n6008) );
  INV_X1 U7577 ( .A(n9532), .ZN(n9378) );
  INV_X1 U7578 ( .A(n9394), .ZN(n9152) );
  OAI22_X1 U7579 ( .A1(n9378), .A2(n6058), .B1(n9152), .B2(n6057), .ZN(n9078)
         );
  INV_X1 U7580 ( .A(n6008), .ZN(n6009) );
  NAND2_X1 U7581 ( .A1(n7319), .A2(n8005), .ZN(n6011) );
  OR2_X1 U7582 ( .A1(n8006), .A2(n7320), .ZN(n6010) );
  NAND2_X1 U7583 ( .A1(n9528), .A2(n6106), .ZN(n6023) );
  INV_X1 U7584 ( .A(n6014), .ZN(n6012) );
  NAND2_X1 U7585 ( .A1(n6012), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6033) );
  INV_X1 U7586 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7587 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  NAND2_X1 U7588 ( .A1(n6033), .A2(n6015), .ZN(n9359) );
  OR2_X1 U7589 ( .A1(n9359), .A2(n6147), .ZN(n6021) );
  INV_X1 U7590 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7591 ( .A1(n7738), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7592 ( .A1(n4313), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6016) );
  OAI211_X1 U7593 ( .C1(n7742), .C2(n6018), .A(n6017), .B(n6016), .ZN(n6019)
         );
  INV_X1 U7594 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7595 ( .A1(n6021), .A2(n6020), .ZN(n9380) );
  NAND2_X1 U7596 ( .A1(n9380), .A2(n6105), .ZN(n6022) );
  NAND2_X1 U7597 ( .A1(n6023), .A2(n6022), .ZN(n6025) );
  XNOR2_X1 U7598 ( .A(n6025), .B(n6024), .ZN(n6028) );
  AND2_X1 U7599 ( .A1(n9380), .A2(n6101), .ZN(n6026) );
  AOI21_X1 U7600 ( .B1(n9528), .B2(n6105), .A(n6026), .ZN(n6027) );
  NAND2_X1 U7601 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  OAI21_X1 U7602 ( .B1(n6028), .B2(n6027), .A(n6029), .ZN(n9125) );
  NAND2_X1 U7603 ( .A1(n7464), .A2(n8005), .ZN(n6031) );
  OR2_X1 U7604 ( .A1(n8006), .A2(n7469), .ZN(n6030) );
  INV_X1 U7605 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7606 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7607 ( .A1(n9346), .A2(n6067), .ZN(n6040) );
  INV_X1 U7608 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7609 ( .A1(n7738), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7610 ( .A1(n5644), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7611 ( .C1(n6037), .C2(n4315), .A(n6036), .B(n6035), .ZN(n6038)
         );
  INV_X1 U7612 ( .A(n6038), .ZN(n6039) );
  OAI22_X1 U7613 ( .A1(n9348), .A2(n6058), .B1(n9176), .B2(n6057), .ZN(n6059)
         );
  NAND2_X1 U7614 ( .A1(n9523), .A2(n6106), .ZN(n6042) );
  NAND2_X1 U7615 ( .A1(n9366), .A2(n6105), .ZN(n6041) );
  NAND2_X1 U7616 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  XNOR2_X1 U7617 ( .A(n6043), .B(n6744), .ZN(n6060) );
  XOR2_X1 U7618 ( .A(n6059), .B(n6060), .Z(n9106) );
  NAND2_X1 U7619 ( .A1(n7516), .A2(n8005), .ZN(n6045) );
  OR2_X1 U7620 ( .A1(n8006), .A2(n7517), .ZN(n6044) );
  INV_X1 U7621 ( .A(n6047), .ZN(n6046) );
  NAND2_X1 U7622 ( .A1(n6046), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6065) );
  INV_X1 U7623 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U7624 ( .A1(n6047), .A2(n9175), .ZN(n6048) );
  NAND2_X1 U7625 ( .A1(n6065), .A2(n6048), .ZN(n9331) );
  INV_X1 U7626 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7627 ( .A1(n7738), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7628 ( .A1(n4313), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6049) );
  OAI211_X1 U7629 ( .C1(n6051), .C2(n7742), .A(n6050), .B(n6049), .ZN(n6052)
         );
  INV_X1 U7630 ( .A(n6052), .ZN(n6053) );
  OAI22_X1 U7631 ( .A1(n9334), .A2(n6055), .B1(n9068), .B2(n6058), .ZN(n6056)
         );
  XNOR2_X1 U7632 ( .A(n6056), .B(n6744), .ZN(n6082) );
  OAI22_X1 U7633 ( .A1(n9334), .A2(n6058), .B1(n9068), .B2(n6057), .ZN(n6081)
         );
  XNOR2_X1 U7634 ( .A(n6082), .B(n6081), .ZN(n9169) );
  NOR2_X1 U7635 ( .A1(n6060), .A2(n6059), .ZN(n9170) );
  NOR2_X1 U7636 ( .A1(n9169), .A2(n9170), .ZN(n6061) );
  NAND2_X1 U7637 ( .A1(n7547), .A2(n8005), .ZN(n6064) );
  OR2_X1 U7638 ( .A1(n8006), .A2(n6062), .ZN(n6063) );
  NAND2_X1 U7639 ( .A1(n9513), .A2(n6106), .ZN(n6075) );
  INV_X1 U7640 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U7641 ( .A1(n6065), .A2(n9067), .ZN(n6066) );
  NAND2_X1 U7642 ( .A1(n9320), .A2(n6067), .ZN(n6073) );
  INV_X1 U7643 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7644 ( .A1(n7738), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7645 ( .A1(n4313), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6068) );
  OAI211_X1 U7646 ( .C1(n6070), .C2(n7742), .A(n6069), .B(n6068), .ZN(n6071)
         );
  INV_X1 U7647 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7648 ( .A1(n9337), .A2(n6105), .ZN(n6074) );
  NAND2_X1 U7649 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  XNOR2_X1 U7650 ( .A(n6076), .B(n6744), .ZN(n6080) );
  NAND2_X1 U7651 ( .A1(n9513), .A2(n6105), .ZN(n6078) );
  NAND2_X1 U7652 ( .A1(n9337), .A2(n6101), .ZN(n6077) );
  NAND2_X1 U7653 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NOR2_X1 U7654 ( .A1(n6080), .A2(n6079), .ZN(n6135) );
  AOI21_X1 U7655 ( .B1(n6080), .B2(n6079), .A(n6135), .ZN(n9063) );
  INV_X1 U7656 ( .A(n9063), .ZN(n6084) );
  NAND2_X1 U7657 ( .A1(n6082), .A2(n6081), .ZN(n9064) );
  INV_X1 U7658 ( .A(n9064), .ZN(n6083) );
  NOR2_X1 U7659 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  INV_X1 U7660 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7555) );
  INV_X1 U7661 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7560) );
  MUX2_X1 U7662 ( .A(n7555), .B(n7560), .S(n8377), .Z(n7721) );
  XNOR2_X1 U7663 ( .A(n7721), .B(SI_28_), .ZN(n7718) );
  NAND2_X1 U7664 ( .A1(n7557), .A2(n8005), .ZN(n6091) );
  OR2_X1 U7665 ( .A1(n8006), .A2(n7560), .ZN(n6090) );
  NAND2_X1 U7666 ( .A1(n9505), .A2(n6105), .ZN(n6103) );
  INV_X1 U7667 ( .A(n6093), .ZN(n6092) );
  NAND2_X1 U7668 ( .A1(n6092), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7750) );
  INV_X1 U7669 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7670 ( .A1(n6093), .A2(n6146), .ZN(n6094) );
  NAND2_X1 U7671 ( .A1(n7750), .A2(n6094), .ZN(n9307) );
  INV_X1 U7672 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7673 ( .A1(n7738), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7674 ( .A1(n4313), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6095) );
  OAI211_X1 U7675 ( .C1(n7742), .C2(n6097), .A(n6096), .B(n6095), .ZN(n6098)
         );
  INV_X1 U7676 ( .A(n6098), .ZN(n6099) );
  NAND2_X1 U7677 ( .A1(n4819), .A2(n6101), .ZN(n6102) );
  NAND2_X1 U7678 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  XNOR2_X1 U7679 ( .A(n6104), .B(n6744), .ZN(n6108) );
  AOI22_X1 U7680 ( .A1(n9505), .A2(n6106), .B1(n6105), .B2(n4819), .ZN(n6107)
         );
  XNOR2_X1 U7681 ( .A(n6108), .B(n6107), .ZN(n6136) );
  INV_X1 U7682 ( .A(n6136), .ZN(n6133) );
  INV_X1 U7683 ( .A(n6135), .ZN(n6132) );
  INV_X1 U7684 ( .A(n7467), .ZN(n6110) );
  NAND2_X1 U7685 ( .A1(n7321), .A2(P1_B_REG_SCAN_IN), .ZN(n6109) );
  OAI22_X1 U7686 ( .A1(n6110), .A2(n6109), .B1(P1_B_REG_SCAN_IN), .B2(n7321), 
        .ZN(n6111) );
  NOR4_X1 U7687 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6115) );
  NOR4_X1 U7688 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6114) );
  NOR4_X1 U7689 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6113) );
  NOR4_X1 U7690 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6112) );
  AND4_X1 U7691 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n6121)
         );
  NOR2_X1 U7692 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .ZN(
        n6119) );
  NOR4_X1 U7693 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6118) );
  NOR4_X1 U7694 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6117) );
  NOR4_X1 U7695 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6116) );
  AND4_X1 U7696 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n6120)
         );
  NAND2_X1 U7697 ( .A1(n6121), .A2(n6120), .ZN(n6638) );
  INV_X1 U7698 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U7699 ( .A1(n6638), .A2(n6122), .ZN(n6123) );
  NAND2_X1 U7700 ( .A1(n7518), .A2(n7321), .ZN(n9603) );
  OAI21_X1 U7701 ( .B1(n9602), .B2(n6123), .A(n9603), .ZN(n6618) );
  NAND2_X1 U7702 ( .A1(n7518), .A2(n7467), .ZN(n6124) );
  NAND2_X1 U7703 ( .A1(n6125), .A2(n6124), .ZN(n6738) );
  NOR2_X1 U7704 ( .A1(n6618), .A2(n6738), .ZN(n6142) );
  NAND2_X1 U7705 ( .A1(n6126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7706 ( .A1(n6142), .A2(n9804), .ZN(n6554) );
  NAND2_X1 U7707 ( .A1(n6129), .A2(n8292), .ZN(n6620) );
  OR2_X1 U7708 ( .A1(n6620), .A2(n9283), .ZN(n6131) );
  INV_X1 U7709 ( .A(n8061), .ZN(n6729) );
  NAND3_X1 U7710 ( .A1(n6134), .A2(n6133), .A3(n4849), .ZN(n6162) );
  NAND3_X1 U7711 ( .A1(n9065), .A2(n9173), .A3(n6136), .ZN(n6161) );
  INV_X1 U7712 ( .A(n6137), .ZN(n6758) );
  INV_X1 U7713 ( .A(n6142), .ZN(n6138) );
  NAND3_X1 U7714 ( .A1(n6758), .A2(n9804), .A3(n6138), .ZN(n6144) );
  AND2_X1 U7715 ( .A1(n8295), .A2(n9283), .ZN(n6139) );
  NAND2_X1 U7716 ( .A1(n6741), .A2(n9804), .ZN(n6616) );
  INV_X1 U7717 ( .A(n6616), .ZN(n6140) );
  AND2_X1 U7718 ( .A1(n6144), .A2(n6140), .ZN(n9646) );
  AND3_X1 U7719 ( .A1(n6741), .A2(n6209), .A3(n6210), .ZN(n6141) );
  OAI21_X1 U7720 ( .B1(n9615), .B2(n6142), .A(n6141), .ZN(n6143) );
  NAND2_X1 U7721 ( .A1(n6143), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6145) );
  OAI22_X1 U7722 ( .A1(n9307), .A2(n9650), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6146), .ZN(n6157) );
  OR2_X1 U7723 ( .A1(n7750), .A2(n6147), .ZN(n6152) );
  INV_X1 U7724 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U7725 ( .A1(n4313), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7726 ( .A1(n5644), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7727 ( .C1(n5709), .C2(n7769), .A(n6149), .B(n6148), .ZN(n6150)
         );
  INV_X1 U7728 ( .A(n6150), .ZN(n6151) );
  NAND2_X1 U7729 ( .A1(n6152), .A2(n6151), .ZN(n9301) );
  INV_X1 U7730 ( .A(n9301), .ZN(n8185) );
  INV_X1 U7731 ( .A(n6554), .ZN(n6153) );
  OR2_X1 U7732 ( .A1(n6727), .A2(n6726), .ZN(n6745) );
  INV_X1 U7733 ( .A(n6745), .ZN(n8348) );
  AND2_X1 U7734 ( .A1(n6153), .A2(n8348), .ZN(n6155) );
  NAND2_X1 U7735 ( .A1(n6155), .A2(n8347), .ZN(n9632) );
  OAI22_X1 U7736 ( .A1(n8185), .A2(n9636), .B1(n7717), .B2(n9632), .ZN(n6156)
         );
  AOI211_X1 U7737 ( .C1(n9505), .C2(n9192), .A(n6157), .B(n6156), .ZN(n6158)
         );
  INV_X1 U7738 ( .A(n6158), .ZN(n6159) );
  NAND3_X1 U7739 ( .A1(n6162), .A2(n6161), .A3(n6160), .ZN(P1_U3218) );
  NAND3_X1 U7740 ( .A1(n6165), .A2(n6164), .A3(n8612), .ZN(n6171) );
  AOI22_X1 U7741 ( .A1(n8682), .A2(n8694), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n6166) );
  OAI21_X1 U7742 ( .B1(n8822), .B2(n8685), .A(n6166), .ZN(n6167) );
  AOI21_X1 U7743 ( .B1(n8793), .B2(n8680), .A(n6167), .ZN(n6168) );
  NAND2_X1 U7744 ( .A1(n6171), .A2(n6170), .ZN(P2_U3242) );
  NAND2_X1 U7745 ( .A1(n7557), .A2(n8370), .ZN(n6173) );
  OR2_X1 U7746 ( .A1(n4317), .A2(n7555), .ZN(n6172) );
  NOR2_X1 U7747 ( .A1(n8776), .A2(n6174), .ZN(n6176) );
  XNOR2_X1 U7748 ( .A(n6176), .B(n6175), .ZN(n6177) );
  XNOR2_X1 U7749 ( .A(n8949), .B(n6177), .ZN(n6190) );
  INV_X1 U7750 ( .A(n6190), .ZN(n6178) );
  NAND2_X1 U7751 ( .A1(n6178), .A2(n8612), .ZN(n6195) );
  INV_X1 U7752 ( .A(n6179), .ZN(n6189) );
  NAND2_X1 U7753 ( .A1(n6196), .A2(n4860), .ZN(n6194) );
  AOI22_X1 U7754 ( .A1(n8623), .A2(n8694), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6188) );
  OR2_X1 U7755 ( .A1(n8040), .A2(n6180), .ZN(n6186) );
  INV_X1 U7756 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7757 ( .A1(n4964), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7758 ( .A1(n4995), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6181) );
  OAI211_X1 U7759 ( .C1(n6183), .C2(n5358), .A(n6182), .B(n6181), .ZN(n6184)
         );
  INV_X1 U7760 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7761 ( .A1(n8682), .A2(n8692), .ZN(n6187) );
  OAI211_X1 U7762 ( .C1(n8633), .C2(n8359), .A(n6188), .B(n6187), .ZN(n6192)
         );
  NOR3_X1 U7763 ( .A1(n6190), .A2(n6189), .A3(n8690), .ZN(n6191) );
  AOI211_X1 U7764 ( .C1(n8688), .C2(n8949), .A(n6192), .B(n6191), .ZN(n6193)
         );
  OAI211_X1 U7765 ( .C1(n6196), .C2(n6195), .A(n6194), .B(n6193), .ZN(P2_U3222) );
  INV_X1 U7766 ( .A(n6210), .ZN(n7246) );
  NOR2_X4 U7767 ( .A1(n6350), .A2(n9888), .ZN(P2_U3966) );
  NAND2_X1 U7768 ( .A1(n4597), .A2(n6198), .ZN(n6199) );
  XNOR2_X1 U7769 ( .A(n6200), .B(n6199), .ZN(n6201) );
  NOR2_X1 U7770 ( .A1(n6201), .A2(n9642), .ZN(n6208) );
  INV_X1 U7771 ( .A(n6202), .ZN(n6940) );
  NOR2_X1 U7772 ( .A1(n9650), .A2(n6940), .ZN(n6207) );
  AND2_X1 U7773 ( .A1(n9192), .A2(n6993), .ZN(n6206) );
  OR2_X1 U7774 ( .A1(n9632), .A2(n6930), .ZN(n6204) );
  AND2_X1 U7775 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9721) );
  INV_X1 U7776 ( .A(n9721), .ZN(n6203) );
  OAI211_X1 U7777 ( .C1(n9636), .C2(n7236), .A(n6204), .B(n6203), .ZN(n6205)
         );
  OR4_X1 U7778 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(P1_U3228)
         );
  NAND2_X1 U7779 ( .A1(n8061), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7780 ( .A1(n6211), .A2(n6210), .ZN(n6313) );
  NAND2_X1 U7781 ( .A1(n6313), .A2(n8002), .ZN(n6212) );
  NAND2_X1 U7782 ( .A1(n6212), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7783 ( .A(n7556), .ZN(n9613) );
  OAI222_X1 U7784 ( .A1(n9609), .A2(n6214), .B1(n9613), .B2(n6220), .C1(
        P1_U3084), .C2(n6213), .ZN(P1_U3351) );
  OAI222_X1 U7785 ( .A1(n9609), .A2(n6216), .B1(n6215), .B2(P1_U3084), .C1(
        n9613), .C2(n6218), .ZN(P1_U3352) );
  OAI222_X1 U7786 ( .A1(n9609), .A2(n6217), .B1(n9613), .B2(n6222), .C1(
        P1_U3084), .C2(n6335), .ZN(P1_U3350) );
  NOR2_X1 U7787 ( .A1(n8001), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9051) );
  INV_X1 U7788 ( .A(n9051), .ZN(n9060) );
  AND2_X1 U7789 ( .A1(n8001), .A2(P2_U3152), .ZN(n7552) );
  INV_X2 U7790 ( .A(n7552), .ZN(n9058) );
  OAI222_X1 U7791 ( .A1(n9060), .A2(n6219), .B1(n9058), .B2(n6218), .C1(n6394), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U7792 ( .A1(n9060), .A2(n6221), .B1(n9058), .B2(n6220), .C1(
        P2_U3152), .C2(n6371), .ZN(P2_U3356) );
  OAI222_X1 U7793 ( .A1(n9060), .A2(n6223), .B1(n9058), .B2(n6222), .C1(
        P2_U3152), .C2(n6471), .ZN(P2_U3355) );
  OAI222_X1 U7794 ( .A1(n9060), .A2(n6224), .B1(n9058), .B2(n6225), .C1(
        P2_U3152), .C2(n6428), .ZN(P2_U3354) );
  OAI222_X1 U7795 ( .A1(n9609), .A2(n6226), .B1(n9613), .B2(n6225), .C1(
        P1_U3084), .C2(n6316), .ZN(P1_U3349) );
  AOI22_X1 U7796 ( .A1(n6489), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9051), .ZN(n6227) );
  OAI21_X1 U7797 ( .B1(n6228), .B2(n9058), .A(n6227), .ZN(P2_U3353) );
  OAI222_X1 U7798 ( .A1(n9609), .A2(n6229), .B1(n9613), .B2(n6228), .C1(
        P1_U3084), .C2(n6315), .ZN(P1_U3348) );
  INV_X1 U7799 ( .A(n6377), .ZN(n6405) );
  INV_X1 U7800 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6234) );
  INV_X1 U7801 ( .A(n6233), .ZN(n6235) );
  INV_X1 U7802 ( .A(n6365), .ZN(n6416) );
  OAI222_X1 U7803 ( .A1(n9060), .A2(n6234), .B1(n9058), .B2(n6235), .C1(
        P2_U3152), .C2(n6416), .ZN(P2_U3351) );
  OAI222_X1 U7804 ( .A1(n9609), .A2(n6236), .B1(n9613), .B2(n6235), .C1(
        P1_U3084), .C2(n6445), .ZN(P1_U3346) );
  NAND2_X1 U7805 ( .A1(n6281), .A2(P2_U3966), .ZN(n6237) );
  OAI21_X1 U7806 ( .B1(P2_U3966), .B2(n4878), .A(n6237), .ZN(P2_U3552) );
  INV_X1 U7807 ( .A(n6238), .ZN(n6240) );
  INV_X1 U7808 ( .A(n9756), .ZN(n6239) );
  OAI222_X1 U7809 ( .A1(n9609), .A2(n7868), .B1(n9613), .B2(n6240), .C1(
        P1_U3084), .C2(n6239), .ZN(P1_U3345) );
  INV_X1 U7810 ( .A(n6511), .ZN(n6520) );
  OAI222_X1 U7811 ( .A1(n9060), .A2(n6241), .B1(n9058), .B2(n6240), .C1(
        P2_U3152), .C2(n6520), .ZN(P2_U3350) );
  INV_X1 U7812 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7813 ( .A1(n6243), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8590) );
  INV_X1 U7814 ( .A(n8590), .ZN(n6245) );
  OAI21_X1 U7815 ( .B1(n9879), .B2(n6245), .A(n6244), .ZN(n6248) );
  NAND2_X1 U7816 ( .A1(n9879), .A2(n6246), .ZN(n6247) );
  INV_X1 U7817 ( .A(n8745), .ZN(n9873) );
  NOR2_X1 U7818 ( .A1(n9873), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7819 ( .A(n6249), .ZN(n6255) );
  INV_X1 U7820 ( .A(n9769), .ZN(n6439) );
  OAI222_X1 U7821 ( .A1(n9613), .A2(n6255), .B1(n6439), .B2(P1_U3084), .C1(
        n6250), .C2(n9609), .ZN(P1_U3344) );
  NAND2_X1 U7822 ( .A1(n4955), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7823 ( .A1(n4995), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7824 ( .A1(n4964), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6251) );
  AND3_X1 U7825 ( .A1(n6253), .A2(n6252), .A3(n6251), .ZN(n8378) );
  NAND2_X1 U7826 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8712), .ZN(n6254) );
  OAI21_X1 U7827 ( .B1(n8378), .B2(n8712), .A(n6254), .ZN(P2_U3582) );
  INV_X1 U7828 ( .A(n6626), .ZN(n6525) );
  OAI222_X1 U7829 ( .A1(n9060), .A2(n6256), .B1(n9058), .B2(n6255), .C1(n6525), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7830 ( .A(n6257), .ZN(n6272) );
  AOI22_X1 U7831 ( .A1(n7047), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9051), .ZN(n6258) );
  OAI21_X1 U7832 ( .B1(n6272), .B2(n9058), .A(n6258), .ZN(P2_U3347) );
  INV_X1 U7833 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6268) );
  OR2_X1 U7834 ( .A1(n6154), .A2(P1_U3084), .ZN(n7558) );
  INV_X1 U7835 ( .A(n6311), .ZN(n9703) );
  NOR2_X1 U7836 ( .A1(n7558), .A2(n9703), .ZN(n6260) );
  INV_X1 U7837 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6261) );
  NAND3_X1 U7838 ( .A1(n9786), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6261), .ZN(
        n6267) );
  NOR2_X1 U7839 ( .A1(n6311), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6262) );
  OR2_X1 U7840 ( .A1(n6154), .A2(n6262), .ZN(n9707) );
  AOI21_X1 U7841 ( .B1(n6261), .B2(n6311), .A(n9707), .ZN(n6263) );
  INV_X1 U7842 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9705) );
  MUX2_X1 U7843 ( .A(n9707), .B(n6263), .S(n9705), .Z(n6265) );
  INV_X1 U7844 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U7845 ( .A1(P1_U3084), .A2(n6561), .ZN(n6264) );
  OAI211_X1 U7846 ( .C1(P1_U3084), .C2(n6265), .A(P1_U3083), .B(n6264), .ZN(
        n6266) );
  OAI211_X1 U7847 ( .C1(n9792), .C2(n6268), .A(n6267), .B(n6266), .ZN(P1_U3241) );
  INV_X1 U7848 ( .A(n6269), .ZN(n6273) );
  INV_X1 U7849 ( .A(n6788), .ZN(n6635) );
  OAI222_X1 U7850 ( .A1(n9060), .A2(n6270), .B1(n9058), .B2(n6273), .C1(n6635), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7851 ( .A(n9777), .ZN(n6677) );
  OAI222_X1 U7852 ( .A1(n9613), .A2(n6272), .B1(n6677), .B2(P1_U3084), .C1(
        n6271), .C2(n9609), .ZN(P1_U3342) );
  INV_X1 U7853 ( .A(n6679), .ZN(n6444) );
  OAI222_X1 U7854 ( .A1(n9609), .A2(n6274), .B1(n6444), .B2(P1_U3084), .C1(
        n9613), .C2(n6273), .ZN(P1_U3343) );
  AND3_X1 U7855 ( .A1(n6806), .A2(n6809), .A3(n6804), .ZN(n6275) );
  INV_X1 U7856 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6298) );
  INV_X1 U7857 ( .A(n6277), .ZN(n6276) );
  NAND2_X1 U7858 ( .A1(n6276), .A2(n8925), .ZN(n8442) );
  NAND2_X1 U7859 ( .A1(n8442), .A2(n8440), .ZN(n6278) );
  NAND2_X1 U7860 ( .A1(n6281), .A2(n6283), .ZN(n6279) );
  NAND2_X1 U7861 ( .A1(n6278), .A2(n6279), .ZN(n6530) );
  OAI21_X1 U7862 ( .B1(n6278), .B2(n6279), .A(n6530), .ZN(n8927) );
  INV_X1 U7863 ( .A(n8927), .ZN(n6296) );
  XNOR2_X1 U7864 ( .A(n6811), .B(n8588), .ZN(n6280) );
  INV_X1 U7865 ( .A(n6281), .ZN(n6282) );
  NAND2_X1 U7866 ( .A1(n6283), .A2(n6282), .ZN(n6884) );
  NAND2_X1 U7867 ( .A1(n8442), .A2(n6884), .ZN(n6541) );
  INV_X1 U7868 ( .A(n8440), .ZN(n6288) );
  INV_X1 U7869 ( .A(n6884), .ZN(n6284) );
  NAND2_X1 U7870 ( .A1(n6278), .A2(n6284), .ZN(n6287) );
  INV_X1 U7871 ( .A(n4312), .ZN(n6286) );
  NAND2_X1 U7872 ( .A1(n6286), .A2(n8433), .ZN(n8381) );
  OAI211_X1 U7873 ( .C1(n6541), .C2(n6288), .A(n6287), .B(n8920), .ZN(n6292)
         );
  NAND2_X1 U7874 ( .A1(n6281), .A2(n8915), .ZN(n6290) );
  NAND2_X1 U7875 ( .A1(n6531), .A2(n8917), .ZN(n6289) );
  NAND2_X1 U7876 ( .A1(n6290), .A2(n6289), .ZN(n6346) );
  INV_X1 U7877 ( .A(n6346), .ZN(n6291) );
  NAND2_X1 U7878 ( .A1(n6292), .A2(n6291), .ZN(n8932) );
  INV_X1 U7879 ( .A(n8932), .ZN(n6295) );
  NAND2_X1 U7880 ( .A1(n6528), .A2(n9892), .ZN(n6988) );
  INV_X1 U7881 ( .A(n6988), .ZN(n6293) );
  AOI21_X1 U7882 ( .B1(n6283), .B2(n8925), .A(n6293), .ZN(n8930) );
  AOI22_X1 U7883 ( .A1(n8930), .A2(n9898), .B1(n9897), .B2(n8925), .ZN(n6294)
         );
  OAI211_X1 U7884 ( .C1(n6296), .C2(n9890), .A(n6295), .B(n6294), .ZN(n6431)
         );
  NAND2_X1 U7885 ( .A1(n9965), .A2(n6431), .ZN(n6297) );
  OAI21_X1 U7886 ( .B1(n9965), .B2(n6298), .A(n6297), .ZN(P2_U3454) );
  NAND2_X1 U7887 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8712), .ZN(n6299) );
  OAI21_X1 U7888 ( .B1(n8864), .B2(n8712), .A(n6299), .ZN(P2_U3575) );
  INV_X1 U7889 ( .A(n6300), .ZN(n6303) );
  INV_X1 U7890 ( .A(n9609), .ZN(n9606) );
  AOI22_X1 U7891 ( .A1(n6774), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9606), .ZN(n6301) );
  OAI21_X1 U7892 ( .B1(n6303), .B2(n9613), .A(n6301), .ZN(P1_U3341) );
  AOI22_X1 U7893 ( .A1(n7087), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9051), .ZN(n6302) );
  OAI21_X1 U7894 ( .B1(n6303), .B2(n9058), .A(n6302), .ZN(P2_U3346) );
  INV_X1 U7895 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6328) );
  NOR2_X1 U7896 ( .A1(n7558), .A2(n6311), .ZN(n6304) );
  NOR2_X1 U7897 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6446), .ZN(n6305) );
  AOI21_X1 U7898 ( .B1(n6446), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6305), .ZN(
        n6310) );
  MUX2_X1 U7899 ( .A(n6937), .B(P1_REG2_REG_4__SCAN_IN), .S(n6316), .Z(n9712)
         );
  NAND2_X1 U7900 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9688) );
  NOR2_X1 U7901 ( .A1(n9688), .A2(n9687), .ZN(n9686) );
  AOI21_X1 U7902 ( .B1(n9682), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9686), .ZN(
        n9697) );
  NAND2_X1 U7903 ( .A1(n9694), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7904 ( .B1(n9694), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6306), .ZN(
        n9696) );
  NAND2_X1 U7905 ( .A1(n6320), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6307) );
  OAI21_X1 U7906 ( .B1(n6320), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6307), .ZN(
        n6330) );
  NAND2_X1 U7907 ( .A1(n9712), .A2(n9713), .ZN(n9711) );
  NAND2_X1 U7908 ( .A1(n6316), .A2(n6937), .ZN(n6308) );
  NAND2_X1 U7909 ( .A1(n9711), .A2(n6308), .ZN(n6309) );
  NAND2_X1 U7910 ( .A1(n6309), .A2(n6310), .ZN(n6448) );
  OAI21_X1 U7911 ( .B1(n6310), .B2(n6309), .A(n6448), .ZN(n6326) );
  NOR2_X1 U7912 ( .A1(n6311), .A2(P1_U3084), .ZN(n7548) );
  AND2_X1 U7913 ( .A1(n7548), .A2(n6154), .ZN(n6312) );
  NAND2_X1 U7914 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n6314) );
  OAI21_X1 U7915 ( .B1(n9264), .B2(n6315), .A(n6314), .ZN(n6325) );
  INV_X1 U7916 ( .A(n6316), .ZN(n9722) );
  INV_X1 U7917 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6317) );
  MUX2_X1 U7918 ( .A(n6317), .B(P1_REG1_REG_4__SCAN_IN), .S(n6316), .Z(n9715)
         );
  NAND2_X1 U7919 ( .A1(n9682), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7920 ( .B1(n9682), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6318), .ZN(
        n9684) );
  NOR3_X1 U7921 ( .A1(n9705), .A2(n6261), .A3(n9684), .ZN(n9683) );
  AOI21_X1 U7922 ( .B1(n9682), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9683), .ZN(
        n9700) );
  XNOR2_X1 U7923 ( .A(n9694), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9699) );
  NOR2_X1 U7924 ( .A1(n9700), .A2(n9699), .ZN(n9698) );
  AOI21_X1 U7925 ( .B1(n9694), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9698), .ZN(
        n6334) );
  NAND2_X1 U7926 ( .A1(n6320), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7927 ( .B1(n6320), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6319), .ZN(
        n6333) );
  NOR2_X1 U7928 ( .A1(n6334), .A2(n6333), .ZN(n6332) );
  AOI21_X1 U7929 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6320), .A(n6332), .ZN(
        n9716) );
  NAND2_X1 U7930 ( .A1(n9715), .A2(n9716), .ZN(n9714) );
  OAI21_X1 U7931 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9722), .A(n9714), .ZN(
        n6323) );
  NAND2_X1 U7932 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6446), .ZN(n6321) );
  OAI21_X1 U7933 ( .B1(n6446), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6321), .ZN(
        n6322) );
  NOR2_X1 U7934 ( .A1(n6323), .A2(n6322), .ZN(n6436) );
  AOI211_X1 U7935 ( .C1(n6323), .C2(n6322), .A(n6436), .B(n9750), .ZN(n6324)
         );
  AOI211_X1 U7936 ( .C1(n9787), .C2(n6326), .A(n6325), .B(n6324), .ZN(n6327)
         );
  OAI21_X1 U7937 ( .B1(n9792), .B2(n6328), .A(n6327), .ZN(P1_U3246) );
  INV_X1 U7938 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6340) );
  AOI211_X1 U7939 ( .C1(n6331), .C2(n6330), .A(n6329), .B(n9763), .ZN(n6338)
         );
  AOI211_X1 U7940 ( .C1(n6334), .C2(n6333), .A(n6332), .B(n9750), .ZN(n6337)
         );
  NAND2_X1 U7941 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6707) );
  OAI21_X1 U7942 ( .B1(n9264), .B2(n6335), .A(n6707), .ZN(n6336) );
  NOR3_X1 U7943 ( .A1(n6338), .A2(n6337), .A3(n6336), .ZN(n6339) );
  OAI21_X1 U7944 ( .B1(n9792), .B2(n6340), .A(n6339), .ZN(P1_U3244) );
  AND2_X1 U7945 ( .A1(n6341), .A2(n9885), .ZN(n6497) );
  INV_X1 U7946 ( .A(n6497), .ZN(n6342) );
  NAND2_X1 U7947 ( .A1(n6342), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6349) );
  OAI21_X1 U7948 ( .B1(n6345), .B2(n6344), .A(n6343), .ZN(n6347) );
  AOI22_X1 U7949 ( .A1(n8612), .A2(n6347), .B1(n8634), .B2(n6346), .ZN(n6348)
         );
  OAI211_X1 U7950 ( .C1(n6528), .C2(n7687), .A(n6349), .B(n6348), .ZN(P2_U3224) );
  OR2_X1 U7951 ( .A1(n4310), .A2(P2_U3152), .ZN(n7553) );
  OAI21_X1 U7952 ( .B1(n6350), .B2(n7553), .A(n8590), .ZN(n6351) );
  NAND2_X1 U7953 ( .A1(n6361), .A2(n4926), .ZN(n6353) );
  NAND2_X1 U7954 ( .A1(n6353), .A2(n8712), .ZN(n6380) );
  AND2_X1 U7955 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8614) );
  INV_X1 U7956 ( .A(n6428), .ZN(n6356) );
  INV_X1 U7957 ( .A(n6471), .ZN(n6354) );
  INV_X1 U7958 ( .A(n6371), .ZN(n6507) );
  INV_X1 U7959 ( .A(n6394), .ZN(n6367) );
  INV_X1 U7960 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9966) );
  XOR2_X1 U7961 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6371), .Z(n6503) );
  NOR2_X1 U7962 ( .A1(n6504), .A2(n6503), .ZN(n6502) );
  MUX2_X1 U7963 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7821), .S(n6471), .Z(n6461)
         );
  NOR2_X1 U7964 ( .A1(n6462), .A2(n6461), .ZN(n6460) );
  AOI21_X1 U7965 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6354), .A(n6460), .ZN(
        n6419) );
  INV_X1 U7966 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6355) );
  MUX2_X1 U7967 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6355), .S(n6428), .Z(n6418)
         );
  NOR2_X1 U7968 ( .A1(n6419), .A2(n6418), .ZN(n6417) );
  NAND2_X1 U7969 ( .A1(n6489), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6357) );
  OAI21_X1 U7970 ( .B1(n6489), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6357), .ZN(
        n6485) );
  XNOR2_X1 U7971 ( .A(n6377), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U7972 ( .A1(n6365), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7973 ( .B1(n6365), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6358), .ZN(
        n6407) );
  NOR2_X1 U7974 ( .A1(n6408), .A2(n6407), .ZN(n6406) );
  XNOR2_X1 U7975 ( .A(n6511), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n6362) );
  AND2_X1 U7976 ( .A1(n4926), .A2(n6359), .ZN(n6360) );
  AOI211_X1 U7977 ( .C1(n6363), .C2(n6362), .A(n7977), .B(n6510), .ZN(n6364)
         );
  AOI211_X1 U7978 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9873), .A(n8614), .B(
        n6364), .ZN(n6384) );
  NAND2_X1 U7979 ( .A1(n6365), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6378) );
  INV_X1 U7980 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6366) );
  MUX2_X1 U7981 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6366), .S(n6365), .Z(n6413)
         );
  INV_X1 U7982 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U7983 ( .A1(n6489), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7984 ( .A1(n6367), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6370) );
  INV_X1 U7985 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7986 ( .A1(n6394), .A2(n6368), .ZN(n6369) );
  NAND4_X1 U7987 ( .A1(n6370), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .A4(n6369), .ZN(n6389) );
  NAND2_X1 U7988 ( .A1(n6389), .A2(n6370), .ZN(n6500) );
  XNOR2_X1 U7989 ( .A(n6371), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6501) );
  AOI22_X1 U7990 ( .A1(n6500), .A2(n6501), .B1(n6507), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n6467) );
  INV_X1 U7991 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7916) );
  MUX2_X1 U7992 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7916), .S(n6471), .Z(n6466)
         );
  NOR2_X1 U7993 ( .A1(n6467), .A2(n6466), .ZN(n6465) );
  NOR2_X1 U7994 ( .A1(n6471), .A2(n7916), .ZN(n6421) );
  MUX2_X1 U7995 ( .A(n4962), .B(P2_REG2_REG_4__SCAN_IN), .S(n6428), .Z(n6372)
         );
  OAI21_X1 U7996 ( .B1(n6465), .B2(n6421), .A(n6372), .ZN(n6424) );
  OAI21_X1 U7997 ( .B1(n4962), .B2(n6428), .A(n6424), .ZN(n6482) );
  INV_X1 U7998 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6373) );
  MUX2_X1 U7999 ( .A(n6373), .B(P2_REG2_REG_5__SCAN_IN), .S(n6489), .Z(n6483)
         );
  INV_X1 U8000 ( .A(n6483), .ZN(n6374) );
  NAND2_X1 U8001 ( .A1(n6482), .A2(n6374), .ZN(n6375) );
  NAND2_X1 U8002 ( .A1(n6376), .A2(n6375), .ZN(n6402) );
  MUX2_X1 U8003 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6835), .S(n6377), .Z(n6401)
         );
  NAND2_X1 U8004 ( .A1(n6402), .A2(n6401), .ZN(n6400) );
  OAI21_X1 U8005 ( .B1(n6835), .B2(n6405), .A(n6400), .ZN(n6412) );
  NAND2_X1 U8006 ( .A1(n6413), .A2(n6412), .ZN(n6411) );
  NAND2_X1 U8007 ( .A1(n6378), .A2(n6411), .ZN(n6382) );
  INV_X1 U8008 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6859) );
  MUX2_X1 U8009 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6859), .S(n6511), .Z(n6381)
         );
  NOR2_X1 U8010 ( .A1(n4310), .A2(n6359), .ZN(n6379) );
  NAND2_X1 U8011 ( .A1(n6382), .A2(n6381), .ZN(n6519) );
  OAI211_X1 U8012 ( .C1(n6382), .C2(n6381), .A(n9867), .B(n6519), .ZN(n6383)
         );
  OAI211_X1 U8013 ( .C1(n9869), .C2(n6520), .A(n6384), .B(n6383), .ZN(P2_U3253) );
  INV_X1 U8014 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7350) );
  NOR2_X1 U8015 ( .A1(n8745), .A2(n7350), .ZN(n6388) );
  NAND2_X1 U8016 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6386) );
  AOI211_X1 U8017 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3152), .A(n6388), .B(
        n6387), .ZN(n6393) );
  AND2_X1 U8018 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6391) );
  MUX2_X1 U8019 ( .A(n6368), .B(P2_REG2_REG_1__SCAN_IN), .S(n6394), .Z(n6390)
         );
  OAI211_X1 U8020 ( .C1(n6391), .C2(n6390), .A(n9867), .B(n6389), .ZN(n6392)
         );
  OAI211_X1 U8021 ( .C1(n9869), .C2(n6394), .A(n6393), .B(n6392), .ZN(P2_U3246) );
  NAND2_X1 U8022 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6648) );
  INV_X1 U8023 ( .A(n6648), .ZN(n6399) );
  AOI211_X1 U8024 ( .C1(n6397), .C2(n6396), .A(n7977), .B(n6395), .ZN(n6398)
         );
  AOI211_X1 U8025 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9873), .A(n6399), .B(
        n6398), .ZN(n6404) );
  OAI211_X1 U8026 ( .C1(n6402), .C2(n6401), .A(n9867), .B(n6400), .ZN(n6403)
         );
  OAI211_X1 U8027 ( .C1(n9869), .C2(n6405), .A(n6404), .B(n6403), .ZN(P2_U3251) );
  NOR2_X1 U8028 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6698), .ZN(n6410) );
  AOI211_X1 U8029 ( .C1(n6408), .C2(n6407), .A(n7977), .B(n6406), .ZN(n6409)
         );
  AOI211_X1 U8030 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9873), .A(n6410), .B(
        n6409), .ZN(n6415) );
  OAI211_X1 U8031 ( .C1(n6413), .C2(n6412), .A(n9867), .B(n6411), .ZN(n6414)
         );
  OAI211_X1 U8032 ( .C1(n9869), .C2(n6416), .A(n6415), .B(n6414), .ZN(P2_U3252) );
  AND2_X1 U8033 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6604) );
  AOI211_X1 U8034 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n7977), .ZN(n6420)
         );
  AOI211_X1 U8035 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9873), .A(n6604), .B(
        n6420), .ZN(n6427) );
  MUX2_X1 U8036 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n4962), .S(n6428), .Z(n6423)
         );
  INV_X1 U8037 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8038 ( .A1(n6423), .A2(n6422), .ZN(n6425) );
  OAI211_X1 U8039 ( .C1(n6465), .C2(n6425), .A(n9867), .B(n6424), .ZN(n6426)
         );
  OAI211_X1 U8040 ( .C1(n9869), .C2(n6428), .A(n6427), .B(n6426), .ZN(P2_U3249) );
  INV_X1 U8041 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8042 ( .A1(n9983), .A2(n6431), .ZN(n6432) );
  OAI21_X1 U8043 ( .B1(n9983), .B2(n6433), .A(n6432), .ZN(P2_U3521) );
  INV_X1 U8044 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6459) );
  INV_X1 U8045 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6434) );
  MUX2_X1 U8046 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6434), .S(n6679), .Z(n6442)
         );
  OR2_X1 U8047 ( .A1(n9769), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6440) );
  XNOR2_X1 U8048 ( .A(n9756), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n9753) );
  OR2_X1 U8049 ( .A1(n9738), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6438) );
  NOR2_X1 U8050 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9738), .ZN(n6435) );
  AOI21_X1 U8051 ( .B1(n9738), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6435), .ZN(
        n9744) );
  INV_X1 U8052 ( .A(n6450), .ZN(n9731) );
  XNOR2_X1 U8053 ( .A(n6450), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9733) );
  AOI21_X1 U8054 ( .B1(n6446), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6436), .ZN(
        n9732) );
  NAND2_X1 U8055 ( .A1(n9733), .A2(n9732), .ZN(n6437) );
  OAI21_X1 U8056 ( .B1(n9731), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6437), .ZN(
        n9743) );
  NAND2_X1 U8057 ( .A1(n9744), .A2(n9743), .ZN(n9742) );
  NAND2_X1 U8058 ( .A1(n6438), .A2(n9742), .ZN(n9752) );
  NOR2_X1 U8059 ( .A1(n9753), .A2(n9752), .ZN(n9751) );
  AOI21_X1 U8060 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9756), .A(n9751), .ZN(
        n9772) );
  INV_X1 U8061 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U8062 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9769), .B1(n6439), .B2(
        n9865), .ZN(n9771) );
  NAND2_X1 U8063 ( .A1(n9772), .A2(n9771), .ZN(n9770) );
  NAND2_X1 U8064 ( .A1(n6440), .A2(n9770), .ZN(n6441) );
  NAND2_X1 U8065 ( .A1(n6442), .A2(n6441), .ZN(n6671) );
  OAI21_X1 U8066 ( .B1(n6442), .B2(n6441), .A(n6671), .ZN(n6457) );
  OR2_X1 U8067 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6443), .ZN(n7392) );
  OAI21_X1 U8068 ( .B1(n9264), .B2(n6444), .A(n7392), .ZN(n6456) );
  XNOR2_X1 U8069 ( .A(n9756), .B(n7257), .ZN(n9758) );
  AOI22_X1 U8070 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9738), .B1(n6445), .B2(
        n7073), .ZN(n9740) );
  OR2_X1 U8071 ( .A1(n6446), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8072 ( .A1(n6448), .A2(n6447), .ZN(n9727) );
  XNOR2_X1 U8073 ( .A(n6450), .B(n6449), .ZN(n9728) );
  NOR2_X1 U8074 ( .A1(n9727), .A2(n9728), .ZN(n9726) );
  OAI21_X1 U8075 ( .B1(n9756), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6451), .ZN(
        n9766) );
  NAND2_X1 U8076 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9769), .ZN(n6452) );
  OAI21_X1 U8077 ( .B1(n9769), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6452), .ZN(
        n9765) );
  NOR2_X1 U8078 ( .A1(n9766), .A2(n9765), .ZN(n9764) );
  XNOR2_X1 U8079 ( .A(n6679), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6453) );
  AOI211_X1 U8080 ( .C1(n6454), .C2(n6453), .A(n6678), .B(n9763), .ZN(n6455)
         );
  AOI211_X1 U8081 ( .C1(n9786), .C2(n6457), .A(n6456), .B(n6455), .ZN(n6458)
         );
  OAI21_X1 U8082 ( .B1(n9792), .B2(n6459), .A(n6458), .ZN(P1_U3251) );
  NOR2_X1 U8083 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6599), .ZN(n6464) );
  AOI211_X1 U8084 ( .C1(n6462), .C2(n6461), .A(n6460), .B(n7977), .ZN(n6463)
         );
  AOI211_X1 U8085 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9873), .A(n6464), .B(
        n6463), .ZN(n6470) );
  AOI211_X1 U8086 ( .C1(n6467), .C2(n6466), .A(n6465), .B(n9871), .ZN(n6468)
         );
  INV_X1 U8087 ( .A(n6468), .ZN(n6469) );
  OAI211_X1 U8088 ( .C1(n9869), .C2(n6471), .A(n6470), .B(n6469), .ZN(P2_U3248) );
  INV_X1 U8089 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6477) );
  XOR2_X1 U8090 ( .A(n6473), .B(n6472), .Z(n6474) );
  AOI22_X1 U8091 ( .A1(n6474), .A2(n8612), .B1(n8623), .B2(n6277), .ZN(n6476)
         );
  INV_X1 U8092 ( .A(n6532), .ZN(n9896) );
  AOI22_X1 U8093 ( .A1(n8682), .A2(n6534), .B1(n8688), .B2(n9896), .ZN(n6475)
         );
  OAI211_X1 U8094 ( .C1(n6497), .C2(n6477), .A(n6476), .B(n6475), .ZN(P2_U3239) );
  INV_X1 U8095 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8096 ( .A1(n6750), .A2(P1_U4006), .ZN(n6478) );
  OAI21_X1 U8097 ( .B1(P1_U4006), .B2(n6479), .A(n6478), .ZN(P1_U3555) );
  INV_X1 U8098 ( .A(n6480), .ZN(n6498) );
  AOI22_X1 U8099 ( .A1(n7170), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9606), .ZN(n6481) );
  OAI21_X1 U8100 ( .B1(n6498), .B2(n9613), .A(n6481), .ZN(P1_U3340) );
  XOR2_X1 U8101 ( .A(n6483), .B(n6482), .Z(n6492) );
  NOR2_X1 U8102 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6568), .ZN(n6488) );
  AOI211_X1 U8103 ( .C1(n6486), .C2(n6485), .A(n7977), .B(n6484), .ZN(n6487)
         );
  AOI211_X1 U8104 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9873), .A(n6488), .B(
        n6487), .ZN(n6491) );
  INV_X1 U8105 ( .A(n9869), .ZN(n8750) );
  NAND2_X1 U8106 ( .A1(n8750), .A2(n6489), .ZN(n6490) );
  OAI211_X1 U8107 ( .C1(n6492), .C2(n9871), .A(n6491), .B(n6490), .ZN(P2_U3250) );
  INV_X1 U8108 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6885) );
  NOR2_X1 U8109 ( .A1(n7687), .A2(n9892), .ZN(n6495) );
  NAND2_X1 U8110 ( .A1(n6281), .A2(n9892), .ZN(n8441) );
  MUX2_X1 U8111 ( .A(n9892), .B(n8441), .S(n8382), .Z(n6493) );
  AOI21_X1 U8112 ( .B1(n6884), .B2(n6493), .A(n8690), .ZN(n6494) );
  AOI211_X1 U8113 ( .C1(n8682), .C2(n6277), .A(n6495), .B(n6494), .ZN(n6496)
         );
  OAI21_X1 U8114 ( .B1(n6497), .B2(n6885), .A(n6496), .ZN(P2_U3234) );
  INV_X1 U8115 ( .A(n7198), .ZN(n7092) );
  OAI222_X1 U8116 ( .A1(n9060), .A2(n6499), .B1(n9058), .B2(n6498), .C1(n7092), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XNOR2_X1 U8117 ( .A(n6501), .B(n6500), .ZN(n6509) );
  INV_X1 U8118 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7349) );
  OAI22_X1 U8119 ( .A1(n8745), .A2(n7349), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6477), .ZN(n6506) );
  AOI211_X1 U8120 ( .C1(n6504), .C2(n6503), .A(n6502), .B(n7977), .ZN(n6505)
         );
  AOI211_X1 U8121 ( .C1(n8750), .C2(n6507), .A(n6506), .B(n6505), .ZN(n6508)
         );
  OAI21_X1 U8122 ( .B1(n6509), .B2(n9871), .A(n6508), .ZN(P2_U3247) );
  NAND2_X1 U8123 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6870) );
  INV_X1 U8124 ( .A(n6870), .ZN(n6516) );
  INV_X1 U8125 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6512) );
  MUX2_X1 U8126 ( .A(n6512), .B(P2_REG1_REG_9__SCAN_IN), .S(n6626), .Z(n6513)
         );
  AOI211_X1 U8127 ( .C1(n6514), .C2(n6513), .A(n7977), .B(n6622), .ZN(n6515)
         );
  AOI211_X1 U8128 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9873), .A(n6516), .B(
        n6515), .ZN(n6524) );
  INV_X1 U8129 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6517) );
  MUX2_X1 U8130 ( .A(n6517), .B(P2_REG2_REG_9__SCAN_IN), .S(n6626), .Z(n6518)
         );
  INV_X1 U8131 ( .A(n6518), .ZN(n6522) );
  OAI21_X1 U8132 ( .B1(n6859), .B2(n6520), .A(n6519), .ZN(n6521) );
  NAND2_X1 U8133 ( .A1(n6522), .A2(n6521), .ZN(n6627) );
  OAI211_X1 U8134 ( .C1(n6522), .C2(n6521), .A(n9867), .B(n6627), .ZN(n6523)
         );
  OAI211_X1 U8135 ( .C1(n9869), .C2(n6525), .A(n6524), .B(n6523), .ZN(P2_U3254) );
  INV_X1 U8136 ( .A(n6526), .ZN(n6551) );
  INV_X1 U8137 ( .A(n9219), .ZN(n9212) );
  OAI222_X1 U8138 ( .A1(n9613), .A2(n6551), .B1(n9212), .B2(P1_U3084), .C1(
        n6527), .C2(n9609), .ZN(P1_U3339) );
  INV_X1 U8139 ( .A(n9030), .ZN(n9947) );
  NAND2_X1 U8140 ( .A1(n6276), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8141 ( .A1(n6530), .A2(n6529), .ZN(n6986) );
  OR2_X1 U8142 ( .A1(n6531), .A2(n6532), .ZN(n8443) );
  NAND2_X1 U8143 ( .A1(n6531), .A2(n6532), .ZN(n8434) );
  AND2_X1 U8144 ( .A1(n8443), .A2(n8434), .ZN(n6542) );
  NAND2_X1 U8145 ( .A1(n6986), .A2(n8383), .ZN(n6985) );
  NAND2_X1 U8146 ( .A1(n6596), .A2(n6532), .ZN(n6533) );
  NAND2_X1 U8147 ( .A1(n6985), .A2(n6533), .ZN(n6535) );
  NAND2_X1 U8148 ( .A1(n6535), .A2(n6540), .ZN(n6580) );
  OR2_X1 U8149 ( .A1(n6535), .A2(n6540), .ZN(n6536) );
  NAND2_X1 U8150 ( .A1(n6580), .A2(n6536), .ZN(n6803) );
  OR2_X1 U8151 ( .A1(n6988), .A2(n9896), .ZN(n6537) );
  INV_X1 U8152 ( .A(n6537), .ZN(n6987) );
  INV_X1 U8153 ( .A(n6958), .ZN(n6538) );
  OAI21_X1 U8154 ( .B1(n6594), .B2(n6987), .A(n6538), .ZN(n6815) );
  OAI22_X1 U8155 ( .A1(n6815), .A2(n9957), .B1(n6594), .B2(n9955), .ZN(n6549)
         );
  INV_X1 U8156 ( .A(n7609), .ZN(n6539) );
  NAND2_X1 U8157 ( .A1(n6803), .A2(n6539), .ZN(n6548) );
  AOI22_X1 U8158 ( .A1(n8915), .A2(n6531), .B1(n8711), .B2(n8917), .ZN(n6547)
         );
  INV_X1 U8159 ( .A(n6540), .ZN(n6543) );
  NAND2_X1 U8160 ( .A1(n6980), .A2(n6542), .ZN(n6981) );
  NAND2_X1 U8161 ( .A1(n6981), .A2(n8443), .ZN(n6544) );
  NAND2_X1 U8162 ( .A1(n6544), .A2(n6543), .ZN(n6582) );
  OAI21_X1 U8163 ( .B1(n6543), .B2(n6544), .A(n6582), .ZN(n6545) );
  NAND2_X1 U8164 ( .A1(n6545), .A2(n8920), .ZN(n6546) );
  NAND3_X1 U8165 ( .A1(n6548), .A2(n6547), .A3(n6546), .ZN(n6818) );
  AOI211_X1 U8166 ( .C1(n9947), .C2(n6803), .A(n6549), .B(n6818), .ZN(n6572)
         );
  NAND2_X1 U8167 ( .A1(n9980), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U8168 ( .B1(n6572), .B2(n9980), .A(n6550), .ZN(P2_U3523) );
  INV_X1 U8169 ( .A(n7418), .ZN(n7196) );
  OAI222_X1 U8170 ( .A1(n9060), .A2(n6552), .B1(n9058), .B2(n6551), .C1(n7196), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8171 ( .A(n6741), .ZN(n6553) );
  OR2_X1 U8172 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U8173 ( .A1(n9181), .A2(n6555), .ZN(n6695) );
  INV_X1 U8174 ( .A(n9636), .ZN(n9188) );
  AOI22_X1 U8175 ( .A1(n9188), .A2(n6717), .B1(n9192), .B2(n6764), .ZN(n6560)
         );
  OAI21_X1 U8176 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(n9704) );
  NAND2_X1 U8177 ( .A1(n9704), .A2(n9173), .ZN(n6559) );
  OAI211_X1 U8178 ( .C1(n6695), .C2(n6561), .A(n6560), .B(n6559), .ZN(P1_U3230) );
  XNOR2_X1 U8179 ( .A(n6563), .B(n6562), .ZN(n6571) );
  NAND2_X1 U8180 ( .A1(n8688), .A2(n6825), .ZN(n6567) );
  OR2_X1 U8181 ( .A1(n6970), .A2(n8863), .ZN(n6565) );
  NAND2_X1 U8182 ( .A1(n8711), .A2(n8915), .ZN(n6564) );
  NAND2_X1 U8183 ( .A1(n6565), .A2(n6564), .ZN(n6584) );
  NAND2_X1 U8184 ( .A1(n8634), .A2(n6584), .ZN(n6566) );
  OAI211_X1 U8185 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6568), .A(n6567), .B(n6566), .ZN(n6569) );
  AOI21_X1 U8186 ( .B1(n8680), .B2(n7099), .A(n6569), .ZN(n6570) );
  OAI21_X1 U8187 ( .B1(n6571), .B2(n8690), .A(n6570), .ZN(P2_U3229) );
  INV_X1 U8188 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6574) );
  OR2_X1 U8189 ( .A1(n6572), .A2(n9963), .ZN(n6573) );
  OAI21_X1 U8190 ( .B1(n9965), .B2(n6574), .A(n6573), .ZN(P2_U3460) );
  INV_X1 U8191 ( .A(n6575), .ZN(n6578) );
  AOI22_X1 U8192 ( .A1(n9249), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9606), .ZN(n6576) );
  OAI21_X1 U8193 ( .B1(n6578), .B2(n9613), .A(n6576), .ZN(P1_U3337) );
  AOI22_X1 U8194 ( .A1(n8720), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9051), .ZN(n6577) );
  OAI21_X1 U8195 ( .B1(n6578), .B2(n9058), .A(n6577), .ZN(P2_U3342) );
  INV_X1 U8196 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8197 ( .A1(n8710), .A2(n7102), .ZN(n8450) );
  NAND2_X1 U8198 ( .A1(n8426), .A2(n8450), .ZN(n8386) );
  INV_X1 U8199 ( .A(n8386), .ZN(n6826) );
  NAND2_X1 U8200 ( .A1(n4829), .A2(n6594), .ZN(n6579) );
  NAND2_X1 U8201 ( .A1(n6580), .A2(n6579), .ZN(n6956) );
  NAND2_X1 U8202 ( .A1(n8711), .A2(n9905), .ZN(n6830) );
  NAND2_X1 U8203 ( .A1(n6595), .A2(n9905), .ZN(n6581) );
  XNOR2_X1 U8204 ( .A(n6826), .B(n6829), .ZN(n7107) );
  INV_X1 U8205 ( .A(n6955), .ZN(n8384) );
  NAND2_X1 U8206 ( .A1(n6831), .A2(n6830), .ZN(n6583) );
  XNOR2_X1 U8207 ( .A(n6583), .B(n8386), .ZN(n6585) );
  AOI21_X1 U8208 ( .B1(n6585), .B2(n8920), .A(n6584), .ZN(n7104) );
  AOI211_X1 U8209 ( .C1(n6825), .C2(n6957), .A(n9957), .B(n4515), .ZN(n7100)
         );
  AOI21_X1 U8210 ( .B1(n9897), .B2(n6825), .A(n7100), .ZN(n6586) );
  OAI211_X1 U8211 ( .C1(n9890), .C2(n7107), .A(n7104), .B(n6586), .ZN(n6589)
         );
  NAND2_X1 U8212 ( .A1(n6589), .A2(n9965), .ZN(n6587) );
  OAI21_X1 U8213 ( .B1(n9965), .B2(n6588), .A(n6587), .ZN(P2_U3466) );
  INV_X1 U8214 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8215 ( .A1(n6589), .A2(n9983), .ZN(n6590) );
  OAI21_X1 U8216 ( .B1(n9983), .B2(n6591), .A(n6590), .ZN(P2_U3525) );
  XNOR2_X1 U8217 ( .A(n6593), .B(n6592), .ZN(n6601) );
  OAI22_X1 U8218 ( .A1(n7687), .A2(n6594), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6599), .ZN(n6598) );
  OAI22_X1 U8219 ( .A1(n6596), .A2(n8685), .B1(n8672), .B2(n6595), .ZN(n6597)
         );
  AOI211_X1 U8220 ( .C1(n8680), .C2(n6599), .A(n6598), .B(n6597), .ZN(n6600)
         );
  OAI21_X1 U8221 ( .B1(n8690), .B2(n6601), .A(n6600), .ZN(P2_U3220) );
  INV_X1 U8222 ( .A(n9905), .ZN(n6605) );
  INV_X1 U8223 ( .A(n8710), .ZN(n6602) );
  OAI22_X1 U8224 ( .A1(n4829), .A2(n8685), .B1(n8672), .B2(n6602), .ZN(n6603)
         );
  AOI211_X1 U8225 ( .C1(n8688), .C2(n6605), .A(n6604), .B(n6603), .ZN(n6611)
         );
  OAI21_X1 U8226 ( .B1(n6608), .B2(n6607), .A(n6606), .ZN(n6609) );
  NAND2_X1 U8227 ( .A1(n6609), .A2(n8612), .ZN(n6610) );
  OAI211_X1 U8228 ( .C1(n8633), .C2(n6959), .A(n6611), .B(n6610), .ZN(P2_U3232) );
  INV_X1 U8229 ( .A(n6612), .ZN(n6614) );
  INV_X1 U8230 ( .A(n7960), .ZN(n7971) );
  OAI222_X1 U8231 ( .A1(n9060), .A2(n6613), .B1(n9058), .B2(n6614), .C1(
        P2_U3152), .C2(n7971), .ZN(P2_U3343) );
  OAI222_X1 U8232 ( .A1(n9609), .A2(n6615), .B1(n9613), .B2(n6614), .C1(
        P1_U3084), .C2(n9234), .ZN(P1_U3338) );
  OAI21_X1 U8233 ( .B1(n9805), .B2(n8332), .A(n6738), .ZN(n6617) );
  INV_X2 U8234 ( .A(n9864), .ZN(n9853) );
  INV_X1 U8235 ( .A(n6764), .ZN(n6721) );
  INV_X1 U8236 ( .A(n6750), .ZN(n6661) );
  NAND2_X1 U8237 ( .A1(n6661), .A2(n6764), .ZN(n6749) );
  NAND2_X1 U8238 ( .A1(n6750), .A2(n6721), .ZN(n8190) );
  NAND2_X1 U8239 ( .A1(n6749), .A2(n8190), .ZN(n8301) );
  INV_X1 U8240 ( .A(n6620), .ZN(n6723) );
  NOR2_X1 U8241 ( .A1(n8348), .A2(n6723), .ZN(n6619) );
  AOI22_X1 U8242 ( .A1(n8301), .A2(n6619), .B1(n9485), .B2(n6717), .ZN(n6767)
         );
  OAI21_X1 U8243 ( .B1(n6721), .B2(n6620), .A(n6767), .ZN(n6643) );
  NAND2_X1 U8244 ( .A1(n6643), .A2(n9853), .ZN(n6621) );
  OAI21_X1 U8245 ( .B1(n9853), .B2(n6261), .A(n6621), .ZN(P1_U3523) );
  INV_X1 U8246 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6623) );
  MUX2_X1 U8247 ( .A(n6623), .B(P2_REG1_REG_10__SCAN_IN), .S(n6788), .Z(n6624)
         );
  NOR2_X1 U8248 ( .A1(n6625), .A2(n6624), .ZN(n6787) );
  AOI211_X1 U8249 ( .C1(n6625), .C2(n6624), .A(n6787), .B(n7977), .ZN(n6637)
         );
  NAND2_X1 U8250 ( .A1(n6626), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U8251 ( .A1(n6628), .A2(n6627), .ZN(n6632) );
  INV_X1 U8252 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6629) );
  MUX2_X1 U8253 ( .A(n6629), .B(P2_REG2_REG_10__SCAN_IN), .S(n6788), .Z(n6630)
         );
  INV_X1 U8254 ( .A(n6630), .ZN(n6631) );
  NAND2_X1 U8255 ( .A1(n6631), .A2(n6632), .ZN(n6783) );
  OAI211_X1 U8256 ( .C1(n6632), .C2(n6631), .A(n9867), .B(n6783), .ZN(n6634)
         );
  AND2_X1 U8257 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6948) );
  AOI21_X1 U8258 ( .B1(n9873), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6948), .ZN(
        n6633) );
  OAI211_X1 U8259 ( .C1(n9869), .C2(n6635), .A(n6634), .B(n6633), .ZN(n6636)
         );
  OR2_X1 U8260 ( .A1(n6637), .A2(n6636), .ZN(P2_U3255) );
  OAI21_X1 U8261 ( .B1(n9602), .B2(P1_D_REG_0__SCAN_IN), .A(n9603), .ZN(n6641)
         );
  INV_X1 U8262 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U8263 ( .A1(n6641), .A2(n6640), .ZN(n6740) );
  NAND2_X1 U8264 ( .A1(n6643), .A2(n9850), .ZN(n6644) );
  OAI21_X1 U8265 ( .B1(n9850), .B2(n6645), .A(n6644), .ZN(P1_U3454) );
  AOI21_X1 U8266 ( .B1(n6647), .B2(n6646), .A(n4401), .ZN(n6652) );
  AOI22_X1 U8267 ( .A1(n8623), .A2(n8710), .B1(n8682), .B2(n8708), .ZN(n6649)
         );
  OAI211_X1 U8268 ( .C1(n9913), .C2(n7687), .A(n6649), .B(n6648), .ZN(n6650)
         );
  AOI21_X1 U8269 ( .B1(n6838), .B2(n8680), .A(n6650), .ZN(n6651) );
  OAI21_X1 U8270 ( .B1(n6652), .B2(n8690), .A(n6651), .ZN(P2_U3241) );
  XNOR2_X1 U8271 ( .A(n6654), .B(n6653), .ZN(n6656) );
  AOI21_X1 U8272 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(n6658) );
  AOI21_X1 U8273 ( .B1(n6659), .B2(n4583), .A(n6658), .ZN(n6665) );
  INV_X1 U8274 ( .A(n6695), .ZN(n6663) );
  NOR2_X1 U8275 ( .A1(n9841), .A2(n6760), .ZN(n9808) );
  AOI22_X1 U8276 ( .A1(n9188), .A2(n9211), .B1(n9808), .B2(n9646), .ZN(n6660)
         );
  OAI21_X1 U8277 ( .B1(n6661), .B2(n9632), .A(n6660), .ZN(n6662) );
  AOI21_X1 U8278 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6663), .A(n6662), .ZN(
        n6664) );
  OAI21_X1 U8279 ( .B1(n6665), .B2(n9642), .A(n6664), .ZN(P1_U3220) );
  INV_X1 U8280 ( .A(n6666), .ZN(n6669) );
  AOI22_X1 U8281 ( .A1(n9266), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9606), .ZN(n6667) );
  OAI21_X1 U8282 ( .B1(n6669), .B2(n9613), .A(n6667), .ZN(P1_U3336) );
  INV_X1 U8283 ( .A(n8732), .ZN(n6668) );
  OAI222_X1 U8284 ( .A1(n9060), .A2(n7863), .B1(n9058), .B2(n6669), .C1(n6668), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8285 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6687) );
  INV_X1 U8286 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U8287 ( .A1(n9777), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n6670), .B2(
        n6677), .ZN(n9783) );
  OAI21_X1 U8288 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6679), .A(n6671), .ZN(
        n9784) );
  NAND2_X1 U8289 ( .A1(n9783), .A2(n9784), .ZN(n9782) );
  OAI21_X1 U8290 ( .B1(n9777), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9782), .ZN(
        n6674) );
  INV_X1 U8291 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8292 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6672), .S(n6774), .Z(n6673)
         );
  NAND2_X1 U8293 ( .A1(n6673), .A2(n6674), .ZN(n6769) );
  OAI21_X1 U8294 ( .B1(n6674), .B2(n6673), .A(n6769), .ZN(n6685) );
  INV_X1 U8295 ( .A(n6774), .ZN(n6676) );
  NAND2_X1 U8296 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6675) );
  OAI21_X1 U8297 ( .B1(n9264), .B2(n6676), .A(n6675), .ZN(n6684) );
  AOI22_X1 U8298 ( .A1(n9777), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n5787), .B2(
        n6677), .ZN(n9780) );
  OAI21_X1 U8299 ( .B1(n9777), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9779), .ZN(
        n6682) );
  NAND2_X1 U8300 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6774), .ZN(n6680) );
  OAI21_X1 U8301 ( .B1(n6774), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6680), .ZN(
        n6681) );
  NOR2_X1 U8302 ( .A1(n6681), .A2(n6682), .ZN(n6773) );
  AOI211_X1 U8303 ( .C1(n6682), .C2(n6681), .A(n6773), .B(n9763), .ZN(n6683)
         );
  AOI211_X1 U8304 ( .C1(n9786), .C2(n6685), .A(n6684), .B(n6683), .ZN(n6686)
         );
  OAI21_X1 U8305 ( .B1(n9792), .B2(n6687), .A(n6686), .ZN(P1_U3253) );
  INV_X1 U8306 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6694) );
  OAI21_X1 U8307 ( .B1(n6689), .B2(n4400), .A(n6688), .ZN(n6690) );
  NAND2_X1 U8308 ( .A1(n6690), .A2(n9173), .ZN(n6693) );
  OAI22_X1 U8309 ( .A1(n6718), .A2(n9632), .B1(n9636), .B2(n6930), .ZN(n6691)
         );
  AOI21_X1 U8310 ( .B1(n9192), .B2(n6876), .A(n6691), .ZN(n6692) );
  OAI211_X1 U8311 ( .C1(n6695), .C2(n6694), .A(n6693), .B(n6692), .ZN(P1_U3235) );
  XNOR2_X1 U8312 ( .A(n6697), .B(n6696), .ZN(n6702) );
  INV_X1 U8313 ( .A(n6975), .ZN(n9920) );
  OAI22_X1 U8314 ( .A1(n7687), .A2(n9920), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6698), .ZN(n6700) );
  OAI22_X1 U8315 ( .A1(n6970), .A2(n8685), .B1(n8672), .B2(n7023), .ZN(n6699)
         );
  AOI211_X1 U8316 ( .C1(n6972), .C2(n8680), .A(n6700), .B(n6699), .ZN(n6701)
         );
  OAI21_X1 U8317 ( .B1(n6702), .B2(n8690), .A(n6701), .ZN(P2_U3215) );
  OAI21_X1 U8318 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6706) );
  NAND2_X1 U8319 ( .A1(n6706), .A2(n9173), .ZN(n6712) );
  INV_X1 U8320 ( .A(n6707), .ZN(n6708) );
  AOI21_X1 U8321 ( .B1(n9160), .B2(n9211), .A(n6708), .ZN(n6709) );
  OAI21_X1 U8322 ( .B1(n6912), .B2(n9636), .A(n6709), .ZN(n6710) );
  AOI21_X1 U8323 ( .B1(n9192), .B2(n6921), .A(n6710), .ZN(n6711) );
  OAI211_X1 U8324 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9650), .A(n6712), .B(
        n6711), .ZN(P1_U3216) );
  INV_X1 U8325 ( .A(n6713), .ZN(n6716) );
  AOI22_X1 U8326 ( .A1(n8749), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9051), .ZN(n6714) );
  OAI21_X1 U8327 ( .B1(n6716), .B2(n9058), .A(n6714), .ZN(P2_U3340) );
  AOI22_X1 U8328 ( .A1(n9276), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9606), .ZN(n6715) );
  OAI21_X1 U8329 ( .B1(n6716), .B2(n9613), .A(n6715), .ZN(P1_U3335) );
  INV_X1 U8330 ( .A(n9805), .ZN(n9848) );
  NAND2_X1 U8331 ( .A1(n6750), .A2(n6764), .ZN(n6737) );
  NAND2_X1 U8332 ( .A1(n6718), .A2(n6760), .ZN(n6719) );
  NAND2_X1 U8333 ( .A1(n6913), .A2(n6876), .ZN(n8193) );
  NAND2_X1 U8334 ( .A1(n9211), .A2(n6896), .ZN(n8195) );
  NAND2_X1 U8335 ( .A1(n6720), .A2(n8303), .ZN(n6898) );
  OAI21_X1 U8336 ( .B1(n6720), .B2(n8303), .A(n6898), .ZN(n6881) );
  OAI21_X1 U8337 ( .B1(n6756), .B2(n6764), .A(n6876), .ZN(n6722) );
  NAND2_X1 U8338 ( .A1(n6918), .A2(n6722), .ZN(n6879) );
  OAI22_X1 U8339 ( .A1(n6879), .A2(n9843), .B1(n6896), .B2(n9841), .ZN(n6733)
         );
  NAND2_X1 U8340 ( .A1(n8350), .A2(n8296), .ZN(n6724) );
  OR2_X1 U8341 ( .A1(n8292), .A2(n8295), .ZN(n8341) );
  INV_X1 U8342 ( .A(n9488), .ZN(n7655) );
  NAND2_X1 U8343 ( .A1(n6747), .A2(n6725), .ZN(n8189) );
  XNOR2_X1 U8344 ( .A(n8189), .B(n8303), .ZN(n6732) );
  NAND2_X1 U8345 ( .A1(n6129), .A2(n9283), .ZN(n6728) );
  MUX2_X1 U8346 ( .A(n6728), .B(n6727), .S(n6726), .Z(n9498) );
  INV_X1 U8347 ( .A(n9498), .ZN(n7476) );
  INV_X1 U8348 ( .A(n9483), .ZN(n7630) );
  OAI22_X1 U8349 ( .A1(n6718), .A2(n7630), .B1(n6930), .B2(n7744), .ZN(n6730)
         );
  AOI21_X1 U8350 ( .B1(n6881), .B2(n7476), .A(n6730), .ZN(n6731) );
  OAI21_X1 U8351 ( .B1(n7655), .B2(n6732), .A(n6731), .ZN(n6875) );
  AOI211_X1 U8352 ( .C1(n9848), .C2(n6881), .A(n6733), .B(n6875), .ZN(n6797)
         );
  NAND2_X1 U8353 ( .A1(n9864), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6734) );
  OAI21_X1 U8354 ( .B1(n6797), .B2(n9864), .A(n6734), .ZN(P1_U3525) );
  OAI21_X1 U8355 ( .B1(n6735), .B2(n6737), .A(n6736), .ZN(n6751) );
  INV_X1 U8356 ( .A(n6751), .ZN(n9806) );
  INV_X1 U8357 ( .A(n6738), .ZN(n6739) );
  NAND2_X1 U8358 ( .A1(n6739), .A2(n9804), .ZN(n9802) );
  NOR2_X1 U8359 ( .A1(n9802), .A2(n6740), .ZN(n6742) );
  NAND2_X1 U8360 ( .A1(n6742), .A2(n6741), .ZN(n6755) );
  NAND2_X1 U8361 ( .A1(n9804), .A2(n8292), .ZN(n6743) );
  NAND2_X1 U8362 ( .A1(n9456), .A2(n8296), .ZN(n7677) );
  INV_X1 U8363 ( .A(n6747), .ZN(n6748) );
  AOI21_X1 U8364 ( .B1(n6735), .B2(n6749), .A(n6748), .ZN(n6754) );
  AOI22_X1 U8365 ( .A1(n9211), .A2(n9485), .B1(n9483), .B2(n6750), .ZN(n6753)
         );
  NAND2_X1 U8366 ( .A1(n6751), .A2(n7476), .ZN(n6752) );
  OAI211_X1 U8367 ( .C1(n6754), .C2(n7655), .A(n6753), .B(n6752), .ZN(n9810)
         );
  NAND2_X1 U8368 ( .A1(n9810), .A2(n9313), .ZN(n6763) );
  NOR2_X2 U8369 ( .A1(n6755), .A2(n8296), .ZN(n9492) );
  XNOR2_X1 U8370 ( .A(n6756), .B(n6764), .ZN(n6757) );
  NOR2_X1 U8371 ( .A1(n6757), .A2(n9843), .ZN(n9807) );
  INV_X2 U8372 ( .A(n7669), .ZN(n9474) );
  AOI22_X1 U8373 ( .A1(n9465), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9474), .ZN(n6759) );
  OAI21_X1 U8374 ( .B1(n6760), .B2(n9477), .A(n6759), .ZN(n6761) );
  AOI21_X1 U8375 ( .B1(n9492), .B2(n9807), .A(n6761), .ZN(n6762) );
  OAI211_X1 U8376 ( .C1(n9806), .C2(n7677), .A(n6763), .B(n6762), .ZN(P1_U3290) );
  AOI22_X1 U8377 ( .A1(n9465), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9474), .ZN(n6766) );
  OAI21_X1 U8378 ( .B1(n9441), .B2(n8017), .A(n6764), .ZN(n6765) );
  OAI211_X1 U8379 ( .C1(n6767), .C2(n9489), .A(n6766), .B(n6765), .ZN(P1_U3291) );
  INV_X1 U8380 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6782) );
  INV_X1 U8381 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6768) );
  MUX2_X1 U8382 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6768), .S(n7170), .Z(n6771)
         );
  OAI21_X1 U8383 ( .B1(n6774), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6769), .ZN(
        n6770) );
  NAND2_X1 U8384 ( .A1(n6771), .A2(n6770), .ZN(n7164) );
  OAI21_X1 U8385 ( .B1(n6771), .B2(n6770), .A(n7164), .ZN(n6780) );
  INV_X1 U8386 ( .A(n7170), .ZN(n6772) );
  NAND2_X1 U8387 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7567) );
  OAI21_X1 U8388 ( .B1(n9264), .B2(n6772), .A(n7567), .ZN(n6779) );
  MUX2_X1 U8389 ( .A(n6775), .B(P1_REG2_REG_13__SCAN_IN), .S(n7170), .Z(n6776)
         );
  AOI211_X1 U8390 ( .C1(n6777), .C2(n6776), .A(n7169), .B(n9763), .ZN(n6778)
         );
  AOI211_X1 U8391 ( .C1(n9786), .C2(n6780), .A(n6779), .B(n6778), .ZN(n6781)
         );
  OAI21_X1 U8392 ( .B1(n9792), .B2(n6782), .A(n6781), .ZN(P1_U3254) );
  NAND2_X1 U8393 ( .A1(n6788), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U8394 ( .A1(n6784), .A2(n6783), .ZN(n6786) );
  INV_X1 U8395 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7119) );
  MUX2_X1 U8396 ( .A(n7119), .B(P2_REG2_REG_11__SCAN_IN), .S(n7047), .Z(n6785)
         );
  NOR2_X1 U8397 ( .A1(n6786), .A2(n6785), .ZN(n7051) );
  AOI21_X1 U8398 ( .B1(n6786), .B2(n6785), .A(n7051), .ZN(n6796) );
  NOR2_X1 U8399 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5107), .ZN(n6793) );
  INV_X1 U8400 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U8401 ( .A(n6789), .B(P2_REG1_REG_11__SCAN_IN), .S(n7047), .Z(n6790)
         );
  AOI211_X1 U8402 ( .C1(n6791), .C2(n6790), .A(n7039), .B(n7977), .ZN(n6792)
         );
  AOI211_X1 U8403 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9873), .A(n6793), .B(
        n6792), .ZN(n6795) );
  NAND2_X1 U8404 ( .A1(n8750), .A2(n7047), .ZN(n6794) );
  OAI211_X1 U8405 ( .C1(n6796), .C2(n9871), .A(n6795), .B(n6794), .ZN(P2_U3256) );
  OR2_X1 U8406 ( .A1(n6797), .A2(n9849), .ZN(n6798) );
  OAI21_X1 U8407 ( .B1(n9850), .B2(n5624), .A(n6798), .ZN(P1_U3460) );
  INV_X1 U8408 ( .A(n6799), .ZN(n6801) );
  OAI222_X1 U8409 ( .A1(n9060), .A2(n6800), .B1(n9058), .B2(n6801), .C1(
        P2_U3152), .C2(n8379), .ZN(P2_U3339) );
  OAI222_X1 U8410 ( .A1(n9609), .A2(n6802), .B1(n9613), .B2(n6801), .C1(n9283), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U8411 ( .A(n6803), .ZN(n6822) );
  NAND3_X1 U8412 ( .A1(n6806), .A2(n6805), .A3(n6804), .ZN(n6807) );
  OR2_X1 U8413 ( .A1(n6811), .A2(n8379), .ZN(n6823) );
  INV_X1 U8414 ( .A(n6823), .ZN(n6812) );
  NAND2_X1 U8415 ( .A1(n8933), .A2(n6812), .ZN(n7619) );
  NOR2_X1 U8416 ( .A1(n8933), .A2(n7916), .ZN(n6817) );
  OAI22_X1 U8417 ( .A1(n8850), .A2(n6815), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8844), .ZN(n6816) );
  AOI211_X1 U8418 ( .C1(n8933), .C2(n6818), .A(n6817), .B(n6816), .ZN(n6821)
         );
  NOR2_X1 U8419 ( .A1(n5516), .A2(n4312), .ZN(n6819) );
  NAND2_X1 U8420 ( .A1(n8926), .A2(n4828), .ZN(n6820) );
  OAI211_X1 U8421 ( .C1(n6822), .C2(n7619), .A(n6821), .B(n6820), .ZN(P2_U3293) );
  NAND2_X1 U8422 ( .A1(n7609), .A2(n6823), .ZN(n6824) );
  NOR2_X1 U8423 ( .A1(n6825), .A2(n8710), .ZN(n6828) );
  NAND2_X1 U8424 ( .A1(n6826), .A2(n8710), .ZN(n6827) );
  NAND2_X1 U8425 ( .A1(n6970), .A2(n6841), .ZN(n8459) );
  INV_X1 U8426 ( .A(n6970), .ZN(n8709) );
  NAND2_X1 U8427 ( .A1(n9913), .A2(n8709), .ZN(n8452) );
  INV_X1 U8428 ( .A(n6833), .ZN(n8387) );
  XNOR2_X1 U8429 ( .A(n6845), .B(n8387), .ZN(n9912) );
  AND2_X1 U8430 ( .A1(n8450), .A2(n6830), .ZN(n8449) );
  OAI21_X1 U8431 ( .B1(n6833), .B2(n6832), .A(n6967), .ZN(n6834) );
  AOI222_X1 U8432 ( .A1(n8920), .A2(n6834), .B1(n8708), .B2(n8917), .C1(n8710), 
        .C2(n8915), .ZN(n9915) );
  MUX2_X1 U8433 ( .A(n6835), .B(n9915), .S(n8933), .Z(n6843) );
  NAND2_X1 U8434 ( .A1(n6836), .A2(n6841), .ZN(n6837) );
  NAND2_X1 U8435 ( .A1(n6971), .A2(n6837), .ZN(n9914) );
  INV_X1 U8436 ( .A(n6838), .ZN(n6839) );
  OAI22_X1 U8437 ( .A1(n8850), .A2(n9914), .B1(n6839), .B2(n8844), .ZN(n6840)
         );
  AOI21_X1 U8438 ( .B1(n8926), .B2(n6841), .A(n6840), .ZN(n6842) );
  OAI211_X1 U8439 ( .C1(n8924), .C2(n9912), .A(n6843), .B(n6842), .ZN(P2_U3290) );
  NAND2_X1 U8440 ( .A1(n9913), .A2(n6970), .ZN(n6844) );
  OR2_X1 U8441 ( .A1(n6975), .A2(n6854), .ZN(n6850) );
  NAND2_X1 U8442 ( .A1(n6975), .A2(n6854), .ZN(n8458) );
  NOR2_X1 U8443 ( .A1(n6975), .A2(n8708), .ZN(n6846) );
  AOI21_X1 U8444 ( .B1(n6966), .B2(n8460), .A(n6846), .ZN(n6847) );
  OR2_X1 U8445 ( .A1(n8615), .A2(n7023), .ZN(n8466) );
  NAND2_X1 U8446 ( .A1(n8615), .A2(n7023), .ZN(n8465) );
  NAND2_X1 U8447 ( .A1(n8466), .A2(n8465), .ZN(n8463) );
  OR2_X1 U8448 ( .A1(n6847), .A2(n8463), .ZN(n6848) );
  NAND2_X1 U8449 ( .A1(n7002), .A2(n6848), .ZN(n9926) );
  INV_X1 U8450 ( .A(n8460), .ZN(n8456) );
  AND2_X1 U8451 ( .A1(n8456), .A2(n8459), .ZN(n6849) );
  NAND2_X1 U8452 ( .A1(n6967), .A2(n6849), .ZN(n6852) );
  AND2_X1 U8453 ( .A1(n6852), .A2(n6850), .ZN(n6853) );
  INV_X1 U8454 ( .A(n8463), .ZN(n8389) );
  INV_X1 U8455 ( .A(n6850), .ZN(n8462) );
  NOR2_X1 U8456 ( .A1(n8462), .A2(n8463), .ZN(n6851) );
  NAND2_X1 U8457 ( .A1(n6852), .A2(n6851), .ZN(n7007) );
  OAI21_X1 U8458 ( .B1(n6853), .B2(n8389), .A(n7007), .ZN(n6856) );
  OAI22_X1 U8459 ( .A1(n6854), .A2(n8861), .B1(n7008), .B2(n8863), .ZN(n6855)
         );
  AOI21_X1 U8460 ( .B1(n6856), .B2(n8920), .A(n6855), .ZN(n6857) );
  OAI21_X1 U8461 ( .B1(n9926), .B2(n7609), .A(n6857), .ZN(n9929) );
  NAND2_X1 U8462 ( .A1(n9929), .A2(n8933), .ZN(n6865) );
  INV_X1 U8463 ( .A(n8616), .ZN(n6858) );
  OAI22_X1 U8464 ( .A1(n8933), .A2(n6859), .B1(n6858), .B2(n8844), .ZN(n6863)
         );
  NOR2_X2 U8465 ( .A1(n6971), .A2(n6975), .ZN(n6860) );
  INV_X1 U8466 ( .A(n8615), .ZN(n9927) );
  OR2_X1 U8467 ( .A1(n6860), .A2(n9927), .ZN(n6861) );
  NAND2_X1 U8468 ( .A1(n7027), .A2(n6861), .ZN(n9928) );
  NOR2_X1 U8469 ( .A1(n8850), .A2(n9928), .ZN(n6862) );
  AOI211_X1 U8470 ( .C1(n8926), .C2(n8615), .A(n6863), .B(n6862), .ZN(n6864)
         );
  OAI211_X1 U8471 ( .C1(n9926), .C2(n7619), .A(n6865), .B(n6864), .ZN(P2_U3288) );
  AOI21_X1 U8472 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6874) );
  NAND2_X1 U8473 ( .A1(n8623), .A2(n8707), .ZN(n6869) );
  OAI211_X1 U8474 ( .C1(n8672), .C2(n7111), .A(n6870), .B(n6869), .ZN(n6871)
         );
  AOI21_X1 U8475 ( .B1(n8688), .B2(n7028), .A(n6871), .ZN(n6873) );
  NAND2_X1 U8476 ( .A1(n8680), .A2(n7031), .ZN(n6872) );
  OAI211_X1 U8477 ( .C1(n6874), .C2(n8690), .A(n6873), .B(n6872), .ZN(P2_U3233) );
  INV_X1 U8478 ( .A(n6875), .ZN(n6883) );
  INV_X1 U8479 ( .A(n7677), .ZN(n7341) );
  INV_X1 U8480 ( .A(n9441), .ZN(n8019) );
  AOI22_X1 U8481 ( .A1(n9465), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9474), .ZN(n6878) );
  NAND2_X1 U8482 ( .A1(n8017), .A2(n6876), .ZN(n6877) );
  OAI211_X1 U8483 ( .C1(n8019), .C2(n6879), .A(n6878), .B(n6877), .ZN(n6880)
         );
  AOI21_X1 U8484 ( .B1(n7341), .B2(n6881), .A(n6880), .ZN(n6882) );
  OAI21_X1 U8485 ( .B1(n6883), .B2(n9489), .A(n6882), .ZN(P1_U3289) );
  NAND2_X1 U8486 ( .A1(n6884), .A2(n8441), .ZN(n9894) );
  INV_X1 U8487 ( .A(n9894), .ZN(n6889) );
  AOI22_X1 U8488 ( .A1(n9894), .A2(n8920), .B1(n8917), .B2(n6277), .ZN(n9891)
         );
  OAI22_X1 U8489 ( .A1(n8931), .A2(n9891), .B1(n6885), .B2(n8844), .ZN(n6886)
         );
  AOI21_X1 U8490 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8931), .A(n6886), .ZN(
        n6888) );
  OAI21_X1 U8491 ( .B1(n8926), .B2(n6814), .A(n6283), .ZN(n6887) );
  OAI211_X1 U8492 ( .C1(n6889), .C2(n8924), .A(n6888), .B(n6887), .ZN(P2_U3296) );
  INV_X1 U8493 ( .A(n8303), .ZN(n6891) );
  INV_X1 U8494 ( .A(n8193), .ZN(n6890) );
  NAND2_X1 U8495 ( .A1(n6930), .A2(n6921), .ZN(n8266) );
  INV_X1 U8496 ( .A(n6930), .ZN(n9210) );
  NAND2_X1 U8497 ( .A1(n9210), .A2(n9811), .ZN(n7057) );
  NAND2_X1 U8498 ( .A1(n6912), .A2(n6993), .ZN(n8267) );
  NAND2_X1 U8499 ( .A1(n9209), .A2(n6941), .ZN(n8268) );
  NAND2_X1 U8500 ( .A1(n8267), .A2(n8268), .ZN(n8304) );
  NAND2_X1 U8501 ( .A1(n7236), .A2(n7132), .ZN(n7147) );
  INV_X1 U8502 ( .A(n7236), .ZN(n9208) );
  NAND2_X1 U8503 ( .A1(n9208), .A2(n9818), .ZN(n8269) );
  OR2_X1 U8504 ( .A1(n6892), .A2(n8306), .ZN(n6893) );
  NAND2_X1 U8505 ( .A1(n7148), .A2(n6893), .ZN(n6895) );
  OAI22_X1 U8506 ( .A1(n7184), .A2(n7744), .B1(n6912), .B2(n7630), .ZN(n6894)
         );
  AOI21_X1 U8507 ( .B1(n6895), .B2(n9488), .A(n6894), .ZN(n9822) );
  NAND2_X1 U8508 ( .A1(n6913), .A2(n6896), .ZN(n6897) );
  NAND2_X1 U8509 ( .A1(n6898), .A2(n6897), .ZN(n6909) );
  NAND2_X1 U8510 ( .A1(n8266), .A2(n7057), .ZN(n8302) );
  NAND2_X1 U8511 ( .A1(n6909), .A2(n8302), .ZN(n6911) );
  NAND2_X1 U8512 ( .A1(n6930), .A2(n9811), .ZN(n6899) );
  NAND2_X1 U8513 ( .A1(n6912), .A2(n6941), .ZN(n6900) );
  INV_X1 U8514 ( .A(n8306), .ZN(n6901) );
  NAND2_X1 U8515 ( .A1(n6903), .A2(n8306), .ZN(n6904) );
  AND2_X1 U8516 ( .A1(n7068), .A2(n6904), .ZN(n9820) );
  NAND2_X1 U8517 ( .A1(n6938), .A2(n9818), .ZN(n7153) );
  OAI211_X1 U8518 ( .C1(n6938), .C2(n9818), .A(n9655), .B(n7153), .ZN(n9817)
         );
  INV_X1 U8519 ( .A(n9492), .ZN(n9306) );
  AOI22_X1 U8520 ( .A1(n9465), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7125), .B2(
        n9474), .ZN(n6906) );
  NAND2_X1 U8521 ( .A1(n8017), .A2(n7132), .ZN(n6905) );
  OAI211_X1 U8522 ( .C1(n9817), .C2(n9306), .A(n6906), .B(n6905), .ZN(n6907)
         );
  AOI21_X1 U8523 ( .B1(n9820), .B2(n9456), .A(n6907), .ZN(n6908) );
  OAI21_X1 U8524 ( .B1(n9822), .B2(n9465), .A(n6908), .ZN(P1_U3286) );
  OR2_X1 U8525 ( .A1(n6909), .A2(n8302), .ZN(n6910) );
  NAND2_X1 U8526 ( .A1(n6911), .A2(n6910), .ZN(n9814) );
  OAI22_X1 U8527 ( .A1(n6913), .A2(n7630), .B1(n6912), .B2(n7744), .ZN(n6914)
         );
  AOI21_X1 U8528 ( .B1(n9814), .B2(n7476), .A(n6914), .ZN(n6917) );
  XNOR2_X1 U8529 ( .A(n8264), .B(n8302), .ZN(n6915) );
  NAND2_X1 U8530 ( .A1(n6915), .A2(n9488), .ZN(n6916) );
  AND2_X1 U8531 ( .A1(n6917), .A2(n6916), .ZN(n9816) );
  NAND2_X1 U8532 ( .A1(n6918), .A2(n6921), .ZN(n6919) );
  NAND2_X1 U8533 ( .A1(n6939), .A2(n6919), .ZN(n9812) );
  AOI22_X1 U8534 ( .A1(n9465), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9474), .B2(
        n6920), .ZN(n6923) );
  NAND2_X1 U8535 ( .A1(n8017), .A2(n6921), .ZN(n6922) );
  OAI211_X1 U8536 ( .C1(n8019), .C2(n9812), .A(n6923), .B(n6922), .ZN(n6924)
         );
  AOI21_X1 U8537 ( .B1(n9814), .B2(n7341), .A(n6924), .ZN(n6925) );
  OAI21_X1 U8538 ( .B1(n9816), .B2(n9489), .A(n6925), .ZN(P1_U3288) );
  INV_X1 U8539 ( .A(n6926), .ZN(n7098) );
  OAI222_X1 U8540 ( .A1(n9613), .A2(n7098), .B1(P1_U3084), .B2(n8295), .C1(
        n6927), .C2(n9609), .ZN(P1_U3333) );
  OAI21_X1 U8541 ( .B1(n6929), .B2(n8304), .A(n6928), .ZN(n6936) );
  INV_X1 U8542 ( .A(n6936), .ZN(n6997) );
  OAI22_X1 U8543 ( .A1(n6930), .A2(n7630), .B1(n7236), .B2(n7744), .ZN(n6935)
         );
  NAND2_X1 U8544 ( .A1(n6931), .A2(n8304), .ZN(n6932) );
  AOI21_X1 U8545 ( .B1(n6933), .B2(n6932), .A(n7655), .ZN(n6934) );
  AOI211_X1 U8546 ( .C1(n7476), .C2(n6936), .A(n6935), .B(n6934), .ZN(n6996)
         );
  MUX2_X1 U8547 ( .A(n6937), .B(n6996), .S(n9313), .Z(n6944) );
  AOI21_X1 U8548 ( .B1(n6993), .B2(n6939), .A(n6938), .ZN(n6994) );
  OAI22_X1 U8549 ( .A1(n9477), .A2(n6941), .B1(n6940), .B2(n7669), .ZN(n6942)
         );
  AOI21_X1 U8550 ( .B1(n6994), .B2(n9441), .A(n6942), .ZN(n6943) );
  OAI211_X1 U8551 ( .C1(n6997), .C2(n7677), .A(n6944), .B(n6943), .ZN(P1_U3287) );
  XNOR2_X1 U8552 ( .A(n6946), .B(n6945), .ZN(n6953) );
  INV_X1 U8553 ( .A(n6947), .ZN(n7012) );
  AOI21_X1 U8554 ( .B1(n8682), .B2(n8704), .A(n6948), .ZN(n6950) );
  INV_X1 U8555 ( .A(n7008), .ZN(n8706) );
  NAND2_X1 U8556 ( .A1(n8623), .A2(n8706), .ZN(n6949) );
  OAI211_X1 U8557 ( .C1(n8633), .C2(n7012), .A(n6950), .B(n6949), .ZN(n6951)
         );
  AOI21_X1 U8558 ( .B1(n8688), .B2(n9941), .A(n6951), .ZN(n6952) );
  OAI21_X1 U8559 ( .B1(n6953), .B2(n8690), .A(n6952), .ZN(P2_U3219) );
  INV_X1 U8560 ( .A(n8924), .ZN(n8928) );
  OAI21_X1 U8561 ( .B1(n6956), .B2(n6955), .A(n6954), .ZN(n9910) );
  OAI21_X1 U8562 ( .B1(n6958), .B2(n9905), .A(n6957), .ZN(n9906) );
  OAI22_X1 U8563 ( .A1(n8850), .A2(n9906), .B1(n6959), .B2(n8844), .ZN(n6960)
         );
  AOI21_X1 U8564 ( .B1(n8928), .B2(n9910), .A(n6960), .ZN(n6965) );
  OAI211_X1 U8565 ( .C1(n8384), .C2(n6961), .A(n6831), .B(n8920), .ZN(n6963)
         );
  AOI22_X1 U8566 ( .A1(n8915), .A2(n6534), .B1(n8710), .B2(n8917), .ZN(n6962)
         );
  AND2_X1 U8567 ( .A1(n6963), .A2(n6962), .ZN(n9907) );
  MUX2_X1 U8568 ( .A(n4962), .B(n9907), .S(n8933), .Z(n6964) );
  OAI211_X1 U8569 ( .C1(n9905), .C2(n8908), .A(n6965), .B(n6964), .ZN(P2_U3292) );
  XNOR2_X1 U8570 ( .A(n6966), .B(n8460), .ZN(n9924) );
  INV_X1 U8571 ( .A(n9924), .ZN(n6979) );
  NAND2_X1 U8572 ( .A1(n6967), .A2(n8459), .ZN(n6968) );
  XNOR2_X1 U8573 ( .A(n6968), .B(n8460), .ZN(n6969) );
  OAI222_X1 U8574 ( .A1(n8863), .A2(n7023), .B1(n8861), .B2(n6970), .C1(n6969), 
        .C2(n8859), .ZN(n9922) );
  XNOR2_X1 U8575 ( .A(n6971), .B(n6975), .ZN(n9921) );
  INV_X1 U8576 ( .A(n6972), .ZN(n6973) );
  OAI22_X1 U8577 ( .A1(n8933), .A2(n6366), .B1(n6973), .B2(n8844), .ZN(n6974)
         );
  AOI21_X1 U8578 ( .B1(n8926), .B2(n6975), .A(n6974), .ZN(n6976) );
  OAI21_X1 U8579 ( .B1(n8850), .B2(n9921), .A(n6976), .ZN(n6977) );
  AOI21_X1 U8580 ( .B1(n9922), .B2(n8933), .A(n6977), .ZN(n6978) );
  OAI21_X1 U8581 ( .B1(n6979), .B2(n8924), .A(n6978), .ZN(P2_U3289) );
  NAND2_X1 U8582 ( .A1(n6982), .A2(n8920), .ZN(n6984) );
  AOI22_X1 U8583 ( .A1(n8915), .A2(n6277), .B1(n6534), .B2(n8917), .ZN(n6983)
         );
  AND2_X1 U8584 ( .A1(n6984), .A2(n6983), .ZN(n9901) );
  OAI21_X1 U8585 ( .B1(n6986), .B2(n8383), .A(n6985), .ZN(n9903) );
  AOI22_X1 U8586 ( .A1(n8928), .A2(n9903), .B1(n8926), .B2(n9896), .ZN(n6992)
         );
  AOI21_X1 U8587 ( .B1(n9896), .B2(n6988), .A(n6987), .ZN(n9899) );
  INV_X1 U8588 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6989) );
  OAI22_X1 U8589 ( .A1(n6989), .A2(n8933), .B1(n6477), .B2(n8844), .ZN(n6990)
         );
  AOI21_X1 U8590 ( .B1(n6814), .B2(n9899), .A(n6990), .ZN(n6991) );
  OAI211_X1 U8591 ( .C1(n8931), .C2(n9901), .A(n6992), .B(n6991), .ZN(P2_U3294) );
  AOI22_X1 U8592 ( .A1(n6994), .A2(n9655), .B1(n6993), .B2(n9615), .ZN(n6995)
         );
  OAI211_X1 U8593 ( .C1(n6997), .C2(n9805), .A(n6996), .B(n6995), .ZN(n6999)
         );
  NAND2_X1 U8594 ( .A1(n6999), .A2(n9853), .ZN(n6998) );
  OAI21_X1 U8595 ( .B1(n9853), .B2(n6317), .A(n6998), .ZN(P1_U3527) );
  NAND2_X1 U8596 ( .A1(n6999), .A2(n9850), .ZN(n7000) );
  OAI21_X1 U8597 ( .B1(n9850), .B2(n5679), .A(n7000), .ZN(P1_U3466) );
  NAND2_X1 U8598 ( .A1(n8615), .A2(n8707), .ZN(n7001) );
  NAND2_X1 U8599 ( .A1(n7028), .A2(n7008), .ZN(n8423) );
  OR2_X1 U8600 ( .A1(n7028), .A2(n8706), .ZN(n7004) );
  NAND2_X1 U8601 ( .A1(n8418), .A2(n8417), .ZN(n7108) );
  NAND2_X1 U8602 ( .A1(n7005), .A2(n8391), .ZN(n7006) );
  NAND2_X1 U8603 ( .A1(n7113), .A2(n7006), .ZN(n9940) );
  NAND2_X1 U8604 ( .A1(n7007), .A2(n8465), .ZN(n7022) );
  NAND2_X1 U8605 ( .A1(n7022), .A2(n8390), .ZN(n7021) );
  NAND2_X1 U8606 ( .A1(n7021), .A2(n8423), .ZN(n7109) );
  XNOR2_X1 U8607 ( .A(n7109), .B(n8391), .ZN(n7010) );
  OAI22_X1 U8608 ( .A1(n7008), .A2(n8861), .B1(n7210), .B2(n8863), .ZN(n7009)
         );
  AOI21_X1 U8609 ( .B1(n7010), .B2(n8920), .A(n7009), .ZN(n7011) );
  OAI21_X1 U8610 ( .B1(n9940), .B2(n7609), .A(n7011), .ZN(n9944) );
  NAND2_X1 U8611 ( .A1(n9944), .A2(n8933), .ZN(n7017) );
  OAI22_X1 U8612 ( .A1(n8933), .A2(n6629), .B1(n7012), .B2(n8844), .ZN(n7015)
         );
  AND2_X1 U8613 ( .A1(n7029), .A2(n9941), .ZN(n7013) );
  OR2_X1 U8614 ( .A1(n7013), .A2(n7116), .ZN(n9943) );
  NOR2_X1 U8615 ( .A1(n9943), .A2(n8850), .ZN(n7014) );
  AOI211_X1 U8616 ( .C1(n8926), .C2(n9941), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI211_X1 U8617 ( .C1(n9940), .C2(n7619), .A(n7017), .B(n7016), .ZN(P2_U3286) );
  INV_X1 U8618 ( .A(n7019), .ZN(n7020) );
  AOI21_X1 U8619 ( .B1(n8390), .B2(n7018), .A(n7020), .ZN(n9933) );
  OAI21_X1 U8620 ( .B1(n8390), .B2(n7022), .A(n7021), .ZN(n7025) );
  OAI22_X1 U8621 ( .A1(n7023), .A2(n8861), .B1(n7111), .B2(n8863), .ZN(n7024)
         );
  AOI21_X1 U8622 ( .B1(n7025), .B2(n8920), .A(n7024), .ZN(n7026) );
  OAI21_X1 U8623 ( .B1(n9933), .B2(n7609), .A(n7026), .ZN(n9936) );
  NAND2_X1 U8624 ( .A1(n9936), .A2(n8933), .ZN(n7036) );
  INV_X1 U8625 ( .A(n7027), .ZN(n7030) );
  INV_X1 U8626 ( .A(n7028), .ZN(n9934) );
  OAI21_X1 U8627 ( .B1(n7030), .B2(n9934), .A(n7029), .ZN(n9935) );
  INV_X1 U8628 ( .A(n9935), .ZN(n7034) );
  AOI22_X1 U8629 ( .A1(n8931), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7031), .B2(
        n8929), .ZN(n7032) );
  OAI21_X1 U8630 ( .B1(n9934), .B2(n8908), .A(n7032), .ZN(n7033) );
  AOI21_X1 U8631 ( .B1(n6814), .B2(n7034), .A(n7033), .ZN(n7035) );
  OAI211_X1 U8632 ( .C1(n9933), .C2(n7619), .A(n7036), .B(n7035), .ZN(P2_U3287) );
  INV_X1 U8633 ( .A(n7037), .ZN(n7146) );
  OAI222_X1 U8634 ( .A1(n9060), .A2(n7038), .B1(n9058), .B2(n7146), .C1(n8409), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8635 ( .A(n7087), .ZN(n7082) );
  NOR2_X1 U8636 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7784), .ZN(n7046) );
  INV_X1 U8637 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9981) );
  MUX2_X1 U8638 ( .A(n9981), .B(P2_REG1_REG_12__SCAN_IN), .S(n7087), .Z(n7042)
         );
  INV_X1 U8639 ( .A(n7042), .ZN(n7040) );
  INV_X1 U8640 ( .A(n7041), .ZN(n7043) );
  NAND2_X1 U8641 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  AOI21_X1 U8642 ( .B1(n7086), .B2(n7044), .A(n7977), .ZN(n7045) );
  AOI211_X1 U8643 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n9873), .A(n7046), .B(
        n7045), .ZN(n7055) );
  NOR2_X1 U8644 ( .A1(n7047), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7052) );
  INV_X1 U8645 ( .A(n7052), .ZN(n7049) );
  INV_X1 U8646 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7218) );
  MUX2_X1 U8647 ( .A(n7218), .B(P2_REG2_REG_12__SCAN_IN), .S(n7087), .Z(n7050)
         );
  NOR2_X1 U8648 ( .A1(n7050), .A2(n7051), .ZN(n7048) );
  NAND2_X1 U8649 ( .A1(n7049), .A2(n7048), .ZN(n7081) );
  OAI21_X1 U8650 ( .B1(n7052), .B2(n7051), .A(n7050), .ZN(n7053) );
  NAND3_X1 U8651 ( .A1(n9867), .A2(n7081), .A3(n7053), .ZN(n7054) );
  OAI211_X1 U8652 ( .C1(n9869), .C2(n7082), .A(n7055), .B(n7054), .ZN(P2_U3257) );
  NAND2_X1 U8653 ( .A1(n7298), .A2(n7078), .ZN(n8067) );
  INV_X1 U8654 ( .A(n7298), .ZN(n9206) );
  NAND2_X1 U8655 ( .A1(n9206), .A2(n9830), .ZN(n8263) );
  NAND2_X1 U8656 ( .A1(n8271), .A2(n8269), .ZN(n7056) );
  NAND2_X1 U8657 ( .A1(n7184), .A2(n7157), .ZN(n8073) );
  NAND2_X1 U8658 ( .A1(n7056), .A2(n8073), .ZN(n7060) );
  AND2_X1 U8659 ( .A1(n8268), .A2(n7057), .ZN(n7058) );
  NAND2_X1 U8660 ( .A1(n7063), .A2(n8276), .ZN(n7062) );
  NAND2_X1 U8661 ( .A1(n8073), .A2(n7147), .ZN(n8265) );
  INV_X1 U8662 ( .A(n8267), .ZN(n7059) );
  OR2_X1 U8663 ( .A1(n8265), .A2(n7059), .ZN(n7061) );
  NAND2_X1 U8664 ( .A1(n7062), .A2(n8197), .ZN(n7064) );
  OAI21_X1 U8665 ( .B1(n8075), .B2(n7064), .A(n4399), .ZN(n7066) );
  OAI22_X1 U8666 ( .A1(n7184), .A2(n7630), .B1(n7251), .B2(n7744), .ZN(n7065)
         );
  AOI21_X1 U8667 ( .B1(n7066), .B2(n9488), .A(n7065), .ZN(n9829) );
  NAND2_X1 U8668 ( .A1(n9208), .A2(n7132), .ZN(n7067) );
  NAND2_X1 U8669 ( .A1(n7184), .A2(n9823), .ZN(n7070) );
  OAI21_X1 U8670 ( .B1(n7071), .B2(n8311), .A(n7250), .ZN(n9833) );
  NAND2_X1 U8671 ( .A1(n9833), .A2(n9456), .ZN(n7080) );
  INV_X1 U8672 ( .A(n7072), .ZN(n7183) );
  OAI22_X1 U8673 ( .A1(n9313), .A2(n7073), .B1(n7183), .B2(n7669), .ZN(n7077)
         );
  INV_X1 U8674 ( .A(n7155), .ZN(n7075) );
  INV_X1 U8675 ( .A(n7258), .ZN(n7074) );
  OAI211_X1 U8676 ( .C1(n9830), .C2(n7075), .A(n7074), .B(n9655), .ZN(n9828)
         );
  NOR2_X1 U8677 ( .A1(n9828), .A2(n9306), .ZN(n7076) );
  AOI211_X1 U8678 ( .C1(n8017), .C2(n7078), .A(n7077), .B(n7076), .ZN(n7079)
         );
  OAI211_X1 U8679 ( .C1(n9465), .C2(n9829), .A(n7080), .B(n7079), .ZN(P1_U3284) );
  OAI21_X1 U8680 ( .B1(n7218), .B2(n7082), .A(n7081), .ZN(n7085) );
  INV_X1 U8681 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7083) );
  AOI22_X1 U8682 ( .A1(n7198), .A2(n7083), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7092), .ZN(n7084) );
  NOR2_X1 U8683 ( .A1(n7085), .A2(n7084), .ZN(n7191) );
  AOI21_X1 U8684 ( .B1(n7085), .B2(n7084), .A(n7191), .ZN(n7097) );
  OAI21_X1 U8685 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7087), .A(n7086), .ZN(
        n7089) );
  INV_X1 U8686 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7778) );
  AOI22_X1 U8687 ( .A1(n7198), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7778), .B2(
        n7092), .ZN(n7088) );
  OAI21_X1 U8688 ( .B1(n7089), .B2(n7088), .A(n7197), .ZN(n7095) );
  INV_X1 U8689 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7091) );
  OAI22_X1 U8690 ( .A1(n8745), .A2(n7091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7090), .ZN(n7094) );
  NOR2_X1 U8691 ( .A1(n9869), .A2(n7092), .ZN(n7093) );
  AOI211_X1 U8692 ( .C1(n9868), .C2(n7095), .A(n7094), .B(n7093), .ZN(n7096)
         );
  OAI21_X1 U8693 ( .B1(n7097), .B2(n9871), .A(n7096), .ZN(P2_U3258) );
  OAI222_X1 U8694 ( .A1(P2_U3152), .A2(n4316), .B1(n9058), .B2(n7098), .C1(
        n7854), .C2(n9060), .ZN(P2_U3338) );
  NOR2_X1 U8695 ( .A1(n8931), .A2(n5290), .ZN(n7956) );
  AOI22_X1 U8696 ( .A1(n7956), .A2(n7100), .B1(n7099), .B2(n8929), .ZN(n7101)
         );
  OAI21_X1 U8697 ( .B1(n7102), .B2(n8908), .A(n7101), .ZN(n7103) );
  INV_X1 U8698 ( .A(n7103), .ZN(n7106) );
  MUX2_X1 U8699 ( .A(n6373), .B(n7104), .S(n8933), .Z(n7105) );
  OAI211_X1 U8700 ( .C1(n7107), .C2(n8924), .A(n7106), .B(n7105), .ZN(P2_U3291) );
  OR2_X1 U8701 ( .A1(n7211), .A2(n7210), .ZN(n8478) );
  NAND2_X1 U8702 ( .A1(n7211), .A2(n7210), .ZN(n8483) );
  NAND2_X1 U8703 ( .A1(n8478), .A2(n8483), .ZN(n8394) );
  XOR2_X1 U8704 ( .A(n7207), .B(n8394), .Z(n7110) );
  OAI222_X1 U8705 ( .A1(n8863), .A2(n7443), .B1(n8861), .B2(n7111), .C1(n8859), 
        .C2(n7110), .ZN(n9951) );
  INV_X1 U8706 ( .A(n9951), .ZN(n7124) );
  NAND2_X1 U8707 ( .A1(n9941), .A2(n8705), .ZN(n7112) );
  NAND2_X1 U8708 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  OAI21_X1 U8709 ( .B1(n7114), .B2(n8394), .A(n7213), .ZN(n7115) );
  INV_X1 U8710 ( .A(n7115), .ZN(n9953) );
  INV_X1 U8711 ( .A(n7211), .ZN(n9949) );
  OR2_X1 U8712 ( .A1(n7116), .A2(n9949), .ZN(n7117) );
  NAND2_X1 U8713 ( .A1(n7215), .A2(n7117), .ZN(n9950) );
  INV_X1 U8714 ( .A(n7142), .ZN(n7118) );
  OAI22_X1 U8715 ( .A1(n8933), .A2(n7119), .B1(n7118), .B2(n8844), .ZN(n7120)
         );
  AOI21_X1 U8716 ( .B1(n8926), .B2(n7211), .A(n7120), .ZN(n7121) );
  OAI21_X1 U8717 ( .B1(n9950), .B2(n8850), .A(n7121), .ZN(n7122) );
  AOI21_X1 U8718 ( .B1(n9953), .B2(n8928), .A(n7122), .ZN(n7123) );
  OAI21_X1 U8719 ( .B1(n7124), .B2(n8931), .A(n7123), .ZN(P2_U3285) );
  INV_X1 U8720 ( .A(n7125), .ZN(n7135) );
  XOR2_X1 U8721 ( .A(n7226), .B(n7225), .Z(n7128) );
  INV_X1 U8722 ( .A(n7126), .ZN(n7127) );
  NAND2_X1 U8723 ( .A1(n7128), .A2(n7127), .ZN(n7224) );
  OAI21_X1 U8724 ( .B1(n7128), .B2(n7127), .A(n7224), .ZN(n7129) );
  NAND2_X1 U8725 ( .A1(n7129), .A2(n9173), .ZN(n7134) );
  AOI22_X1 U8726 ( .A1(n9160), .A2(n9209), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3084), .ZN(n7130) );
  OAI21_X1 U8727 ( .B1(n7184), .B2(n9636), .A(n7130), .ZN(n7131) );
  AOI21_X1 U8728 ( .B1(n9192), .B2(n7132), .A(n7131), .ZN(n7133) );
  OAI211_X1 U8729 ( .C1(n9650), .C2(n7135), .A(n7134), .B(n7133), .ZN(P1_U3225) );
  XNOR2_X1 U8730 ( .A(n7137), .B(n7136), .ZN(n7144) );
  NOR2_X1 U8731 ( .A1(n7687), .A2(n9949), .ZN(n7141) );
  NAND2_X1 U8732 ( .A1(n8682), .A2(n8703), .ZN(n7139) );
  NAND2_X1 U8733 ( .A1(n8623), .A2(n8705), .ZN(n7138) );
  OAI211_X1 U8734 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5107), .A(n7139), .B(n7138), .ZN(n7140) );
  AOI211_X1 U8735 ( .C1(n8680), .C2(n7142), .A(n7141), .B(n7140), .ZN(n7143)
         );
  OAI21_X1 U8736 ( .B1(n7144), .B2(n8690), .A(n7143), .ZN(P2_U3238) );
  OAI222_X1 U8737 ( .A1(n9613), .A2(n7146), .B1(P1_U3084), .B2(n8292), .C1(
        n7145), .C2(n9609), .ZN(P1_U3332) );
  NAND2_X1 U8738 ( .A1(n7148), .A2(n7147), .ZN(n8070) );
  XOR2_X1 U8739 ( .A(n8305), .B(n8070), .Z(n7152) );
  OAI21_X1 U8740 ( .B1(n4398), .B2(n7069), .A(n7149), .ZN(n9827) );
  OAI22_X1 U8741 ( .A1(n7298), .A2(n7744), .B1(n7236), .B2(n7630), .ZN(n7150)
         );
  AOI21_X1 U8742 ( .B1(n9827), .B2(n7476), .A(n7150), .ZN(n7151) );
  OAI21_X1 U8743 ( .B1(n7152), .B2(n7655), .A(n7151), .ZN(n9825) );
  INV_X1 U8744 ( .A(n9825), .ZN(n7162) );
  NAND2_X1 U8745 ( .A1(n7153), .A2(n7157), .ZN(n7154) );
  NAND2_X1 U8746 ( .A1(n7155), .A2(n7154), .ZN(n9824) );
  AOI22_X1 U8747 ( .A1(n9489), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7156), .B2(
        n9474), .ZN(n7159) );
  NAND2_X1 U8748 ( .A1(n8017), .A2(n7157), .ZN(n7158) );
  OAI211_X1 U8749 ( .C1(n9824), .C2(n8019), .A(n7159), .B(n7158), .ZN(n7160)
         );
  AOI21_X1 U8750 ( .B1(n9827), .B2(n7341), .A(n7160), .ZN(n7161) );
  OAI21_X1 U8751 ( .B1(n7162), .B2(n9489), .A(n7161), .ZN(P1_U3285) );
  INV_X1 U8752 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7177) );
  INV_X1 U8753 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7163) );
  MUX2_X1 U8754 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7163), .S(n9219), .Z(n7166)
         );
  OAI21_X1 U8755 ( .B1(n7170), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7164), .ZN(
        n7165) );
  NAND2_X1 U8756 ( .A1(n7166), .A2(n7165), .ZN(n9218) );
  OAI21_X1 U8757 ( .B1(n7166), .B2(n7165), .A(n9218), .ZN(n7175) );
  NOR2_X1 U8758 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7167), .ZN(n7641) );
  INV_X1 U8759 ( .A(n7641), .ZN(n7168) );
  OAI21_X1 U8760 ( .B1(n9264), .B2(n9212), .A(n7168), .ZN(n7174) );
  INV_X1 U8761 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7171) );
  NOR2_X1 U8762 ( .A1(n7171), .A2(n7172), .ZN(n9214) );
  AOI211_X1 U8763 ( .C1(n7172), .C2(n7171), .A(n9214), .B(n9763), .ZN(n7173)
         );
  AOI211_X1 U8764 ( .C1(n9786), .C2(n7175), .A(n7174), .B(n7173), .ZN(n7176)
         );
  OAI21_X1 U8765 ( .B1(n9792), .B2(n7177), .A(n7176), .ZN(P1_U3255) );
  XNOR2_X1 U8766 ( .A(n7179), .B(n7178), .ZN(n7180) );
  XNOR2_X1 U8767 ( .A(n7181), .B(n7180), .ZN(n7182) );
  NAND2_X1 U8768 ( .A1(n7182), .A2(n9173), .ZN(n7190) );
  NOR2_X1 U8769 ( .A1(n9650), .A2(n7183), .ZN(n7188) );
  OR2_X1 U8770 ( .A1(n9632), .A2(n7184), .ZN(n7186) );
  NOR2_X1 U8771 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5611), .ZN(n9737) );
  INV_X1 U8772 ( .A(n9737), .ZN(n7185) );
  OAI211_X1 U8773 ( .C1(n9636), .C2(n7251), .A(n7186), .B(n7185), .ZN(n7187)
         );
  NOR2_X1 U8774 ( .A1(n7188), .A2(n7187), .ZN(n7189) );
  OAI211_X1 U8775 ( .C1(n9830), .C2(n9181), .A(n7190), .B(n7189), .ZN(P1_U3211) );
  NOR2_X1 U8776 ( .A1(n7198), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7192) );
  NOR2_X1 U8777 ( .A1(n7192), .A2(n7191), .ZN(n7195) );
  INV_X1 U8778 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7193) );
  AOI22_X1 U8779 ( .A1(n7418), .A2(n7193), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7196), .ZN(n7194) );
  NOR2_X1 U8780 ( .A1(n7195), .A2(n7194), .ZN(n7414) );
  AOI21_X1 U8781 ( .B1(n7195), .B2(n7194), .A(n7414), .ZN(n7206) );
  AOI22_X1 U8782 ( .A1(n7418), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n4421), .B2(
        n7196), .ZN(n7200) );
  OAI21_X1 U8783 ( .B1(n7200), .B2(n7199), .A(n7417), .ZN(n7201) );
  NAND2_X1 U8784 ( .A1(n7201), .A2(n9868), .ZN(n7205) );
  INV_X1 U8785 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8786 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7496) );
  OAI21_X1 U8787 ( .B1(n8745), .B2(n7202), .A(n7496), .ZN(n7203) );
  AOI21_X1 U8788 ( .B1(n8750), .B2(n7418), .A(n7203), .ZN(n7204) );
  OAI211_X1 U8789 ( .C1(n7206), .C2(n9871), .A(n7205), .B(n7204), .ZN(P2_U3259) );
  NAND2_X1 U8790 ( .A1(n7207), .A2(n8483), .ZN(n7208) );
  NAND2_X1 U8791 ( .A1(n7270), .A2(n7443), .ZN(n8484) );
  NAND2_X1 U8792 ( .A1(n4348), .A2(n8484), .ZN(n8395) );
  XOR2_X1 U8793 ( .A(n7436), .B(n8395), .Z(n7209) );
  OAI222_X1 U8794 ( .A1(n8863), .A2(n7430), .B1(n8861), .B2(n7210), .C1(n8859), 
        .C2(n7209), .ZN(n9959) );
  INV_X1 U8795 ( .A(n9959), .ZN(n7223) );
  NAND2_X1 U8796 ( .A1(n7211), .A2(n8704), .ZN(n7212) );
  OAI21_X1 U8797 ( .B1(n7214), .B2(n8395), .A(n7429), .ZN(n9961) );
  OR2_X2 U8798 ( .A1(n7215), .A2(n7270), .ZN(n7449) );
  NAND2_X1 U8799 ( .A1(n7215), .A2(n7270), .ZN(n7216) );
  NAND2_X1 U8800 ( .A1(n7449), .A2(n7216), .ZN(n9958) );
  INV_X1 U8801 ( .A(n7217), .ZN(n7268) );
  OAI22_X1 U8802 ( .A1(n8933), .A2(n7218), .B1(n7268), .B2(n8844), .ZN(n7219)
         );
  AOI21_X1 U8803 ( .B1(n8926), .B2(n7270), .A(n7219), .ZN(n7220) );
  OAI21_X1 U8804 ( .B1(n9958), .B2(n8850), .A(n7220), .ZN(n7221) );
  AOI21_X1 U8805 ( .B1(n9961), .B2(n8928), .A(n7221), .ZN(n7222) );
  OAI21_X1 U8806 ( .B1(n7223), .B2(n8931), .A(n7222), .ZN(P2_U3284) );
  OAI21_X1 U8807 ( .B1(n7226), .B2(n7225), .A(n7224), .ZN(n7230) );
  XNOR2_X1 U8808 ( .A(n7228), .B(n7227), .ZN(n7229) );
  XNOR2_X1 U8809 ( .A(n7230), .B(n7229), .ZN(n7231) );
  NAND2_X1 U8810 ( .A1(n7231), .A2(n9173), .ZN(n7240) );
  NOR2_X1 U8811 ( .A1(n9650), .A2(n7232), .ZN(n7238) );
  OR2_X1 U8812 ( .A1(n9636), .A2(n7298), .ZN(n7235) );
  INV_X1 U8813 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7233) );
  NOR2_X1 U8814 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7233), .ZN(n9730) );
  INV_X1 U8815 ( .A(n9730), .ZN(n7234) );
  OAI211_X1 U8816 ( .C1(n9632), .C2(n7236), .A(n7235), .B(n7234), .ZN(n7237)
         );
  NOR2_X1 U8817 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  OAI211_X1 U8818 ( .C1(n9823), .C2(n9181), .A(n7240), .B(n7239), .ZN(P1_U3237) );
  INV_X1 U8819 ( .A(n7241), .ZN(n8020) );
  OAI222_X1 U8820 ( .A1(n9609), .A2(n7242), .B1(n9613), .B2(n8020), .C1(n6129), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U8821 ( .A1(n7245), .A2(n7552), .ZN(n7243) );
  OAI211_X1 U8822 ( .C1(n7244), .C2(n9060), .A(n7243), .B(n8590), .ZN(P2_U3335) );
  NAND2_X1 U8823 ( .A1(n7245), .A2(n7556), .ZN(n7247) );
  NAND2_X1 U8824 ( .A1(n7246), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8352) );
  OAI211_X1 U8825 ( .C1(n7248), .C2(n9609), .A(n7247), .B(n8352), .ZN(P1_U3330) );
  NAND2_X1 U8826 ( .A1(n7298), .A2(n9830), .ZN(n7249) );
  NAND2_X1 U8827 ( .A1(n7251), .A2(n7275), .ZN(n8080) );
  NAND2_X1 U8828 ( .A1(n9835), .A2(n9205), .ZN(n8218) );
  NAND2_X1 U8829 ( .A1(n7274), .A2(n8308), .ZN(n7252) );
  NAND2_X1 U8830 ( .A1(n7326), .A2(n7252), .ZN(n9834) );
  XNOR2_X1 U8831 ( .A(n7280), .B(n8308), .ZN(n7254) );
  INV_X1 U8832 ( .A(n9204), .ZN(n7391) );
  OAI22_X1 U8833 ( .A1(n7391), .A2(n7744), .B1(n7298), .B2(n7630), .ZN(n7253)
         );
  AOI21_X1 U8834 ( .B1(n7254), .B2(n9488), .A(n7253), .ZN(n7255) );
  OAI21_X1 U8835 ( .B1(n9834), .B2(n9498), .A(n7255), .ZN(n9837) );
  NAND2_X1 U8836 ( .A1(n9837), .A2(n9313), .ZN(n7263) );
  INV_X1 U8837 ( .A(n7256), .ZN(n7297) );
  OAI22_X1 U8838 ( .A1(n9313), .A2(n7257), .B1(n7297), .B2(n7669), .ZN(n7261)
         );
  NOR2_X1 U8839 ( .A1(n7258), .A2(n9835), .ZN(n7259) );
  OR2_X1 U8840 ( .A1(n7335), .A2(n7259), .ZN(n9836) );
  NOR2_X1 U8841 ( .A1(n9836), .A2(n8019), .ZN(n7260) );
  AOI211_X1 U8842 ( .C1(n8017), .C2(n7275), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI211_X1 U8843 ( .C1(n9834), .C2(n7677), .A(n7263), .B(n7262), .ZN(P1_U3283) );
  XNOR2_X1 U8844 ( .A(n7264), .B(n7265), .ZN(n7272) );
  AOI22_X1 U8845 ( .A1(n8682), .A2(n8702), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7267) );
  NAND2_X1 U8846 ( .A1(n8623), .A2(n8704), .ZN(n7266) );
  OAI211_X1 U8847 ( .C1(n8633), .C2(n7268), .A(n7267), .B(n7266), .ZN(n7269)
         );
  AOI21_X1 U8848 ( .B1(n8688), .B2(n7270), .A(n7269), .ZN(n7271) );
  OAI21_X1 U8849 ( .B1(n7272), .B2(n8690), .A(n7271), .ZN(P2_U3226) );
  OR2_X1 U8850 ( .A1(n8308), .A2(n4380), .ZN(n7273) );
  NOR2_X1 U8851 ( .A1(n7274), .A2(n7273), .ZN(n7278) );
  NAND2_X1 U8852 ( .A1(n9205), .A2(n7275), .ZN(n7325) );
  AND2_X1 U8853 ( .A1(n4858), .A2(n7325), .ZN(n7276) );
  NOR2_X1 U8854 ( .A1(n4380), .A2(n7276), .ZN(n7277) );
  NAND2_X1 U8855 ( .A1(n9616), .A2(n7378), .ZN(n8085) );
  NAND2_X1 U8856 ( .A1(n8204), .A2(n8085), .ZN(n7307) );
  NOR2_X1 U8857 ( .A1(n9616), .A2(n9203), .ZN(n7279) );
  OR2_X1 U8858 ( .A1(n9582), .A2(n9202), .ZN(n7470) );
  NAND2_X1 U8859 ( .A1(n9582), .A2(n9202), .ZN(n7472) );
  AND2_X1 U8860 ( .A1(n7470), .A2(n7472), .ZN(n8078) );
  XNOR2_X1 U8861 ( .A(n7471), .B(n8078), .ZN(n9584) );
  NAND2_X1 U8862 ( .A1(n7280), .A2(n8218), .ZN(n7281) );
  NAND2_X1 U8863 ( .A1(n7281), .A2(n8080), .ZN(n7328) );
  OR2_X1 U8864 ( .A1(n7391), .A2(n7337), .ZN(n8082) );
  NAND2_X1 U8865 ( .A1(n7337), .A2(n7391), .ZN(n8081) );
  NAND2_X1 U8866 ( .A1(n8082), .A2(n8081), .ZN(n8310) );
  OR2_X1 U8867 ( .A1(n8310), .A2(n7307), .ZN(n7282) );
  OR2_X1 U8868 ( .A1(n7307), .A2(n8082), .ZN(n7283) );
  AND2_X2 U8869 ( .A1(n7284), .A2(n7283), .ZN(n7308) );
  INV_X1 U8870 ( .A(n8078), .ZN(n8313) );
  XNOR2_X1 U8871 ( .A(n7474), .B(n8313), .ZN(n7285) );
  OAI222_X1 U8872 ( .A1(n7744), .A2(n7570), .B1(n7630), .B2(n7378), .C1(n7285), 
        .C2(n7655), .ZN(n9580) );
  INV_X1 U8873 ( .A(n9582), .ZN(n7413) );
  INV_X1 U8874 ( .A(n7337), .ZN(n9842) );
  INV_X1 U8875 ( .A(n7481), .ZN(n7287) );
  AOI211_X1 U8876 ( .C1(n9582), .C2(n7313), .A(n9843), .B(n7287), .ZN(n9581)
         );
  NAND2_X1 U8877 ( .A1(n9581), .A2(n9492), .ZN(n7289) );
  AOI22_X1 U8878 ( .A1(n9489), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7410), .B2(
        n9474), .ZN(n7288) );
  OAI211_X1 U8879 ( .C1(n7413), .C2(n9477), .A(n7289), .B(n7288), .ZN(n7290)
         );
  AOI21_X1 U8880 ( .B1(n9580), .B2(n9313), .A(n7290), .ZN(n7291) );
  OAI21_X1 U8881 ( .B1(n9584), .B2(n9494), .A(n7291), .ZN(P1_U3280) );
  XNOR2_X1 U8882 ( .A(n7293), .B(n7292), .ZN(n7294) );
  XNOR2_X1 U8883 ( .A(n7295), .B(n7294), .ZN(n7296) );
  NAND2_X1 U8884 ( .A1(n7296), .A2(n9173), .ZN(n7305) );
  NOR2_X1 U8885 ( .A1(n9650), .A2(n7297), .ZN(n7303) );
  OR2_X1 U8886 ( .A1(n9632), .A2(n7298), .ZN(n7301) );
  INV_X1 U8887 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7299) );
  NOR2_X1 U8888 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7299), .ZN(n9755) );
  INV_X1 U8889 ( .A(n9755), .ZN(n7300) );
  OAI211_X1 U8890 ( .C1(n9636), .C2(n7391), .A(n7301), .B(n7300), .ZN(n7302)
         );
  NOR2_X1 U8891 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  OAI211_X1 U8892 ( .C1(n9835), .C2(n9181), .A(n7305), .B(n7304), .ZN(P1_U3219) );
  XNOR2_X1 U8893 ( .A(n7306), .B(n7307), .ZN(n9620) );
  OR2_X1 U8894 ( .A1(n7328), .A2(n8310), .ZN(n7329) );
  NAND2_X1 U8895 ( .A1(n7329), .A2(n8082), .ZN(n7309) );
  INV_X1 U8896 ( .A(n7307), .ZN(n8314) );
  OAI211_X1 U8897 ( .C1(n7309), .C2(n8314), .A(n7308), .B(n9488), .ZN(n7311)
         );
  AOI22_X1 U8898 ( .A1(n9483), .A2(n9204), .B1(n9202), .B2(n9485), .ZN(n7310)
         );
  NAND2_X1 U8899 ( .A1(n7311), .A2(n7310), .ZN(n7312) );
  AOI21_X1 U8900 ( .B1(n9620), .B2(n7476), .A(n7312), .ZN(n9622) );
  AOI21_X1 U8901 ( .B1(n4397), .B2(n9616), .A(n9843), .ZN(n7314) );
  NAND2_X1 U8902 ( .A1(n7314), .A2(n7313), .ZN(n9618) );
  AOI22_X1 U8903 ( .A1(n9489), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7389), .B2(
        n9474), .ZN(n7316) );
  NAND2_X1 U8904 ( .A1(n9616), .A2(n8017), .ZN(n7315) );
  OAI211_X1 U8905 ( .C1(n9618), .C2(n9306), .A(n7316), .B(n7315), .ZN(n7317)
         );
  AOI21_X1 U8906 ( .B1(n9620), .B2(n7341), .A(n7317), .ZN(n7318) );
  OAI21_X1 U8907 ( .B1(n9622), .B2(n9489), .A(n7318), .ZN(P1_U3281) );
  INV_X1 U8908 ( .A(n7319), .ZN(n7323) );
  OAI222_X1 U8909 ( .A1(n9613), .A2(n7323), .B1(P1_U3084), .B2(n7321), .C1(
        n7320), .C2(n9609), .ZN(P1_U3329) );
  OAI222_X1 U8910 ( .A1(n7324), .A2(P2_U3152), .B1(n9058), .B2(n7323), .C1(
        n7322), .C2(n9060), .ZN(P2_U3334) );
  NAND2_X1 U8911 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
  XNOR2_X1 U8912 ( .A(n7327), .B(n8310), .ZN(n7334) );
  AOI22_X1 U8913 ( .A1(n9483), .A2(n9205), .B1(n9203), .B2(n9485), .ZN(n7333)
         );
  INV_X1 U8914 ( .A(n7328), .ZN(n7331) );
  INV_X1 U8915 ( .A(n8310), .ZN(n7330) );
  OAI211_X1 U8916 ( .C1(n7331), .C2(n7330), .A(n7329), .B(n9488), .ZN(n7332)
         );
  OAI211_X1 U8917 ( .C1(n7334), .C2(n9498), .A(n7333), .B(n7332), .ZN(n9845)
         );
  INV_X1 U8918 ( .A(n9845), .ZN(n7343) );
  INV_X1 U8919 ( .A(n7334), .ZN(n9847) );
  OR2_X1 U8920 ( .A1(n7335), .A2(n9842), .ZN(n7336) );
  NAND2_X1 U8921 ( .A1(n4397), .A2(n7336), .ZN(n9844) );
  AOI22_X1 U8922 ( .A1(n9489), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7380), .B2(
        n9474), .ZN(n7339) );
  NAND2_X1 U8923 ( .A1(n8017), .A2(n7337), .ZN(n7338) );
  OAI211_X1 U8924 ( .C1(n9844), .C2(n8019), .A(n7339), .B(n7338), .ZN(n7340)
         );
  AOI21_X1 U8925 ( .B1(n9847), .B2(n7341), .A(n7340), .ZN(n7342) );
  OAI21_X1 U8926 ( .B1(n7343), .B2(n9489), .A(n7342), .ZN(P1_U3282) );
  INV_X1 U8927 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U8928 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7344) );
  AOI21_X1 U8929 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n7344), .ZN(n9990) );
  NOR2_X1 U8930 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7345) );
  AOI21_X1 U8931 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7345), .ZN(n9993) );
  NOR2_X1 U8932 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7346) );
  AOI21_X1 U8933 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7346), .ZN(n9996) );
  NOR2_X1 U8934 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7347) );
  AOI21_X1 U8935 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7347), .ZN(n9999) );
  NOR2_X1 U8936 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7348) );
  AOI21_X1 U8937 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7348), .ZN(n10002) );
  AOI22_X1 U8938 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9725), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n7918), .ZN(n10031) );
  NAND2_X1 U8939 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7354) );
  XOR2_X1 U8940 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10029) );
  NAND2_X1 U8941 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7352) );
  AOI22_X1 U8942 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n7349), .B2(n7867), .ZN(n10027) );
  AOI21_X1 U8943 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9984) );
  NAND3_X1 U8944 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9986) );
  OAI21_X1 U8945 ( .B1(n9984), .B2(n7350), .A(n9986), .ZN(n10026) );
  NAND2_X1 U8946 ( .A1(n10027), .A2(n10026), .ZN(n7351) );
  NAND2_X1 U8947 ( .A1(n7352), .A2(n7351), .ZN(n10028) );
  NAND2_X1 U8948 ( .A1(n10029), .A2(n10028), .ZN(n7353) );
  NAND2_X1 U8949 ( .A1(n7354), .A2(n7353), .ZN(n10030) );
  NOR2_X1 U8950 ( .A1(n10031), .A2(n10030), .ZN(n7355) );
  AOI21_X1 U8951 ( .B1(n7918), .B2(n9725), .A(n7355), .ZN(n7356) );
  NOR2_X1 U8952 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7356), .ZN(n10015) );
  AND2_X1 U8953 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7356), .ZN(n10014) );
  NOR2_X1 U8954 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10014), .ZN(n7357) );
  NAND2_X1 U8955 ( .A1(n7358), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7360) );
  XOR2_X1 U8956 ( .A(n7358), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10013) );
  NAND2_X1 U8957 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10013), .ZN(n7359) );
  NAND2_X1 U8958 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  NAND2_X1 U8959 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7361), .ZN(n7363) );
  XOR2_X1 U8960 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7361), .Z(n10025) );
  NAND2_X1 U8961 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10025), .ZN(n7362) );
  NAND2_X1 U8962 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  NAND2_X1 U8963 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7364), .ZN(n7366) );
  XOR2_X1 U8964 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7364), .Z(n10024) );
  NAND2_X1 U8965 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10024), .ZN(n7365) );
  NAND2_X1 U8966 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  AND2_X1 U8967 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7367), .ZN(n7368) );
  INV_X1 U8968 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10023) );
  XNOR2_X1 U8969 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7367), .ZN(n10022) );
  NOR2_X1 U8970 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  NAND2_X1 U8971 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7369) );
  OAI21_X1 U8972 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7369), .ZN(n10010) );
  NAND2_X1 U8973 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7370) );
  OAI21_X1 U8974 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7370), .ZN(n10007) );
  NOR2_X1 U8975 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7371) );
  AOI21_X1 U8976 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7371), .ZN(n10004) );
  NAND2_X1 U8977 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  NAND2_X1 U8978 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  NAND2_X1 U8979 ( .A1(n9999), .A2(n9998), .ZN(n9997) );
  OAI21_X1 U8980 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9997), .ZN(n9995) );
  NAND2_X1 U8981 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OAI21_X1 U8982 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9994), .ZN(n9992) );
  NAND2_X1 U8983 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  OAI21_X1 U8984 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9991), .ZN(n9989) );
  NAND2_X1 U8985 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  NOR2_X1 U8986 ( .A1(n10019), .A2(n10018), .ZN(n7372) );
  NAND2_X1 U8987 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  OAI21_X1 U8988 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7372), .A(n10017), .ZN(
        n7374) );
  XNOR2_X1 U8989 ( .A(n4413), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7373) );
  XNOR2_X1 U8990 ( .A(n7374), .B(n7373), .ZN(ADD_1071_U4) );
  NAND2_X1 U8991 ( .A1(n7400), .A2(n7375), .ZN(n7384) );
  OAI21_X1 U8992 ( .B1(n7375), .B2(n7400), .A(n7384), .ZN(n7376) );
  NAND2_X1 U8993 ( .A1(n7376), .A2(n9173), .ZN(n7382) );
  AND2_X1 U8994 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9768) );
  AOI21_X1 U8995 ( .B1(n9160), .B2(n9205), .A(n9768), .ZN(n7377) );
  OAI21_X1 U8996 ( .B1(n7378), .B2(n9636), .A(n7377), .ZN(n7379) );
  AOI21_X1 U8997 ( .B1(n7380), .B2(n9164), .A(n7379), .ZN(n7381) );
  OAI211_X1 U8998 ( .C1(n9842), .C2(n9181), .A(n7382), .B(n7381), .ZN(P1_U3229) );
  NAND2_X1 U8999 ( .A1(n7384), .A2(n7383), .ZN(n7388) );
  NAND2_X1 U9000 ( .A1(n7386), .A2(n7385), .ZN(n7387) );
  XNOR2_X1 U9001 ( .A(n7388), .B(n7387), .ZN(n7398) );
  INV_X1 U9002 ( .A(n7389), .ZN(n7390) );
  NOR2_X1 U9003 ( .A1(n9650), .A2(n7390), .ZN(n7395) );
  INV_X1 U9004 ( .A(n9202), .ZN(n7475) );
  OR2_X1 U9005 ( .A1(n7391), .A2(n9632), .ZN(n7393) );
  OAI211_X1 U9006 ( .C1(n9636), .C2(n7475), .A(n7393), .B(n7392), .ZN(n7394)
         );
  NOR2_X1 U9007 ( .A1(n7395), .A2(n7394), .ZN(n7397) );
  NAND2_X1 U9008 ( .A1(n9616), .A2(n9192), .ZN(n7396) );
  OAI211_X1 U9009 ( .C1(n7398), .C2(n9642), .A(n7397), .B(n7396), .ZN(P1_U3215) );
  NAND2_X1 U9010 ( .A1(n7400), .A2(n7399), .ZN(n7405) );
  NAND2_X1 U9011 ( .A1(n7405), .A2(n7401), .ZN(n7403) );
  AOI21_X1 U9012 ( .B1(n7403), .B2(n7402), .A(n9642), .ZN(n7407) );
  NAND2_X1 U9013 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  NAND2_X1 U9014 ( .A1(n7407), .A2(n7406), .ZN(n7412) );
  AND2_X1 U9015 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9776) );
  AOI21_X1 U9016 ( .B1(n9160), .B2(n9203), .A(n9776), .ZN(n7408) );
  OAI21_X1 U9017 ( .B1(n7570), .B2(n9636), .A(n7408), .ZN(n7409) );
  AOI21_X1 U9018 ( .B1(n7410), .B2(n9164), .A(n7409), .ZN(n7411) );
  OAI211_X1 U9019 ( .C1(n7413), .C2(n9181), .A(n7412), .B(n7411), .ZN(P1_U3234) );
  NOR2_X1 U9020 ( .A1(n7418), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7415) );
  NOR2_X1 U9021 ( .A1(n7415), .A2(n7414), .ZN(n7959) );
  XNOR2_X1 U9022 ( .A(n7959), .B(n7960), .ZN(n7416) );
  NOR2_X1 U9023 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7416), .ZN(n7961) );
  AOI21_X1 U9024 ( .B1(n7416), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7961), .ZN(
        n7427) );
  XNOR2_X1 U9025 ( .A(n7970), .B(n7971), .ZN(n7419) );
  INV_X1 U9026 ( .A(n7419), .ZN(n7422) );
  INV_X1 U9027 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7420) );
  NOR2_X1 U9028 ( .A1(n7420), .A2(n7419), .ZN(n7972) );
  INV_X1 U9029 ( .A(n7972), .ZN(n7421) );
  OAI211_X1 U9030 ( .C1(n7422), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9868), .B(
        n7421), .ZN(n7426) );
  AND2_X1 U9031 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7424) );
  NOR2_X1 U9032 ( .A1(n9869), .A2(n7971), .ZN(n7423) );
  AOI211_X1 U9033 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9873), .A(n7424), .B(
        n7423), .ZN(n7425) );
  OAI211_X1 U9034 ( .C1(n7427), .C2(n9871), .A(n7426), .B(n7425), .ZN(P2_U3260) );
  NAND2_X1 U9035 ( .A1(n9020), .A2(n7600), .ZN(n8493) );
  NAND2_X1 U9036 ( .A1(n8494), .A2(n8493), .ZN(n7510) );
  NAND2_X1 U9037 ( .A1(n9956), .A2(n7443), .ZN(n7428) );
  OR2_X1 U9038 ( .A1(n9025), .A2(n7430), .ZN(n8487) );
  NAND2_X1 U9039 ( .A1(n9025), .A2(n7430), .ZN(n8480) );
  NAND2_X1 U9040 ( .A1(n9025), .A2(n8702), .ZN(n7431) );
  INV_X1 U9041 ( .A(n7504), .ZN(n7432) );
  AOI21_X1 U9042 ( .B1(n8498), .B2(n7433), .A(n7432), .ZN(n9024) );
  INV_X1 U9043 ( .A(n7448), .ZN(n7434) );
  INV_X1 U9044 ( .A(n9020), .ZN(n7497) );
  AOI21_X1 U9045 ( .B1(n9020), .B2(n7434), .A(n7505), .ZN(n9021) );
  AOI22_X1 U9046 ( .A1(n8931), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7500), .B2(
        n8929), .ZN(n7435) );
  OAI21_X1 U9047 ( .B1(n7497), .B2(n8908), .A(n7435), .ZN(n7439) );
  XNOR2_X1 U9048 ( .A(n7511), .B(n8498), .ZN(n7437) );
  AOI222_X1 U9049 ( .A1(n8920), .A2(n7437), .B1(n8700), .B2(n8917), .C1(n8702), 
        .C2(n8915), .ZN(n9023) );
  NOR2_X1 U9050 ( .A1(n9023), .A2(n8931), .ZN(n7438) );
  AOI211_X1 U9051 ( .C1(n9021), .C2(n6814), .A(n7439), .B(n7438), .ZN(n7440)
         );
  OAI21_X1 U9052 ( .B1(n9024), .B2(n8924), .A(n7440), .ZN(P2_U3282) );
  OAI21_X1 U9053 ( .B1(n8489), .B2(n7442), .A(n7441), .ZN(n7447) );
  OAI22_X1 U9054 ( .A1(n7443), .A2(n8861), .B1(n7600), .B2(n8863), .ZN(n7446)
         );
  OAI21_X1 U9055 ( .B1(n4393), .B2(n8396), .A(n7444), .ZN(n9029) );
  NOR2_X1 U9056 ( .A1(n9029), .A2(n7609), .ZN(n7445) );
  AOI211_X1 U9057 ( .C1(n8920), .C2(n7447), .A(n7446), .B(n7445), .ZN(n9028)
         );
  AOI21_X1 U9058 ( .B1(n9025), .B2(n7449), .A(n7448), .ZN(n9026) );
  INV_X1 U9059 ( .A(n9025), .ZN(n7451) );
  AOI22_X1 U9060 ( .A1(n8931), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7534), .B2(
        n8929), .ZN(n7450) );
  OAI21_X1 U9061 ( .B1(n7451), .B2(n8908), .A(n7450), .ZN(n7453) );
  NOR2_X1 U9062 ( .A1(n9029), .A2(n7619), .ZN(n7452) );
  AOI211_X1 U9063 ( .C1(n9026), .C2(n6814), .A(n7453), .B(n7452), .ZN(n7454)
         );
  OAI21_X1 U9064 ( .B1(n9028), .B2(n8931), .A(n7454), .ZN(P2_U3283) );
  XNOR2_X1 U9065 ( .A(n7457), .B(n7456), .ZN(n7458) );
  XNOR2_X1 U9066 ( .A(n7455), .B(n7458), .ZN(n7463) );
  AOI22_X1 U9067 ( .A1(n9188), .A2(n9200), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7460) );
  NAND2_X1 U9068 ( .A1(n9164), .A2(n7484), .ZN(n7459) );
  OAI211_X1 U9069 ( .C1(n7475), .C2(n9632), .A(n7460), .B(n7459), .ZN(n7461)
         );
  AOI21_X1 U9070 ( .B1(n9574), .B2(n9192), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9071 ( .B1(n7463), .B2(n9642), .A(n7462), .ZN(P1_U3222) );
  INV_X1 U9072 ( .A(n7464), .ZN(n7468) );
  OAI222_X1 U9073 ( .A1(n9060), .A2(n7466), .B1(n9058), .B2(n7468), .C1(n7465), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9074 ( .A1(n9609), .A2(n7469), .B1(n9613), .B2(n7468), .C1(n7467), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U9075 ( .A1(n7471), .A2(n7470), .ZN(n7473) );
  NAND2_X1 U9076 ( .A1(n7473), .A2(n7472), .ZN(n7526) );
  OR2_X1 U9077 ( .A1(n9574), .A2(n7570), .ZN(n8095) );
  NAND2_X1 U9078 ( .A1(n9574), .A2(n7570), .ZN(n8100) );
  NAND2_X1 U9079 ( .A1(n8095), .A2(n8100), .ZN(n7525) );
  XNOR2_X1 U9080 ( .A(n7526), .B(n8315), .ZN(n7477) );
  INV_X1 U9081 ( .A(n7477), .ZN(n9577) );
  NAND2_X1 U9082 ( .A1(n9582), .A2(n7475), .ZN(n8099) );
  OR2_X1 U9083 ( .A1(n9582), .A2(n7475), .ZN(n8094) );
  XNOR2_X1 U9084 ( .A(n7519), .B(n8315), .ZN(n7480) );
  NAND2_X1 U9085 ( .A1(n7477), .A2(n7476), .ZN(n7479) );
  AOI22_X1 U9086 ( .A1(n9483), .A2(n9202), .B1(n9200), .B2(n9485), .ZN(n7478)
         );
  OAI211_X1 U9087 ( .C1(n7655), .C2(n7480), .A(n7479), .B(n7478), .ZN(n9579)
         );
  NAND2_X1 U9088 ( .A1(n9579), .A2(n9313), .ZN(n7490) );
  INV_X1 U9089 ( .A(n7529), .ZN(n7483) );
  AOI21_X1 U9090 ( .B1(n7481), .B2(n9574), .A(n9843), .ZN(n7482) );
  NAND2_X1 U9091 ( .A1(n7483), .A2(n7482), .ZN(n9575) );
  INV_X1 U9092 ( .A(n9575), .ZN(n7488) );
  INV_X1 U9093 ( .A(n9574), .ZN(n7486) );
  AOI22_X1 U9094 ( .A1(n9489), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7484), .B2(
        n9474), .ZN(n7485) );
  OAI21_X1 U9095 ( .B1(n7486), .B2(n9477), .A(n7485), .ZN(n7487) );
  AOI21_X1 U9096 ( .B1(n7488), .B2(n9492), .A(n7487), .ZN(n7489) );
  OAI211_X1 U9097 ( .C1(n9577), .C2(n7677), .A(n7490), .B(n7489), .ZN(P1_U3279) );
  INV_X1 U9098 ( .A(n7491), .ZN(n7492) );
  AOI21_X1 U9099 ( .B1(n7494), .B2(n7493), .A(n7492), .ZN(n7502) );
  NAND2_X1 U9100 ( .A1(n8623), .A2(n8702), .ZN(n7495) );
  OAI211_X1 U9101 ( .C1(n8672), .C2(n8499), .A(n7496), .B(n7495), .ZN(n7499)
         );
  NOR2_X1 U9102 ( .A1(n7497), .A2(n7687), .ZN(n7498) );
  AOI211_X1 U9103 ( .C1(n8680), .C2(n7500), .A(n7499), .B(n7498), .ZN(n7501)
         );
  OAI21_X1 U9104 ( .B1(n7502), .B2(n8690), .A(n7501), .ZN(P2_U3217) );
  INV_X1 U9105 ( .A(n7600), .ZN(n8701) );
  OR2_X1 U9106 ( .A1(n9020), .A2(n8701), .ZN(n7503) );
  XNOR2_X1 U9107 ( .A(n9015), .B(n8700), .ZN(n8397) );
  XNOR2_X1 U9108 ( .A(n7576), .B(n8397), .ZN(n9019) );
  INV_X1 U9109 ( .A(n7505), .ZN(n7507) );
  INV_X1 U9110 ( .A(n9015), .ZN(n7509) );
  NAND2_X1 U9111 ( .A1(n7505), .A2(n7509), .ZN(n7616) );
  INV_X1 U9112 ( .A(n7616), .ZN(n7506) );
  AOI21_X1 U9113 ( .B1(n9015), .B2(n7507), .A(n7506), .ZN(n9016) );
  AOI22_X1 U9114 ( .A1(n8931), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7597), .B2(
        n8929), .ZN(n7508) );
  OAI21_X1 U9115 ( .B1(n7509), .B2(n8908), .A(n7508), .ZN(n7514) );
  INV_X1 U9116 ( .A(n8397), .ZN(n8503) );
  XNOR2_X1 U9117 ( .A(n7581), .B(n8503), .ZN(n7512) );
  INV_X1 U9118 ( .A(n8646), .ZN(n8699) );
  AOI222_X1 U9119 ( .A1(n8920), .A2(n7512), .B1(n8699), .B2(n8917), .C1(n8701), 
        .C2(n8915), .ZN(n9018) );
  NOR2_X1 U9120 ( .A1(n9018), .A2(n8931), .ZN(n7513) );
  AOI211_X1 U9121 ( .C1(n9016), .C2(n6814), .A(n7514), .B(n7513), .ZN(n7515)
         );
  OAI21_X1 U9122 ( .B1(n8924), .B2(n9019), .A(n7515), .ZN(P2_U3281) );
  INV_X1 U9123 ( .A(n7516), .ZN(n7545) );
  OAI222_X1 U9124 ( .A1(n9613), .A2(n7545), .B1(P1_U3084), .B2(n7518), .C1(
        n7517), .C2(n9609), .ZN(P1_U3327) );
  INV_X1 U9125 ( .A(n7522), .ZN(n7520) );
  INV_X1 U9126 ( .A(n8095), .ZN(n8101) );
  INV_X1 U9127 ( .A(n9200), .ZN(n7644) );
  OR2_X1 U9128 ( .A1(n7622), .A2(n7644), .ZN(n8093) );
  NAND2_X1 U9129 ( .A1(n7622), .A2(n7644), .ZN(n8065) );
  NAND2_X1 U9130 ( .A1(n8093), .A2(n8065), .ZN(n8317) );
  OAI21_X1 U9131 ( .B1(n7520), .B2(n8101), .A(n8317), .ZN(n7523) );
  NOR2_X1 U9132 ( .A1(n8317), .A2(n8101), .ZN(n7521) );
  NAND2_X1 U9133 ( .A1(n7522), .A2(n7521), .ZN(n7625) );
  NAND2_X1 U9134 ( .A1(n7523), .A2(n7625), .ZN(n7524) );
  AOI222_X1 U9135 ( .A1(n9488), .A2(n7524), .B1(n9199), .B2(n9485), .C1(n9201), 
        .C2(n9483), .ZN(n9672) );
  NAND2_X1 U9136 ( .A1(n9574), .A2(n9201), .ZN(n7527) );
  XOR2_X1 U9137 ( .A(n7624), .B(n8317), .Z(n9675) );
  NAND2_X1 U9138 ( .A1(n9675), .A2(n9456), .ZN(n7533) );
  INV_X1 U9139 ( .A(n7572), .ZN(n7528) );
  OAI22_X1 U9140 ( .A1(n9313), .A2(n6775), .B1(n7528), .B2(n7669), .ZN(n7531)
         );
  NAND2_X1 U9141 ( .A1(n7529), .A2(n9673), .ZN(n7649) );
  OAI211_X1 U9142 ( .C1(n7529), .C2(n9673), .A(n7649), .B(n9655), .ZN(n9671)
         );
  NOR2_X1 U9143 ( .A1(n9671), .A2(n9306), .ZN(n7530) );
  AOI211_X1 U9144 ( .C1(n8017), .C2(n7622), .A(n7531), .B(n7530), .ZN(n7532)
         );
  OAI211_X1 U9145 ( .C1(n9465), .C2(n9672), .A(n7533), .B(n7532), .ZN(P1_U3278) );
  INV_X1 U9146 ( .A(n7534), .ZN(n7538) );
  NOR2_X1 U9147 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7090), .ZN(n7535) );
  AOI21_X1 U9148 ( .B1(n8682), .B2(n8701), .A(n7535), .ZN(n7537) );
  NAND2_X1 U9149 ( .A1(n8623), .A2(n8703), .ZN(n7536) );
  OAI211_X1 U9150 ( .C1(n8633), .C2(n7538), .A(n7537), .B(n7536), .ZN(n7543)
         );
  XNOR2_X1 U9151 ( .A(n7539), .B(n7540), .ZN(n7541) );
  NOR2_X1 U9152 ( .A1(n7541), .A2(n8690), .ZN(n7542) );
  AOI211_X1 U9153 ( .C1(n8688), .C2(n9025), .A(n7543), .B(n7542), .ZN(n7544)
         );
  INV_X1 U9154 ( .A(n7544), .ZN(P2_U3236) );
  OAI222_X1 U9155 ( .A1(n7546), .A2(P2_U3152), .B1(n9058), .B2(n7545), .C1(
        n7762), .C2(n9060), .ZN(P2_U3332) );
  INV_X1 U9156 ( .A(n7547), .ZN(n7550) );
  AOI21_X1 U9157 ( .B1(n9606), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7548), .ZN(
        n7549) );
  OAI21_X1 U9158 ( .B1(n7550), .B2(n9613), .A(n7549), .ZN(P1_U3326) );
  OAI222_X1 U9159 ( .A1(n9060), .A2(n7551), .B1(n9058), .B2(n7550), .C1(n6359), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U9160 ( .A1(n7557), .A2(n7552), .ZN(n7554) );
  OAI211_X1 U9161 ( .C1(n9060), .C2(n7555), .A(n7554), .B(n7553), .ZN(P2_U3330) );
  NAND2_X1 U9162 ( .A1(n7557), .A2(n7556), .ZN(n7559) );
  OAI211_X1 U9163 ( .C1(n9609), .C2(n7560), .A(n7559), .B(n7558), .ZN(P1_U3325) );
  NOR2_X1 U9164 ( .A1(n7561), .A2(n4590), .ZN(n7566) );
  AOI21_X1 U9165 ( .B1(n7564), .B2(n7563), .A(n7562), .ZN(n7565) );
  OAI21_X1 U9166 ( .B1(n7566), .B2(n7565), .A(n9173), .ZN(n7574) );
  INV_X1 U9167 ( .A(n7567), .ZN(n7568) );
  AOI21_X1 U9168 ( .B1(n9188), .B2(n9199), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9169 ( .B1(n7570), .B2(n9632), .A(n7569), .ZN(n7571) );
  AOI21_X1 U9170 ( .B1(n7572), .B2(n9164), .A(n7571), .ZN(n7573) );
  OAI211_X1 U9171 ( .C1(n9673), .C2(n9181), .A(n7574), .B(n7573), .ZN(P1_U3232) );
  NAND2_X1 U9172 ( .A1(n9007), .A2(n8686), .ZN(n8413) );
  NOR2_X1 U9173 ( .A1(n9015), .A2(n8700), .ZN(n7575) );
  NAND2_X1 U9174 ( .A1(n9010), .A2(n8646), .ZN(n8505) );
  NAND2_X1 U9175 ( .A1(n7606), .A2(n7605), .ZN(n7608) );
  NAND2_X1 U9176 ( .A1(n9010), .A2(n8699), .ZN(n7577) );
  INV_X1 U9177 ( .A(n7941), .ZN(n7578) );
  AOI21_X1 U9178 ( .B1(n8507), .B2(n7579), .A(n7578), .ZN(n9009) );
  NAND2_X1 U9179 ( .A1(n9015), .A2(n8499), .ZN(n7580) );
  NAND2_X1 U9180 ( .A1(n7581), .A2(n7580), .ZN(n7583) );
  OR2_X1 U9181 ( .A1(n9015), .A2(n8499), .ZN(n7582) );
  INV_X1 U9182 ( .A(n8505), .ZN(n7584) );
  OAI211_X1 U9183 ( .C1(n4394), .C2(n8507), .A(n8911), .B(n8920), .ZN(n7586)
         );
  OR2_X1 U9184 ( .A1(n8646), .A2(n8861), .ZN(n7585) );
  OAI211_X1 U9185 ( .C1(n7948), .C2(n8863), .A(n7586), .B(n7585), .ZN(n9005)
         );
  INV_X1 U9186 ( .A(n9007), .ZN(n7590) );
  OR2_X1 U9187 ( .A1(n7616), .A2(n9010), .ZN(n7587) );
  NOR2_X2 U9188 ( .A1(n7587), .A2(n9007), .ZN(n8903) );
  AOI211_X1 U9189 ( .C1(n9007), .C2(n7587), .A(n9957), .B(n8903), .ZN(n9006)
         );
  NAND2_X1 U9190 ( .A1(n9006), .A2(n7956), .ZN(n7589) );
  AOI22_X1 U9191 ( .A1(n8931), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8643), .B2(
        n8929), .ZN(n7588) );
  OAI211_X1 U9192 ( .C1(n7590), .C2(n8908), .A(n7589), .B(n7588), .ZN(n7591)
         );
  AOI21_X1 U9193 ( .B1(n9005), .B2(n8933), .A(n7591), .ZN(n7592) );
  OAI21_X1 U9194 ( .B1(n9009), .B2(n8924), .A(n7592), .ZN(P2_U3279) );
  NAND2_X1 U9195 ( .A1(n7594), .A2(n7593), .ZN(n7596) );
  XNOR2_X1 U9196 ( .A(n7596), .B(n7595), .ZN(n7603) );
  NAND2_X1 U9197 ( .A1(n8680), .A2(n7597), .ZN(n7599) );
  AOI22_X1 U9198 ( .A1(n8682), .A2(n8699), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n7598) );
  OAI211_X1 U9199 ( .C1(n7600), .C2(n8685), .A(n7599), .B(n7598), .ZN(n7601)
         );
  AOI21_X1 U9200 ( .B1(n8688), .B2(n9015), .A(n7601), .ZN(n7602) );
  OAI21_X1 U9201 ( .B1(n7603), .B2(n8690), .A(n7602), .ZN(P2_U3243) );
  XNOR2_X1 U9202 ( .A(n7604), .B(n7605), .ZN(n7612) );
  OAI22_X1 U9203 ( .A1(n8499), .A2(n8861), .B1(n8686), .B2(n8863), .ZN(n7611)
         );
  OR2_X1 U9204 ( .A1(n7606), .A2(n7605), .ZN(n7607) );
  NAND2_X1 U9205 ( .A1(n7608), .A2(n7607), .ZN(n9014) );
  NOR2_X1 U9206 ( .A1(n9014), .A2(n7609), .ZN(n7610) );
  AOI211_X1 U9207 ( .C1(n8920), .C2(n7612), .A(n7611), .B(n7610), .ZN(n9013)
         );
  INV_X1 U9208 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7614) );
  INV_X1 U9209 ( .A(n7684), .ZN(n7613) );
  OAI22_X1 U9210 ( .A1(n8933), .A2(n7614), .B1(n7613), .B2(n8844), .ZN(n7615)
         );
  AOI21_X1 U9211 ( .B1(n9010), .B2(n8926), .A(n7615), .ZN(n7618) );
  INV_X1 U9212 ( .A(n9010), .ZN(n7688) );
  XNOR2_X1 U9213 ( .A(n7616), .B(n7688), .ZN(n9011) );
  NAND2_X1 U9214 ( .A1(n9011), .A2(n6814), .ZN(n7617) );
  OAI211_X1 U9215 ( .C1(n9014), .C2(n7619), .A(n7618), .B(n7617), .ZN(n7620)
         );
  INV_X1 U9216 ( .A(n7620), .ZN(n7621) );
  OAI21_X1 U9217 ( .B1(n9013), .B2(n8931), .A(n7621), .ZN(P2_U3280) );
  AND2_X1 U9218 ( .A1(n7622), .A2(n9200), .ZN(n7623) );
  OR2_X1 U9219 ( .A1(n9193), .A2(n9631), .ZN(n8110) );
  NAND2_X1 U9220 ( .A1(n9193), .A2(n9631), .ZN(n8222) );
  NAND2_X1 U9221 ( .A1(n8110), .A2(n8222), .ZN(n8320) );
  NAND2_X1 U9222 ( .A1(n7662), .A2(n8320), .ZN(n7696) );
  NAND2_X1 U9223 ( .A1(n9193), .A2(n9198), .ZN(n7694) );
  NAND2_X1 U9224 ( .A1(n7696), .A2(n7694), .ZN(n9467) );
  OR2_X1 U9225 ( .A1(n7689), .A2(n7665), .ZN(n8112) );
  NAND2_X1 U9226 ( .A1(n7689), .A2(n7665), .ZN(n9479) );
  NAND2_X1 U9227 ( .A1(n8112), .A2(n9479), .ZN(n9466) );
  XNOR2_X1 U9228 ( .A(n9467), .B(n9466), .ZN(n9656) );
  NAND2_X1 U9229 ( .A1(n7625), .A2(n8065), .ZN(n7656) );
  XNOR2_X1 U9230 ( .A(n9570), .B(n9186), .ZN(n8319) );
  OR2_X2 U9231 ( .A1(n7656), .A2(n8319), .ZN(n7653) );
  OR2_X1 U9232 ( .A1(n9570), .A2(n9186), .ZN(n8103) );
  INV_X1 U9233 ( .A(n9466), .ZN(n8322) );
  NAND3_X1 U9234 ( .A1(n7627), .A2(n8222), .A3(n9466), .ZN(n7628) );
  AND2_X1 U9235 ( .A1(n9480), .A2(n7628), .ZN(n7629) );
  OAI222_X1 U9236 ( .A1(n7744), .A2(n9635), .B1(n7630), .B2(n9631), .C1(n7655), 
        .C2(n7629), .ZN(n9657) );
  AOI211_X1 U9237 ( .C1(n7689), .C2(n4330), .A(n9843), .B(n7749), .ZN(n9658)
         );
  NAND2_X1 U9238 ( .A1(n9658), .A2(n9492), .ZN(n7634) );
  AOI22_X1 U9239 ( .A1(n9465), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7632), .B2(
        n9474), .ZN(n7633) );
  OAI211_X1 U9240 ( .C1(n9638), .C2(n9477), .A(n7634), .B(n7633), .ZN(n7635)
         );
  AOI21_X1 U9241 ( .B1(n9657), .B2(n9313), .A(n7635), .ZN(n7636) );
  OAI21_X1 U9242 ( .B1(n9656), .B2(n9494), .A(n7636), .ZN(P1_U3275) );
  NAND2_X1 U9243 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  XOR2_X1 U9244 ( .A(n7640), .B(n7639), .Z(n7647) );
  AOI21_X1 U9245 ( .B1(n9188), .B2(n9198), .A(n7641), .ZN(n7643) );
  NAND2_X1 U9246 ( .A1(n9164), .A2(n7650), .ZN(n7642) );
  OAI211_X1 U9247 ( .C1(n7644), .C2(n9632), .A(n7643), .B(n7642), .ZN(n7645)
         );
  AOI21_X1 U9248 ( .B1(n9570), .B2(n9192), .A(n7645), .ZN(n7646) );
  OAI21_X1 U9249 ( .B1(n7647), .B2(n9642), .A(n7646), .ZN(P1_U3213) );
  XOR2_X1 U9250 ( .A(n7648), .B(n8319), .Z(n9573) );
  AOI211_X1 U9251 ( .C1(n9570), .C2(n7649), .A(n9843), .B(n7631), .ZN(n9569)
         );
  AOI22_X1 U9252 ( .A1(n9489), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7650), .B2(
        n9474), .ZN(n7651) );
  OAI21_X1 U9253 ( .B1(n7652), .B2(n9477), .A(n7651), .ZN(n7660) );
  NOR2_X1 U9254 ( .A1(n9631), .A2(n7744), .ZN(n7658) );
  INV_X1 U9255 ( .A(n7653), .ZN(n7654) );
  AOI211_X1 U9256 ( .C1(n8319), .C2(n7656), .A(n7655), .B(n7654), .ZN(n7657)
         );
  AOI211_X1 U9257 ( .C1(n9483), .C2(n9200), .A(n7658), .B(n7657), .ZN(n9572)
         );
  NOR2_X1 U9258 ( .A1(n9572), .A2(n9489), .ZN(n7659) );
  AOI211_X1 U9259 ( .C1(n9492), .C2(n9569), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI21_X1 U9260 ( .B1(n9494), .B2(n9573), .A(n7661), .ZN(P1_U3277) );
  XNOR2_X1 U9261 ( .A(n7662), .B(n8320), .ZN(n9662) );
  XNOR2_X1 U9262 ( .A(n7663), .B(n8320), .ZN(n7667) );
  NAND2_X1 U9263 ( .A1(n9199), .A2(n9483), .ZN(n7664) );
  OAI21_X1 U9264 ( .B1(n7665), .B2(n7744), .A(n7664), .ZN(n7666) );
  AOI21_X1 U9265 ( .B1(n7667), .B2(n9488), .A(n7666), .ZN(n9667) );
  OAI21_X1 U9266 ( .B1(n9662), .B2(n9498), .A(n9667), .ZN(n7668) );
  NAND2_X1 U9267 ( .A1(n7668), .A2(n9313), .ZN(n7676) );
  OAI22_X1 U9268 ( .A1(n9313), .A2(n7670), .B1(n9190), .B2(n7669), .ZN(n7674)
         );
  NAND2_X1 U9269 ( .A1(n7671), .A2(n9193), .ZN(n7672) );
  NAND2_X1 U9270 ( .A1(n4330), .A2(n7672), .ZN(n9664) );
  NOR2_X1 U9271 ( .A1(n9664), .A2(n8019), .ZN(n7673) );
  AOI211_X1 U9272 ( .C1(n8017), .C2(n9193), .A(n7674), .B(n7673), .ZN(n7675)
         );
  OAI211_X1 U9273 ( .C1(n9662), .C2(n7677), .A(n7676), .B(n7675), .ZN(P1_U3276) );
  OAI21_X1 U9274 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  NAND2_X1 U9275 ( .A1(n7681), .A2(n8612), .ZN(n7686) );
  NAND2_X1 U9276 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U9277 ( .A1(n8623), .A2(n8700), .ZN(n7682) );
  OAI211_X1 U9278 ( .C1(n8672), .C2(n8686), .A(n8717), .B(n7682), .ZN(n7683)
         );
  AOI21_X1 U9279 ( .B1(n7684), .B2(n8680), .A(n7683), .ZN(n7685) );
  OAI211_X1 U9280 ( .C1(n7688), .C2(n7687), .A(n7686), .B(n7685), .ZN(P2_U3228) );
  INV_X1 U9281 ( .A(n9505), .ZN(n9310) );
  OR2_X1 U9282 ( .A1(n9552), .A2(n9162), .ZN(n8236) );
  NAND2_X1 U9283 ( .A1(n9552), .A2(n9162), .ZN(n8231) );
  NAND2_X1 U9284 ( .A1(n8236), .A2(n8231), .ZN(n9430) );
  INV_X1 U9285 ( .A(n9430), .ZN(n9435) );
  NAND2_X1 U9286 ( .A1(n9560), .A2(n9486), .ZN(n7693) );
  OR2_X1 U9287 ( .A1(n9560), .A2(n9119), .ZN(n8126) );
  NAND2_X1 U9288 ( .A1(n9560), .A2(n9119), .ZN(n8122) );
  INV_X1 U9289 ( .A(n9452), .ZN(n7692) );
  OR2_X1 U9290 ( .A1(n9565), .A2(n9446), .ZN(n7698) );
  INV_X1 U9291 ( .A(n7698), .ZN(n7691) );
  NAND2_X1 U9292 ( .A1(n7689), .A2(n9484), .ZN(n9468) );
  NAND2_X1 U9293 ( .A1(n9565), .A2(n9446), .ZN(n8115) );
  AND2_X1 U9294 ( .A1(n9468), .A2(n8115), .ZN(n7690) );
  OR2_X1 U9295 ( .A1(n7692), .A2(n9450), .ZN(n9454) );
  AND2_X1 U9296 ( .A1(n7694), .A2(n7697), .ZN(n7695) );
  NAND2_X1 U9297 ( .A1(n7696), .A2(n7695), .ZN(n7702) );
  INV_X1 U9298 ( .A(n7697), .ZN(n7700) );
  AND2_X1 U9299 ( .A1(n9466), .A2(n7698), .ZN(n9449) );
  AND2_X1 U9300 ( .A1(n9449), .A2(n9452), .ZN(n9427) );
  AND2_X1 U9301 ( .A1(n9427), .A2(n9430), .ZN(n7699) );
  OR2_X1 U9302 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  NAND2_X1 U9303 ( .A1(n9552), .A2(n9447), .ZN(n7703) );
  OR2_X1 U9304 ( .A1(n9548), .A2(n9437), .ZN(n7704) );
  NAND2_X1 U9305 ( .A1(n9548), .A2(n9437), .ZN(n7705) );
  AND2_X1 U9306 ( .A1(n9543), .A2(n9422), .ZN(n7706) );
  OR2_X1 U9307 ( .A1(n9543), .A2(n9422), .ZN(n7707) );
  NOR2_X1 U9308 ( .A1(n9537), .A2(n9409), .ZN(n7710) );
  NAND2_X1 U9309 ( .A1(n9537), .A2(n9409), .ZN(n7709) );
  AND2_X1 U9310 ( .A1(n9532), .A2(n9394), .ZN(n7711) );
  NAND2_X1 U9311 ( .A1(n9528), .A2(n9380), .ZN(n7712) );
  NAND2_X1 U9312 ( .A1(n9523), .A2(n9176), .ZN(n8249) );
  OR2_X1 U9313 ( .A1(n9523), .A2(n9366), .ZN(n7713) );
  INV_X1 U9314 ( .A(n7714), .ZN(n9328) );
  NAND2_X1 U9315 ( .A1(n9334), .A2(n9352), .ZN(n8254) );
  NAND2_X1 U9316 ( .A1(n9517), .A2(n9068), .ZN(n9322) );
  NAND2_X1 U9317 ( .A1(n9328), .A2(n7715), .ZN(n9327) );
  NAND2_X1 U9318 ( .A1(n9517), .A2(n9352), .ZN(n7716) );
  NAND2_X1 U9319 ( .A1(n9513), .A2(n7717), .ZN(n8183) );
  NAND2_X1 U9320 ( .A1(n9505), .A2(n9071), .ZN(n8184) );
  INV_X1 U9321 ( .A(SI_28_), .ZN(n7720) );
  NAND2_X1 U9322 ( .A1(n7721), .A2(n7720), .ZN(n7984) );
  NAND2_X1 U9323 ( .A1(n7987), .A2(n7984), .ZN(n7723) );
  INV_X1 U9324 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9059) );
  INV_X1 U9325 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9610) );
  MUX2_X1 U9326 ( .A(n9059), .B(n9610), .S(n8377), .Z(n7989) );
  XNOR2_X1 U9327 ( .A(n7989), .B(SI_29_), .ZN(n7722) );
  NAND2_X1 U9328 ( .A1(n9056), .A2(n8005), .ZN(n7725) );
  OR2_X1 U9329 ( .A1(n8006), .A2(n9610), .ZN(n7724) );
  XOR2_X1 U9330 ( .A(n9301), .B(n9499), .Z(n8329) );
  NAND2_X1 U9331 ( .A1(n9565), .A2(n9635), .ZN(n8300) );
  AND2_X1 U9332 ( .A1(n8300), .A2(n9479), .ZN(n7727) );
  NAND2_X1 U9333 ( .A1(n9480), .A2(n7727), .ZN(n9444) );
  OR2_X1 U9334 ( .A1(n9565), .A2(n9635), .ZN(n9443) );
  AND2_X1 U9335 ( .A1(n8126), .A2(n9443), .ZN(n8234) );
  NAND2_X1 U9336 ( .A1(n9444), .A2(n8234), .ZN(n7728) );
  NAND2_X1 U9337 ( .A1(n7728), .A2(n8122), .ZN(n9436) );
  NAND2_X1 U9338 ( .A1(n9436), .A2(n9435), .ZN(n7729) );
  NAND2_X1 U9339 ( .A1(n7729), .A2(n8231), .ZN(n9421) );
  INV_X1 U9340 ( .A(n9437), .ZN(n9090) );
  OR2_X1 U9341 ( .A1(n9548), .A2(n9090), .ZN(n8299) );
  NAND2_X1 U9342 ( .A1(n9421), .A2(n8299), .ZN(n7730) );
  NAND2_X1 U9343 ( .A1(n9548), .A2(n9090), .ZN(n8298) );
  OR2_X1 U9344 ( .A1(n9543), .A2(n9136), .ZN(n8239) );
  NAND2_X1 U9345 ( .A1(n9543), .A2(n9136), .ZN(n9390) );
  INV_X1 U9346 ( .A(n9409), .ZN(n9101) );
  AND2_X1 U9347 ( .A1(n9537), .A2(n9101), .ZN(n8145) );
  INV_X1 U9348 ( .A(n9390), .ZN(n7731) );
  OR2_X1 U9349 ( .A1(n8145), .A2(n7731), .ZN(n8201) );
  INV_X1 U9350 ( .A(n8201), .ZN(n7732) );
  OR2_X1 U9351 ( .A1(n9537), .A2(n9101), .ZN(n8241) );
  OR2_X1 U9352 ( .A1(n9532), .A2(n9152), .ZN(n8139) );
  NAND2_X1 U9353 ( .A1(n9532), .A2(n9152), .ZN(n8245) );
  NAND2_X1 U9354 ( .A1(n8139), .A2(n8245), .ZN(n9371) );
  INV_X1 U9355 ( .A(n9380), .ZN(n9110) );
  OR2_X1 U9356 ( .A1(n9528), .A2(n9110), .ZN(n8142) );
  NAND2_X1 U9357 ( .A1(n9528), .A2(n9110), .ZN(n9349) );
  NAND2_X2 U9358 ( .A1(n9364), .A2(n9365), .ZN(n9363) );
  INV_X1 U9359 ( .A(n9349), .ZN(n8251) );
  NOR2_X1 U9360 ( .A1(n9342), .A2(n8251), .ZN(n7734) );
  INV_X1 U9361 ( .A(n9322), .ZN(n8181) );
  NOR2_X1 U9362 ( .A1(n9315), .A2(n8181), .ZN(n8152) );
  INV_X1 U9363 ( .A(n8286), .ZN(n7735) );
  INV_X1 U9364 ( .A(n9298), .ZN(n7736) );
  OAI21_X1 U9365 ( .B1(n9299), .B2(n7736), .A(n8179), .ZN(n7737) );
  INV_X1 U9366 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U9367 ( .A1(n4313), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U9368 ( .A1(n7738), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7739) );
  OAI211_X1 U9369 ( .C1(n7742), .C2(n7741), .A(n7740), .B(n7739), .ZN(n9197)
         );
  AND2_X1 U9370 ( .A1(n9703), .A2(P1_B_REG_SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9371 ( .A1(n7744), .A2(n7743), .ZN(n8015) );
  NAND2_X1 U9372 ( .A1(n9197), .A2(n8015), .ZN(n7745) );
  AOI21_X2 U9373 ( .B1(n7748), .B2(n9488), .A(n7747), .ZN(n9502) );
  NOR2_X1 U9374 ( .A1(n9502), .A2(n9489), .ZN(n7756) );
  NAND2_X1 U9375 ( .A1(n7749), .A2(n9478), .ZN(n9471) );
  INV_X1 U9376 ( .A(n9548), .ZN(n9419) );
  AOI21_X1 U9377 ( .B1(n9499), .B2(n9305), .A(n9289), .ZN(n9500) );
  INV_X1 U9378 ( .A(n9499), .ZN(n8173) );
  INV_X1 U9379 ( .A(n7750), .ZN(n7751) );
  AOI22_X1 U9380 ( .A1(n7751), .A2(n9474), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9489), .ZN(n7752) );
  OAI21_X1 U9381 ( .B1(n8173), .B2(n9477), .A(n7752), .ZN(n7753) );
  OAI21_X1 U9382 ( .B1(n9503), .B2(n9494), .A(n7757), .ZN(n7939) );
  INV_X1 U9383 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7821) );
  INV_X1 U9384 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U9385 ( .A1(n7821), .A2(keyinput20), .B1(n9793), .B2(keyinput7), 
        .ZN(n7758) );
  OAI221_X1 U9386 ( .B1(n7821), .B2(keyinput20), .C1(n9793), .C2(keyinput7), 
        .A(n7758), .ZN(n7767) );
  AOI22_X1 U9387 ( .A1(n7778), .A2(keyinput42), .B1(n7760), .B2(keyinput39), 
        .ZN(n7759) );
  OAI221_X1 U9388 ( .B1(n7778), .B2(keyinput42), .C1(n7760), .C2(keyinput39), 
        .A(n7759), .ZN(n7766) );
  AOI22_X1 U9389 ( .A1(n7762), .A2(keyinput58), .B1(n5579), .B2(keyinput31), 
        .ZN(n7761) );
  OAI221_X1 U9390 ( .B1(n7762), .B2(keyinput58), .C1(n5579), .C2(keyinput31), 
        .A(n7761), .ZN(n7765) );
  INV_X1 U9391 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9680) );
  INV_X1 U9392 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U9393 ( .A1(n9680), .A2(keyinput13), .B1(n9795), .B2(keyinput26), 
        .ZN(n7763) );
  OAI221_X1 U9394 ( .B1(n9680), .B2(keyinput13), .C1(n9795), .C2(keyinput26), 
        .A(n7763), .ZN(n7764) );
  OR4_X1 U9395 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7764), .ZN(n7909) );
  AOI22_X1 U9396 ( .A1(n7769), .A2(keyinput82), .B1(n6037), .B2(keyinput127), 
        .ZN(n7768) );
  OAI221_X1 U9397 ( .B1(n7769), .B2(keyinput82), .C1(n6037), .C2(keyinput127), 
        .A(n7768), .ZN(n7776) );
  INV_X1 U9398 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7772) );
  AOI22_X1 U9399 ( .A1(n7772), .A2(keyinput89), .B1(n7771), .B2(keyinput123), 
        .ZN(n7770) );
  OAI221_X1 U9400 ( .B1(n7772), .B2(keyinput89), .C1(n7771), .C2(keyinput123), 
        .A(n7770), .ZN(n7775) );
  AOI22_X1 U9401 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput108), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput88), .ZN(n7773) );
  OAI221_X1 U9402 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput108), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput88), .A(n7773), .ZN(n7774) );
  NOR3_X1 U9403 ( .A1(n7776), .A2(n7775), .A3(n7774), .ZN(n7794) );
  INV_X1 U9404 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U9405 ( .A1(n9880), .A2(keyinput69), .B1(keyinput106), .B2(n7778), 
        .ZN(n7777) );
  OAI221_X1 U9406 ( .B1(n9880), .B2(keyinput69), .C1(n7778), .C2(keyinput106), 
        .A(n7777), .ZN(n7781) );
  AOI22_X1 U9407 ( .A1(n6768), .A2(keyinput109), .B1(P1_U3084), .B2(
        keyinput112), .ZN(n7779) );
  OAI221_X1 U9408 ( .B1(n6768), .B2(keyinput109), .C1(P1_U3084), .C2(
        keyinput112), .A(n7779), .ZN(n7780) );
  NOR2_X1 U9409 ( .A1(n7781), .A2(n7780), .ZN(n7793) );
  INV_X1 U9410 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10012) );
  INV_X1 U9411 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U9412 ( .A1(n10012), .A2(keyinput119), .B1(n9881), .B2(keyinput99), 
        .ZN(n7782) );
  OAI221_X1 U9413 ( .B1(n10012), .B2(keyinput119), .C1(n9881), .C2(keyinput99), 
        .A(n7782), .ZN(n7786) );
  AOI22_X1 U9414 ( .A1(n7784), .A2(keyinput124), .B1(n5567), .B2(keyinput101), 
        .ZN(n7783) );
  OAI221_X1 U9415 ( .B1(n7784), .B2(keyinput124), .C1(n5567), .C2(keyinput101), 
        .A(n7783), .ZN(n7785) );
  NOR2_X1 U9416 ( .A1(n7786), .A2(n7785), .ZN(n7792) );
  AOI22_X1 U9417 ( .A1(n6512), .A2(keyinput98), .B1(n9680), .B2(keyinput77), 
        .ZN(n7787) );
  OAI221_X1 U9418 ( .B1(n6512), .B2(keyinput98), .C1(n9680), .C2(keyinput77), 
        .A(n7787), .ZN(n7790) );
  INV_X1 U9419 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U9420 ( .A1(n7867), .A2(keyinput116), .B1(n9794), .B2(keyinput120), 
        .ZN(n7788) );
  OAI221_X1 U9421 ( .B1(n7867), .B2(keyinput116), .C1(n9794), .C2(keyinput120), 
        .A(n7788), .ZN(n7789) );
  NOR2_X1 U9422 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  AND4_X1 U9423 ( .A1(n7794), .A2(n7793), .A3(n7792), .A4(n7791), .ZN(n7852)
         );
  OAI22_X1 U9424 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput118), .B1(
        keyinput64), .B2(P1_D_REG_2__SCAN_IN), .ZN(n7795) );
  AOI221_X1 U9425 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput118), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput64), .A(n7795), .ZN(n7802) );
  OAI22_X1 U9426 ( .A1(SI_21_), .A2(keyinput86), .B1(P2_REG2_REG_8__SCAN_IN), 
        .B2(keyinput74), .ZN(n7796) );
  AOI221_X1 U9427 ( .B1(SI_21_), .B2(keyinput86), .C1(keyinput74), .C2(
        P2_REG2_REG_8__SCAN_IN), .A(n7796), .ZN(n7801) );
  OAI22_X1 U9428 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput68), .B1(
        P2_IR_REG_22__SCAN_IN), .B2(keyinput67), .ZN(n7797) );
  AOI221_X1 U9429 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput68), .C1(
        keyinput67), .C2(P2_IR_REG_22__SCAN_IN), .A(n7797), .ZN(n7800) );
  OAI22_X1 U9430 ( .A1(P1_D_REG_19__SCAN_IN), .A2(keyinput90), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(keyinput104), .ZN(n7798) );
  AOI221_X1 U9431 ( .B1(P1_D_REG_19__SCAN_IN), .B2(keyinput90), .C1(
        keyinput104), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7798), .ZN(n7799) );
  NAND4_X1 U9432 ( .A1(n7802), .A2(n7801), .A3(n7800), .A4(n7799), .ZN(n7807)
         );
  AOI22_X1 U9433 ( .A1(n7913), .A2(keyinput111), .B1(keyinput73), .B2(n5611), 
        .ZN(n7803) );
  OAI221_X1 U9434 ( .B1(n7913), .B2(keyinput111), .C1(n5611), .C2(keyinput73), 
        .A(n7803), .ZN(n7806) );
  INV_X1 U9435 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n7883) );
  AOI22_X1 U9436 ( .A1(n9079), .A2(keyinput105), .B1(keyinput87), .B2(n7883), 
        .ZN(n7804) );
  OAI221_X1 U9437 ( .B1(n9079), .B2(keyinput105), .C1(n7883), .C2(keyinput87), 
        .A(n7804), .ZN(n7805) );
  NOR3_X1 U9438 ( .A1(n7807), .A2(n7806), .A3(n7805), .ZN(n7851) );
  OAI22_X1 U9439 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput95), .B1(keyinput80), .B2(P2_IR_REG_15__SCAN_IN), .ZN(n7808) );
  AOI221_X1 U9440 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput95), .C1(
        P2_IR_REG_15__SCAN_IN), .C2(keyinput80), .A(n7808), .ZN(n7815) );
  OAI22_X1 U9441 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(keyinput114), .B1(
        P2_REG2_REG_23__SCAN_IN), .B2(keyinput107), .ZN(n7809) );
  AOI221_X1 U9442 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(keyinput114), .C1(
        keyinput107), .C2(P2_REG2_REG_23__SCAN_IN), .A(n7809), .ZN(n7814) );
  OAI22_X1 U9443 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput91), .B1(
        P2_REG0_REG_25__SCAN_IN), .B2(keyinput100), .ZN(n7810) );
  AOI221_X1 U9444 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput91), .C1(
        keyinput100), .C2(P2_REG0_REG_25__SCAN_IN), .A(n7810), .ZN(n7813) );
  OAI22_X1 U9445 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput78), .B1(SI_5_), 
        .B2(keyinput103), .ZN(n7811) );
  AOI221_X1 U9446 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput78), .C1(
        keyinput103), .C2(SI_5_), .A(n7811), .ZN(n7812) );
  NAND4_X1 U9447 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n7830)
         );
  INV_X1 U9448 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7911) );
  AOI22_X1 U9449 ( .A1(n7911), .A2(keyinput110), .B1(keyinput117), .B2(n9725), 
        .ZN(n7816) );
  OAI221_X1 U9450 ( .B1(n7911), .B2(keyinput110), .C1(n9725), .C2(keyinput117), 
        .A(n7816), .ZN(n7829) );
  XNOR2_X1 U9451 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput83), .ZN(n7820) );
  XNOR2_X1 U9452 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput81), .ZN(n7819) );
  XNOR2_X1 U9453 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput72), .ZN(n7818) );
  XNOR2_X1 U9454 ( .A(keyinput113), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7817) );
  AND4_X1 U9455 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n7827)
         );
  XNOR2_X1 U9456 ( .A(keyinput92), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n7826) );
  XNOR2_X1 U9457 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput85), .ZN(n7823) );
  XNOR2_X1 U9458 ( .A(keyinput84), .B(n7821), .ZN(n7822) );
  NOR2_X1 U9459 ( .A1(n7823), .A2(n7822), .ZN(n7825) );
  XNOR2_X1 U9460 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput96), .ZN(n7824) );
  NAND4_X1 U9461 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7824), .ZN(n7828)
         );
  NOR3_X1 U9462 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(n7850) );
  OAI22_X1 U9463 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(keyinput66), .B1(keyinput76), .B2(P2_REG0_REG_13__SCAN_IN), .ZN(n7831) );
  AOI221_X1 U9464 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(keyinput66), .C1(
        P2_REG0_REG_13__SCAN_IN), .C2(keyinput76), .A(n7831), .ZN(n7838) );
  OAI22_X1 U9465 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput94), .B1(
        keyinput126), .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n7832) );
  AOI221_X1 U9466 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput94), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput126), .A(n7832), .ZN(n7837) );
  OAI22_X1 U9467 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput115), .B1(keyinput121), .B2(P1_D_REG_3__SCAN_IN), .ZN(n7833) );
  AOI221_X1 U9468 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput115), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput121), .A(n7833), .ZN(n7836) );
  OAI22_X1 U9469 ( .A1(P1_D_REG_7__SCAN_IN), .A2(keyinput65), .B1(keyinput79), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n7834) );
  AOI221_X1 U9470 ( .B1(P1_D_REG_7__SCAN_IN), .B2(keyinput65), .C1(
        P2_REG2_REG_16__SCAN_IN), .C2(keyinput79), .A(n7834), .ZN(n7835) );
  NAND4_X1 U9471 ( .A1(n7838), .A2(n7837), .A3(n7836), .A4(n7835), .ZN(n7848)
         );
  OAI22_X1 U9472 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(keyinput93), .B1(
        keyinput70), .B2(P2_REG1_REG_22__SCAN_IN), .ZN(n7839) );
  AOI221_X1 U9473 ( .B1(P1_REG0_REG_18__SCAN_IN), .B2(keyinput93), .C1(
        P2_REG1_REG_22__SCAN_IN), .C2(keyinput70), .A(n7839), .ZN(n7846) );
  OAI22_X1 U9474 ( .A1(P1_D_REG_28__SCAN_IN), .A2(keyinput71), .B1(
        P2_REG0_REG_24__SCAN_IN), .B2(keyinput97), .ZN(n7840) );
  AOI221_X1 U9475 ( .B1(P1_D_REG_28__SCAN_IN), .B2(keyinput71), .C1(keyinput97), .C2(P2_REG0_REG_24__SCAN_IN), .A(n7840), .ZN(n7845) );
  OAI22_X1 U9476 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput122), .B1(
        keyinput75), .B2(P2_IR_REG_10__SCAN_IN), .ZN(n7841) );
  AOI221_X1 U9477 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput122), .C1(
        P2_IR_REG_10__SCAN_IN), .C2(keyinput75), .A(n7841), .ZN(n7844) );
  OAI22_X1 U9478 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput125), .B1(
        keyinput102), .B2(P1_REG0_REG_22__SCAN_IN), .ZN(n7842) );
  AOI221_X1 U9479 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput125), .C1(
        P1_REG0_REG_22__SCAN_IN), .C2(keyinput102), .A(n7842), .ZN(n7843) );
  NAND4_X1 U9480 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n7847)
         );
  NOR2_X1 U9481 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  NAND4_X1 U9482 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n7878)
         );
  AOI22_X1 U9483 ( .A1(n7854), .A2(keyinput50), .B1(keyinput16), .B2(n4882), 
        .ZN(n7853) );
  OAI221_X1 U9484 ( .B1(n7854), .B2(keyinput50), .C1(n4882), .C2(keyinput16), 
        .A(n7853), .ZN(n7860) );
  XNOR2_X1 U9485 ( .A(n9794), .B(keyinput56), .ZN(n7859) );
  XNOR2_X1 U9486 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput19), .ZN(n7857) );
  XNOR2_X1 U9487 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput32), .ZN(n7856) );
  XNOR2_X1 U9488 ( .A(keyinput2), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7855) );
  NAND3_X1 U9489 ( .A1(n7857), .A2(n7856), .A3(n7855), .ZN(n7858) );
  NOR3_X1 U9490 ( .A1(n7860), .A2(n7859), .A3(n7858), .ZN(n7877) );
  INV_X1 U9491 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9796) );
  INV_X1 U9492 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U9493 ( .A1(n9796), .A2(keyinput1), .B1(keyinput57), .B2(n9799), 
        .ZN(n7861) );
  OAI221_X1 U9494 ( .B1(n9796), .B2(keyinput1), .C1(n9799), .C2(keyinput57), 
        .A(n7861), .ZN(n7865) );
  AOI22_X1 U9495 ( .A1(n7863), .A2(keyinput54), .B1(keyinput4), .B2(n5754), 
        .ZN(n7862) );
  OAI221_X1 U9496 ( .B1(n7863), .B2(keyinput54), .C1(n5754), .C2(keyinput4), 
        .A(n7862), .ZN(n7864) );
  NOR2_X1 U9497 ( .A1(n7865), .A2(n7864), .ZN(n7876) );
  AOI22_X1 U9498 ( .A1(n7868), .A2(keyinput61), .B1(keyinput52), .B2(n7867), 
        .ZN(n7866) );
  OAI221_X1 U9499 ( .B1(n7868), .B2(keyinput61), .C1(n7867), .C2(keyinput52), 
        .A(n7866), .ZN(n7874) );
  INV_X1 U9500 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U9501 ( .A1(n9797), .A2(keyinput51), .B1(keyinput62), .B2(n9966), 
        .ZN(n7869) );
  OAI221_X1 U9502 ( .B1(n9797), .B2(keyinput51), .C1(n9966), .C2(keyinput62), 
        .A(n7869), .ZN(n7873) );
  INV_X1 U9503 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9948) );
  AOI22_X1 U9504 ( .A1(n9948), .A2(keyinput30), .B1(keyinput6), .B2(n7871), 
        .ZN(n7870) );
  OAI221_X1 U9505 ( .B1(n9948), .B2(keyinput30), .C1(n7871), .C2(keyinput6), 
        .A(n7870), .ZN(n7872) );
  NOR3_X1 U9506 ( .A1(n7874), .A2(n7873), .A3(n7872), .ZN(n7875) );
  NAND4_X1 U9507 ( .A1(n7878), .A2(n7877), .A3(n7876), .A4(n7875), .ZN(n7908)
         );
  AOI22_X1 U9508 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput36), .B1(
        P2_IR_REG_10__SCAN_IN), .B2(keyinput11), .ZN(n7879) );
  OAI221_X1 U9509 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput36), .C1(
        P2_IR_REG_10__SCAN_IN), .C2(keyinput11), .A(n7879), .ZN(n7887) );
  AOI22_X1 U9510 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput18), .B1(
        P1_REG2_REG_7__SCAN_IN), .B2(keyinput49), .ZN(n7880) );
  OAI221_X1 U9511 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput18), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(keyinput49), .A(n7880), .ZN(n7886) );
  AOI22_X1 U9512 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput44), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput24), .ZN(n7881) );
  OAI221_X1 U9513 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput44), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput24), .A(n7881), .ZN(n7885) );
  AOI22_X1 U9514 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput33), .B1(n7883), 
        .B2(keyinput23), .ZN(n7882) );
  OAI221_X1 U9515 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput33), .C1(n7883), 
        .C2(keyinput23), .A(n7882), .ZN(n7884) );
  NOR4_X1 U9516 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n7906)
         );
  AOI22_X1 U9517 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(keyinput55), .B1(SI_4_), 
        .B2(keyinput59), .ZN(n7888) );
  OAI221_X1 U9518 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(keyinput55), .C1(SI_4_), 
        .C2(keyinput59), .A(n7888), .ZN(n7895) );
  AOI22_X1 U9519 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput43), .B1(
        P2_IR_REG_21__SCAN_IN), .B2(keyinput8), .ZN(n7889) );
  OAI221_X1 U9520 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput43), .C1(
        P2_IR_REG_21__SCAN_IN), .C2(keyinput8), .A(n7889), .ZN(n7894) );
  AOI22_X1 U9521 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput10), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput37), .ZN(n7890) );
  OAI221_X1 U9522 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput10), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput37), .A(n7890), .ZN(n7893) );
  AOI22_X1 U9523 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput60), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput35), .ZN(n7891) );
  OAI221_X1 U9524 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput60), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput35), .A(n7891), .ZN(n7892) );
  NOR4_X1 U9525 ( .A1(n7895), .A2(n7894), .A3(n7893), .A4(n7892), .ZN(n7905)
         );
  AOI22_X1 U9526 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput48), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput17), .ZN(n7896) );
  OAI221_X1 U9527 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput48), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput17), .A(n7896), .ZN(n7903) );
  AOI22_X1 U9528 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(keyinput15), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput27), .ZN(n7897) );
  OAI221_X1 U9529 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(keyinput15), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput27), .A(n7897), .ZN(n7902) );
  AOI22_X1 U9530 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput21), .B1(
        P1_REG1_REG_13__SCAN_IN), .B2(keyinput45), .ZN(n7898) );
  OAI221_X1 U9531 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput21), .C1(
        P1_REG1_REG_13__SCAN_IN), .C2(keyinput45), .A(n7898), .ZN(n7901) );
  AOI22_X1 U9532 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(keyinput25), .B1(
        P1_REG0_REG_18__SCAN_IN), .B2(keyinput29), .ZN(n7899) );
  OAI221_X1 U9533 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG0_REG_18__SCAN_IN), .C2(keyinput29), .A(n7899), .ZN(n7900) );
  NOR4_X1 U9534 ( .A1(n7903), .A2(n7902), .A3(n7901), .A4(n7900), .ZN(n7904)
         );
  NAND3_X1 U9535 ( .A1(n7906), .A2(n7905), .A3(n7904), .ZN(n7907) );
  NOR3_X1 U9536 ( .A1(n7909), .A2(n7908), .A3(n7907), .ZN(n7937) );
  AOI22_X1 U9537 ( .A1(n9079), .A2(keyinput41), .B1(keyinput46), .B2(n7911), 
        .ZN(n7910) );
  OAI221_X1 U9538 ( .B1(n9079), .B2(keyinput41), .C1(n7911), .C2(keyinput46), 
        .A(n7910), .ZN(n7923) );
  AOI22_X1 U9539 ( .A1(n7914), .A2(keyinput14), .B1(keyinput47), .B2(n7913), 
        .ZN(n7912) );
  OAI221_X1 U9540 ( .B1(n7914), .B2(keyinput14), .C1(n7913), .C2(keyinput47), 
        .A(n7912), .ZN(n7922) );
  AOI22_X1 U9541 ( .A1(n7916), .A2(keyinput28), .B1(n6037), .B2(keyinput63), 
        .ZN(n7915) );
  OAI221_X1 U9542 ( .B1(n7916), .B2(keyinput28), .C1(n6037), .C2(keyinput63), 
        .A(n7915), .ZN(n7921) );
  AOI22_X1 U9543 ( .A1(n7919), .A2(keyinput22), .B1(keyinput40), .B2(n7918), 
        .ZN(n7917) );
  OAI221_X1 U9544 ( .B1(n7919), .B2(keyinput22), .C1(n7918), .C2(keyinput40), 
        .A(n7917), .ZN(n7920) );
  NOR4_X1 U9545 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n7936)
         );
  INV_X1 U9546 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7925) );
  AOI22_X1 U9547 ( .A1(n9725), .A2(keyinput53), .B1(n7925), .B2(keyinput38), 
        .ZN(n7924) );
  OAI221_X1 U9548 ( .B1(n9725), .B2(keyinput53), .C1(n7925), .C2(keyinput38), 
        .A(n7924), .ZN(n7934) );
  INV_X1 U9549 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U9550 ( .A1(n7927), .A2(keyinput3), .B1(n9800), .B2(keyinput0), 
        .ZN(n7926) );
  OAI221_X1 U9551 ( .B1(n7927), .B2(keyinput3), .C1(n9800), .C2(keyinput0), 
        .A(n7926), .ZN(n7933) );
  AOI22_X1 U9552 ( .A1(n9880), .A2(keyinput5), .B1(n5611), .B2(keyinput9), 
        .ZN(n7928) );
  OAI221_X1 U9553 ( .B1(n9880), .B2(keyinput5), .C1(n5611), .C2(keyinput9), 
        .A(n7928), .ZN(n7932) );
  INV_X1 U9554 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7930) );
  AOI22_X1 U9555 ( .A1(n7930), .A2(keyinput12), .B1(keyinput34), .B2(n6512), 
        .ZN(n7929) );
  OAI221_X1 U9556 ( .B1(n7930), .B2(keyinput12), .C1(n6512), .C2(keyinput34), 
        .A(n7929), .ZN(n7931) );
  NOR4_X1 U9557 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n7935)
         );
  NAND3_X1 U9558 ( .A1(n7937), .A2(n7936), .A3(n7935), .ZN(n7938) );
  XNOR2_X1 U9559 ( .A(n7939), .B(n7938), .ZN(P1_U3355) );
  OR2_X1 U9560 ( .A1(n9007), .A2(n8916), .ZN(n7940) );
  NOR2_X1 U9561 ( .A1(n9000), .A2(n8698), .ZN(n7942) );
  OR2_X1 U9562 ( .A1(n8996), .A2(n8661), .ZN(n8522) );
  NAND2_X1 U9563 ( .A1(n8996), .A2(n8661), .ZN(n8526) );
  XNOR2_X1 U9564 ( .A(n8024), .B(n8401), .ZN(n8999) );
  INV_X1 U9565 ( .A(n9000), .ZN(n8909) );
  AND2_X2 U9566 ( .A1(n8909), .A2(n8903), .ZN(n8904) );
  INV_X1 U9567 ( .A(n8904), .ZN(n7944) );
  INV_X1 U9568 ( .A(n8996), .ZN(n7947) );
  INV_X1 U9569 ( .A(n8892), .ZN(n7943) );
  AOI211_X1 U9570 ( .C1(n8996), .C2(n7944), .A(n9957), .B(n7943), .ZN(n8995)
         );
  INV_X1 U9571 ( .A(n8606), .ZN(n7945) );
  AOI22_X1 U9572 ( .A1(n8931), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n7945), .B2(
        n8929), .ZN(n7946) );
  OAI21_X1 U9573 ( .B1(n7947), .B2(n8908), .A(n7946), .ZN(n7955) );
  OR2_X1 U9574 ( .A1(n9000), .A2(n7948), .ZN(n8511) );
  NAND2_X1 U9575 ( .A1(n9000), .A2(n7948), .ZN(n8524) );
  AND2_X1 U9576 ( .A1(n8910), .A2(n8914), .ZN(n7949) );
  NAND2_X1 U9577 ( .A1(n7950), .A2(n7952), .ZN(n8044) );
  OAI21_X1 U9578 ( .B1(n7952), .B2(n7950), .A(n7951), .ZN(n7953) );
  AOI222_X1 U9579 ( .A1(n8920), .A2(n7953), .B1(n8881), .B2(n8917), .C1(n8698), 
        .C2(n8915), .ZN(n8998) );
  NOR2_X1 U9580 ( .A1(n8998), .A2(n8931), .ZN(n7954) );
  AOI211_X1 U9581 ( .C1(n8995), .C2(n7956), .A(n7955), .B(n7954), .ZN(n7957)
         );
  OAI21_X1 U9582 ( .B1(n8924), .B2(n8999), .A(n7957), .ZN(P2_U3277) );
  NAND2_X1 U9583 ( .A1(n8732), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7964) );
  XOR2_X1 U9584 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8732), .Z(n8728) );
  NAND2_X1 U9585 ( .A1(n8720), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7963) );
  OR2_X1 U9586 ( .A1(n8720), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7958) );
  AND2_X1 U9587 ( .A1(n7958), .A2(n7963), .ZN(n8722) );
  NOR2_X1 U9588 ( .A1(n7960), .A2(n7959), .ZN(n7962) );
  NOR2_X1 U9589 ( .A1(n7962), .A2(n7961), .ZN(n8723) );
  NAND2_X1 U9590 ( .A1(n8722), .A2(n8723), .ZN(n8721) );
  NAND2_X1 U9591 ( .A1(n7963), .A2(n8721), .ZN(n8729) );
  NAND2_X1 U9592 ( .A1(n8728), .A2(n8729), .ZN(n8727) );
  NAND2_X1 U9593 ( .A1(n7964), .A2(n8727), .ZN(n7965) );
  NOR2_X1 U9594 ( .A1(n7965), .A2(n8749), .ZN(n7967) );
  AOI21_X1 U9595 ( .B1(n8749), .B2(n7965), .A(n7967), .ZN(n7966) );
  INV_X1 U9596 ( .A(n7966), .ZN(n8742) );
  NOR2_X1 U9597 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8742), .ZN(n8741) );
  NOR2_X1 U9598 ( .A1(n8741), .A2(n7967), .ZN(n7968) );
  XOR2_X1 U9599 ( .A(n7968), .B(P2_REG2_REG_19__SCAN_IN), .Z(n7981) );
  INV_X1 U9600 ( .A(n7981), .ZN(n7978) );
  INV_X1 U9601 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7969) );
  XNOR2_X1 U9602 ( .A(n8749), .B(n7969), .ZN(n8744) );
  XNOR2_X1 U9603 ( .A(n8732), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8735) );
  OR2_X1 U9604 ( .A1(n8720), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7974) );
  XOR2_X1 U9605 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8720), .Z(n8714) );
  NOR2_X1 U9606 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  NOR2_X1 U9607 ( .A1(n8749), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7975) );
  AOI21_X1 U9608 ( .B1(n8744), .B2(n8743), .A(n7975), .ZN(n7976) );
  XNOR2_X1 U9609 ( .A(n7976), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U9610 ( .A1(n9868), .A2(n7979), .ZN(n7980) );
  NAND2_X1 U9611 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n7982) );
  INV_X1 U9612 ( .A(SI_29_), .ZN(n7983) );
  AND2_X1 U9613 ( .A1(n7989), .A2(n7983), .ZN(n7986) );
  INV_X1 U9614 ( .A(n7984), .ZN(n7985) );
  NOR2_X1 U9615 ( .A1(n7986), .A2(n7985), .ZN(n7988) );
  NAND2_X1 U9616 ( .A1(n7988), .A2(n7987), .ZN(n7992) );
  INV_X1 U9617 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U9618 ( .A1(n7990), .A2(SI_29_), .ZN(n7991) );
  NAND2_X1 U9619 ( .A1(n7992), .A2(n7991), .ZN(n7995) );
  MUX2_X1 U9620 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8001), .Z(n7994) );
  INV_X1 U9621 ( .A(n8004), .ZN(n7993) );
  NAND2_X1 U9622 ( .A1(n7993), .A2(SI_30_), .ZN(n7997) );
  NAND2_X1 U9623 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND2_X1 U9624 ( .A1(n7997), .A2(n7996), .ZN(n8000) );
  MUX2_X1 U9625 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8001), .Z(n7998) );
  XNOR2_X1 U9626 ( .A(n7998), .B(SI_31_), .ZN(n7999) );
  MUX2_X1 U9627 ( .A(n9048), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8001), .Z(n8003) );
  NAND2_X1 U9628 ( .A1(n8371), .A2(n8005), .ZN(n8008) );
  INV_X1 U9629 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8367) );
  OR2_X1 U9630 ( .A1(n8006), .A2(n8367), .ZN(n8007) );
  INV_X1 U9631 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8009) );
  NOR2_X1 U9632 ( .A1(n9313), .A2(n8009), .ZN(n8016) );
  NAND2_X1 U9633 ( .A1(n5644), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8014) );
  OR2_X1 U9634 ( .A1(n4314), .A2(n8009), .ZN(n8013) );
  INV_X1 U9635 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8011) );
  OR2_X1 U9636 ( .A1(n5709), .A2(n8011), .ZN(n8012) );
  NAND2_X1 U9637 ( .A1(n9196), .A2(n8015), .ZN(n9651) );
  NOR2_X1 U9638 ( .A1(n9651), .A2(n9489), .ZN(n9292) );
  AOI211_X1 U9639 ( .C1(n9495), .C2(n8017), .A(n8016), .B(n9292), .ZN(n8018)
         );
  OAI21_X1 U9640 ( .B1(n9497), .B2(n8019), .A(n8018), .ZN(P1_U3261) );
  OAI222_X1 U9641 ( .A1(n9060), .A2(n8021), .B1(n9058), .B2(n8020), .C1(
        P2_U3152), .C2(n5519), .ZN(P2_U3336) );
  AND2_X1 U9642 ( .A1(n8996), .A2(n8918), .ZN(n8023) );
  NAND2_X1 U9643 ( .A1(n8990), .A2(n8025), .ZN(n8527) );
  NAND2_X1 U9644 ( .A1(n8528), .A2(n8527), .ZN(n8889) );
  OR2_X1 U9645 ( .A1(n8046), .A2(n4341), .ZN(n8029) );
  NAND2_X1 U9646 ( .A1(n8985), .A2(n8897), .ZN(n8027) );
  NAND2_X1 U9647 ( .A1(n8990), .A2(n8881), .ZN(n8870) );
  OR2_X1 U9648 ( .A1(n4341), .A2(n8870), .ZN(n8026) );
  AND2_X1 U9649 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  NAND2_X1 U9650 ( .A1(n8980), .A2(n8837), .ZN(n8533) );
  NAND2_X1 U9651 ( .A1(n8834), .A2(n8533), .ZN(n8860) );
  OR2_X1 U9652 ( .A1(n8848), .A2(n8864), .ZN(n8519) );
  NAND2_X1 U9653 ( .A1(n8848), .A2(n8864), .ZN(n8541) );
  NAND2_X1 U9654 ( .A1(n8519), .A2(n8541), .ZN(n8518) );
  INV_X1 U9655 ( .A(n8518), .ZN(n8833) );
  OR2_X1 U9656 ( .A1(n8968), .A2(n8838), .ZN(n8543) );
  NAND2_X1 U9657 ( .A1(n8968), .A2(n8838), .ZN(n8542) );
  NAND2_X1 U9658 ( .A1(n8543), .A2(n8542), .ZN(n8820) );
  INV_X1 U9659 ( .A(n8838), .ZN(n8697) );
  XNOR2_X1 U9660 ( .A(n8965), .B(n8822), .ZN(n8802) );
  NAND2_X1 U9661 ( .A1(n8039), .A2(n8695), .ZN(n8552) );
  NAND2_X1 U9662 ( .A1(n8961), .A2(n8775), .ZN(n8555) );
  XNOR2_X1 U9663 ( .A(n8954), .B(n8694), .ZN(n8554) );
  INV_X1 U9664 ( .A(n8554), .ZN(n8774) );
  NAND2_X1 U9665 ( .A1(n8768), .A2(n8774), .ZN(n8767) );
  NAND2_X1 U9666 ( .A1(n8767), .A2(n8032), .ZN(n8362) );
  NAND2_X1 U9667 ( .A1(n8949), .A2(n8776), .ZN(n8563) );
  NAND2_X1 U9668 ( .A1(n8033), .A2(n8776), .ZN(n8034) );
  NAND2_X1 U9669 ( .A1(n8363), .A2(n8034), .ZN(n8038) );
  NAND2_X1 U9670 ( .A1(n9056), .A2(n8370), .ZN(n8036) );
  OR2_X1 U9671 ( .A1(n4947), .A2(n9059), .ZN(n8035) );
  INV_X1 U9672 ( .A(n8942), .ZN(n8043) );
  INV_X1 U9673 ( .A(n8051), .ZN(n8566) );
  NAND2_X1 U9674 ( .A1(n8567), .A2(n8566), .ZN(n8407) );
  INV_X1 U9675 ( .A(n8407), .ZN(n8565) );
  INV_X1 U9676 ( .A(n8968), .ZN(n8818) );
  INV_X1 U9677 ( .A(n8985), .ZN(n8877) );
  NOR2_X2 U9678 ( .A1(n8848), .A2(n8854), .ZN(n8842) );
  NAND2_X1 U9679 ( .A1(n8818), .A2(n8842), .ZN(n8813) );
  NOR2_X2 U9680 ( .A1(n8813), .A2(n8965), .ZN(n8806) );
  NAND2_X1 U9681 ( .A1(n8039), .A2(n8806), .ZN(n8790) );
  NOR2_X2 U9682 ( .A1(n8954), .A2(n8790), .ZN(n8770) );
  AOI21_X1 U9683 ( .B1(n8942), .B2(n8356), .A(n8761), .ZN(n8943) );
  INV_X1 U9684 ( .A(n8040), .ZN(n8041) );
  AOI22_X1 U9685 ( .A1(n8931), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8041), .B2(
        n8929), .ZN(n8042) );
  OAI21_X1 U9686 ( .B1(n8043), .B2(n8908), .A(n8042), .ZN(n8059) );
  NAND2_X1 U9687 ( .A1(n8044), .A2(n8526), .ZN(n8896) );
  INV_X1 U9688 ( .A(n8896), .ZN(n8047) );
  AOI21_X1 U9689 ( .B1(n8047), .B2(n8046), .A(n8045), .ZN(n8879) );
  OR2_X1 U9690 ( .A1(n8985), .A2(n8862), .ZN(n8529) );
  NAND2_X1 U9691 ( .A1(n8985), .A2(n8862), .ZN(n8532) );
  INV_X1 U9692 ( .A(n8834), .ZN(n8049) );
  NOR2_X1 U9693 ( .A1(n8518), .A2(n8049), .ZN(n8537) );
  INV_X1 U9694 ( .A(n8541), .ZN(n8821) );
  OR2_X1 U9695 ( .A1(n8822), .A2(n8965), .ZN(n8550) );
  OAI21_X1 U9696 ( .B1(n8803), .B2(n8802), .A(n8550), .ZN(n8787) );
  INV_X1 U9697 ( .A(n8694), .ZN(n8789) );
  INV_X1 U9698 ( .A(n8562), .ZN(n8050) );
  AOI21_X1 U9699 ( .B1(n8354), .B2(n8405), .A(n8050), .ZN(n8052) );
  NAND2_X1 U9700 ( .A1(n8369), .A2(n8567), .ZN(n8057) );
  AOI21_X1 U9701 ( .B1(n8052), .B2(n8407), .A(n8859), .ZN(n8056) );
  INV_X1 U9702 ( .A(P2_B_REG_SCAN_IN), .ZN(n8053) );
  NOR2_X1 U9703 ( .A1(n6359), .A2(n8053), .ZN(n8054) );
  OR2_X1 U9704 ( .A1(n8863), .A2(n8054), .ZN(n8754) );
  OAI22_X1 U9705 ( .A1(n8776), .A2(n8861), .B1(n8378), .B2(n8754), .ZN(n8055)
         );
  NOR2_X1 U9706 ( .A1(n8945), .A2(n8931), .ZN(n8058) );
  AOI211_X2 U9707 ( .C1(n6814), .C2(n8943), .A(n8059), .B(n8058), .ZN(n8060)
         );
  OAI21_X1 U9708 ( .B1(n8947), .B2(n8924), .A(n8060), .ZN(P2_U3267) );
  NOR2_X1 U9709 ( .A1(n9495), .A2(n8062), .ZN(n8342) );
  NAND2_X1 U9710 ( .A1(n8340), .A2(n8296), .ZN(n8336) );
  NOR3_X1 U9711 ( .A1(n8342), .A2(n8061), .A3(n8336), .ZN(n8346) );
  NAND2_X1 U9712 ( .A1(n9495), .A2(n8062), .ZN(n8259) );
  INV_X1 U9713 ( .A(n9197), .ZN(n8258) );
  NOR2_X1 U9714 ( .A1(n9290), .A2(n8258), .ZN(n8330) );
  NAND2_X1 U9715 ( .A1(n9495), .A2(n8330), .ZN(n8063) );
  NAND2_X1 U9716 ( .A1(n8259), .A2(n8063), .ZN(n8164) );
  NAND2_X1 U9717 ( .A1(n9197), .A2(n9196), .ZN(n8064) );
  NAND2_X1 U9718 ( .A1(n9290), .A2(n8064), .ZN(n8289) );
  NAND2_X1 U9719 ( .A1(n9570), .A2(n9186), .ZN(n8105) );
  NAND2_X1 U9720 ( .A1(n8105), .A2(n8065), .ZN(n8221) );
  NAND2_X1 U9721 ( .A1(n8070), .A2(n8168), .ZN(n8066) );
  NAND3_X1 U9722 ( .A1(n8066), .A2(n8075), .A3(n8305), .ZN(n8069) );
  NAND2_X1 U9723 ( .A1(n8080), .A2(n8067), .ZN(n8209) );
  INV_X1 U9724 ( .A(n8168), .ZN(n8171) );
  NAND2_X1 U9725 ( .A1(n8209), .A2(n8171), .ZN(n8068) );
  NAND2_X1 U9726 ( .A1(n8069), .A2(n8068), .ZN(n8072) );
  OR3_X1 U9727 ( .A1(n8070), .A2(n8168), .A3(n8209), .ZN(n8071) );
  NAND2_X1 U9728 ( .A1(n8072), .A2(n8071), .ZN(n8088) );
  AND2_X1 U9729 ( .A1(n8204), .A2(n8082), .ZN(n8229) );
  AND2_X1 U9730 ( .A1(n8085), .A2(n8081), .ZN(n8203) );
  AND2_X1 U9731 ( .A1(n8218), .A2(n8263), .ZN(n8077) );
  MUX2_X1 U9732 ( .A(n8073), .B(n8271), .S(n8168), .Z(n8074) );
  INV_X1 U9733 ( .A(n8074), .ZN(n8076) );
  NAND2_X1 U9734 ( .A1(n8076), .A2(n8075), .ZN(n8087) );
  AND4_X1 U9735 ( .A1(n8229), .A2(n8203), .A3(n8077), .A4(n8087), .ZN(n8079)
         );
  AOI21_X1 U9736 ( .B1(n8088), .B2(n8079), .A(n8078), .ZN(n8092) );
  AOI21_X1 U9737 ( .B1(n8081), .B2(n8080), .A(n8171), .ZN(n8084) );
  AOI21_X1 U9738 ( .B1(n8082), .B2(n8218), .A(n8168), .ZN(n8083) );
  AOI22_X1 U9739 ( .A1(n8229), .A2(n8084), .B1(n8203), .B2(n8083), .ZN(n8091)
         );
  NAND2_X1 U9740 ( .A1(n8100), .A2(n8085), .ZN(n8086) );
  NAND2_X1 U9741 ( .A1(n8086), .A2(n8168), .ZN(n8090) );
  NAND4_X1 U9742 ( .A1(n8088), .A2(n8171), .A3(n8203), .A4(n8087), .ZN(n8089)
         );
  NAND4_X1 U9743 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n8098)
         );
  AND2_X1 U9744 ( .A1(n8103), .A2(n8093), .ZN(n8104) );
  NAND2_X1 U9745 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  NAND2_X1 U9746 ( .A1(n8096), .A2(n8100), .ZN(n8220) );
  NAND3_X1 U9747 ( .A1(n8098), .A2(n8104), .A3(n8220), .ZN(n8097) );
  OR2_X1 U9748 ( .A1(n8098), .A2(n4617), .ZN(n8102) );
  NAND2_X1 U9749 ( .A1(n8100), .A2(n8099), .ZN(n8202) );
  INV_X1 U9750 ( .A(n8320), .ZN(n8109) );
  NAND2_X1 U9751 ( .A1(n8221), .A2(n8103), .ZN(n8107) );
  INV_X1 U9752 ( .A(n8104), .ZN(n8106) );
  NAND2_X1 U9753 ( .A1(n8106), .A2(n8105), .ZN(n8219) );
  MUX2_X1 U9754 ( .A(n8107), .B(n8219), .S(n8171), .Z(n8108) );
  AND2_X1 U9755 ( .A1(n9479), .A2(n8222), .ZN(n8111) );
  AND2_X1 U9756 ( .A1(n8112), .A2(n8110), .ZN(n8227) );
  MUX2_X1 U9757 ( .A(n8111), .B(n8227), .S(n8168), .Z(n8114) );
  MUX2_X1 U9758 ( .A(n8112), .B(n9479), .S(n8168), .Z(n8113) );
  OAI21_X1 U9759 ( .B1(n9446), .B2(n8168), .A(n8115), .ZN(n8117) );
  NAND2_X1 U9760 ( .A1(n8122), .A2(n8300), .ZN(n8212) );
  AND2_X1 U9761 ( .A1(n8212), .A2(n8171), .ZN(n8116) );
  AOI21_X1 U9762 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n8125) );
  OAI21_X1 U9763 ( .B1(n8119), .B2(n9565), .A(n8234), .ZN(n8120) );
  NAND2_X1 U9764 ( .A1(n8120), .A2(n8168), .ZN(n8121) );
  NAND2_X1 U9765 ( .A1(n8125), .A2(n8121), .ZN(n8124) );
  AND2_X1 U9766 ( .A1(n8231), .A2(n8122), .ZN(n8233) );
  NAND2_X1 U9767 ( .A1(n8124), .A2(n8233), .ZN(n8123) );
  NAND2_X1 U9768 ( .A1(n8123), .A2(n8236), .ZN(n8131) );
  NAND3_X1 U9769 ( .A1(n8124), .A2(n9162), .A3(n8126), .ZN(n8129) );
  INV_X1 U9770 ( .A(n8125), .ZN(n8127) );
  AOI21_X1 U9771 ( .B1(n8127), .B2(n8126), .A(n9162), .ZN(n8128) );
  AOI21_X1 U9772 ( .B1(n8129), .B2(n4483), .A(n8128), .ZN(n8130) );
  MUX2_X1 U9773 ( .A(n8131), .B(n8130), .S(n8171), .Z(n8132) );
  AND2_X1 U9774 ( .A1(n9408), .A2(n8299), .ZN(n8133) );
  OAI21_X1 U9775 ( .B1(n8298), .B2(n8168), .A(n8241), .ZN(n8138) );
  NAND2_X1 U9776 ( .A1(n9349), .A2(n8245), .ZN(n8143) );
  INV_X1 U9777 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9778 ( .A1(n8134), .A2(n9390), .ZN(n8135) );
  AOI21_X1 U9779 ( .B1(n8135), .B2(n8241), .A(n8168), .ZN(n8136) );
  NOR2_X1 U9780 ( .A1(n8143), .A2(n8136), .ZN(n8137) );
  NAND2_X1 U9781 ( .A1(n8142), .A2(n8139), .ZN(n8248) );
  NAND2_X1 U9782 ( .A1(n8248), .A2(n8171), .ZN(n8140) );
  NAND2_X1 U9783 ( .A1(n8141), .A2(n8140), .ZN(n8153) );
  NAND2_X1 U9784 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  AND2_X1 U9785 ( .A1(n8249), .A2(n8144), .ZN(n8284) );
  NAND2_X1 U9786 ( .A1(n8145), .A2(n8171), .ZN(n8147) );
  NAND4_X1 U9787 ( .A1(n9349), .A2(n9378), .A3(n8168), .A4(n9394), .ZN(n8146)
         );
  OAI211_X1 U9788 ( .C1(n8248), .C2(n8147), .A(n8253), .B(n8146), .ZN(n8148)
         );
  INV_X1 U9789 ( .A(n8148), .ZN(n8149) );
  OAI211_X1 U9790 ( .C1(n8284), .C2(n8168), .A(n8254), .B(n8149), .ZN(n8150)
         );
  INV_X1 U9791 ( .A(n8150), .ZN(n8151) );
  AOI21_X1 U9792 ( .B1(n8254), .B2(n8253), .A(n8168), .ZN(n8154) );
  NAND2_X1 U9793 ( .A1(n8154), .A2(n9322), .ZN(n8156) );
  NAND4_X1 U9794 ( .A1(n8254), .A2(n9176), .A3(n8168), .A4(n9523), .ZN(n8155)
         );
  OAI211_X1 U9795 ( .C1(n8171), .C2(n9322), .A(n8156), .B(n8155), .ZN(n8157)
         );
  NAND2_X1 U9796 ( .A1(n8157), .A2(n9323), .ZN(n8159) );
  MUX2_X1 U9797 ( .A(n8286), .B(n8183), .S(n8168), .Z(n8158) );
  MUX2_X1 U9798 ( .A(n8179), .B(n8184), .S(n8171), .Z(n8160) );
  INV_X1 U9799 ( .A(n8165), .ZN(n8161) );
  INV_X1 U9800 ( .A(n8164), .ZN(n8294) );
  OAI21_X1 U9801 ( .B1(n8161), .B2(n8185), .A(n8294), .ZN(n8170) );
  INV_X1 U9802 ( .A(n8259), .ZN(n8331) );
  MUX2_X1 U9803 ( .A(n8185), .B(n8173), .S(n8171), .Z(n8162) );
  NAND2_X1 U9804 ( .A1(n8289), .A2(n8162), .ZN(n8163) );
  NOR2_X1 U9805 ( .A1(n8164), .A2(n8163), .ZN(n8176) );
  NAND3_X1 U9806 ( .A1(n8176), .A2(n8179), .A3(n8172), .ZN(n8167) );
  NAND2_X1 U9807 ( .A1(n8165), .A2(n9499), .ZN(n8166) );
  OAI211_X1 U9808 ( .C1(n8331), .C2(n8289), .A(n8167), .B(n8166), .ZN(n8169)
         );
  MUX2_X1 U9809 ( .A(n8170), .B(n8169), .S(n8168), .Z(n8178) );
  NAND3_X1 U9810 ( .A1(n8172), .A2(n8171), .A3(n8184), .ZN(n8174) );
  NAND3_X1 U9811 ( .A1(n8174), .A2(n8173), .A3(n8185), .ZN(n8175) );
  AND2_X1 U9812 ( .A1(n8176), .A2(n8175), .ZN(n8177) );
  OR2_X1 U9813 ( .A1(n9499), .A2(n8185), .ZN(n8180) );
  AND2_X1 U9814 ( .A1(n8180), .A2(n8179), .ZN(n8188) );
  NAND2_X1 U9815 ( .A1(n8286), .A2(n8181), .ZN(n8182) );
  NAND3_X1 U9816 ( .A1(n8184), .A2(n8183), .A3(n8182), .ZN(n8187) );
  AND2_X1 U9817 ( .A1(n9499), .A2(n8185), .ZN(n8186) );
  AOI21_X1 U9818 ( .B1(n8188), .B2(n8187), .A(n8186), .ZN(n8288) );
  INV_X1 U9819 ( .A(n8188), .ZN(n8291) );
  INV_X1 U9820 ( .A(n8189), .ZN(n8194) );
  NAND3_X1 U9821 ( .A1(n8191), .A2(n8190), .A3(n8332), .ZN(n8192) );
  NAND3_X1 U9822 ( .A1(n8194), .A2(n8193), .A3(n8192), .ZN(n8196) );
  AOI21_X1 U9823 ( .B1(n8196), .B2(n8195), .A(n4621), .ZN(n8199) );
  INV_X1 U9824 ( .A(n8276), .ZN(n8198) );
  OAI21_X1 U9825 ( .B1(n8199), .B2(n8198), .A(n8197), .ZN(n8216) );
  AND2_X1 U9826 ( .A1(n8239), .A2(n4475), .ZN(n8200) );
  NOR2_X1 U9827 ( .A1(n8201), .A2(n8200), .ZN(n8244) );
  INV_X1 U9828 ( .A(n8221), .ZN(n8208) );
  INV_X1 U9829 ( .A(n8202), .ZN(n8207) );
  INV_X1 U9830 ( .A(n8203), .ZN(n8205) );
  NAND2_X1 U9831 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  NAND4_X1 U9832 ( .A1(n8222), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8228)
         );
  NOR2_X1 U9833 ( .A1(n8228), .A2(n8209), .ZN(n8210) );
  NAND2_X1 U9834 ( .A1(n8231), .A2(n8210), .ZN(n8213) );
  INV_X1 U9835 ( .A(n9479), .ZN(n8211) );
  OR2_X1 U9836 ( .A1(n8212), .A2(n8211), .ZN(n8217) );
  NOR2_X1 U9837 ( .A1(n8213), .A2(n8217), .ZN(n8214) );
  AND2_X1 U9838 ( .A1(n8244), .A2(n8214), .ZN(n8277) );
  INV_X1 U9839 ( .A(n8277), .ZN(n8215) );
  AOI21_X1 U9840 ( .B1(n8263), .B2(n8216), .A(n8215), .ZN(n8247) );
  INV_X1 U9841 ( .A(n8217), .ZN(n8232) );
  INV_X1 U9842 ( .A(n8228), .ZN(n8225) );
  INV_X1 U9843 ( .A(n8218), .ZN(n8224) );
  OAI21_X1 U9844 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8223) );
  AOI22_X1 U9845 ( .A1(n8225), .A2(n8224), .B1(n8223), .B2(n8222), .ZN(n8226)
         );
  OAI211_X1 U9846 ( .C1(n8229), .C2(n8228), .A(n8227), .B(n8226), .ZN(n8230)
         );
  NAND3_X1 U9847 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(n8238) );
  INV_X1 U9848 ( .A(n8233), .ZN(n8235) );
  OR2_X1 U9849 ( .A1(n8235), .A2(n8234), .ZN(n8237) );
  AND4_X1 U9850 ( .A1(n8299), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n8240)
         );
  NAND2_X1 U9851 ( .A1(n8240), .A2(n8239), .ZN(n8243) );
  INV_X1 U9852 ( .A(n8241), .ZN(n8242) );
  AOI21_X1 U9853 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8281) );
  INV_X1 U9854 ( .A(n8281), .ZN(n8246) );
  OAI21_X1 U9855 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8252) );
  INV_X1 U9856 ( .A(n8248), .ZN(n8280) );
  INV_X1 U9857 ( .A(n8249), .ZN(n8250) );
  AOI211_X1 U9858 ( .C1(n8252), .C2(n8280), .A(n8251), .B(n8250), .ZN(n8256)
         );
  AND2_X1 U9859 ( .A1(n8254), .A2(n8253), .ZN(n8287) );
  INV_X1 U9860 ( .A(n8287), .ZN(n8255) );
  OR4_X1 U9861 ( .A1(n8291), .A2(n9315), .A3(n8256), .A4(n8255), .ZN(n8257) );
  AOI21_X1 U9862 ( .B1(n8288), .B2(n8257), .A(n8330), .ZN(n8261) );
  AOI21_X1 U9863 ( .B1(n8258), .B2(n9290), .A(n8342), .ZN(n8334) );
  INV_X1 U9864 ( .A(n8334), .ZN(n8260) );
  OAI21_X1 U9865 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8262) );
  XNOR2_X1 U9866 ( .A(n8262), .B(n9283), .ZN(n8339) );
  INV_X1 U9867 ( .A(n8263), .ZN(n8279) );
  INV_X1 U9868 ( .A(n8265), .ZN(n8274) );
  NAND2_X1 U9869 ( .A1(n8267), .A2(n8266), .ZN(n8270) );
  NAND3_X1 U9870 ( .A1(n8270), .A2(n8269), .A3(n8268), .ZN(n8273) );
  INV_X1 U9871 ( .A(n8271), .ZN(n8272) );
  AOI21_X1 U9872 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8275) );
  AOI21_X1 U9873 ( .B1(n4477), .B2(n8276), .A(n8275), .ZN(n8278) );
  OAI21_X1 U9874 ( .B1(n8279), .B2(n8278), .A(n8277), .ZN(n8282) );
  NAND3_X1 U9875 ( .A1(n8282), .A2(n8281), .A3(n8280), .ZN(n8283) );
  NAND2_X1 U9876 ( .A1(n8284), .A2(n8283), .ZN(n8285) );
  NAND3_X1 U9877 ( .A1(n8287), .A2(n8286), .A3(n8285), .ZN(n8290) );
  OAI211_X1 U9878 ( .C1(n8291), .C2(n8290), .A(n8289), .B(n8288), .ZN(n8293)
         );
  AOI211_X1 U9879 ( .C1(n8294), .C2(n8293), .A(n8292), .B(n8342), .ZN(n8297)
         );
  OR3_X1 U9880 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n8337) );
  INV_X1 U9881 ( .A(n9365), .ZN(n8326) );
  NAND2_X1 U9882 ( .A1(n8299), .A2(n8298), .ZN(n9420) );
  NOR4_X1 U9883 ( .A1(n6735), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n8307)
         );
  NAND4_X1 U9884 ( .A1(n8307), .A2(n8306), .A3(n4780), .A4(n8305), .ZN(n8312)
         );
  INV_X1 U9885 ( .A(n8308), .ZN(n8309) );
  NOR4_X1 U9886 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n8316)
         );
  NAND4_X1 U9887 ( .A1(n8316), .A2(n8315), .A3(n8314), .A4(n8313), .ZN(n8318)
         );
  NOR4_X1 U9888 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n8321)
         );
  NAND3_X1 U9889 ( .A1(n9481), .A2(n8322), .A3(n8321), .ZN(n8323) );
  NOR4_X1 U9890 ( .A1(n9420), .A2(n9430), .A3(n9452), .A4(n8323), .ZN(n8324)
         );
  XNOR2_X1 U9891 ( .A(n9537), .B(n9409), .ZN(n9392) );
  NAND4_X1 U9892 ( .A1(n7733), .A2(n9408), .A3(n8324), .A4(n9392), .ZN(n8325)
         );
  NOR4_X1 U9893 ( .A1(n7715), .A2(n9342), .A3(n8326), .A4(n8325), .ZN(n8327)
         );
  NAND3_X1 U9894 ( .A1(n8327), .A2(n9298), .A3(n9323), .ZN(n8328) );
  NOR4_X1 U9895 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n8333)
         );
  AOI21_X1 U9896 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8335) );
  MUX2_X1 U9897 ( .A(n8337), .B(n8336), .S(n8335), .Z(n8338) );
  OAI21_X1 U9898 ( .B1(n8340), .B2(n8339), .A(n8338), .ZN(n8344) );
  NOR4_X1 U9899 ( .A1(n8345), .A2(n8350), .A3(n8342), .A4(n8341), .ZN(n8343)
         );
  AOI211_X1 U9900 ( .C1(n8346), .C2(n8345), .A(n8344), .B(n8343), .ZN(n8353)
         );
  NAND4_X1 U9901 ( .A1(n8348), .A2(n9804), .A3(n8347), .A4(n9703), .ZN(n8349)
         );
  OAI211_X1 U9902 ( .C1(n8350), .C2(n8352), .A(n8349), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8351) );
  OAI21_X1 U9903 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(P1_U3240) );
  XNOR2_X1 U9904 ( .A(n8354), .B(n8559), .ZN(n8355) );
  AOI222_X1 U9905 ( .A1(n8920), .A2(n8355), .B1(n8692), .B2(n8917), .C1(n8694), 
        .C2(n8915), .ZN(n8952) );
  INV_X1 U9906 ( .A(n8770), .ZN(n8358) );
  INV_X1 U9907 ( .A(n8356), .ZN(n8357) );
  AOI21_X1 U9908 ( .B1(n8949), .B2(n8358), .A(n8357), .ZN(n8950) );
  INV_X1 U9909 ( .A(n8359), .ZN(n8360) );
  AOI22_X1 U9910 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n8931), .B1(n8360), .B2(
        n8929), .ZN(n8361) );
  OAI21_X1 U9911 ( .B1(n8033), .B2(n8908), .A(n8361), .ZN(n8364) );
  OAI21_X1 U9912 ( .B1(n8931), .B2(n8952), .A(n8365), .ZN(P2_U3268) );
  INV_X1 U9913 ( .A(n8371), .ZN(n9054) );
  OAI222_X1 U9914 ( .A1(n9609), .A2(n8367), .B1(n9613), .B2(n9054), .C1(
        P1_U3084), .C2(n8366), .ZN(P1_U3323) );
  NAND2_X1 U9915 ( .A1(n8371), .A2(n8370), .ZN(n8373) );
  INV_X1 U9916 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9055) );
  OR2_X1 U9917 ( .A1(n4947), .A2(n9055), .ZN(n8372) );
  INV_X1 U9918 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U9919 ( .A1(n4995), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U9920 ( .A1(n4964), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8374) );
  OAI211_X1 U9921 ( .C1(n5358), .C2(n8376), .A(n8375), .B(n8374), .ZN(n8755)
         );
  NAND2_X1 U9922 ( .A1(n9627), .A2(n8378), .ZN(n8569) );
  XNOR2_X1 U9923 ( .A(n8380), .B(n8379), .ZN(n8584) );
  NAND2_X1 U9924 ( .A1(n8572), .A2(n4857), .ZN(n8411) );
  INV_X1 U9925 ( .A(n8914), .ZN(n8400) );
  NOR4_X1 U9926 ( .A1(n9894), .A2(n6278), .A3(n8383), .A4(n4312), .ZN(n8385)
         );
  NAND3_X1 U9927 ( .A1(n8385), .A2(n8384), .A3(n6543), .ZN(n8388) );
  NOR4_X1 U9928 ( .A1(n8388), .A2(n8460), .A3(n8387), .A4(n8386), .ZN(n8392)
         );
  NAND4_X1 U9929 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n8393)
         );
  NOR4_X1 U9930 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n8398)
         );
  NAND4_X1 U9931 ( .A1(n8504), .A2(n8498), .A3(n8398), .A4(n8397), .ZN(n8399)
         );
  NOR4_X1 U9932 ( .A1(n8401), .A2(n8400), .A3(n4311), .A4(n8399), .ZN(n8402)
         );
  NAND4_X1 U9933 ( .A1(n8048), .A2(n8880), .A3(n8046), .A4(n8402), .ZN(n8403)
         );
  NOR4_X1 U9934 ( .A1(n8788), .A2(n8820), .A3(n8518), .A4(n8403), .ZN(n8404)
         );
  INV_X1 U9935 ( .A(n8802), .ZN(n8545) );
  NAND4_X1 U9936 ( .A1(n8405), .A2(n8404), .A3(n8554), .A4(n8545), .ZN(n8406)
         );
  NOR4_X1 U9937 ( .A1(n8411), .A2(n4356), .A3(n8407), .A4(n8406), .ZN(n8408)
         );
  XOR2_X1 U9938 ( .A(n8408), .B(n5290), .Z(n8410) );
  AOI22_X1 U9939 ( .A1(n8410), .A2(n8409), .B1(n8580), .B2(n4312), .ZN(n8577)
         );
  NAND3_X1 U9940 ( .A1(n5519), .A2(n5290), .A3(n8433), .ZN(n8570) );
  MUX2_X1 U9941 ( .A(n4356), .B(n8411), .S(n8570), .Z(n8575) );
  AND2_X1 U9942 ( .A1(n8965), .A2(n8822), .ZN(n8412) );
  OAI21_X1 U9943 ( .B1(n8788), .B2(n8412), .A(n8570), .ZN(n8549) );
  NAND2_X1 U9944 ( .A1(n8511), .A2(n8910), .ZN(n8415) );
  INV_X1 U9945 ( .A(n8413), .ZN(n8414) );
  INV_X1 U9946 ( .A(n8570), .ZN(n8556) );
  MUX2_X1 U9947 ( .A(n8415), .B(n8414), .S(n8556), .Z(n8416) );
  INV_X1 U9948 ( .A(n8416), .ZN(n8510) );
  NAND2_X1 U9949 ( .A1(n8483), .A2(n8417), .ZN(n8421) );
  OAI211_X1 U9950 ( .C1(n8472), .C2(n8419), .A(n8478), .B(n8418), .ZN(n8420)
         );
  MUX2_X1 U9951 ( .A(n8421), .B(n8420), .S(n8570), .Z(n8422) );
  INV_X1 U9952 ( .A(n8422), .ZN(n8477) );
  INV_X1 U9953 ( .A(n8423), .ZN(n8475) );
  NAND2_X1 U9954 ( .A1(n8426), .A2(n8424), .ZN(n8427) );
  INV_X1 U9955 ( .A(n8449), .ZN(n8425) );
  MUX2_X1 U9956 ( .A(n8427), .B(n8425), .S(n8570), .Z(n8451) );
  NAND2_X1 U9957 ( .A1(n8451), .A2(n8426), .ZN(n8432) );
  INV_X1 U9958 ( .A(n8427), .ZN(n8429) );
  NAND2_X1 U9959 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  INV_X1 U9960 ( .A(n8459), .ZN(n8430) );
  AOI21_X1 U9961 ( .B1(n8432), .B2(n8431), .A(n8430), .ZN(n8439) );
  AND2_X1 U9962 ( .A1(n8441), .A2(n8433), .ZN(n8435) );
  OAI211_X1 U9963 ( .C1(n8435), .C2(n6541), .A(n8434), .B(n8440), .ZN(n8436)
         );
  NAND3_X1 U9964 ( .A1(n8436), .A2(n8443), .A3(n8570), .ZN(n8437) );
  NAND2_X1 U9965 ( .A1(n8437), .A2(n6543), .ZN(n8438) );
  OAI22_X1 U9966 ( .A1(n8439), .A2(n8556), .B1(n8438), .B2(n8451), .ZN(n8447)
         );
  NAND2_X1 U9967 ( .A1(n8441), .A2(n8440), .ZN(n8444) );
  NAND3_X1 U9968 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8445) );
  NAND3_X1 U9969 ( .A1(n8445), .A2(n8556), .A3(n8434), .ZN(n8446) );
  NAND3_X1 U9970 ( .A1(n8447), .A2(n8452), .A3(n8446), .ZN(n8457) );
  AOI22_X1 U9971 ( .A1(n8451), .A2(n8450), .B1(n8449), .B2(n8448), .ZN(n8454)
         );
  INV_X1 U9972 ( .A(n8452), .ZN(n8453) );
  OAI21_X1 U9973 ( .B1(n8454), .B2(n8453), .A(n8556), .ZN(n8455) );
  NAND3_X1 U9974 ( .A1(n8457), .A2(n8456), .A3(n8455), .ZN(n8471) );
  OAI21_X1 U9975 ( .B1(n8460), .B2(n8459), .A(n8458), .ZN(n8461) );
  MUX2_X1 U9976 ( .A(n8462), .B(n8461), .S(n8556), .Z(n8464) );
  NOR2_X1 U9977 ( .A1(n8464), .A2(n8463), .ZN(n8470) );
  INV_X1 U9978 ( .A(n8465), .ZN(n8468) );
  INV_X1 U9979 ( .A(n8466), .ZN(n8467) );
  MUX2_X1 U9980 ( .A(n8468), .B(n8467), .S(n8556), .Z(n8469) );
  AOI21_X1 U9981 ( .B1(n8471), .B2(n8470), .A(n8469), .ZN(n8474) );
  INV_X1 U9982 ( .A(n8472), .ZN(n8473) );
  OAI21_X1 U9983 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8476) );
  NAND2_X1 U9984 ( .A1(n8477), .A2(n8476), .ZN(n8485) );
  NAND3_X1 U9985 ( .A1(n8485), .A2(n4348), .A3(n8478), .ZN(n8479) );
  NAND2_X1 U9986 ( .A1(n8479), .A2(n8484), .ZN(n8482) );
  INV_X1 U9987 ( .A(n8480), .ZN(n8481) );
  AOI21_X1 U9988 ( .B1(n8482), .B2(n8489), .A(n8481), .ZN(n8492) );
  NAND3_X1 U9989 ( .A1(n8485), .A2(n8484), .A3(n8483), .ZN(n8486) );
  NAND2_X1 U9990 ( .A1(n8486), .A2(n4348), .ZN(n8490) );
  INV_X1 U9991 ( .A(n8487), .ZN(n8488) );
  AOI21_X1 U9992 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8491) );
  INV_X1 U9993 ( .A(n8493), .ZN(n8496) );
  INV_X1 U9994 ( .A(n8494), .ZN(n8495) );
  MUX2_X1 U9995 ( .A(n8496), .B(n8495), .S(n8556), .Z(n8497) );
  NAND2_X1 U9996 ( .A1(n8700), .A2(n8556), .ZN(n8501) );
  NAND2_X1 U9997 ( .A1(n8499), .A2(n8570), .ZN(n8500) );
  MUX2_X1 U9998 ( .A(n8501), .B(n8500), .S(n9015), .Z(n8502) );
  MUX2_X1 U9999 ( .A(n4352), .B(n8505), .S(n8570), .Z(n8506) );
  NAND3_X1 U10000 ( .A1(n8508), .A2(n8507), .A3(n8506), .ZN(n8509) );
  NAND3_X1 U10001 ( .A1(n8510), .A2(n8509), .A3(n8524), .ZN(n8525) );
  NAND2_X1 U10002 ( .A1(n8525), .A2(n8511), .ZN(n8512) );
  NAND2_X1 U10003 ( .A1(n8512), .A2(n8526), .ZN(n8513) );
  NAND3_X1 U10004 ( .A1(n8513), .A2(n8528), .A3(n8522), .ZN(n8514) );
  NAND3_X1 U10005 ( .A1(n8514), .A2(n8532), .A3(n8527), .ZN(n8515) );
  NAND2_X1 U10006 ( .A1(n8515), .A2(n8529), .ZN(n8517) );
  NAND2_X1 U10007 ( .A1(n8834), .A2(n8556), .ZN(n8516) );
  INV_X1 U10008 ( .A(n8519), .ZN(n8520) );
  INV_X1 U10009 ( .A(n8521), .ZN(n8536) );
  INV_X1 U10010 ( .A(n8522), .ZN(n8523) );
  AOI21_X1 U10011 ( .B1(n8525), .B2(n8524), .A(n8523), .ZN(n8531) );
  NAND2_X1 U10012 ( .A1(n8527), .A2(n8526), .ZN(n8530) );
  OAI211_X1 U10013 ( .C1(n8531), .C2(n8530), .A(n8529), .B(n8528), .ZN(n8534)
         );
  NAND3_X1 U10014 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n8535) );
  NAND3_X1 U10015 ( .A1(n8537), .A2(n8536), .A3(n8535), .ZN(n8539) );
  INV_X1 U10016 ( .A(n8542), .ZN(n8538) );
  AOI21_X1 U10017 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n8547) );
  AOI21_X1 U10018 ( .B1(n8542), .B2(n8541), .A(n8556), .ZN(n8546) );
  OR2_X1 U10019 ( .A1(n8543), .A2(n8556), .ZN(n8544) );
  OAI211_X1 U10020 ( .C1(n8547), .C2(n8546), .A(n8545), .B(n8544), .ZN(n8548)
         );
  NAND2_X1 U10021 ( .A1(n8549), .A2(n8548), .ZN(n8553) );
  AOI21_X1 U10022 ( .B1(n8552), .B2(n8550), .A(n8570), .ZN(n8551) );
  OAI21_X1 U10023 ( .B1(n8555), .B2(n8570), .A(n8554), .ZN(n8561) );
  AND2_X1 U10024 ( .A1(n8954), .A2(n8789), .ZN(n8557) );
  MUX2_X1 U10025 ( .A(n8557), .B(n4372), .S(n8556), .Z(n8558) );
  NOR2_X1 U10026 ( .A1(n8559), .A2(n8558), .ZN(n8560) );
  MUX2_X1 U10027 ( .A(n8563), .B(n8562), .S(n8570), .Z(n8564) );
  MUX2_X1 U10028 ( .A(n8567), .B(n8566), .S(n8570), .Z(n8568) );
  MUX2_X1 U10029 ( .A(n8572), .B(n8571), .S(n8570), .Z(n8573) );
  OAI21_X1 U10030 ( .B1(n8575), .B2(n8574), .A(n8573), .ZN(n8576) );
  AND2_X1 U10031 ( .A1(n8576), .A2(n4316), .ZN(n8578) );
  INV_X1 U10032 ( .A(n8578), .ZN(n8581) );
  NOR3_X1 U10033 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n8582) );
  INV_X1 U10034 ( .A(n6359), .ZN(n8585) );
  NAND3_X1 U10035 ( .A1(n8586), .A2(n8585), .A3(n8915), .ZN(n8587) );
  OAI211_X1 U10036 ( .C1(n8588), .C2(n8590), .A(n8587), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8589) );
  NAND2_X1 U10037 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  XOR2_X1 U10038 ( .A(n8594), .B(n8593), .Z(n8599) );
  AOI22_X1 U10039 ( .A1(n8682), .A2(n8697), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8596) );
  NAND2_X1 U10040 ( .A1(n8623), .A2(n8882), .ZN(n8595) );
  OAI211_X1 U10041 ( .C1(n8633), .C2(n8845), .A(n8596), .B(n8595), .ZN(n8597)
         );
  AOI21_X1 U10042 ( .B1(n8848), .B2(n8688), .A(n8597), .ZN(n8598) );
  OAI21_X1 U10043 ( .B1(n8599), .B2(n8690), .A(n8598), .ZN(P2_U3218) );
  NAND2_X1 U10044 ( .A1(n8601), .A2(n8600), .ZN(n8603) );
  XOR2_X1 U10045 ( .A(n8603), .B(n8602), .Z(n8609) );
  AOI22_X1 U10046 ( .A1(n8623), .A2(n8698), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8605) );
  NAND2_X1 U10047 ( .A1(n8682), .A2(n8881), .ZN(n8604) );
  OAI211_X1 U10048 ( .C1(n8633), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8607)
         );
  AOI21_X1 U10049 ( .B1(n8996), .B2(n8688), .A(n8607), .ZN(n8608) );
  OAI21_X1 U10050 ( .B1(n8609), .B2(n8690), .A(n8608), .ZN(P2_U3221) );
  XOR2_X1 U10051 ( .A(n8611), .B(n8610), .Z(n8613) );
  NAND2_X1 U10052 ( .A1(n8613), .A2(n8612), .ZN(n8620) );
  AOI21_X1 U10053 ( .B1(n8688), .B2(n8615), .A(n8614), .ZN(n8619) );
  AOI22_X1 U10054 ( .A1(n8623), .A2(n8708), .B1(n8682), .B2(n8706), .ZN(n8618)
         );
  NAND2_X1 U10055 ( .A1(n8680), .A2(n8616), .ZN(n8617) );
  NAND4_X1 U10056 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(
        P2_U3223) );
  XNOR2_X1 U10057 ( .A(n8621), .B(n8622), .ZN(n8628) );
  AOI22_X1 U10058 ( .A1(n8682), .A2(n8882), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8625) );
  NAND2_X1 U10059 ( .A1(n8623), .A2(n8881), .ZN(n8624) );
  OAI211_X1 U10060 ( .C1(n8633), .C2(n8874), .A(n8625), .B(n8624), .ZN(n8626)
         );
  AOI21_X1 U10061 ( .B1(n8985), .B2(n8688), .A(n8626), .ZN(n8627) );
  OAI21_X1 U10062 ( .B1(n8628), .B2(n8690), .A(n8627), .ZN(P2_U3225) );
  XNOR2_X1 U10063 ( .A(n8631), .B(n8630), .ZN(n8632) );
  XNOR2_X1 U10064 ( .A(n8629), .B(n8632), .ZN(n8640) );
  NOR2_X1 U10065 ( .A1(n8633), .A2(n8807), .ZN(n8638) );
  INV_X1 U10066 ( .A(n8634), .ZN(n8636) );
  AOI22_X1 U10067 ( .A1(n8695), .A2(n8917), .B1(n8697), .B2(n8915), .ZN(n8804)
         );
  OAI22_X1 U10068 ( .A1(n8636), .A2(n8804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8635), .ZN(n8637) );
  AOI211_X1 U10069 ( .C1(n8965), .C2(n8688), .A(n8638), .B(n8637), .ZN(n8639)
         );
  OAI21_X1 U10070 ( .B1(n8640), .B2(n8690), .A(n8639), .ZN(P2_U3227) );
  XNOR2_X1 U10071 ( .A(n8642), .B(n8641), .ZN(n8649) );
  NAND2_X1 U10072 ( .A1(n8680), .A2(n8643), .ZN(n8645) );
  AOI22_X1 U10073 ( .A1(n8682), .A2(n8698), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8644) );
  OAI211_X1 U10074 ( .C1(n8646), .C2(n8685), .A(n8645), .B(n8644), .ZN(n8647)
         );
  AOI21_X1 U10075 ( .B1(n9007), .B2(n8688), .A(n8647), .ZN(n8648) );
  OAI21_X1 U10076 ( .B1(n8649), .B2(n8690), .A(n8648), .ZN(P2_U3230) );
  XNOR2_X1 U10077 ( .A(n8650), .B(n8651), .ZN(n8656) );
  NAND2_X1 U10078 ( .A1(n8680), .A2(n8816), .ZN(n8653) );
  AOI22_X1 U10079 ( .A1(n8682), .A2(n8696), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8652) );
  OAI211_X1 U10080 ( .C1(n8864), .C2(n8685), .A(n8653), .B(n8652), .ZN(n8654)
         );
  AOI21_X1 U10081 ( .B1(n8968), .B2(n8688), .A(n8654), .ZN(n8655) );
  OAI21_X1 U10082 ( .B1(n8656), .B2(n8690), .A(n8655), .ZN(P2_U3231) );
  XNOR2_X1 U10083 ( .A(n8658), .B(n8657), .ZN(n8664) );
  NAND2_X1 U10084 ( .A1(n8680), .A2(n8893), .ZN(n8660) );
  AOI22_X1 U10085 ( .A1(n8682), .A2(n8897), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8659) );
  OAI211_X1 U10086 ( .C1(n8661), .C2(n8685), .A(n8660), .B(n8659), .ZN(n8662)
         );
  AOI21_X1 U10087 ( .B1(n8990), .B2(n8688), .A(n8662), .ZN(n8663) );
  OAI21_X1 U10088 ( .B1(n8664), .B2(n8690), .A(n8663), .ZN(P2_U3235) );
  NAND2_X1 U10089 ( .A1(n8666), .A2(n8665), .ZN(n8670) );
  XOR2_X1 U10090 ( .A(n8668), .B(n8667), .Z(n8669) );
  XNOR2_X1 U10091 ( .A(n8670), .B(n8669), .ZN(n8677) );
  NOR2_X1 U10092 ( .A1(n8685), .A2(n8862), .ZN(n8674) );
  OAI22_X1 U10093 ( .A1(n8672), .A2(n8864), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8671), .ZN(n8673) );
  AOI211_X1 U10094 ( .C1(n8680), .C2(n8856), .A(n8674), .B(n8673), .ZN(n8676)
         );
  NAND2_X1 U10095 ( .A1(n8980), .A2(n8688), .ZN(n8675) );
  OAI211_X1 U10096 ( .C1(n8677), .C2(n8690), .A(n8676), .B(n8675), .ZN(
        P2_U3237) );
  XNOR2_X1 U10097 ( .A(n8679), .B(n8678), .ZN(n8691) );
  NAND2_X1 U10098 ( .A1(n8680), .A2(n8906), .ZN(n8684) );
  NOR2_X1 U10099 ( .A1(n8681), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8747) );
  AOI21_X1 U10100 ( .B1(n8682), .B2(n8918), .A(n8747), .ZN(n8683) );
  OAI211_X1 U10101 ( .C1(n8686), .C2(n8685), .A(n8684), .B(n8683), .ZN(n8687)
         );
  AOI21_X1 U10102 ( .B1(n9000), .B2(n8688), .A(n8687), .ZN(n8689) );
  OAI21_X1 U10103 ( .B1(n8691), .B2(n8690), .A(n8689), .ZN(P2_U3240) );
  MUX2_X1 U10104 ( .A(n8755), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8712), .Z(
        P2_U3583) );
  MUX2_X1 U10105 ( .A(n8692), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8712), .Z(
        P2_U3581) );
  MUX2_X1 U10106 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8693), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10107 ( .A(n8694), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8712), .Z(
        P2_U3579) );
  MUX2_X1 U10108 ( .A(n8695), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8712), .Z(
        P2_U3578) );
  MUX2_X1 U10109 ( .A(n8696), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8712), .Z(
        P2_U3577) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8697), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10111 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8882), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10112 ( .A(n8897), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8712), .Z(
        P2_U3573) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8881), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8918), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8698), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8916), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8699), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10118 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8700), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8701), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8702), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10121 ( .A(n8703), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8712), .Z(
        P2_U3564) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8704), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8705), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10124 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8706), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10125 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8707), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10126 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8708), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10127 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8709), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10128 ( .A(n8710), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8712), .Z(
        P2_U3557) );
  MUX2_X1 U10129 ( .A(n8711), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8712), .Z(
        P2_U3556) );
  MUX2_X1 U10130 ( .A(n6534), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8712), .Z(
        P2_U3555) );
  MUX2_X1 U10131 ( .A(n6531), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8712), .Z(
        P2_U3554) );
  MUX2_X1 U10132 ( .A(n6277), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8712), .Z(
        P2_U3553) );
  OAI21_X1 U10133 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8716) );
  NAND2_X1 U10134 ( .A1(n8716), .A2(n9868), .ZN(n8726) );
  INV_X1 U10135 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8718) );
  OAI21_X1 U10136 ( .B1(n8745), .B2(n8718), .A(n8717), .ZN(n8719) );
  AOI21_X1 U10137 ( .B1(n8750), .B2(n8720), .A(n8719), .ZN(n8725) );
  OAI211_X1 U10138 ( .C1(n8723), .C2(n8722), .A(n9867), .B(n8721), .ZN(n8724)
         );
  NAND3_X1 U10139 ( .A1(n8726), .A2(n8725), .A3(n8724), .ZN(P2_U3261) );
  OAI211_X1 U10140 ( .C1(n8729), .C2(n8728), .A(n9867), .B(n8727), .ZN(n8740)
         );
  NOR2_X1 U10141 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8730), .ZN(n8731) );
  AOI21_X1 U10142 ( .B1(n9873), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8731), .ZN(
        n8739) );
  NAND2_X1 U10143 ( .A1(n8750), .A2(n8732), .ZN(n8738) );
  AOI21_X1 U10144 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8736) );
  NAND2_X1 U10145 ( .A1(n9868), .A2(n8736), .ZN(n8737) );
  NAND4_X1 U10146 ( .A1(n8740), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(
        P2_U3262) );
  AOI21_X1 U10147 ( .B1(n8742), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8741), .ZN(
        n8753) );
  XNOR2_X1 U10148 ( .A(n8744), .B(n8743), .ZN(n8748) );
  NOR2_X1 U10149 ( .A1(n8745), .A2(n10019), .ZN(n8746) );
  AOI211_X1 U10150 ( .C1(n9868), .C2(n8748), .A(n8747), .B(n8746), .ZN(n8752)
         );
  NAND2_X1 U10151 ( .A1(n8750), .A2(n8749), .ZN(n8751) );
  OAI211_X1 U10152 ( .C1(n8753), .C2(n9871), .A(n8752), .B(n8751), .ZN(
        P2_U3263) );
  INV_X1 U10153 ( .A(n9627), .ZN(n8762) );
  INV_X1 U10154 ( .A(n8754), .ZN(n8756) );
  NAND2_X1 U10155 ( .A1(n8756), .A2(n8755), .ZN(n8939) );
  INV_X1 U10156 ( .A(n8939), .ZN(n9626) );
  NAND2_X1 U10157 ( .A1(n8933), .A2(n9626), .ZN(n8763) );
  NAND2_X1 U10158 ( .A1(n8931), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8757) );
  OAI211_X1 U10159 ( .C1(n8941), .C2(n8908), .A(n8763), .B(n8757), .ZN(n8758)
         );
  AOI21_X1 U10160 ( .B1(n8938), .B2(n6814), .A(n8758), .ZN(n8759) );
  INV_X1 U10161 ( .A(n8759), .ZN(P2_U3265) );
  OAI21_X1 U10162 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n9624) );
  INV_X1 U10163 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8764) );
  OAI21_X1 U10164 ( .B1(n8933), .B2(n8764), .A(n8763), .ZN(n8765) );
  AOI21_X1 U10165 ( .B1(n9627), .B2(n8926), .A(n8765), .ZN(n8766) );
  OAI21_X1 U10166 ( .B1(n9624), .B2(n8850), .A(n8766), .ZN(P2_U3266) );
  OAI21_X1 U10167 ( .B1(n8768), .B2(n8774), .A(n8767), .ZN(n8769) );
  INV_X1 U10168 ( .A(n8769), .ZN(n8958) );
  AOI21_X1 U10169 ( .B1(n8954), .B2(n8790), .A(n8770), .ZN(n8955) );
  AOI22_X1 U10170 ( .A1(n8931), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8771), .B2(
        n8929), .ZN(n8772) );
  OAI21_X1 U10171 ( .B1(n8773), .B2(n8908), .A(n8772), .ZN(n8781) );
  AOI21_X1 U10172 ( .B1(n4362), .B2(n8774), .A(n8859), .ZN(n8779) );
  OAI22_X1 U10173 ( .A1(n8776), .A2(n8863), .B1(n8775), .B2(n8861), .ZN(n8777)
         );
  AOI21_X1 U10174 ( .B1(n8779), .B2(n8778), .A(n8777), .ZN(n8957) );
  NOR2_X1 U10175 ( .A1(n8957), .A2(n8931), .ZN(n8780) );
  AOI211_X1 U10176 ( .C1(n8955), .C2(n6814), .A(n8781), .B(n8780), .ZN(n8782)
         );
  OAI21_X1 U10177 ( .B1(n8958), .B2(n8924), .A(n8782), .ZN(P2_U3269) );
  OAI21_X1 U10178 ( .B1(n8784), .B2(n8788), .A(n8783), .ZN(n8785) );
  INV_X1 U10179 ( .A(n8785), .ZN(n8962) );
  INV_X1 U10180 ( .A(n8806), .ZN(n8792) );
  INV_X1 U10181 ( .A(n8790), .ZN(n8791) );
  AOI211_X1 U10182 ( .C1(n8961), .C2(n8792), .A(n9957), .B(n8791), .ZN(n8960)
         );
  INV_X1 U10183 ( .A(n8960), .ZN(n8795) );
  INV_X1 U10184 ( .A(n8793), .ZN(n8794) );
  OAI22_X1 U10185 ( .A1(n8795), .A2(n5290), .B1(n8844), .B2(n8794), .ZN(n8796)
         );
  OAI21_X1 U10186 ( .B1(n8959), .B2(n8796), .A(n8933), .ZN(n8798) );
  AOI22_X1 U10187 ( .A1(n8961), .A2(n8926), .B1(n8931), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U10188 ( .C1(n8962), .C2(n8924), .A(n8798), .B(n8797), .ZN(
        P2_U3270) );
  OAI21_X1 U10189 ( .B1(n8800), .B2(n8802), .A(n8799), .ZN(n8801) );
  INV_X1 U10190 ( .A(n8801), .ZN(n8967) );
  XNOR2_X1 U10191 ( .A(n8803), .B(n8802), .ZN(n8805) );
  OAI21_X1 U10192 ( .B1(n8805), .B2(n8859), .A(n8804), .ZN(n8963) );
  AOI211_X1 U10193 ( .C1(n8965), .C2(n8813), .A(n9957), .B(n8806), .ZN(n8964)
         );
  INV_X1 U10194 ( .A(n8964), .ZN(n8808) );
  OAI22_X1 U10195 ( .A1(n8808), .A2(n5290), .B1(n8844), .B2(n8807), .ZN(n8809)
         );
  OAI21_X1 U10196 ( .B1(n8963), .B2(n8809), .A(n8933), .ZN(n8811) );
  AOI22_X1 U10197 ( .A1(n8965), .A2(n8926), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8931), .ZN(n8810) );
  OAI211_X1 U10198 ( .C1(n8967), .C2(n8924), .A(n8811), .B(n8810), .ZN(
        P2_U3271) );
  XNOR2_X1 U10199 ( .A(n8812), .B(n8820), .ZN(n8972) );
  INV_X1 U10200 ( .A(n8842), .ZN(n8815) );
  INV_X1 U10201 ( .A(n8813), .ZN(n8814) );
  AOI21_X1 U10202 ( .B1(n8968), .B2(n8815), .A(n8814), .ZN(n8969) );
  AOI22_X1 U10203 ( .A1(n8931), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8816), .B2(
        n8929), .ZN(n8817) );
  OAI21_X1 U10204 ( .B1(n8818), .B2(n8908), .A(n8817), .ZN(n8827) );
  NOR2_X1 U10205 ( .A1(n8819), .A2(n8859), .ZN(n8825) );
  OAI21_X1 U10206 ( .B1(n8835), .B2(n8821), .A(n8820), .ZN(n8824) );
  OAI22_X1 U10207 ( .A1(n8822), .A2(n8863), .B1(n8864), .B2(n8861), .ZN(n8823)
         );
  AOI21_X1 U10208 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8971) );
  NOR2_X1 U10209 ( .A1(n8971), .A2(n8931), .ZN(n8826) );
  AOI211_X1 U10210 ( .C1(n8969), .C2(n6814), .A(n8827), .B(n8826), .ZN(n8828)
         );
  OAI21_X1 U10211 ( .B1(n8924), .B2(n8972), .A(n8828), .ZN(P2_U3272) );
  NAND2_X1 U10212 ( .A1(n8829), .A2(n8833), .ZN(n8830) );
  NAND2_X1 U10213 ( .A1(n8831), .A2(n8830), .ZN(n8973) );
  AOI21_X1 U10214 ( .B1(n8832), .B2(n8834), .A(n8833), .ZN(n8836) );
  OAI21_X1 U10215 ( .B1(n8836), .B2(n8835), .A(n8920), .ZN(n8841) );
  OAI22_X1 U10216 ( .A1(n8838), .A2(n8863), .B1(n8837), .B2(n8861), .ZN(n8839)
         );
  INV_X1 U10217 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U10218 ( .A1(n8841), .A2(n8840), .ZN(n8977) );
  AND2_X1 U10219 ( .A1(n8848), .A2(n8854), .ZN(n8843) );
  OR2_X1 U10220 ( .A1(n8843), .A2(n8842), .ZN(n8975) );
  OAI22_X1 U10221 ( .A1(n8933), .A2(n8846), .B1(n8845), .B2(n8844), .ZN(n8847)
         );
  AOI21_X1 U10222 ( .B1(n8848), .B2(n8926), .A(n8847), .ZN(n8849) );
  OAI21_X1 U10223 ( .B1(n8975), .B2(n8850), .A(n8849), .ZN(n8851) );
  AOI21_X1 U10224 ( .B1(n8977), .B2(n8933), .A(n8851), .ZN(n8852) );
  OAI21_X1 U10225 ( .B1(n8973), .B2(n8924), .A(n8852), .ZN(P2_U3273) );
  XNOR2_X1 U10226 ( .A(n8853), .B(n8860), .ZN(n8984) );
  INV_X1 U10227 ( .A(n8854), .ZN(n8855) );
  AOI21_X1 U10228 ( .B1(n8980), .B2(n8872), .A(n8855), .ZN(n8981) );
  AOI22_X1 U10229 ( .A1(n8931), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8856), .B2(
        n8929), .ZN(n8857) );
  OAI21_X1 U10230 ( .B1(n4519), .B2(n8908), .A(n8857), .ZN(n8868) );
  AOI21_X1 U10231 ( .B1(n8858), .B2(n8860), .A(n8859), .ZN(n8866) );
  OAI22_X1 U10232 ( .A1(n8864), .A2(n8863), .B1(n8862), .B2(n8861), .ZN(n8865)
         );
  AOI21_X1 U10233 ( .B1(n8866), .B2(n8832), .A(n8865), .ZN(n8983) );
  NOR2_X1 U10234 ( .A1(n8983), .A2(n8931), .ZN(n8867) );
  AOI211_X1 U10235 ( .C1(n8981), .C2(n6814), .A(n8868), .B(n8867), .ZN(n8869)
         );
  OAI21_X1 U10236 ( .B1(n8924), .B2(n8984), .A(n8869), .ZN(P2_U3274) );
  OR2_X1 U10237 ( .A1(n8887), .A2(n8046), .ZN(n8888) );
  NAND2_X1 U10238 ( .A1(n8888), .A2(n8870), .ZN(n8871) );
  XOR2_X1 U10239 ( .A(n8871), .B(n8880), .Z(n8989) );
  INV_X1 U10240 ( .A(n8872), .ZN(n8873) );
  AOI21_X1 U10241 ( .B1(n8985), .B2(n4521), .A(n8873), .ZN(n8986) );
  INV_X1 U10242 ( .A(n8874), .ZN(n8875) );
  AOI22_X1 U10243 ( .A1(n8931), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8875), .B2(
        n8929), .ZN(n8876) );
  OAI21_X1 U10244 ( .B1(n8877), .B2(n8908), .A(n8876), .ZN(n8885) );
  OAI21_X1 U10245 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8883) );
  AOI222_X1 U10246 ( .A1(n8920), .A2(n8883), .B1(n8882), .B2(n8917), .C1(n8881), .C2(n8915), .ZN(n8988) );
  NOR2_X1 U10247 ( .A1(n8988), .A2(n8931), .ZN(n8884) );
  AOI211_X1 U10248 ( .C1(n8986), .C2(n6814), .A(n8885), .B(n8884), .ZN(n8886)
         );
  OAI21_X1 U10249 ( .B1(n8924), .B2(n8989), .A(n8886), .ZN(P2_U3275) );
  INV_X1 U10250 ( .A(n8887), .ZN(n8890) );
  OAI21_X1 U10251 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8994) );
  AOI21_X1 U10252 ( .B1(n8990), .B2(n8892), .A(n8891), .ZN(n8991) );
  INV_X1 U10253 ( .A(n8990), .ZN(n8895) );
  AOI22_X1 U10254 ( .A1(n8931), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8893), .B2(
        n8929), .ZN(n8894) );
  OAI21_X1 U10255 ( .B1(n8895), .B2(n8908), .A(n8894), .ZN(n8900) );
  XNOR2_X1 U10256 ( .A(n8896), .B(n8046), .ZN(n8898) );
  AOI222_X1 U10257 ( .A1(n8920), .A2(n8898), .B1(n8897), .B2(n8917), .C1(n8918), .C2(n8915), .ZN(n8993) );
  NOR2_X1 U10258 ( .A1(n8993), .A2(n8931), .ZN(n8899) );
  AOI211_X1 U10259 ( .C1(n8991), .C2(n6814), .A(n8900), .B(n8899), .ZN(n8901)
         );
  OAI21_X1 U10260 ( .B1(n8924), .B2(n8994), .A(n8901), .ZN(P2_U3276) );
  XNOR2_X1 U10261 ( .A(n8902), .B(n8914), .ZN(n9004) );
  INV_X1 U10262 ( .A(n8903), .ZN(n8905) );
  AOI21_X1 U10263 ( .B1(n9000), .B2(n8905), .A(n8904), .ZN(n9001) );
  AOI22_X1 U10264 ( .A1(n8931), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8906), .B2(
        n8929), .ZN(n8907) );
  OAI21_X1 U10265 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n8922) );
  AND2_X1 U10266 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  OAI21_X1 U10267 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8919) );
  AOI222_X1 U10268 ( .A1(n8920), .A2(n8919), .B1(n8918), .B2(n8917), .C1(n8916), .C2(n8915), .ZN(n9003) );
  NOR2_X1 U10269 ( .A1(n9003), .A2(n8931), .ZN(n8921) );
  AOI211_X1 U10270 ( .C1(n9001), .C2(n6814), .A(n8922), .B(n8921), .ZN(n8923)
         );
  OAI21_X1 U10271 ( .B1(n9004), .B2(n8924), .A(n8923), .ZN(P2_U3278) );
  AOI22_X1 U10272 ( .A1(n8928), .A2(n8927), .B1(n8926), .B2(n8925), .ZN(n8937)
         );
  AOI22_X1 U10273 ( .A1(n6814), .A2(n8930), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8929), .ZN(n8936) );
  NAND2_X1 U10274 ( .A1(n8931), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U10275 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND4_X1 U10276 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), .ZN(
        P2_U3295) );
  NAND2_X1 U10277 ( .A1(n8938), .A2(n9898), .ZN(n8940) );
  OAI211_X1 U10278 ( .C1(n9955), .C2(n8941), .A(n8940), .B(n8939), .ZN(n9031)
         );
  MUX2_X1 U10279 ( .A(n9031), .B(P2_REG1_REG_31__SCAN_IN), .S(n9980), .Z(
        P2_U3551) );
  AOI22_X1 U10280 ( .A1(n8943), .A2(n9898), .B1(n9897), .B2(n8942), .ZN(n8944)
         );
  INV_X1 U10281 ( .A(n8948), .ZN(n8953) );
  AOI22_X1 U10282 ( .A1(n8950), .A2(n9898), .B1(n9897), .B2(n8949), .ZN(n8951)
         );
  OAI211_X1 U10283 ( .C1(n9890), .C2(n8953), .A(n8952), .B(n8951), .ZN(n9032)
         );
  MUX2_X1 U10284 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9032), .S(n9983), .Z(
        P2_U3548) );
  AOI22_X1 U10285 ( .A1(n8955), .A2(n9898), .B1(n9897), .B2(n8954), .ZN(n8956)
         );
  OAI211_X1 U10286 ( .C1(n9890), .C2(n8958), .A(n8957), .B(n8956), .ZN(n9033)
         );
  MUX2_X1 U10287 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9033), .S(n9983), .Z(
        P2_U3547) );
  MUX2_X1 U10288 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9034), .S(n9983), .Z(
        P2_U3546) );
  AOI211_X1 U10289 ( .C1(n9897), .C2(n8965), .A(n8964), .B(n8963), .ZN(n8966)
         );
  OAI21_X1 U10290 ( .B1(n9890), .B2(n8967), .A(n8966), .ZN(n9035) );
  MUX2_X1 U10291 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9035), .S(n9983), .Z(
        P2_U3545) );
  AOI22_X1 U10292 ( .A1(n8969), .A2(n9898), .B1(n9897), .B2(n8968), .ZN(n8970)
         );
  OAI211_X1 U10293 ( .C1(n8972), .C2(n9890), .A(n8971), .B(n8970), .ZN(n9036)
         );
  MUX2_X1 U10294 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9036), .S(n9983), .Z(
        P2_U3544) );
  OR2_X1 U10295 ( .A1(n8973), .A2(n9890), .ZN(n8979) );
  OAI22_X1 U10296 ( .A1(n8975), .A2(n9957), .B1(n8974), .B2(n9955), .ZN(n8976)
         );
  NOR2_X1 U10297 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  NAND2_X1 U10298 ( .A1(n8979), .A2(n8978), .ZN(n9037) );
  MUX2_X1 U10299 ( .A(n9037), .B(P2_REG1_REG_23__SCAN_IN), .S(n9980), .Z(
        P2_U3543) );
  AOI22_X1 U10300 ( .A1(n8981), .A2(n9898), .B1(n9897), .B2(n8980), .ZN(n8982)
         );
  OAI211_X1 U10301 ( .C1(n8984), .C2(n9890), .A(n8983), .B(n8982), .ZN(n9038)
         );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9038), .S(n9983), .Z(
        P2_U3542) );
  AOI22_X1 U10303 ( .A1(n8986), .A2(n9898), .B1(n9897), .B2(n8985), .ZN(n8987)
         );
  OAI211_X1 U10304 ( .C1(n8989), .C2(n9890), .A(n8988), .B(n8987), .ZN(n9039)
         );
  MUX2_X1 U10305 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9039), .S(n9983), .Z(
        P2_U3541) );
  AOI22_X1 U10306 ( .A1(n8991), .A2(n9898), .B1(n9897), .B2(n8990), .ZN(n8992)
         );
  OAI211_X1 U10307 ( .C1(n8994), .C2(n9890), .A(n8993), .B(n8992), .ZN(n9040)
         );
  MUX2_X1 U10308 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9040), .S(n9983), .Z(
        P2_U3540) );
  AOI21_X1 U10309 ( .B1(n9897), .B2(n8996), .A(n8995), .ZN(n8997) );
  OAI211_X1 U10310 ( .C1(n9890), .C2(n8999), .A(n8998), .B(n8997), .ZN(n9041)
         );
  MUX2_X1 U10311 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9041), .S(n9983), .Z(
        P2_U3539) );
  AOI22_X1 U10312 ( .A1(n9001), .A2(n9898), .B1(n9897), .B2(n9000), .ZN(n9002)
         );
  OAI211_X1 U10313 ( .C1(n9890), .C2(n9004), .A(n9003), .B(n9002), .ZN(n9042)
         );
  MUX2_X1 U10314 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9042), .S(n9983), .Z(
        P2_U3538) );
  AOI211_X1 U10315 ( .C1(n9897), .C2(n9007), .A(n9006), .B(n9005), .ZN(n9008)
         );
  OAI21_X1 U10316 ( .B1(n9009), .B2(n9890), .A(n9008), .ZN(n9043) );
  MUX2_X1 U10317 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9043), .S(n9983), .Z(
        P2_U3537) );
  AOI22_X1 U10318 ( .A1(n9011), .A2(n9898), .B1(n9897), .B2(n9010), .ZN(n9012)
         );
  OAI211_X1 U10319 ( .C1(n9030), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9044)
         );
  MUX2_X1 U10320 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9044), .S(n9983), .Z(
        P2_U3536) );
  AOI22_X1 U10321 ( .A1(n9016), .A2(n9898), .B1(n9897), .B2(n9015), .ZN(n9017)
         );
  OAI211_X1 U10322 ( .C1(n9890), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9045)
         );
  MUX2_X1 U10323 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9045), .S(n9983), .Z(
        P2_U3535) );
  AOI22_X1 U10324 ( .A1(n9021), .A2(n9898), .B1(n9897), .B2(n9020), .ZN(n9022)
         );
  OAI211_X1 U10325 ( .C1(n9024), .C2(n9890), .A(n9023), .B(n9022), .ZN(n9046)
         );
  MUX2_X1 U10326 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9046), .S(n9983), .Z(
        P2_U3534) );
  AOI22_X1 U10327 ( .A1(n9026), .A2(n9898), .B1(n9897), .B2(n9025), .ZN(n9027)
         );
  OAI211_X1 U10328 ( .C1(n9030), .C2(n9029), .A(n9028), .B(n9027), .ZN(n9047)
         );
  MUX2_X1 U10329 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9047), .S(n9983), .Z(
        P2_U3533) );
  MUX2_X1 U10330 ( .A(n9031), .B(P2_REG0_REG_31__SCAN_IN), .S(n9963), .Z(
        P2_U3519) );
  MUX2_X1 U10331 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9032), .S(n9965), .Z(
        P2_U3516) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9033), .S(n9965), .Z(
        P2_U3515) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9034), .S(n9965), .Z(
        P2_U3514) );
  MUX2_X1 U10334 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9035), .S(n9965), .Z(
        P2_U3513) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9036), .S(n9965), .Z(
        P2_U3512) );
  MUX2_X1 U10336 ( .A(n9037), .B(P2_REG0_REG_23__SCAN_IN), .S(n9963), .Z(
        P2_U3511) );
  MUX2_X1 U10337 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9038), .S(n9965), .Z(
        P2_U3510) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9039), .S(n9965), .Z(
        P2_U3509) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9040), .S(n9965), .Z(
        P2_U3508) );
  MUX2_X1 U10340 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9041), .S(n9965), .Z(
        P2_U3507) );
  MUX2_X1 U10341 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9042), .S(n9965), .Z(
        P2_U3505) );
  MUX2_X1 U10342 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9043), .S(n9965), .Z(
        P2_U3502) );
  MUX2_X1 U10343 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9044), .S(n9965), .Z(
        P2_U3499) );
  MUX2_X1 U10344 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9045), .S(n9965), .Z(
        P2_U3496) );
  MUX2_X1 U10345 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9046), .S(n9965), .Z(
        P2_U3493) );
  MUX2_X1 U10346 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9047), .S(n9965), .Z(
        P2_U3490) );
  INV_X1 U10347 ( .A(n9048), .ZN(n9608) );
  NOR4_X1 U10348 ( .A1(n4560), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9049), .A4(
        P2_U3152), .ZN(n9050) );
  AOI21_X1 U10349 ( .B1(n9051), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9050), .ZN(
        n9052) );
  OAI21_X1 U10350 ( .B1(n9608), .B2(n9058), .A(n9052), .ZN(P2_U3327) );
  OAI222_X1 U10351 ( .A1(n9060), .A2(n9055), .B1(n9058), .B2(n9054), .C1(
        P2_U3152), .C2(n9053), .ZN(P2_U3328) );
  INV_X1 U10352 ( .A(n9056), .ZN(n9612) );
  OAI222_X1 U10353 ( .A1(n9060), .A2(n9059), .B1(n9058), .B2(n9612), .C1(n9057), .C2(P2_U3152), .ZN(P2_U3329) );
  INV_X1 U10354 ( .A(n9061), .ZN(n9062) );
  MUX2_X1 U10355 ( .A(n9062), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI21_X1 U10356 ( .B1(n9172), .B2(n9064), .A(n9063), .ZN(n9066) );
  OAI21_X1 U10357 ( .B1(n9066), .B2(n9065), .A(n9173), .ZN(n9074) );
  OAI22_X1 U10358 ( .A1(n9068), .A2(n9632), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9067), .ZN(n9069) );
  AOI21_X1 U10359 ( .B1(n9320), .B2(n9164), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10360 ( .B1(n9071), .B2(n9636), .A(n9070), .ZN(n9072) );
  AOI21_X1 U10361 ( .B1(n9513), .B2(n9192), .A(n9072), .ZN(n9073) );
  NAND2_X1 U10362 ( .A1(n9074), .A2(n9073), .ZN(P1_U3212) );
  NAND2_X1 U10363 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  XOR2_X1 U10364 ( .A(n9078), .B(n9077), .Z(n9084) );
  OAI22_X1 U10365 ( .A1(n9110), .A2(n9636), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9079), .ZN(n9080) );
  AOI21_X1 U10366 ( .B1(n9160), .B2(n9409), .A(n9080), .ZN(n9081) );
  OAI21_X1 U10367 ( .B1(n9650), .B2(n9375), .A(n9081), .ZN(n9082) );
  AOI21_X1 U10368 ( .B1(n9532), .B2(n9192), .A(n9082), .ZN(n9083) );
  OAI21_X1 U10369 ( .B1(n9084), .B2(n9642), .A(n9083), .ZN(P1_U3214) );
  XNOR2_X1 U10370 ( .A(n9086), .B(n9085), .ZN(n9087) );
  XNOR2_X1 U10371 ( .A(n9088), .B(n9087), .ZN(n9094) );
  NAND2_X1 U10372 ( .A1(n9160), .A2(n9486), .ZN(n9089) );
  NAND2_X1 U10373 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9286) );
  OAI211_X1 U10374 ( .C1(n9090), .C2(n9636), .A(n9089), .B(n9286), .ZN(n9092)
         );
  NOR2_X1 U10375 ( .A1(n4483), .A2(n9181), .ZN(n9091) );
  AOI211_X1 U10376 ( .C1(n9433), .C2(n9164), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI21_X1 U10377 ( .B1(n9094), .B2(n9642), .A(n9093), .ZN(P1_U3217) );
  NAND2_X1 U10378 ( .A1(n9143), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U10379 ( .A1(n9097), .A2(n9098), .ZN(n9096) );
  OAI21_X1 U10380 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9099) );
  NAND2_X1 U10381 ( .A1(n9099), .A2(n9173), .ZN(n9104) );
  AOI22_X1 U10382 ( .A1(n9160), .A2(n9437), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9100) );
  OAI21_X1 U10383 ( .B1(n9101), .B2(n9636), .A(n9100), .ZN(n9102) );
  AOI21_X1 U10384 ( .B1(n9403), .B2(n9164), .A(n9102), .ZN(n9103) );
  OAI211_X1 U10385 ( .C1(n9405), .C2(n9181), .A(n9104), .B(n9103), .ZN(
        P1_U3221) );
  OAI21_X1 U10386 ( .B1(n9106), .B2(n9105), .A(n9168), .ZN(n9107) );
  NAND2_X1 U10387 ( .A1(n9107), .A2(n9173), .ZN(n9113) );
  NAND2_X1 U10388 ( .A1(n9352), .A2(n9188), .ZN(n9109) );
  NAND2_X1 U10389 ( .A1(P1_U3084), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9108) );
  OAI211_X1 U10390 ( .C1(n9110), .C2(n9632), .A(n9109), .B(n9108), .ZN(n9111)
         );
  AOI21_X1 U10391 ( .B1(n9346), .B2(n9164), .A(n9111), .ZN(n9112) );
  OAI211_X1 U10392 ( .C1(n9348), .C2(n9181), .A(n9113), .B(n9112), .ZN(
        P1_U3223) );
  OAI21_X1 U10393 ( .B1(n9116), .B2(n9114), .A(n9115), .ZN(n9117) );
  NAND2_X1 U10394 ( .A1(n9117), .A2(n9173), .ZN(n9122) );
  NAND2_X1 U10395 ( .A1(n9160), .A2(n9484), .ZN(n9118) );
  NAND2_X1 U10396 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9253) );
  OAI211_X1 U10397 ( .C1(n9119), .C2(n9636), .A(n9118), .B(n9253), .ZN(n9120)
         );
  AOI21_X1 U10398 ( .B1(n9475), .B2(n9164), .A(n9120), .ZN(n9121) );
  OAI211_X1 U10399 ( .C1(n9478), .C2(n9181), .A(n9122), .B(n9121), .ZN(
        P1_U3226) );
  INV_X1 U10400 ( .A(n9123), .ZN(n9124) );
  AOI21_X1 U10401 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9131) );
  NAND2_X1 U10402 ( .A1(n9366), .A2(n9188), .ZN(n9128) );
  AOI22_X1 U10403 ( .A1(n9160), .A2(n9394), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9127) );
  OAI211_X1 U10404 ( .C1(n9650), .C2(n9359), .A(n9128), .B(n9127), .ZN(n9129)
         );
  AOI21_X1 U10405 ( .B1(n9528), .B2(n9192), .A(n9129), .ZN(n9130) );
  OAI21_X1 U10406 ( .B1(n9131), .B2(n9642), .A(n9130), .ZN(P1_U3227) );
  INV_X1 U10407 ( .A(n9143), .ZN(n9132) );
  AOI21_X1 U10408 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9141) );
  OAI22_X1 U10409 ( .A1(n9636), .A2(n9136), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9135), .ZN(n9137) );
  AOI21_X1 U10410 ( .B1(n9160), .B2(n9447), .A(n9137), .ZN(n9138) );
  OAI21_X1 U10411 ( .B1(n9650), .B2(n9416), .A(n9138), .ZN(n9139) );
  AOI21_X1 U10412 ( .B1(n9548), .B2(n9192), .A(n9139), .ZN(n9140) );
  OAI21_X1 U10413 ( .B1(n9141), .B2(n9642), .A(n9140), .ZN(P1_U3231) );
  NAND2_X1 U10414 ( .A1(n9143), .A2(n9142), .ZN(n9145) );
  NAND2_X1 U10415 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U10416 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  XOR2_X1 U10417 ( .A(n9149), .B(n9148), .Z(n9155) );
  AOI22_X1 U10418 ( .A1(n9160), .A2(n9422), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9151) );
  NAND2_X1 U10419 ( .A1(n9164), .A2(n9387), .ZN(n9150) );
  OAI211_X1 U10420 ( .C1(n9152), .C2(n9636), .A(n9151), .B(n9150), .ZN(n9153)
         );
  AOI21_X1 U10421 ( .B1(n9537), .B2(n9192), .A(n9153), .ZN(n9154) );
  OAI21_X1 U10422 ( .B1(n9155), .B2(n9642), .A(n9154), .ZN(P1_U3233) );
  XNOR2_X1 U10423 ( .A(n9157), .B(n9156), .ZN(n9158) );
  XNOR2_X1 U10424 ( .A(n9159), .B(n9158), .ZN(n9167) );
  NAND2_X1 U10425 ( .A1(n9160), .A2(n9446), .ZN(n9161) );
  NAND2_X1 U10426 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9262) );
  OAI211_X1 U10427 ( .C1(n9162), .C2(n9636), .A(n9161), .B(n9262), .ZN(n9163)
         );
  AOI21_X1 U10428 ( .B1(n9459), .B2(n9164), .A(n9163), .ZN(n9166) );
  NAND2_X1 U10429 ( .A1(n9560), .A2(n9192), .ZN(n9165) );
  OAI211_X1 U10430 ( .C1(n9167), .C2(n9642), .A(n9166), .B(n9165), .ZN(
        P1_U3236) );
  INV_X1 U10431 ( .A(n9168), .ZN(n9171) );
  OAI21_X1 U10432 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9174) );
  NAND3_X1 U10433 ( .A1(n9174), .A2(n9173), .A3(n9172), .ZN(n9180) );
  NOR2_X1 U10434 ( .A1(n9331), .A2(n9650), .ZN(n9178) );
  OAI22_X1 U10435 ( .A1(n9176), .A2(n9632), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9175), .ZN(n9177) );
  AOI211_X1 U10436 ( .C1(n9337), .C2(n9188), .A(n9178), .B(n9177), .ZN(n9179)
         );
  OAI211_X1 U10437 ( .C1(n9334), .C2(n9181), .A(n9180), .B(n9179), .ZN(
        P1_U3238) );
  NAND2_X1 U10438 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  XOR2_X1 U10439 ( .A(n9185), .B(n9184), .Z(n9195) );
  AND2_X1 U10440 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9222) );
  NOR2_X1 U10441 ( .A1(n9632), .A2(n9186), .ZN(n9187) );
  AOI211_X1 U10442 ( .C1(n9188), .C2(n9484), .A(n9222), .B(n9187), .ZN(n9189)
         );
  OAI21_X1 U10443 ( .B1(n9650), .B2(n9190), .A(n9189), .ZN(n9191) );
  AOI21_X1 U10444 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9194) );
  OAI21_X1 U10445 ( .B1(n9195), .B2(n9642), .A(n9194), .ZN(P1_U3239) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9196), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9197), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9301), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n4819), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9337), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9352), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9366), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9380), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9394), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9409), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9422), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9437), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9447), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9486), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9446), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9484), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9198), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9199), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9200), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9201), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9202), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9203), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9204), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9205), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9206), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9207), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9208), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9209), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9210), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9211), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6717), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U10477 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9226) );
  NOR2_X1 U10478 ( .A1(n9213), .A2(n9212), .ZN(n9215) );
  NOR2_X1 U10479 ( .A1(n9215), .A2(n9214), .ZN(n9227) );
  XNOR2_X1 U10480 ( .A(n9227), .B(n9234), .ZN(n9216) );
  NOR2_X1 U10481 ( .A1(n7670), .A2(n9216), .ZN(n9228) );
  AOI211_X1 U10482 ( .C1(n9216), .C2(n7670), .A(n9228), .B(n9763), .ZN(n9217)
         );
  INV_X1 U10483 ( .A(n9217), .ZN(n9225) );
  OAI21_X1 U10484 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9219), .A(n9218), .ZN(
        n9233) );
  XNOR2_X1 U10485 ( .A(n9234), .B(n9233), .ZN(n9220) );
  INV_X1 U10486 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9670) );
  NOR2_X1 U10487 ( .A1(n9670), .A2(n9220), .ZN(n9235) );
  AOI211_X1 U10488 ( .C1(n9220), .C2(n9670), .A(n9235), .B(n9750), .ZN(n9221)
         );
  AOI211_X1 U10489 ( .C1(n9778), .C2(n9223), .A(n9222), .B(n9221), .ZN(n9224)
         );
  OAI211_X1 U10490 ( .C1(n9792), .C2(n9226), .A(n9225), .B(n9224), .ZN(
        P1_U3256) );
  NOR2_X1 U10491 ( .A1(n9227), .A2(n9234), .ZN(n9229) );
  NOR2_X1 U10492 ( .A1(n9229), .A2(n9228), .ZN(n9232) );
  NAND2_X1 U10493 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9249), .ZN(n9230) );
  OAI21_X1 U10494 ( .B1(n9249), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9230), .ZN(
        n9231) );
  NOR2_X1 U10495 ( .A1(n9232), .A2(n9231), .ZN(n9248) );
  AOI211_X1 U10496 ( .C1(n9232), .C2(n9231), .A(n9248), .B(n9763), .ZN(n9244)
         );
  NOR2_X1 U10497 ( .A1(n9234), .A2(n9233), .ZN(n9236) );
  NOR2_X1 U10498 ( .A1(n9236), .A2(n9235), .ZN(n9239) );
  INV_X1 U10499 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9237) );
  MUX2_X1 U10500 ( .A(n9237), .B(P1_REG1_REG_16__SCAN_IN), .S(n9249), .Z(n9238) );
  NOR2_X1 U10501 ( .A1(n9239), .A2(n9238), .ZN(n9245) );
  AOI211_X1 U10502 ( .C1(n9239), .C2(n9238), .A(n9245), .B(n9750), .ZN(n9243)
         );
  INV_X1 U10503 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U10504 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U10505 ( .A1(n9778), .A2(n9249), .ZN(n9240) );
  OAI211_X1 U10506 ( .C1(n9792), .C2(n9241), .A(n9633), .B(n9240), .ZN(n9242)
         );
  OR3_X1 U10507 ( .A1(n9244), .A2(n9243), .A3(n9242), .ZN(P1_U3257) );
  AOI21_X1 U10508 ( .B1(n9249), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9245), .ZN(
        n9247) );
  XNOR2_X1 U10509 ( .A(n9266), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9246) );
  NOR2_X1 U10510 ( .A1(n9247), .A2(n9246), .ZN(n9259) );
  AOI211_X1 U10511 ( .C1(n9247), .C2(n9246), .A(n9259), .B(n9750), .ZN(n9257)
         );
  AOI21_X1 U10512 ( .B1(n9249), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9248), .ZN(
        n9252) );
  INV_X1 U10513 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9250) );
  MUX2_X1 U10514 ( .A(n9250), .B(P1_REG2_REG_17__SCAN_IN), .S(n9266), .Z(n9251) );
  NOR2_X1 U10515 ( .A1(n9252), .A2(n9251), .ZN(n9265) );
  AOI211_X1 U10516 ( .C1(n9252), .C2(n9251), .A(n9265), .B(n9763), .ZN(n9256)
         );
  INV_X1 U10517 ( .A(n9266), .ZN(n9254) );
  OAI21_X1 U10518 ( .B1(n9264), .B2(n9254), .A(n9253), .ZN(n9255) );
  NOR3_X1 U10519 ( .A1(n9257), .A2(n9256), .A3(n9255), .ZN(n9258) );
  OAI21_X1 U10520 ( .B1(n9792), .B2(n7911), .A(n9258), .ZN(P1_U3258) );
  INV_X1 U10521 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9273) );
  XOR2_X1 U10522 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9276), .Z(n9261) );
  AOI21_X1 U10523 ( .B1(n9266), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9259), .ZN(
        n9260) );
  NAND2_X1 U10524 ( .A1(n9261), .A2(n9260), .ZN(n9275) );
  OAI21_X1 U10525 ( .B1(n9261), .B2(n9260), .A(n9275), .ZN(n9271) );
  INV_X1 U10526 ( .A(n9276), .ZN(n9263) );
  OAI21_X1 U10527 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9270) );
  XNOR2_X1 U10528 ( .A(n9276), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9267) );
  AOI211_X1 U10529 ( .C1(n9268), .C2(n9267), .A(n9274), .B(n9763), .ZN(n9269)
         );
  AOI211_X1 U10530 ( .C1(n9786), .C2(n9271), .A(n9270), .B(n9269), .ZN(n9272)
         );
  OAI21_X1 U10531 ( .B1(n9792), .B2(n9273), .A(n9272), .ZN(P1_U3259) );
  NAND2_X1 U10532 ( .A1(n9282), .A2(n9787), .ZN(n9280) );
  OAI21_X1 U10533 ( .B1(n9276), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9275), .ZN(
        n9278) );
  INV_X1 U10534 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9277) );
  XNOR2_X1 U10535 ( .A(n9278), .B(n9277), .ZN(n9281) );
  AOI21_X1 U10536 ( .B1(n9281), .B2(n9786), .A(n9778), .ZN(n9279) );
  NAND2_X1 U10537 ( .A1(n9280), .A2(n9279), .ZN(n9285) );
  OAI22_X1 U10538 ( .A1(n9282), .A2(n9763), .B1(n9281), .B2(n9750), .ZN(n9284)
         );
  MUX2_X1 U10539 ( .A(n9285), .B(n9284), .S(n9283), .Z(n9288) );
  OAI21_X1 U10540 ( .B1(n9792), .B2(n4877), .A(n9286), .ZN(n9287) );
  XNOR2_X1 U10541 ( .A(n9290), .B(n9289), .ZN(n9654) );
  NAND2_X1 U10542 ( .A1(n9654), .A2(n9441), .ZN(n9294) );
  AND2_X1 U10543 ( .A1(n9489), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9291) );
  NOR2_X1 U10544 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  OAI211_X1 U10545 ( .C1(n9652), .C2(n9477), .A(n9294), .B(n9293), .ZN(
        P1_U3262) );
  NAND2_X1 U10546 ( .A1(n9295), .A2(n9298), .ZN(n9296) );
  NAND2_X1 U10547 ( .A1(n9297), .A2(n9296), .ZN(n9504) );
  XNOR2_X1 U10548 ( .A(n9299), .B(n9298), .ZN(n9300) );
  NAND2_X1 U10549 ( .A1(n9300), .A2(n9488), .ZN(n9303) );
  AOI22_X1 U10550 ( .A1(n9337), .A2(n9483), .B1(n9485), .B2(n9301), .ZN(n9302)
         );
  NAND2_X1 U10551 ( .A1(n9303), .A2(n9302), .ZN(n9509) );
  NAND2_X1 U10552 ( .A1(n9505), .A2(n9317), .ZN(n9304) );
  NAND3_X1 U10553 ( .A1(n9305), .A2(n9655), .A3(n9304), .ZN(n9507) );
  NOR2_X1 U10554 ( .A1(n9507), .A2(n9306), .ZN(n9312) );
  INV_X1 U10555 ( .A(n9307), .ZN(n9308) );
  AOI22_X1 U10556 ( .A1(n9308), .A2(n9474), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9465), .ZN(n9309) );
  OAI21_X1 U10557 ( .B1(n9310), .B2(n9477), .A(n9309), .ZN(n9311) );
  AOI211_X1 U10558 ( .C1(n9509), .C2(n9313), .A(n9312), .B(n9311), .ZN(n9314)
         );
  OAI21_X1 U10559 ( .B1(n9504), .B2(n9494), .A(n9314), .ZN(P1_U3263) );
  XNOR2_X1 U10560 ( .A(n9316), .B(n9315), .ZN(n9516) );
  INV_X1 U10561 ( .A(n9329), .ZN(n9319) );
  INV_X1 U10562 ( .A(n9317), .ZN(n9318) );
  AOI211_X1 U10563 ( .C1(n9513), .C2(n9319), .A(n9843), .B(n9318), .ZN(n9512)
         );
  AOI22_X1 U10564 ( .A1(n9320), .A2(n9474), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9465), .ZN(n9321) );
  OAI21_X1 U10565 ( .B1(n4821), .B2(n9477), .A(n9321), .ZN(n9326) );
  XNOR2_X1 U10566 ( .A(n9324), .B(n9323), .ZN(n9325) );
  OAI21_X1 U10567 ( .B1(n9328), .B2(n7715), .A(n9327), .ZN(n9521) );
  INV_X1 U10568 ( .A(n9344), .ZN(n9330) );
  AOI21_X1 U10569 ( .B1(n9517), .B2(n9330), .A(n9329), .ZN(n9518) );
  INV_X1 U10570 ( .A(n9331), .ZN(n9332) );
  AOI22_X1 U10571 ( .A1(n9332), .A2(n9474), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9465), .ZN(n9333) );
  OAI21_X1 U10572 ( .B1(n9334), .B2(n9477), .A(n9333), .ZN(n9340) );
  OAI21_X1 U10573 ( .B1(n4355), .B2(n9336), .A(n9335), .ZN(n9338) );
  AOI222_X1 U10574 ( .A1(n9488), .A2(n9338), .B1(n9337), .B2(n9485), .C1(n9366), .C2(n9483), .ZN(n9520) );
  NOR2_X1 U10575 ( .A1(n9520), .A2(n9489), .ZN(n9339) );
  AOI211_X1 U10576 ( .C1(n9518), .C2(n9441), .A(n9340), .B(n9339), .ZN(n9341)
         );
  OAI21_X1 U10577 ( .B1(n9494), .B2(n9521), .A(n9341), .ZN(P1_U3265) );
  XNOR2_X1 U10578 ( .A(n9343), .B(n9342), .ZN(n9526) );
  INV_X1 U10579 ( .A(n9358), .ZN(n9345) );
  AOI211_X1 U10580 ( .C1(n9523), .C2(n9345), .A(n9843), .B(n9344), .ZN(n9522)
         );
  AOI22_X1 U10581 ( .A1(n9346), .A2(n9474), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9465), .ZN(n9347) );
  OAI21_X1 U10582 ( .B1(n9348), .B2(n9477), .A(n9347), .ZN(n9355) );
  NAND2_X1 U10583 ( .A1(n9363), .A2(n9349), .ZN(n9351) );
  XNOR2_X1 U10584 ( .A(n9351), .B(n9350), .ZN(n9353) );
  AOI222_X1 U10585 ( .A1(n9488), .A2(n9353), .B1(n9352), .B2(n9485), .C1(n9380), .C2(n9483), .ZN(n9525) );
  NOR2_X1 U10586 ( .A1(n9525), .A2(n9489), .ZN(n9354) );
  AOI211_X1 U10587 ( .C1(n9522), .C2(n9492), .A(n9355), .B(n9354), .ZN(n9356)
         );
  OAI21_X1 U10588 ( .B1(n9494), .B2(n9526), .A(n9356), .ZN(P1_U3266) );
  XNOR2_X1 U10589 ( .A(n9357), .B(n9365), .ZN(n9531) );
  AOI211_X1 U10590 ( .C1(n9528), .C2(n9373), .A(n9843), .B(n9358), .ZN(n9527)
         );
  INV_X1 U10591 ( .A(n9528), .ZN(n9362) );
  INV_X1 U10592 ( .A(n9359), .ZN(n9360) );
  AOI22_X1 U10593 ( .A1(n9360), .A2(n9474), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9465), .ZN(n9361) );
  OAI21_X1 U10594 ( .B1(n9362), .B2(n9477), .A(n9361), .ZN(n9369) );
  OAI21_X1 U10595 ( .B1(n9365), .B2(n9364), .A(n9363), .ZN(n9367) );
  AOI222_X1 U10596 ( .A1(n9488), .A2(n9367), .B1(n9366), .B2(n9485), .C1(n9394), .C2(n9483), .ZN(n9530) );
  NOR2_X1 U10597 ( .A1(n9530), .A2(n9465), .ZN(n9368) );
  AOI211_X1 U10598 ( .C1(n9527), .C2(n9492), .A(n9369), .B(n9368), .ZN(n9370)
         );
  OAI21_X1 U10599 ( .B1(n9531), .B2(n9494), .A(n9370), .ZN(P1_U3267) );
  XNOR2_X1 U10600 ( .A(n9372), .B(n9371), .ZN(n9536) );
  INV_X1 U10601 ( .A(n9373), .ZN(n9374) );
  AOI21_X1 U10602 ( .B1(n9532), .B2(n9386), .A(n9374), .ZN(n9533) );
  INV_X1 U10603 ( .A(n9375), .ZN(n9376) );
  AOI22_X1 U10604 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n9489), .B1(n9376), .B2(
        n9474), .ZN(n9377) );
  OAI21_X1 U10605 ( .B1(n9378), .B2(n9477), .A(n9377), .ZN(n9383) );
  OAI21_X1 U10606 ( .B1(n4863), .B2(n7733), .A(n9379), .ZN(n9381) );
  AOI222_X1 U10607 ( .A1(n9488), .A2(n9381), .B1(n9380), .B2(n9485), .C1(n9409), .C2(n9483), .ZN(n9535) );
  NOR2_X1 U10608 ( .A1(n9535), .A2(n9489), .ZN(n9382) );
  AOI211_X1 U10609 ( .C1(n9533), .C2(n9441), .A(n9383), .B(n9382), .ZN(n9384)
         );
  OAI21_X1 U10610 ( .B1(n9494), .B2(n9536), .A(n9384), .ZN(P1_U3268) );
  XNOR2_X1 U10611 ( .A(n9385), .B(n9392), .ZN(n9541) );
  AOI21_X1 U10612 ( .B1(n9537), .B2(n9401), .A(n4484), .ZN(n9538) );
  INV_X1 U10613 ( .A(n9537), .ZN(n9389) );
  AOI22_X1 U10614 ( .A1(n9465), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9387), .B2(
        n9474), .ZN(n9388) );
  OAI21_X1 U10615 ( .B1(n9389), .B2(n9477), .A(n9388), .ZN(n9397) );
  INV_X1 U10616 ( .A(n9392), .ZN(n9393) );
  NAND2_X1 U10617 ( .A1(n9406), .A2(n9390), .ZN(n9391) );
  MUX2_X1 U10618 ( .A(n9393), .B(n9392), .S(n9391), .Z(n9395) );
  AOI222_X1 U10619 ( .A1(n9488), .A2(n9395), .B1(n9394), .B2(n9485), .C1(n9422), .C2(n9483), .ZN(n9540) );
  NOR2_X1 U10620 ( .A1(n9540), .A2(n9489), .ZN(n9396) );
  AOI211_X1 U10621 ( .C1(n9538), .C2(n9441), .A(n9397), .B(n9396), .ZN(n9398)
         );
  OAI21_X1 U10622 ( .B1(n9494), .B2(n9541), .A(n9398), .ZN(P1_U3269) );
  XOR2_X1 U10623 ( .A(n9399), .B(n9408), .Z(n9546) );
  INV_X1 U10624 ( .A(n9400), .ZN(n9402) );
  AOI211_X1 U10625 ( .C1(n9543), .C2(n9402), .A(n9843), .B(n4481), .ZN(n9542)
         );
  AOI22_X1 U10626 ( .A1(n9465), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9403), .B2(
        n9474), .ZN(n9404) );
  OAI21_X1 U10627 ( .B1(n9405), .B2(n9477), .A(n9404), .ZN(n9412) );
  OAI21_X1 U10628 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9410) );
  AOI222_X1 U10629 ( .A1(n9488), .A2(n9410), .B1(n9437), .B2(n9483), .C1(n9409), .C2(n9485), .ZN(n9545) );
  NOR2_X1 U10630 ( .A1(n9545), .A2(n9489), .ZN(n9411) );
  AOI211_X1 U10631 ( .C1(n9542), .C2(n9492), .A(n9412), .B(n9411), .ZN(n9413)
         );
  OAI21_X1 U10632 ( .B1(n9546), .B2(n9494), .A(n9413), .ZN(P1_U3270) );
  XNOR2_X1 U10633 ( .A(n9414), .B(n9420), .ZN(n9551) );
  INV_X1 U10634 ( .A(n9432), .ZN(n9415) );
  AOI211_X1 U10635 ( .C1(n9548), .C2(n9415), .A(n9843), .B(n9400), .ZN(n9547)
         );
  INV_X1 U10636 ( .A(n9416), .ZN(n9417) );
  AOI22_X1 U10637 ( .A1(n9465), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9417), .B2(
        n9474), .ZN(n9418) );
  OAI21_X1 U10638 ( .B1(n9419), .B2(n9477), .A(n9418), .ZN(n9425) );
  XOR2_X1 U10639 ( .A(n9421), .B(n9420), .Z(n9423) );
  AOI222_X1 U10640 ( .A1(n9488), .A2(n9423), .B1(n9422), .B2(n9485), .C1(n9447), .C2(n9483), .ZN(n9550) );
  NOR2_X1 U10641 ( .A1(n9550), .A2(n9489), .ZN(n9424) );
  AOI211_X1 U10642 ( .C1(n9547), .C2(n9492), .A(n9425), .B(n9424), .ZN(n9426)
         );
  OAI21_X1 U10643 ( .B1(n9494), .B2(n9551), .A(n9426), .ZN(P1_U3271) );
  NAND2_X1 U10644 ( .A1(n9467), .A2(n9427), .ZN(n9455) );
  NAND2_X1 U10645 ( .A1(n9455), .A2(n9428), .ZN(n9431) );
  OAI21_X1 U10646 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9556) );
  AOI21_X1 U10647 ( .B1(n9552), .B2(n9457), .A(n9432), .ZN(n9553) );
  AOI22_X1 U10648 ( .A1(n9489), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9433), .B2(
        n9474), .ZN(n9434) );
  OAI21_X1 U10649 ( .B1(n4483), .B2(n9477), .A(n9434), .ZN(n9440) );
  XNOR2_X1 U10650 ( .A(n9436), .B(n9435), .ZN(n9438) );
  AOI222_X1 U10651 ( .A1(n9488), .A2(n9438), .B1(n9437), .B2(n9485), .C1(n9486), .C2(n9483), .ZN(n9555) );
  NOR2_X1 U10652 ( .A1(n9555), .A2(n9489), .ZN(n9439) );
  AOI211_X1 U10653 ( .C1(n9553), .C2(n9441), .A(n9440), .B(n9439), .ZN(n9442)
         );
  OAI21_X1 U10654 ( .B1(n9494), .B2(n9556), .A(n9442), .ZN(P1_U3272) );
  NAND2_X1 U10655 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  XNOR2_X1 U10656 ( .A(n9445), .B(n9452), .ZN(n9448) );
  AOI222_X1 U10657 ( .A1(n9488), .A2(n9448), .B1(n9447), .B2(n9485), .C1(n9446), .C2(n9483), .ZN(n9562) );
  NAND2_X1 U10658 ( .A1(n9467), .A2(n9449), .ZN(n9451) );
  NAND2_X1 U10659 ( .A1(n9451), .A2(n9450), .ZN(n9453) );
  OR2_X1 U10660 ( .A1(n9453), .A2(n9452), .ZN(n9558) );
  AND2_X1 U10661 ( .A1(n9455), .A2(n9454), .ZN(n9557) );
  NAND3_X1 U10662 ( .A1(n9558), .A2(n9557), .A3(n9456), .ZN(n9464) );
  INV_X1 U10663 ( .A(n9457), .ZN(n9458) );
  AOI211_X1 U10664 ( .C1(n9560), .C2(n9471), .A(n9843), .B(n9458), .ZN(n9559)
         );
  INV_X1 U10665 ( .A(n9560), .ZN(n9461) );
  AOI22_X1 U10666 ( .A1(n9489), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9459), .B2(
        n9474), .ZN(n9460) );
  OAI21_X1 U10667 ( .B1(n9461), .B2(n9477), .A(n9460), .ZN(n9462) );
  AOI21_X1 U10668 ( .B1(n9559), .B2(n9492), .A(n9462), .ZN(n9463) );
  OAI211_X1 U10669 ( .C1(n9465), .C2(n9562), .A(n9464), .B(n9463), .ZN(
        P1_U3273) );
  NAND2_X1 U10670 ( .A1(n9467), .A2(n9466), .ZN(n9469) );
  NAND2_X1 U10671 ( .A1(n9469), .A2(n9468), .ZN(n9470) );
  XOR2_X1 U10672 ( .A(n9481), .B(n9470), .Z(n9568) );
  INV_X1 U10673 ( .A(n7749), .ZN(n9473) );
  INV_X1 U10674 ( .A(n9471), .ZN(n9472) );
  AOI211_X1 U10675 ( .C1(n9565), .C2(n9473), .A(n9843), .B(n9472), .ZN(n9564)
         );
  AOI22_X1 U10676 ( .A1(n9489), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9475), .B2(
        n9474), .ZN(n9476) );
  OAI21_X1 U10677 ( .B1(n9478), .B2(n9477), .A(n9476), .ZN(n9491) );
  NAND2_X1 U10678 ( .A1(n9480), .A2(n9479), .ZN(n9482) );
  XNOR2_X1 U10679 ( .A(n9482), .B(n9481), .ZN(n9487) );
  AOI222_X1 U10680 ( .A1(n9488), .A2(n9487), .B1(n9486), .B2(n9485), .C1(n9484), .C2(n9483), .ZN(n9567) );
  NOR2_X1 U10681 ( .A1(n9567), .A2(n9489), .ZN(n9490) );
  AOI211_X1 U10682 ( .C1(n9564), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9493)
         );
  OAI21_X1 U10683 ( .B1(n9494), .B2(n9568), .A(n9493), .ZN(P1_U3274) );
  NAND2_X1 U10684 ( .A1(n9495), .A2(n9615), .ZN(n9496) );
  OAI211_X1 U10685 ( .C1(n9497), .C2(n9843), .A(n9651), .B(n9496), .ZN(n9585)
         );
  MUX2_X1 U10686 ( .A(n9585), .B(P1_REG1_REG_31__SCAN_IN), .S(n9864), .Z(
        P1_U3554) );
  AOI22_X1 U10687 ( .A1(n9500), .A2(n9655), .B1(n9499), .B2(n9615), .ZN(n9501)
         );
  OAI211_X1 U10688 ( .C1(n9503), .C2(n9661), .A(n9502), .B(n9501), .ZN(n9586)
         );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9586), .S(n9853), .Z(
        P1_U3552) );
  NAND2_X1 U10690 ( .A1(n9505), .A2(n9615), .ZN(n9506) );
  NAND2_X1 U10691 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  NOR2_X1 U10692 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U10693 ( .A1(n9511), .A2(n9510), .ZN(n9587) );
  MUX2_X1 U10694 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9587), .S(n9853), .Z(
        P1_U3551) );
  AOI21_X1 U10695 ( .B1(n9513), .B2(n9615), .A(n9512), .ZN(n9514) );
  OAI211_X1 U10696 ( .C1(n9516), .C2(n9661), .A(n9515), .B(n9514), .ZN(n9588)
         );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9588), .S(n9853), .Z(
        P1_U3550) );
  AOI22_X1 U10698 ( .A1(n9518), .A2(n9655), .B1(n9517), .B2(n9615), .ZN(n9519)
         );
  OAI211_X1 U10699 ( .C1(n9521), .C2(n9661), .A(n9520), .B(n9519), .ZN(n9589)
         );
  MUX2_X1 U10700 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9589), .S(n9853), .Z(
        P1_U3549) );
  AOI21_X1 U10701 ( .B1(n9523), .B2(n9615), .A(n9522), .ZN(n9524) );
  OAI211_X1 U10702 ( .C1(n9526), .C2(n9661), .A(n9525), .B(n9524), .ZN(n9590)
         );
  MUX2_X1 U10703 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9590), .S(n9853), .Z(
        P1_U3548) );
  AOI21_X1 U10704 ( .B1(n9528), .B2(n9615), .A(n9527), .ZN(n9529) );
  OAI211_X1 U10705 ( .C1(n9531), .C2(n9661), .A(n9530), .B(n9529), .ZN(n9591)
         );
  MUX2_X1 U10706 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9591), .S(n9853), .Z(
        P1_U3547) );
  AOI22_X1 U10707 ( .A1(n9533), .A2(n9655), .B1(n9532), .B2(n9615), .ZN(n9534)
         );
  OAI211_X1 U10708 ( .C1(n9536), .C2(n9661), .A(n9535), .B(n9534), .ZN(n9592)
         );
  MUX2_X1 U10709 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9592), .S(n9853), .Z(
        P1_U3546) );
  AOI22_X1 U10710 ( .A1(n9538), .A2(n9655), .B1(n9537), .B2(n9615), .ZN(n9539)
         );
  OAI211_X1 U10711 ( .C1(n9541), .C2(n9661), .A(n9540), .B(n9539), .ZN(n9593)
         );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9593), .S(n9853), .Z(
        P1_U3545) );
  AOI21_X1 U10713 ( .B1(n9543), .B2(n9615), .A(n9542), .ZN(n9544) );
  OAI211_X1 U10714 ( .C1(n9546), .C2(n9661), .A(n9545), .B(n9544), .ZN(n9594)
         );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9594), .S(n9853), .Z(
        P1_U3544) );
  AOI21_X1 U10716 ( .B1(n9548), .B2(n9615), .A(n9547), .ZN(n9549) );
  OAI211_X1 U10717 ( .C1(n9551), .C2(n9661), .A(n9550), .B(n9549), .ZN(n9595)
         );
  MUX2_X1 U10718 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9595), .S(n9853), .Z(
        P1_U3543) );
  AOI22_X1 U10719 ( .A1(n9553), .A2(n9655), .B1(n9552), .B2(n9615), .ZN(n9554)
         );
  OAI211_X1 U10720 ( .C1(n9556), .C2(n9661), .A(n9555), .B(n9554), .ZN(n9596)
         );
  MUX2_X1 U10721 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9596), .S(n9853), .Z(
        P1_U3542) );
  INV_X1 U10722 ( .A(n9661), .ZN(n9832) );
  NAND3_X1 U10723 ( .A1(n9558), .A2(n9557), .A3(n9832), .ZN(n9563) );
  AOI21_X1 U10724 ( .B1(n9560), .B2(n9615), .A(n9559), .ZN(n9561) );
  NAND3_X1 U10725 ( .A1(n9563), .A2(n9562), .A3(n9561), .ZN(n9597) );
  MUX2_X1 U10726 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9597), .S(n9853), .Z(
        P1_U3541) );
  AOI21_X1 U10727 ( .B1(n9565), .B2(n9615), .A(n9564), .ZN(n9566) );
  OAI211_X1 U10728 ( .C1(n9568), .C2(n9661), .A(n9567), .B(n9566), .ZN(n9598)
         );
  MUX2_X1 U10729 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9598), .S(n9853), .Z(
        P1_U3540) );
  AOI21_X1 U10730 ( .B1(n9570), .B2(n9615), .A(n9569), .ZN(n9571) );
  OAI211_X1 U10731 ( .C1(n9573), .C2(n9661), .A(n9572), .B(n9571), .ZN(n9599)
         );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9599), .S(n9853), .Z(
        P1_U3537) );
  NAND2_X1 U10733 ( .A1(n9574), .A2(n9615), .ZN(n9576) );
  OAI211_X1 U10734 ( .C1(n9577), .C2(n9805), .A(n9576), .B(n9575), .ZN(n9578)
         );
  OR2_X1 U10735 ( .A1(n9579), .A2(n9578), .ZN(n9600) );
  MUX2_X1 U10736 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9600), .S(n9853), .Z(
        P1_U3535) );
  AOI211_X1 U10737 ( .C1(n9582), .C2(n9615), .A(n9581), .B(n9580), .ZN(n9583)
         );
  OAI21_X1 U10738 ( .B1(n9661), .B2(n9584), .A(n9583), .ZN(n9601) );
  MUX2_X1 U10739 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9601), .S(n9853), .Z(
        P1_U3534) );
  MUX2_X1 U10740 ( .A(n9585), .B(P1_REG0_REG_31__SCAN_IN), .S(n9849), .Z(
        P1_U3522) );
  MUX2_X1 U10741 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9586), .S(n9850), .Z(
        P1_U3520) );
  MUX2_X1 U10742 ( .A(n9587), .B(P1_REG0_REG_28__SCAN_IN), .S(n9849), .Z(
        P1_U3519) );
  MUX2_X1 U10743 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9588), .S(n9850), .Z(
        P1_U3518) );
  MUX2_X1 U10744 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9589), .S(n9850), .Z(
        P1_U3517) );
  MUX2_X1 U10745 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9590), .S(n9850), .Z(
        P1_U3516) );
  MUX2_X1 U10746 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9591), .S(n9850), .Z(
        P1_U3515) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9592), .S(n9850), .Z(
        P1_U3514) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9593), .S(n9850), .Z(
        P1_U3513) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9594), .S(n9850), .Z(
        P1_U3512) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9595), .S(n9850), .Z(
        P1_U3511) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9596), .S(n9850), .Z(
        P1_U3510) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9597), .S(n9850), .Z(
        P1_U3508) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9598), .S(n9850), .Z(
        P1_U3505) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9599), .S(n9850), .Z(
        P1_U3496) );
  MUX2_X1 U10755 ( .A(n9600), .B(P1_REG0_REG_12__SCAN_IN), .S(n9849), .Z(
        P1_U3490) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9601), .S(n9850), .Z(
        P1_U3487) );
  MUX2_X1 U10757 ( .A(P1_D_REG_0__SCAN_IN), .B(n9603), .S(n9801), .Z(P1_U3440)
         );
  NOR4_X1 U10758 ( .A1(n9604), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5557), .ZN(n9605) );
  AOI21_X1 U10759 ( .B1(n9606), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9605), .ZN(
        n9607) );
  OAI21_X1 U10760 ( .B1(n9608), .B2(n9613), .A(n9607), .ZN(P1_U3322) );
  OAI222_X1 U10761 ( .A1(n9613), .A2(n9612), .B1(n9611), .B2(P1_U3084), .C1(
        n9610), .C2(n9609), .ZN(P1_U3324) );
  MUX2_X1 U10762 ( .A(n9614), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NAND2_X1 U10763 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  NAND2_X1 U10764 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U10765 ( .B1(n9620), .B2(n9848), .A(n9619), .ZN(n9621) );
  AND2_X1 U10766 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  AOI22_X1 U10767 ( .A1(n9850), .A2(n9623), .B1(n5772), .B2(n9849), .ZN(
        P1_U3484) );
  AOI22_X1 U10768 ( .A1(n9853), .A2(n9623), .B1(n6434), .B2(n9864), .ZN(
        P1_U3533) );
  NOR2_X1 U10769 ( .A1(n9624), .A2(n9957), .ZN(n9625) );
  INV_X1 U10770 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9628) );
  AOI22_X1 U10771 ( .A1(n9983), .A2(n9630), .B1(n9628), .B2(n9980), .ZN(
        P2_U3550) );
  INV_X1 U10772 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U10773 ( .A1(n9965), .A2(n9630), .B1(n9629), .B2(n9963), .ZN(
        P2_U3518) );
  OR2_X1 U10774 ( .A1(n9632), .A2(n9631), .ZN(n9634) );
  OAI211_X1 U10775 ( .C1(n9636), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9637)
         );
  INV_X1 U10776 ( .A(n9637), .ZN(n9648) );
  NOR2_X1 U10777 ( .A1(n9638), .A2(n9841), .ZN(n9659) );
  NAND2_X1 U10778 ( .A1(n9639), .A2(n9182), .ZN(n9641) );
  NAND2_X1 U10779 ( .A1(n9641), .A2(n9640), .ZN(n9643) );
  AOI21_X1 U10780 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9645) );
  AOI21_X1 U10781 ( .B1(n9646), .B2(n9659), .A(n9645), .ZN(n9647) );
  OAI211_X1 U10782 ( .C1(n9650), .C2(n9649), .A(n9648), .B(n9647), .ZN(
        P1_U3224) );
  OAI21_X1 U10783 ( .B1(n9652), .B2(n9841), .A(n9651), .ZN(n9653) );
  AOI21_X1 U10784 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9677) );
  AOI22_X1 U10785 ( .A1(n9853), .A2(n9677), .B1(n7741), .B2(n9864), .ZN(
        P1_U3553) );
  NOR2_X1 U10786 ( .A1(n9656), .A2(n9661), .ZN(n9660) );
  NOR4_X1 U10787 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n9678)
         );
  AOI22_X1 U10788 ( .A1(n9853), .A2(n9678), .B1(n9237), .B2(n9864), .ZN(
        P1_U3539) );
  OR2_X1 U10789 ( .A1(n9662), .A2(n9661), .ZN(n9669) );
  OAI22_X1 U10790 ( .A1(n9664), .A2(n9843), .B1(n9663), .B2(n9841), .ZN(n9665)
         );
  INV_X1 U10791 ( .A(n9665), .ZN(n9666) );
  AND2_X1 U10792 ( .A1(n9667), .A2(n9666), .ZN(n9668) );
  AOI22_X1 U10793 ( .A1(n9853), .A2(n9679), .B1(n9670), .B2(n9864), .ZN(
        P1_U3538) );
  OAI211_X1 U10794 ( .C1(n9673), .C2(n9841), .A(n9672), .B(n9671), .ZN(n9674)
         );
  AOI21_X1 U10795 ( .B1(n9675), .B2(n9832), .A(n9674), .ZN(n9681) );
  AOI22_X1 U10796 ( .A1(n9853), .A2(n9681), .B1(n6768), .B2(n9864), .ZN(
        P1_U3536) );
  INV_X1 U10797 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U10798 ( .A1(n9850), .A2(n9677), .B1(n9676), .B2(n9849), .ZN(
        P1_U3521) );
  AOI22_X1 U10799 ( .A1(n9850), .A2(n9678), .B1(n5593), .B2(n9849), .ZN(
        P1_U3502) );
  AOI22_X1 U10800 ( .A1(n9850), .A2(n9679), .B1(n5875), .B2(n9849), .ZN(
        P1_U3499) );
  AOI22_X1 U10801 ( .A1(n9850), .A2(n9681), .B1(n9680), .B2(n9849), .ZN(
        P1_U3493) );
  XNOR2_X1 U10802 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10803 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U10804 ( .A1(n9778), .A2(n9682), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9692) );
  INV_X1 U10805 ( .A(n9792), .ZN(n9760) );
  NAND2_X1 U10806 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9685) );
  AOI211_X1 U10807 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9750), .ZN(n9690)
         );
  AOI211_X1 U10808 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9763), .ZN(n9689)
         );
  AOI211_X1 U10809 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9760), .A(n9690), .B(
        n9689), .ZN(n9691) );
  NAND2_X1 U10810 ( .A1(n9692), .A2(n9691), .ZN(P1_U3242) );
  AOI22_X1 U10811 ( .A1(n9778), .A2(n9694), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n9710) );
  AOI211_X1 U10812 ( .C1(n9697), .C2(n9696), .A(n9695), .B(n9763), .ZN(n9702)
         );
  AOI211_X1 U10813 ( .C1(n9700), .C2(n9699), .A(n9698), .B(n9750), .ZN(n9701)
         );
  AOI211_X1 U10814 ( .C1(n9760), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9702), .B(
        n9701), .ZN(n9709) );
  MUX2_X1 U10815 ( .A(n9704), .B(n9705), .S(n9703), .Z(n9708) );
  NAND2_X1 U10816 ( .A1(n9707), .A2(n9705), .ZN(n9706) );
  OAI211_X1 U10817 ( .C1(n9708), .C2(n9707), .A(P1_U4006), .B(n9706), .ZN(
        n9719) );
  NAND3_X1 U10818 ( .A1(n9710), .A2(n9709), .A3(n9719), .ZN(P1_U3243) );
  OAI21_X1 U10819 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9718) );
  OAI21_X1 U10820 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9717) );
  AOI22_X1 U10821 ( .A1(n9787), .A2(n9718), .B1(n9786), .B2(n9717), .ZN(n9724)
         );
  INV_X1 U10822 ( .A(n9719), .ZN(n9720) );
  AOI211_X1 U10823 ( .C1(n9778), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9723)
         );
  OAI211_X1 U10824 ( .C1(n9725), .C2(n9792), .A(n9724), .B(n9723), .ZN(
        P1_U3245) );
  AOI211_X1 U10825 ( .C1(n9728), .C2(n9727), .A(n9726), .B(n9763), .ZN(n9729)
         );
  AOI211_X1 U10826 ( .C1(n9778), .C2(n9731), .A(n9730), .B(n9729), .ZN(n9736)
         );
  XNOR2_X1 U10827 ( .A(n9733), .B(n9732), .ZN(n9734) );
  AOI22_X1 U10828 ( .A1(n9760), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9786), .B2(
        n9734), .ZN(n9735) );
  NAND2_X1 U10829 ( .A1(n9736), .A2(n9735), .ZN(P1_U3247) );
  INV_X1 U10830 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9749) );
  AOI21_X1 U10831 ( .B1(n9778), .B2(n9738), .A(n9737), .ZN(n9748) );
  OAI21_X1 U10832 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9746) );
  OAI21_X1 U10833 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(n9745) );
  AOI22_X1 U10834 ( .A1(n9787), .A2(n9746), .B1(n9786), .B2(n9745), .ZN(n9747)
         );
  OAI211_X1 U10835 ( .C1(n9792), .C2(n9749), .A(n9748), .B(n9747), .ZN(
        P1_U3248) );
  AOI211_X1 U10836 ( .C1(n9753), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9754)
         );
  AOI211_X1 U10837 ( .C1(n9778), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9762)
         );
  XNOR2_X1 U10838 ( .A(n9758), .B(n9757), .ZN(n9759) );
  AOI22_X1 U10839 ( .A1(n9760), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9787), .B2(
        n9759), .ZN(n9761) );
  NAND2_X1 U10840 ( .A1(n9762), .A2(n9761), .ZN(P1_U3249) );
  AOI211_X1 U10841 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9767)
         );
  AOI211_X1 U10842 ( .C1(n9778), .C2(n9769), .A(n9768), .B(n9767), .ZN(n9775)
         );
  OAI21_X1 U10843 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9773) );
  NAND2_X1 U10844 ( .A1(n9786), .A2(n9773), .ZN(n9774) );
  OAI211_X1 U10845 ( .C1(n10023), .C2(n9792), .A(n9775), .B(n9774), .ZN(
        P1_U3250) );
  INV_X1 U10846 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9791) );
  AOI21_X1 U10847 ( .B1(n9778), .B2(n9777), .A(n9776), .ZN(n9790) );
  OAI21_X1 U10848 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9788) );
  OAI21_X1 U10849 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9785) );
  AOI22_X1 U10850 ( .A1(n9788), .A2(n9787), .B1(n9786), .B2(n9785), .ZN(n9789)
         );
  OAI211_X1 U10851 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n9789), .ZN(
        P1_U3252) );
  AND2_X1 U10852 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9798), .ZN(P1_U3292) );
  AND2_X1 U10853 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9798), .ZN(P1_U3293) );
  AND2_X1 U10854 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9798), .ZN(P1_U3294) );
  NOR2_X1 U10855 ( .A1(n9801), .A2(n9793), .ZN(P1_U3295) );
  AND2_X1 U10856 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9798), .ZN(P1_U3296) );
  AND2_X1 U10857 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9798), .ZN(P1_U3297) );
  AND2_X1 U10858 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9798), .ZN(P1_U3298) );
  AND2_X1 U10859 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9798), .ZN(P1_U3299) );
  AND2_X1 U10860 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9798), .ZN(P1_U3300) );
  NOR2_X1 U10861 ( .A1(n9801), .A2(n9794), .ZN(P1_U3301) );
  AND2_X1 U10862 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9798), .ZN(P1_U3302) );
  AND2_X1 U10863 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9798), .ZN(P1_U3303) );
  NOR2_X1 U10864 ( .A1(n9801), .A2(n9795), .ZN(P1_U3304) );
  AND2_X1 U10865 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9798), .ZN(P1_U3305) );
  AND2_X1 U10866 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9798), .ZN(P1_U3306) );
  AND2_X1 U10867 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9798), .ZN(P1_U3307) );
  AND2_X1 U10868 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9798), .ZN(P1_U3308) );
  AND2_X1 U10869 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9798), .ZN(P1_U3309) );
  AND2_X1 U10870 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9798), .ZN(P1_U3310) );
  AND2_X1 U10871 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9798), .ZN(P1_U3311) );
  AND2_X1 U10872 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9798), .ZN(P1_U3312) );
  AND2_X1 U10873 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9798), .ZN(P1_U3313) );
  AND2_X1 U10874 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9798), .ZN(P1_U3314) );
  AND2_X1 U10875 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9798), .ZN(P1_U3315) );
  NOR2_X1 U10876 ( .A1(n9801), .A2(n9796), .ZN(P1_U3316) );
  AND2_X1 U10877 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9798), .ZN(P1_U3317) );
  NOR2_X1 U10878 ( .A1(n9801), .A2(n9797), .ZN(P1_U3318) );
  AND2_X1 U10879 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9798), .ZN(P1_U3319) );
  NOR2_X1 U10880 ( .A1(n9801), .A2(n9799), .ZN(P1_U3320) );
  NOR2_X1 U10881 ( .A1(n9801), .A2(n9800), .ZN(P1_U3321) );
  INV_X1 U10882 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9803) );
  OAI21_X1 U10883 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(P1_U3441) );
  NOR2_X1 U10884 ( .A1(n9806), .A2(n9805), .ZN(n9809) );
  NOR4_X1 U10885 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n9852)
         );
  AOI22_X1 U10886 ( .A1(n9850), .A2(n9852), .B1(n5635), .B2(n9849), .ZN(
        P1_U3457) );
  OAI22_X1 U10887 ( .A1(n9812), .A2(n9843), .B1(n9811), .B2(n9841), .ZN(n9813)
         );
  AOI21_X1 U10888 ( .B1(n9814), .B2(n9848), .A(n9813), .ZN(n9815) );
  AND2_X1 U10889 ( .A1(n9816), .A2(n9815), .ZN(n9855) );
  AOI22_X1 U10890 ( .A1(n9850), .A2(n9855), .B1(n5661), .B2(n9849), .ZN(
        P1_U3463) );
  OAI21_X1 U10891 ( .B1(n9818), .B2(n9841), .A(n9817), .ZN(n9819) );
  AOI21_X1 U10892 ( .B1(n9820), .B2(n9832), .A(n9819), .ZN(n9821) );
  AND2_X1 U10893 ( .A1(n9822), .A2(n9821), .ZN(n9857) );
  AOI22_X1 U10894 ( .A1(n9850), .A2(n9857), .B1(n5710), .B2(n9849), .ZN(
        P1_U3469) );
  OAI22_X1 U10895 ( .A1(n9824), .A2(n9843), .B1(n9823), .B2(n9841), .ZN(n9826)
         );
  AOI211_X1 U10896 ( .C1(n9848), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9859)
         );
  AOI22_X1 U10897 ( .A1(n9850), .A2(n9859), .B1(n5697), .B2(n9849), .ZN(
        P1_U3472) );
  OAI211_X1 U10898 ( .C1(n9830), .C2(n9841), .A(n9829), .B(n9828), .ZN(n9831)
         );
  AOI21_X1 U10899 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9861) );
  AOI22_X1 U10900 ( .A1(n9850), .A2(n9861), .B1(n5613), .B2(n9849), .ZN(
        P1_U3475) );
  INV_X1 U10901 ( .A(n9834), .ZN(n9839) );
  OAI22_X1 U10902 ( .A1(n9836), .A2(n9843), .B1(n9835), .B2(n9841), .ZN(n9838)
         );
  AOI211_X1 U10903 ( .C1(n9848), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9863)
         );
  INV_X1 U10904 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10905 ( .A1(n9850), .A2(n9863), .B1(n9840), .B2(n9849), .ZN(
        P1_U3478) );
  OAI22_X1 U10906 ( .A1(n9844), .A2(n9843), .B1(n9842), .B2(n9841), .ZN(n9846)
         );
  AOI211_X1 U10907 ( .C1(n9848), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9866)
         );
  AOI22_X1 U10908 ( .A1(n9850), .A2(n9866), .B1(n5754), .B2(n9849), .ZN(
        P1_U3481) );
  INV_X1 U10909 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10910 ( .A1(n9853), .A2(n9852), .B1(n9851), .B2(n9864), .ZN(
        P1_U3524) );
  INV_X1 U10911 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10912 ( .A1(n9853), .A2(n9855), .B1(n9854), .B2(n9864), .ZN(
        P1_U3526) );
  INV_X1 U10913 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U10914 ( .A1(n9853), .A2(n9857), .B1(n9856), .B2(n9864), .ZN(
        P1_U3528) );
  INV_X1 U10915 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10916 ( .A1(n9853), .A2(n9859), .B1(n9858), .B2(n9864), .ZN(
        P1_U3529) );
  INV_X1 U10917 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U10918 ( .A1(n9853), .A2(n9861), .B1(n9860), .B2(n9864), .ZN(
        P1_U3530) );
  INV_X1 U10919 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U10920 ( .A1(n9853), .A2(n9863), .B1(n9862), .B2(n9864), .ZN(
        P1_U3531) );
  AOI22_X1 U10921 ( .A1(n9853), .A2(n9866), .B1(n9865), .B2(n9864), .ZN(
        P1_U3532) );
  AOI22_X1 U10922 ( .A1(n9867), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9868), .ZN(n9877) );
  NAND2_X1 U10923 ( .A1(n9868), .A2(n9966), .ZN(n9870) );
  OAI211_X1 U10924 ( .C1(n9871), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9870), .B(
        n9869), .ZN(n9872) );
  INV_X1 U10925 ( .A(n9872), .ZN(n9875) );
  AOI22_X1 U10926 ( .A1(n9873), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9874) );
  OAI221_X1 U10927 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9877), .C1(n9876), .C2(
        n9875), .A(n9874), .ZN(P2_U3245) );
  AND2_X1 U10928 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9882), .ZN(P2_U3297) );
  AND2_X1 U10929 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9882), .ZN(P2_U3298) );
  AND2_X1 U10930 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9882), .ZN(P2_U3299) );
  INV_X1 U10931 ( .A(n9882), .ZN(n9886) );
  NOR2_X1 U10932 ( .A1(n9886), .A2(n9880), .ZN(P2_U3300) );
  AND2_X1 U10933 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9882), .ZN(P2_U3301) );
  AND2_X1 U10934 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9882), .ZN(P2_U3302) );
  AND2_X1 U10935 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9882), .ZN(P2_U3303) );
  AND2_X1 U10936 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9882), .ZN(P2_U3304) );
  AND2_X1 U10937 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9882), .ZN(P2_U3305) );
  AND2_X1 U10938 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9882), .ZN(P2_U3306) );
  AND2_X1 U10939 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9882), .ZN(P2_U3307) );
  AND2_X1 U10940 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9882), .ZN(P2_U3308) );
  AND2_X1 U10941 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9882), .ZN(P2_U3309) );
  AND2_X1 U10942 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9882), .ZN(P2_U3310) );
  AND2_X1 U10943 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9882), .ZN(P2_U3311) );
  AND2_X1 U10944 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9882), .ZN(P2_U3312) );
  AND2_X1 U10945 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9882), .ZN(P2_U3313) );
  AND2_X1 U10946 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9882), .ZN(P2_U3314) );
  AND2_X1 U10947 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9882), .ZN(P2_U3315) );
  AND2_X1 U10948 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9882), .ZN(P2_U3316) );
  AND2_X1 U10949 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9882), .ZN(P2_U3317) );
  AND2_X1 U10950 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9882), .ZN(P2_U3318) );
  AND2_X1 U10951 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9882), .ZN(P2_U3319) );
  NOR2_X1 U10952 ( .A1(n9886), .A2(n9881), .ZN(P2_U3320) );
  AND2_X1 U10953 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9882), .ZN(P2_U3321) );
  AND2_X1 U10954 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9882), .ZN(P2_U3322) );
  AND2_X1 U10955 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9882), .ZN(P2_U3323) );
  AND2_X1 U10956 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9882), .ZN(P2_U3324) );
  AND2_X1 U10957 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9882), .ZN(P2_U3325) );
  AND2_X1 U10958 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9882), .ZN(P2_U3326) );
  AOI22_X1 U10959 ( .A1(n9885), .A2(n9884), .B1(n9883), .B2(n9882), .ZN(
        P2_U3437) );
  OAI22_X1 U10960 ( .A1(n9888), .A2(n9887), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n9886), .ZN(n9889) );
  INV_X1 U10961 ( .A(n9889), .ZN(P2_U3438) );
  OAI21_X1 U10962 ( .B1(n9892), .B2(n5516), .A(n9891), .ZN(n9893) );
  AOI21_X1 U10963 ( .B1(n9894), .B2(n9962), .A(n9893), .ZN(n9967) );
  INV_X1 U10964 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U10965 ( .A1(n9965), .A2(n9967), .B1(n9895), .B2(n9963), .ZN(
        P2_U3451) );
  AOI22_X1 U10966 ( .A1(n9899), .A2(n9898), .B1(n9897), .B2(n9896), .ZN(n9900)
         );
  NAND2_X1 U10967 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  AOI21_X1 U10968 ( .B1(n9962), .B2(n9903), .A(n9902), .ZN(n9969) );
  INV_X1 U10969 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10970 ( .A1(n9965), .A2(n9969), .B1(n9904), .B2(n9963), .ZN(
        P2_U3457) );
  OAI22_X1 U10971 ( .A1(n9906), .A2(n9957), .B1(n9905), .B2(n9955), .ZN(n9909)
         );
  INV_X1 U10972 ( .A(n9907), .ZN(n9908) );
  AOI211_X1 U10973 ( .C1(n9962), .C2(n9910), .A(n9909), .B(n9908), .ZN(n9970)
         );
  INV_X1 U10974 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10975 ( .A1(n9965), .A2(n9970), .B1(n9911), .B2(n9963), .ZN(
        P2_U3463) );
  INV_X1 U10976 ( .A(n9912), .ZN(n9918) );
  OAI22_X1 U10977 ( .A1(n9914), .A2(n9957), .B1(n9913), .B2(n9955), .ZN(n9917)
         );
  INV_X1 U10978 ( .A(n9915), .ZN(n9916) );
  AOI211_X1 U10979 ( .C1(n9918), .C2(n9962), .A(n9917), .B(n9916), .ZN(n9972)
         );
  INV_X1 U10980 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10981 ( .A1(n9965), .A2(n9972), .B1(n9919), .B2(n9963), .ZN(
        P2_U3469) );
  OAI22_X1 U10982 ( .A1(n9921), .A2(n9957), .B1(n9920), .B2(n9955), .ZN(n9923)
         );
  AOI211_X1 U10983 ( .C1(n9962), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9974)
         );
  INV_X1 U10984 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U10985 ( .A1(n9965), .A2(n9974), .B1(n9925), .B2(n9963), .ZN(
        P2_U3472) );
  INV_X1 U10986 ( .A(n9926), .ZN(n9931) );
  OAI22_X1 U10987 ( .A1(n9928), .A2(n9957), .B1(n9927), .B2(n9955), .ZN(n9930)
         );
  AOI211_X1 U10988 ( .C1(n9947), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9976)
         );
  INV_X1 U10989 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U10990 ( .A1(n9965), .A2(n9976), .B1(n9932), .B2(n9963), .ZN(
        P2_U3475) );
  INV_X1 U10991 ( .A(n9933), .ZN(n9938) );
  OAI22_X1 U10992 ( .A1(n9935), .A2(n9957), .B1(n9934), .B2(n9955), .ZN(n9937)
         );
  AOI211_X1 U10993 ( .C1(n9947), .C2(n9938), .A(n9937), .B(n9936), .ZN(n9977)
         );
  INV_X1 U10994 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U10995 ( .A1(n9965), .A2(n9977), .B1(n9939), .B2(n9963), .ZN(
        P2_U3478) );
  INV_X1 U10996 ( .A(n9940), .ZN(n9946) );
  INV_X1 U10997 ( .A(n9941), .ZN(n9942) );
  OAI22_X1 U10998 ( .A1(n9943), .A2(n9957), .B1(n9942), .B2(n9955), .ZN(n9945)
         );
  AOI211_X1 U10999 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9978)
         );
  AOI22_X1 U11000 ( .A1(n9965), .A2(n9978), .B1(n9948), .B2(n9963), .ZN(
        P2_U3481) );
  OAI22_X1 U11001 ( .A1(n9950), .A2(n9957), .B1(n9949), .B2(n9955), .ZN(n9952)
         );
  AOI211_X1 U11002 ( .C1(n9953), .C2(n9962), .A(n9952), .B(n9951), .ZN(n9979)
         );
  INV_X1 U11003 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11004 ( .A1(n9965), .A2(n9979), .B1(n9954), .B2(n9963), .ZN(
        P2_U3484) );
  OAI22_X1 U11005 ( .A1(n9958), .A2(n9957), .B1(n9956), .B2(n9955), .ZN(n9960)
         );
  AOI211_X1 U11006 ( .C1(n9962), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9982)
         );
  INV_X1 U11007 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11008 ( .A1(n9965), .A2(n9982), .B1(n9964), .B2(n9963), .ZN(
        P2_U3487) );
  AOI22_X1 U11009 ( .A1(n9983), .A2(n9967), .B1(n9966), .B2(n9980), .ZN(
        P2_U3520) );
  INV_X1 U11010 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9968) );
  AOI22_X1 U11011 ( .A1(n9983), .A2(n9969), .B1(n9968), .B2(n9980), .ZN(
        P2_U3522) );
  AOI22_X1 U11012 ( .A1(n9983), .A2(n9970), .B1(n6355), .B2(n9980), .ZN(
        P2_U3524) );
  INV_X1 U11013 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11014 ( .A1(n9983), .A2(n9972), .B1(n9971), .B2(n9980), .ZN(
        P2_U3526) );
  INV_X1 U11015 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U11016 ( .A1(n9983), .A2(n9974), .B1(n9973), .B2(n9980), .ZN(
        P2_U3527) );
  INV_X1 U11017 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U11018 ( .A1(n9983), .A2(n9976), .B1(n9975), .B2(n9980), .ZN(
        P2_U3528) );
  AOI22_X1 U11019 ( .A1(n9983), .A2(n9977), .B1(n6512), .B2(n9980), .ZN(
        P2_U3529) );
  AOI22_X1 U11020 ( .A1(n9983), .A2(n9978), .B1(n6623), .B2(n9980), .ZN(
        P2_U3530) );
  AOI22_X1 U11021 ( .A1(n9983), .A2(n9979), .B1(n6789), .B2(n9980), .ZN(
        P2_U3531) );
  AOI22_X1 U11022 ( .A1(n9983), .A2(n9982), .B1(n9981), .B2(n9980), .ZN(
        P2_U3532) );
  INV_X1 U11023 ( .A(n9984), .ZN(n9985) );
  NAND2_X1 U11024 ( .A1(n9986), .A2(n9985), .ZN(n9987) );
  XNOR2_X1 U11025 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9987), .ZN(ADD_1071_U5) );
  XOR2_X1 U11026 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11027 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(ADD_1071_U56) );
  OAI21_X1 U11028 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(ADD_1071_U57) );
  OAI21_X1 U11029 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(ADD_1071_U58) );
  OAI21_X1 U11030 ( .B1(n9999), .B2(n9998), .A(n9997), .ZN(ADD_1071_U59) );
  OAI21_X1 U11031 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(ADD_1071_U60) );
  OAI21_X1 U11032 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(ADD_1071_U61) );
  AOI21_X1 U11033 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(ADD_1071_U62) );
  AOI21_X1 U11034 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11035 ( .A(n10013), .B(n10012), .ZN(ADD_1071_U50) );
  NOR2_X1 U11036 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  XOR2_X1 U11037 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10016), .Z(ADD_1071_U51) );
  OAI21_X1 U11038 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  XNOR2_X1 U11039 ( .A(n10020), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11040 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(ADD_1071_U47) );
  XOR2_X1 U11041 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10024), .Z(ADD_1071_U48) );
  XOR2_X1 U11042 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10025), .Z(ADD_1071_U49) );
  XOR2_X1 U11043 ( .A(n10027), .B(n10026), .Z(ADD_1071_U54) );
  XOR2_X1 U11044 ( .A(n10029), .B(n10028), .Z(ADD_1071_U53) );
  XNOR2_X1 U11045 ( .A(n10031), .B(n10030), .ZN(ADD_1071_U52) );
  INV_X1 U4821 ( .A(n8010), .ZN(n4313) );
  CLKBUF_X1 U4837 ( .A(n8010), .Z(n4314) );
  CLKBUF_X1 U4848 ( .A(n5530), .Z(n4310) );
  CLKBUF_X1 U4861 ( .A(n8010), .Z(n4315) );
  CLKBUF_X1 U4867 ( .A(n5518), .Z(n4316) );
endmodule

