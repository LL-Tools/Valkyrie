

module b20_C_SARLock_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4416, n4417, n4418, n4419, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401;

  OAI21_X1 U4923 ( .B1(n6929), .B2(n6931), .A(n6930), .ZN(n7098) );
  INV_X1 U4924 ( .A(n6776), .ZN(n4419) );
  INV_X2 U4925 ( .A(n6776), .ZN(n7808) );
  INV_X2 U4926 ( .A(n5880), .ZN(n6844) );
  INV_X1 U4927 ( .A(n5148), .ZN(n5352) );
  INV_X1 U4928 ( .A(n6973), .ZN(n5722) );
  INV_X1 U4929 ( .A(n6127), .ZN(n6139) );
  CLKBUF_X2 U4930 ( .A(n6501), .Z(n4417) );
  INV_X1 U4931 ( .A(n7696), .ZN(n7812) );
  NAND2_X1 U4932 ( .A1(n6739), .A2(n6740), .ZN(n6746) );
  INV_X1 U4933 ( .A(n7826), .ZN(n7807) );
  INV_X1 U4934 ( .A(n5377), .ZN(n5429) );
  AOI211_X1 U4935 ( .C1(n4416), .C2(n5009), .A(n9778), .B(n7588), .ZN(n7463)
         );
  INV_X1 U4936 ( .A(n7335), .ZN(n6659) );
  INV_X1 U4937 ( .A(n5376), .ZN(n5428) );
  NAND2_X1 U4939 ( .A1(n9770), .A2(n5848), .ZN(n9769) );
  NAND2_X1 U4940 ( .A1(n7699), .A2(n9928), .ZN(n7453) );
  INV_X1 U4941 ( .A(n9299), .ZN(n7699) );
  NAND2_X1 U4942 ( .A1(n5381), .A2(n10021), .ZN(n5167) );
  INV_X1 U4943 ( .A(n5953), .ZN(n7968) );
  AOI211_X1 U4945 ( .C1(n8183), .C2(n10191), .A(n8182), .B(n8181), .ZN(n8184)
         );
  NAND2_X2 U4946 ( .A1(n9644), .A2(n4996), .ZN(n9647) );
  NAND2_X2 U4947 ( .A1(n4955), .A2(n4954), .ZN(n9644) );
  NAND4_X4 U4948 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n6777)
         );
  OAI22_X2 U4949 ( .A1(n7553), .A2(n6294), .B1(n8688), .B2(n7906), .ZN(n8684)
         );
  NAND2_X2 U4950 ( .A1(n6293), .A2(n6292), .ZN(n7553) );
  AOI211_X2 U4951 ( .C1(n7854), .C2(n7853), .A(n7847), .B(n7852), .ZN(n7861)
         );
  OAI21_X2 U4952 ( .B1(n9226), .B2(n7705), .A(n7704), .ZN(n9204) );
  OAI211_X1 U4953 ( .C1(n5143), .C2(n6411), .A(n5213), .B(n5212), .ZN(n9299)
         );
  NOR2_X2 U4954 ( .A1(n6823), .A2(n6824), .ZN(n6875) );
  INV_X1 U4955 ( .A(n10184), .ZN(n4418) );
  OAI211_X1 U4956 ( .C1(n6429), .C2(n10050), .A(n5207), .B(n5206), .ZN(n10184)
         );
  INV_X1 U4957 ( .A(n6741), .ZN(n8767) );
  NAND2_X1 U4958 ( .A1(n5408), .A2(n5407), .ZN(n6665) );
  CLKBUF_X2 U4959 ( .A(n5943), .Z(n4423) );
  INV_X1 U4960 ( .A(n5904), .ZN(n5907) );
  NAND2_X1 U4961 ( .A1(n5903), .A2(n5902), .ZN(n8869) );
  CLKBUF_X1 U4962 ( .A(n5167), .Z(n6429) );
  MUX2_X1 U4963 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5901), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5903) );
  OR2_X1 U4964 ( .A1(n4424), .A2(n9038), .ZN(n5012) );
  NOR2_X1 U4965 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5168) );
  AND2_X1 U4966 ( .A1(n9531), .A2(n9530), .ZN(n9540) );
  AND2_X1 U4967 ( .A1(n8197), .A2(n8196), .ZN(n8204) );
  AND2_X1 U4968 ( .A1(n4545), .A2(n4544), .ZN(n9193) );
  NAND2_X1 U4969 ( .A1(n9595), .A2(n4448), .ZN(n9594) );
  OR2_X1 U4970 ( .A1(n9325), .A2(n9324), .ZN(n4545) );
  NAND2_X1 U4971 ( .A1(n9236), .A2(n7785), .ZN(n9188) );
  AOI21_X1 U4972 ( .B1(n4634), .B2(n4633), .A(n4630), .ZN(n7967) );
  NAND2_X1 U4973 ( .A1(n4550), .A2(n4554), .ZN(n9214) );
  NAND2_X1 U4974 ( .A1(n8629), .A2(n4738), .ZN(n8736) );
  NAND2_X1 U4975 ( .A1(n9691), .A2(n5856), .ZN(n9676) );
  AOI21_X1 U4976 ( .B1(n9814), .B2(n10280), .A(n9813), .ZN(n4948) );
  OR2_X1 U4977 ( .A1(n8188), .A2(n8168), .ZN(n9515) );
  NAND2_X1 U4978 ( .A1(n7744), .A2(n7743), .ZN(n4537) );
  OR2_X1 U4979 ( .A1(n8169), .A2(n4518), .ZN(n4533) );
  OR2_X1 U4980 ( .A1(n8189), .A2(n4519), .ZN(n4534) );
  AND2_X1 U4981 ( .A1(n4539), .A2(n4538), .ZN(n7741) );
  NAND2_X1 U4982 ( .A1(n9740), .A2(n5853), .ZN(n9723) );
  OAI21_X1 U4983 ( .B1(n7303), .B2(n4784), .A(n4783), .ZN(n6293) );
  INV_X1 U4984 ( .A(n4779), .ZN(n4783) );
  OAI21_X1 U4985 ( .B1(n4781), .B2(n4780), .A(n8014), .ZN(n4779) );
  OR2_X1 U4986 ( .A1(n7191), .A2(n4867), .ZN(n4866) );
  AOI21_X1 U4987 ( .B1(n7292), .B2(n7291), .A(n4998), .ZN(n7293) );
  AND2_X1 U4988 ( .A1(n5234), .A2(n5233), .ZN(n8118) );
  NAND2_X1 U4989 ( .A1(n6050), .A2(n6049), .ZN(n7633) );
  NAND2_X1 U4990 ( .A1(n4620), .A2(n4619), .ZN(n5218) );
  NAND2_X1 U4991 ( .A1(n4548), .A2(n4547), .ZN(n7483) );
  AOI21_X1 U4992 ( .B1(n7092), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6773), .ZN(
        n6775) );
  OAI211_X1 U4993 ( .C1(n6429), .C2(n6398), .A(n5182), .B(n5181), .ZN(n7381)
         );
  NAND2_X1 U4994 ( .A1(n4994), .A2(n4993), .ZN(n6890) );
  AND4_X1 U4995 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n6997)
         );
  INV_X4 U4997 ( .A(n7679), .ZN(n4982) );
  AND2_X1 U4998 ( .A1(n7017), .A2(n6665), .ZN(n6660) );
  INV_X2 U4999 ( .A(n9394), .ZN(P1_U3973) );
  NAND2_X1 U5000 ( .A1(n6659), .A2(n7281), .ZN(n6663) );
  NAND2_X2 U5001 ( .A1(n6318), .A2(n6417), .ZN(n6385) );
  NOR2_X1 U5002 ( .A1(n8117), .A2(n7637), .ZN(n5408) );
  XNOR2_X1 U5003 ( .A(n5386), .B(n5385), .ZN(n8049) );
  INV_X2 U5004 ( .A(n6414), .ZN(n8489) );
  NOR2_X1 U5005 ( .A1(n4719), .A2(n4723), .ZN(n4718) );
  INV_X1 U5006 ( .A(n5185), .ZN(n4723) );
  AND2_X1 U5007 ( .A1(n5029), .A2(n5028), .ZN(n5154) );
  NAND2_X1 U5008 ( .A1(n5367), .A2(n5366), .ZN(n7281) );
  NAND2_X1 U5009 ( .A1(n5364), .A2(n5409), .ZN(n7538) );
  XNOR2_X1 U5010 ( .A(n5359), .B(n5358), .ZN(n7335) );
  AND2_X1 U5011 ( .A1(n5044), .A2(n5043), .ZN(n5185) );
  NAND2_X1 U5012 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5359) );
  AND2_X1 U5013 ( .A1(n5034), .A2(n5033), .ZN(n5165) );
  NAND2_X1 U5014 ( .A1(n5902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5899) );
  AND2_X1 U5015 ( .A1(n6271), .A2(n4433), .ZN(n5914) );
  INV_X2 U5016 ( .A(n10013), .ZN(n8174) );
  OR2_X1 U5017 ( .A1(n6436), .A2(n6697), .ZN(n6464) );
  INV_X2 U5018 ( .A(n9175), .ZN(n8874) );
  NAND2_X1 U5019 ( .A1(n4778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6332) );
  AND2_X1 U5020 ( .A1(n5127), .A2(n4939), .ZN(n4938) );
  OAI211_X1 U5021 ( .C1(n5925), .C2(n4884), .A(n5937), .B(n4883), .ZN(n6501)
         );
  NOR2_X1 U5022 ( .A1(n5887), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4574) );
  NAND4_X1 U5023 ( .A1(n5886), .A2(n5885), .A3(n5998), .A4(n5959), .ZN(n5887)
         );
  AND4_X1 U5024 ( .A1(n5219), .A2(n5126), .A3(n5230), .A4(n5225), .ZN(n5127)
         );
  AND2_X1 U5025 ( .A1(n4953), .A2(n8881), .ZN(n5149) );
  INV_X1 U5026 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4727) );
  INV_X1 U5027 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6103) );
  INV_X1 U5028 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5230) );
  NOR2_X1 U5029 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5885) );
  INV_X1 U5030 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5128) );
  INV_X1 U5031 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5998) );
  NOR2_X1 U5032 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4952) );
  NOR2_X1 U5033 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4990) );
  INV_X1 U5034 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6046) );
  NOR2_X1 U5035 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5126) );
  NOR2_X1 U5036 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5219) );
  INV_X4 U5037 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5038 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5039 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6104) );
  AND2_X1 U5040 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6909) );
  NAND2_X2 U5041 ( .A1(n9769), .A2(n4440), .ZN(n9736) );
  OAI22_X2 U5042 ( .A1(n8588), .A2(n8595), .B1(n8596), .B2(n8605), .ZN(n8576)
         );
  BUF_X2 U5043 ( .A(n5941), .Z(n4421) );
  XNOR2_X2 U5044 ( .A(n5370), .B(n5133), .ZN(n5381) );
  NAND2_X2 U5045 ( .A1(n4692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  NAND2_X4 U5046 ( .A1(n6665), .A2(n4812), .ZN(n6776) );
  CLKBUF_X1 U5047 ( .A(n5943), .Z(n4422) );
  AND2_X1 U5048 ( .A1(n5904), .A2(n8869), .ZN(n5943) );
  AND2_X1 U5049 ( .A1(n4887), .A2(n4888), .ZN(n4424) );
  AND2_X1 U5050 ( .A1(n4887), .A2(n4888), .ZN(n4425) );
  INV_X8 U5051 ( .A(n6392), .ZN(n5928) );
  INV_X1 U5052 ( .A(n7696), .ZN(n4426) );
  AND2_X1 U5053 ( .A1(n8791), .A2(n8258), .ZN(n7960) );
  OR2_X1 U5054 ( .A1(n8803), .A2(n8561), .ZN(n5003) );
  OR2_X1 U5055 ( .A1(n8842), .A2(n8276), .ZN(n7923) );
  XNOR2_X1 U5056 ( .A(n5336), .B(n5335), .ZN(n5339) );
  OR2_X1 U5057 ( .A1(n5288), .A2(n5287), .ZN(n4629) );
  NAND2_X1 U5058 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5913) );
  INV_X1 U5059 ( .A(n6746), .ZN(n8106) );
  NAND2_X1 U5060 ( .A1(n8785), .A2(n8526), .ZN(n6312) );
  INV_X1 U5061 ( .A(n5708), .ZN(n5697) );
  INV_X1 U5062 ( .A(n5711), .ZN(n5695) );
  MUX2_X1 U5063 ( .A(n7851), .B(n7850), .S(n7973), .Z(n7852) );
  NOR2_X1 U5064 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  INV_X1 U5065 ( .A(n8568), .ZN(n4852) );
  AND2_X1 U5066 ( .A1(n4849), .A2(n4640), .ZN(n4846) );
  NAND2_X1 U5067 ( .A1(n4847), .A2(n4850), .ZN(n4640) );
  INV_X1 U5068 ( .A(n7956), .ZN(n4849) );
  INV_X1 U5069 ( .A(n7959), .ZN(n4843) );
  NAND2_X1 U5070 ( .A1(n7760), .A2(n9272), .ZN(n4559) );
  AND2_X1 U5071 ( .A1(n4509), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U5072 ( .A1(n5090), .A2(n5296), .ZN(n4908) );
  AOI21_X1 U5073 ( .B1(n7411), .B2(n7410), .A(n7409), .ZN(n7412) );
  INV_X1 U5074 ( .A(n7629), .ZN(n4963) );
  INV_X1 U5075 ( .A(n6764), .ZN(n4978) );
  OR2_X1 U5076 ( .A1(n7675), .A2(n6266), .ZN(n7985) );
  NOR2_X1 U5077 ( .A1(n8785), .A2(n8336), .ZN(n7963) );
  OR2_X1 U5078 ( .A1(n8803), .A2(n8285), .ZN(n7996) );
  NOR2_X1 U5079 ( .A1(n6304), .A2(n6305), .ZN(n4774) );
  NOR2_X1 U5080 ( .A1(n4767), .A2(n5887), .ZN(n4766) );
  AND2_X1 U5081 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  NAND2_X1 U5082 ( .A1(n9636), .A2(n9666), .ZN(n4601) );
  AND2_X1 U5083 ( .A1(n9629), .A2(n8151), .ZN(n4947) );
  NOR2_X1 U5084 ( .A1(n9725), .A2(n9747), .ZN(n4603) );
  NOR2_X1 U5085 ( .A1(n9804), .A2(n10257), .ZN(n4605) );
  XNOR2_X1 U5086 ( .A(n6777), .B(n5469), .ZN(n6837) );
  AND2_X1 U5087 ( .A1(n8159), .A2(n8158), .ZN(n4956) );
  NAND2_X1 U5088 ( .A1(n9563), .A2(n9576), .ZN(n8158) );
  OR2_X1 U5089 ( .A1(n9956), .A2(n9566), .ZN(n8156) );
  NAND2_X1 U5090 ( .A1(n9650), .A2(n9664), .ZN(n5776) );
  NOR2_X1 U5091 ( .A1(n9395), .A2(n8056), .ZN(n6962) );
  NAND2_X1 U5092 ( .A1(n5117), .A2(n5116), .ZN(n5327) );
  AND2_X1 U5093 ( .A1(n5122), .A2(n5121), .ZN(n5328) );
  NAND2_X1 U5094 ( .A1(n4905), .A2(n4626), .ZN(n4625) );
  INV_X1 U5095 ( .A(n5307), .ZN(n4626) );
  NAND2_X1 U5096 ( .A1(n4453), .A2(n4827), .ZN(n4826) );
  AND2_X1 U5097 ( .A1(n5129), .A2(n4828), .ZN(n4827) );
  INV_X1 U5098 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5129) );
  INV_X1 U5099 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U5100 ( .A1(n4629), .A2(n5089), .ZN(n5299) );
  NAND2_X1 U5101 ( .A1(n4925), .A2(n4923), .ZN(n5288) );
  INV_X1 U5102 ( .A(n4924), .ZN(n4923) );
  OAI21_X1 U5103 ( .B1(n4928), .B2(n5084), .A(n5083), .ZN(n4924) );
  NAND2_X1 U5104 ( .A1(n4636), .A2(n9032), .ZN(n5072) );
  NAND2_X1 U5105 ( .A1(n4932), .A2(n4931), .ZN(n4636) );
  INV_X1 U5106 ( .A(n4933), .ZN(n4931) );
  AND2_X1 U5107 ( .A1(n5214), .A2(n4450), .ZN(n4619) );
  OR2_X1 U5108 ( .A1(n8263), .A2(n8659), .ZN(n4586) );
  NAND2_X1 U5109 ( .A1(n4969), .A2(n4967), .ZN(n8262) );
  AND2_X1 U5110 ( .A1(n4968), .A2(n4492), .ZN(n4967) );
  NAND2_X1 U5111 ( .A1(n8215), .A2(n4445), .ZN(n4969) );
  NAND2_X1 U5112 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  OR2_X1 U5113 ( .A1(n8098), .A2(n8545), .ZN(n8099) );
  OAI21_X1 U5114 ( .B1(n4736), .B2(n8037), .A(n4431), .ZN(n4734) );
  AND2_X1 U5115 ( .A1(n8036), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5116 ( .A1(n4477), .A2(n8034), .ZN(n4737) );
  AND2_X1 U5117 ( .A1(n7967), .A2(n7966), .ZN(n7978) );
  NAND2_X1 U5118 ( .A1(n7085), .A2(n6284), .ZN(n4810) );
  NAND2_X1 U5119 ( .A1(n4740), .A2(n4741), .ZN(n8514) );
  AOI21_X1 U5120 ( .B1(n4473), .B2(n4743), .A(n4436), .ZN(n4741) );
  AOI21_X1 U5121 ( .B1(n4804), .B2(n4806), .A(n4803), .ZN(n4802) );
  NOR2_X1 U5122 ( .A1(n8797), .A2(n8545), .ZN(n4803) );
  NAND2_X1 U5123 ( .A1(n8809), .A2(n8307), .ZN(n8550) );
  OR2_X1 U5124 ( .A1(n6309), .A2(n8307), .ZN(n5002) );
  AOI21_X1 U5125 ( .B1(n4755), .B2(n4758), .A(n4754), .ZN(n4753) );
  INV_X1 U5126 ( .A(n5952), .ZN(n7677) );
  INV_X1 U5127 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4979) );
  OR2_X1 U5128 ( .A1(n9238), .A2(n4818), .ZN(n4817) );
  INV_X1 U5129 ( .A(n6663), .ZN(n4812) );
  AND4_X1 U5130 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n9631)
         );
  AND2_X1 U5131 ( .A1(n9705), .A2(n5854), .ZN(n4949) );
  OR2_X1 U5132 ( .A1(n9804), .A2(n10274), .ZN(n9771) );
  NAND2_X1 U5133 ( .A1(n6672), .A2(n10005), .ZN(n6952) );
  AND2_X1 U5134 ( .A1(n7610), .A2(n5844), .ZN(n4951) );
  INV_X1 U5135 ( .A(n5143), .ZN(n5293) );
  INV_X1 U5136 ( .A(n6429), .ZN(n5292) );
  OAI21_X1 U5137 ( .B1(n9556), .B2(n8143), .A(n8142), .ZN(n9541) );
  AOI21_X1 U5138 ( .B1(n4430), .B2(n4667), .A(n4502), .ZN(n4663) );
  NAND2_X1 U5139 ( .A1(n4602), .A2(n9699), .ZN(n4682) );
  INV_X1 U5140 ( .A(n4683), .ZN(n4681) );
  OAI21_X1 U5141 ( .B1(n5339), .B2(n5338), .A(n5337), .ZN(n5346) );
  OR2_X1 U5142 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  INV_X1 U5143 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4813) );
  INV_X1 U5144 ( .A(n10156), .ZN(n10175) );
  AOI21_X1 U5145 ( .B1(n10014), .B2(n5352), .A(n5351), .ZN(n9514) );
  OAI21_X1 U5146 ( .B1(n7845), .B2(n4856), .A(n4854), .ZN(n7849) );
  NAND2_X1 U5147 ( .A1(n4857), .A2(n8034), .ZN(n4856) );
  NAND2_X1 U5148 ( .A1(n7846), .A2(n4855), .ZN(n4854) );
  AOI21_X1 U5149 ( .B1(n4833), .B2(n7868), .A(n4832), .ZN(n4836) );
  OAI21_X1 U5150 ( .B1(n4835), .B2(n4834), .A(n7862), .ZN(n4833) );
  NAND2_X1 U5151 ( .A1(n7875), .A2(n7874), .ZN(n4531) );
  NOR2_X1 U5152 ( .A1(n7873), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U5153 ( .A1(n4694), .A2(n4458), .ZN(n4693) );
  OAI21_X1 U5154 ( .B1(n4700), .B2(n4469), .A(n4699), .ZN(n4698) );
  NOR2_X1 U5155 ( .A1(n8695), .A2(n7909), .ZN(n4862) );
  OAI21_X1 U5156 ( .B1(n4464), .B2(n4526), .A(n9705), .ZN(n5639) );
  OAI21_X1 U5157 ( .B1(n5607), .B2(n6845), .A(n5611), .ZN(n4526) );
  INV_X1 U5158 ( .A(n9613), .ZN(n4726) );
  AND3_X1 U5159 ( .A1(n7939), .A2(n7929), .A3(n7937), .ZN(n7932) );
  NAND2_X1 U5160 ( .A1(n7950), .A2(n7977), .ZN(n4638) );
  NAND2_X1 U5161 ( .A1(n8161), .A2(n6845), .ZN(n4715) );
  AND2_X1 U5162 ( .A1(n7458), .A2(n5527), .ZN(n5739) );
  AOI21_X1 U5163 ( .B1(n4842), .B2(n4840), .A(n8524), .ZN(n4635) );
  NOR2_X1 U5164 ( .A1(n4845), .A2(n4843), .ZN(n4842) );
  INV_X1 U5165 ( .A(n4846), .ZN(n4845) );
  OR2_X1 U5166 ( .A1(n4844), .A2(n4843), .ZN(n4841) );
  AOI21_X1 U5167 ( .B1(n4846), .B2(n4460), .A(n4805), .ZN(n4844) );
  OR2_X1 U5168 ( .A1(n4847), .A2(n4851), .ZN(n4639) );
  INV_X1 U5169 ( .A(n7965), .ZN(n4631) );
  INV_X1 U5170 ( .A(n6885), .ZN(n4797) );
  AND2_X1 U5171 ( .A1(n4559), .A2(n9264), .ZN(n4555) );
  NAND2_X1 U5172 ( .A1(n4507), .A2(n4559), .ZN(n4554) );
  OAI21_X1 U5173 ( .B1(n8114), .B2(n4912), .A(n4910), .ZN(n5767) );
  INV_X1 U5174 ( .A(n5343), .ZN(n4912) );
  AND2_X1 U5175 ( .A1(n5760), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U5176 ( .A1(n5343), .A2(n5148), .ZN(n4911) );
  OAI21_X1 U5177 ( .B1(n9604), .B2(n9842), .A(n8137), .ZN(n8138) );
  OR2_X1 U5178 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  INV_X1 U5179 ( .A(n5122), .ZN(n4901) );
  INV_X1 U5180 ( .A(n4900), .ZN(n4899) );
  OAI21_X1 U5181 ( .B1(n5328), .B2(n4901), .A(n5332), .ZN(n4900) );
  NOR2_X1 U5182 ( .A1(n8297), .A2(n4981), .ZN(n4980) );
  INV_X1 U5183 ( .A(n5000), .ZN(n4981) );
  OR2_X1 U5184 ( .A1(n8034), .A2(n8037), .ZN(n6736) );
  NAND2_X1 U5185 ( .A1(n4445), .A2(n8216), .ZN(n4968) );
  INV_X1 U5186 ( .A(n6765), .ZN(n6762) );
  NAND2_X1 U5187 ( .A1(n7045), .A2(n4535), .ZN(n7170) );
  NAND2_X1 U5188 ( .A1(n4536), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4535) );
  AND2_X1 U5189 ( .A1(n6193), .A2(n9010), .ZN(n6195) );
  OR2_X1 U5190 ( .A1(n8596), .A2(n8579), .ZN(n7943) );
  OR2_X1 U5191 ( .A1(n7633), .A2(n7599), .ZN(n7898) );
  INV_X1 U5192 ( .A(n6290), .ZN(n4789) );
  OR2_X1 U5193 ( .A1(n8251), .A2(n8085), .ZN(n7945) );
  NOR2_X1 U5194 ( .A1(n7919), .A2(n7844), .ZN(n4759) );
  OR2_X1 U5195 ( .A1(n8848), .A2(n8672), .ZN(n7916) );
  NAND2_X1 U5196 ( .A1(n8485), .A2(n8037), .ZN(n6739) );
  NAND2_X1 U5197 ( .A1(n6044), .A2(n4428), .ZN(n6105) );
  INV_X1 U5198 ( .A(n7785), .ZN(n4818) );
  INV_X1 U5199 ( .A(n7691), .ZN(n4822) );
  NAND2_X1 U5200 ( .A1(n4546), .A2(n4457), .ZN(n7282) );
  NAND2_X1 U5201 ( .A1(n7821), .A2(n7483), .ZN(n4546) );
  AND2_X1 U5202 ( .A1(n5714), .A2(n5427), .ZN(n5869) );
  OR2_X1 U5203 ( .A1(n9814), .A2(n9548), .ZN(n8161) );
  OR2_X1 U5204 ( .A1(n9563), .A2(n9956), .ZN(n4607) );
  OR2_X1 U5205 ( .A1(n9914), .A2(n10276), .ZN(n5851) );
  OR2_X1 U5206 ( .A1(n10004), .A2(n5406), .ZN(n6672) );
  INV_X1 U5207 ( .A(n4672), .ZN(n4671) );
  OAI21_X1 U5208 ( .B1(n7583), .B2(n4673), .A(n8120), .ZN(n4672) );
  INV_X1 U5209 ( .A(n7608), .ZN(n4673) );
  OR2_X1 U5210 ( .A1(n10257), .A2(n9794), .ZN(n9790) );
  INV_X1 U5211 ( .A(n7281), .ZN(n6673) );
  OR2_X1 U5212 ( .A1(n8188), .A2(n9528), .ZN(n5828) );
  OR2_X1 U5213 ( .A1(n9946), .A2(n9527), .ZN(n8160) );
  NOR2_X1 U5214 ( .A1(n9598), .A2(n9956), .ZN(n9581) );
  OR2_X1 U5215 ( .A1(n9838), .A2(n9842), .ZN(n8155) );
  OR2_X1 U5216 ( .A1(n9665), .A2(n4599), .ZN(n9619) );
  INV_X1 U5217 ( .A(n4601), .ZN(n4600) );
  NAND2_X1 U5218 ( .A1(n6392), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4942) );
  NOR2_X1 U5219 ( .A1(n4959), .A2(n5132), .ZN(n4958) );
  NAND2_X1 U5220 ( .A1(n4960), .A2(n5410), .ZN(n4959) );
  INV_X1 U5221 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U5222 ( .A1(n4891), .A2(n4889), .ZN(n5324) );
  AOI21_X1 U5223 ( .B1(n4893), .B2(n4895), .A(n4890), .ZN(n4889) );
  INV_X1 U5224 ( .A(n5111), .ZN(n4890) );
  AND2_X1 U5225 ( .A1(n5111), .A2(n5110), .ZN(n5320) );
  NAND2_X1 U5226 ( .A1(n4915), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5227 ( .A1(n5205), .A2(n5052), .ZN(n4611) );
  NOR2_X1 U5228 ( .A1(n4618), .A2(n4614), .ZN(n4613) );
  INV_X1 U5229 ( .A(n5052), .ZN(n4614) );
  NOR2_X1 U5230 ( .A1(n4616), .A2(n4914), .ZN(n4615) );
  NAND2_X1 U5231 ( .A1(n4619), .A2(n4617), .ZN(n4616) );
  NOR2_X1 U5232 ( .A1(n5223), .A2(n4920), .ZN(n4919) );
  INV_X1 U5233 ( .A(n5059), .ZN(n4920) );
  XNOR2_X1 U5234 ( .A(n5060), .B(SI_11_), .ZN(n5223) );
  OR2_X1 U5235 ( .A1(n5204), .A2(n5205), .ZN(n4608) );
  XNOR2_X1 U5236 ( .A(n5049), .B(SI_8_), .ZN(n5205) );
  NAND2_X1 U5237 ( .A1(n5193), .A2(n5048), .ZN(n5204) );
  INV_X1 U5238 ( .A(n5177), .ZN(n4719) );
  INV_X1 U5239 ( .A(n5039), .ZN(n4722) );
  INV_X1 U5240 ( .A(SI_7_), .ZN(n9071) );
  OAI21_X1 U5241 ( .B1(n5928), .B2(n5024), .A(n5023), .ZN(n5025) );
  OR2_X1 U5242 ( .A1(n8103), .A2(n8102), .ZN(n5007) );
  OR2_X1 U5243 ( .A1(n8082), .A2(n8605), .ZN(n8083) );
  XNOR2_X1 U5244 ( .A(n6890), .B(n6746), .ZN(n6758) );
  INV_X1 U5245 ( .A(n7338), .ZN(n4589) );
  NAND2_X1 U5246 ( .A1(n4592), .A2(n7338), .ZN(n4590) );
  INV_X1 U5247 ( .A(n7442), .ZN(n7425) );
  OR2_X1 U5248 ( .A1(n7597), .A2(n4963), .ZN(n4962) );
  OAI21_X1 U5249 ( .B1(n7597), .B2(n4474), .A(n8688), .ZN(n4965) );
  INV_X1 U5250 ( .A(n4578), .ZN(n4577) );
  OAI21_X1 U5251 ( .B1(n4980), .B2(n4579), .A(n8247), .ZN(n4578) );
  INV_X1 U5252 ( .A(n8083), .ZN(n4579) );
  NAND2_X1 U5253 ( .A1(n4520), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U5254 ( .A1(n7595), .A2(n7596), .ZN(n4573) );
  OAI21_X1 U5255 ( .B1(n4586), .B2(n4584), .A(n8271), .ZN(n4583) );
  NOR2_X1 U5256 ( .A1(n4974), .A2(n4588), .ZN(n4592) );
  INV_X1 U5257 ( .A(n7008), .ZN(n4588) );
  INV_X1 U5258 ( .A(n6323), .ZN(n6260) );
  NAND2_X1 U5259 ( .A1(n4881), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U5260 ( .A1(n6496), .A2(n6517), .ZN(n6525) );
  OR2_X1 U5261 ( .A1(n6541), .A2(n4459), .ZN(n4561) );
  OAI21_X1 U5262 ( .B1(n6875), .B2(n6873), .A(n6874), .ZN(n7045) );
  NOR2_X1 U5263 ( .A1(n6862), .A2(n6808), .ZN(n4567) );
  INV_X1 U5264 ( .A(n4569), .ZN(n4563) );
  NOR2_X1 U5265 ( .A1(n7046), .A2(n6863), .ZN(n4568) );
  NOR2_X1 U5266 ( .A1(n9174), .A2(n7448), .ZN(n4867) );
  NAND2_X1 U5267 ( .A1(n7517), .A2(n7518), .ZN(n7519) );
  NAND2_X1 U5268 ( .A1(n7519), .A2(n7520), .ZN(n8372) );
  OAI22_X1 U5269 ( .A1(n8505), .A2(n6257), .B1(n6328), .B2(n8779), .ZN(n7990)
         );
  NAND2_X1 U5270 ( .A1(n6165), .A2(n9031), .ZN(n6175) );
  INV_X1 U5271 ( .A(n6166), .ZN(n6165) );
  OR2_X1 U5272 ( .A1(n6155), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6166) );
  OR2_X1 U5273 ( .A1(n6073), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6084) );
  OR2_X1 U5274 ( .A1(n6051), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U5275 ( .A1(n7898), .A2(n7900), .ZN(n8014) );
  NAND2_X1 U5276 ( .A1(n4792), .A2(n4786), .ZN(n4784) );
  NAND2_X1 U5277 ( .A1(n7303), .A2(n4788), .ZN(n4782) );
  OR2_X1 U5278 ( .A1(n7490), .A2(n7442), .ZN(n7881) );
  OR2_X1 U5279 ( .A1(n6024), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6037) );
  AND4_X1 U5280 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n7623)
         );
  INV_X1 U5281 ( .A(n5991), .ZN(n5990) );
  INV_X1 U5282 ( .A(n8007), .ZN(n6286) );
  AND2_X1 U5283 ( .A1(n7223), .A2(n7884), .ZN(n8007) );
  AOI21_X1 U5284 ( .B1(n8514), .B2(n7961), .A(n7963), .ZN(n8505) );
  XNOR2_X1 U5285 ( .A(n8779), .B(n8517), .ZN(n8506) );
  AOI21_X1 U5286 ( .B1(n4746), .B2(n4745), .A(n4744), .ZN(n4743) );
  INV_X1 U5287 ( .A(n4750), .ZN(n4745) );
  INV_X1 U5288 ( .A(n7957), .ZN(n4744) );
  NAND2_X1 U5289 ( .A1(n4480), .A2(n5003), .ZN(n4806) );
  INV_X1 U5290 ( .A(n5002), .ZN(n4807) );
  NOR2_X1 U5291 ( .A1(n7951), .A2(n4751), .ZN(n4750) );
  INV_X1 U5292 ( .A(n7949), .ZN(n4751) );
  OR2_X1 U5293 ( .A1(n7951), .A2(n7950), .ZN(n4749) );
  AND2_X1 U5294 ( .A1(n7996), .A2(n7995), .ZN(n8553) );
  OR2_X1 U5295 ( .A1(n8815), .A2(n8560), .ZN(n6308) );
  NAND2_X1 U5296 ( .A1(n6303), .A2(n4777), .ZN(n4775) );
  OAI211_X1 U5297 ( .C1(n4774), .C2(n6303), .A(n4771), .B(n4769), .ZN(n4773)
         );
  NAND2_X1 U5298 ( .A1(n6133), .A2(n6132), .ZN(n8629) );
  AND4_X1 U5299 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n8647)
         );
  OR2_X1 U5300 ( .A1(n6731), .A2(n7973), .ZN(n8673) );
  AND2_X1 U5301 ( .A1(n7923), .A2(n7925), .ZN(n8645) );
  AOI21_X1 U5302 ( .B1(n4757), .B2(n4759), .A(n4756), .ZN(n4755) );
  INV_X1 U5303 ( .A(n4761), .ZN(n4757) );
  INV_X1 U5304 ( .A(n7916), .ZN(n4756) );
  INV_X1 U5305 ( .A(n4759), .ZN(n4758) );
  NOR2_X1 U5306 ( .A1(n4762), .A2(n7915), .ZN(n4761) );
  INV_X1 U5307 ( .A(n7911), .ZN(n4762) );
  INV_X1 U5308 ( .A(n8671), .ZN(n8687) );
  INV_X1 U5309 ( .A(n8673), .ZN(n8685) );
  NAND2_X1 U5310 ( .A1(n6317), .A2(n6316), .ZN(n8690) );
  AND2_X1 U5311 ( .A1(n6361), .A2(n6594), .ZN(n6577) );
  INV_X1 U5312 ( .A(n8764), .ZN(n8766) );
  NAND2_X1 U5313 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  INV_X1 U5314 ( .A(n8879), .ZN(n6342) );
  INV_X1 U5315 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6336) );
  INV_X1 U5316 ( .A(n5887), .ZN(n4763) );
  NOR2_X1 U5317 ( .A1(n4767), .A2(n5950), .ZN(n4764) );
  NAND2_X1 U5318 ( .A1(n6135), .A2(n5890), .ZN(n6136) );
  INV_X1 U5319 ( .A(n9914), .ZN(n8122) );
  OAI22_X1 U5320 ( .A1(n6785), .A2(n6776), .B1(n4426), .B2(n8056), .ZN(n6773)
         );
  OR2_X1 U5321 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  AND2_X1 U5322 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  OR2_X1 U5323 ( .A1(n7793), .A2(n9191), .ZN(n7796) );
  NAND2_X1 U5324 ( .A1(n4452), .A2(n4818), .ZN(n4816) );
  INV_X1 U5325 ( .A(n7791), .ZN(n9189) );
  NOR2_X1 U5326 ( .A1(n7311), .A2(n4543), .ZN(n7294) );
  AND2_X1 U5327 ( .A1(n7286), .A2(n7285), .ZN(n4543) );
  NAND3_X1 U5328 ( .A1(n4537), .A2(n7746), .A3(n7745), .ZN(n9365) );
  INV_X1 U5329 ( .A(n9367), .ZN(n7745) );
  AND2_X1 U5330 ( .A1(n6832), .A2(n6659), .ZN(n6842) );
  OAI21_X1 U5331 ( .B1(n5833), .B2(n5722), .A(n5723), .ZN(n5724) );
  INV_X1 U5332 ( .A(n8049), .ZN(n5407) );
  NAND2_X1 U5333 ( .A1(n10084), .A2(n10085), .ZN(n4649) );
  NAND2_X1 U5334 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5335 ( .A1(n10091), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5336 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  INV_X1 U5337 ( .A(n10097), .ZN(n4646) );
  NOR2_X1 U5338 ( .A1(n10041), .A2(n4643), .ZN(n10057) );
  NOR2_X1 U5339 ( .A1(n6613), .A2(n5497), .ZN(n4643) );
  NOR2_X1 U5340 ( .A1(n10057), .A2(n4524), .ZN(n10056) );
  AND2_X1 U5341 ( .A1(n8161), .A2(n5727), .ZN(n9532) );
  NAND2_X1 U5342 ( .A1(n9573), .A2(n8157), .ZN(n9560) );
  AND4_X1 U5343 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n9576)
         );
  NAND2_X1 U5344 ( .A1(n9594), .A2(n8155), .ZN(n9574) );
  AND2_X1 U5345 ( .A1(n5777), .A2(n5776), .ZN(n8151) );
  AND2_X1 U5346 ( .A1(n8149), .A2(n5857), .ZN(n4954) );
  AND4_X1 U5347 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n9664)
         );
  NAND2_X1 U5348 ( .A1(n9723), .A2(n9722), .ZN(n4950) );
  AND4_X1 U5349 ( .A1(n5592), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(n9712)
         );
  NOR2_X1 U5350 ( .A1(n9776), .A2(n9914), .ZN(n9762) );
  AOI21_X1 U5351 ( .B1(n9798), .B2(n9797), .A(n4997), .ZN(n9775) );
  NAND2_X1 U5352 ( .A1(n5843), .A2(n5742), .ZN(n7578) );
  NOR2_X1 U5353 ( .A1(n7478), .A2(n7483), .ZN(n7477) );
  XNOR2_X1 U5354 ( .A(n9391), .B(n7275), .ZN(n7268) );
  INV_X1 U5355 ( .A(n9393), .ZN(n7102) );
  NAND2_X1 U5356 ( .A1(n5470), .A2(n6964), .ZN(n6836) );
  AND2_X1 U5357 ( .A1(n5377), .A2(n5376), .ZN(n5479) );
  OR2_X1 U5358 ( .A1(n5490), .A2(n5457), .ZN(n5458) );
  AND2_X1 U5359 ( .A1(n5413), .A2(n10007), .ZN(n6670) );
  NOR2_X1 U5360 ( .A1(n9532), .A2(n4687), .ZN(n4686) );
  INV_X1 U5361 ( .A(n8145), .ZN(n4687) );
  OAI21_X1 U5362 ( .B1(n9572), .B2(n8141), .A(n8140), .ZN(n9556) );
  AND2_X1 U5363 ( .A1(n9610), .A2(n8130), .ZN(n9590) );
  NOR2_X1 U5364 ( .A1(n9967), .A2(n9631), .ZN(n9591) );
  AOI21_X1 U5365 ( .B1(n9674), .B2(n8127), .A(n8126), .ZN(n9660) );
  AND2_X1 U5366 ( .A1(n4512), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5367 ( .A1(n4678), .A2(n4677), .ZN(n4680) );
  INV_X1 U5368 ( .A(n4680), .ZN(n9719) );
  INV_X1 U5369 ( .A(n10234), .ZN(n10275) );
  INV_X1 U5370 ( .A(n9929), .ZN(n10273) );
  INV_X1 U5371 ( .A(n6403), .ZN(n4549) );
  AND2_X1 U5372 ( .A1(n10235), .A2(n5880), .ZN(n10280) );
  AND2_X1 U5373 ( .A1(n7335), .A2(n7538), .ZN(n10235) );
  INV_X1 U5374 ( .A(n9927), .ZN(n10283) );
  XNOR2_X1 U5375 ( .A(n5346), .B(n5345), .ZN(n8114) );
  NAND2_X1 U5376 ( .A1(n4898), .A2(n5122), .ZN(n5331) );
  XNOR2_X1 U5377 ( .A(n5327), .B(n5328), .ZN(n8875) );
  XNOR2_X1 U5378 ( .A(n5319), .B(n5320), .ZN(n7647) );
  NAND2_X1 U5379 ( .A1(n4892), .A2(n5107), .ZN(n5319) );
  NAND2_X1 U5380 ( .A1(n5316), .A2(n5315), .ZN(n4892) );
  INV_X1 U5381 ( .A(n4624), .ZN(n4623) );
  OR2_X1 U5382 ( .A1(n5288), .A2(n4513), .ZN(n4621) );
  OAI21_X1 U5383 ( .B1(n4625), .B2(n4627), .A(n5096), .ZN(n4624) );
  AND2_X1 U5384 ( .A1(n5101), .A2(n5100), .ZN(n5311) );
  NAND2_X1 U5385 ( .A1(n4622), .A2(n4905), .ZN(n5308) );
  NAND2_X1 U5386 ( .A1(n4629), .A2(n4627), .ZN(n4622) );
  NAND2_X1 U5387 ( .A1(n4903), .A2(n4902), .ZN(n5304) );
  NAND2_X1 U5388 ( .A1(n5090), .A2(n5296), .ZN(n4902) );
  NAND2_X1 U5389 ( .A1(n4825), .A2(n4938), .ZN(n5284) );
  AND2_X1 U5390 ( .A1(n4921), .A2(n4928), .ZN(n5283) );
  INV_X1 U5391 ( .A(n4927), .ZN(n4922) );
  INV_X1 U5392 ( .A(n4636), .ZN(n5262) );
  NAND2_X1 U5393 ( .A1(n5245), .A2(n5069), .ZN(n5252) );
  NAND2_X1 U5394 ( .A1(n5243), .A2(n5242), .ZN(n5245) );
  NAND2_X1 U5395 ( .A1(n5064), .A2(n5063), .ZN(n5235) );
  NAND2_X1 U5396 ( .A1(n5218), .A2(n4919), .ZN(n4916) );
  AND2_X1 U5397 ( .A1(n5059), .A2(n5058), .ZN(n5214) );
  NAND3_X1 U5398 ( .A1(n4988), .A2(n4987), .A3(n5007), .ZN(n8207) );
  INV_X1 U5399 ( .A(n8206), .ZN(n4987) );
  OAI21_X1 U5400 ( .B1(n8072), .B2(n8071), .A(n8070), .ZN(n8215) );
  AOI21_X1 U5401 ( .B1(n8322), .B2(n8323), .A(n4503), .ZN(n8232) );
  NAND2_X1 U5402 ( .A1(n8232), .A2(n8231), .ZN(n8230) );
  AND2_X1 U5403 ( .A1(n6234), .A2(n6233), .ZN(n8258) );
  NAND2_X1 U5404 ( .A1(n6123), .A2(n6122), .ZN(n8631) );
  AND2_X1 U5405 ( .A1(n6211), .A2(n6210), .ZN(n8307) );
  INV_X1 U5406 ( .A(n8526), .ZN(n8336) );
  AOI21_X1 U5407 ( .B1(n4735), .B2(n4525), .A(n4734), .ZN(n8039) );
  INV_X1 U5408 ( .A(n8258), .ZN(n8535) );
  NAND2_X1 U5409 ( .A1(n6222), .A2(n6221), .ZN(n8545) );
  INV_X1 U5410 ( .A(n8307), .ZN(n8570) );
  XNOR2_X1 U5411 ( .A(n6858), .B(n6828), .ZN(n6860) );
  NAND2_X1 U5412 ( .A1(n6059), .A2(n6058), .ZN(n7906) );
  NAND2_X1 U5413 ( .A1(n7803), .A2(n7802), .ZN(n9255) );
  NAND2_X1 U5414 ( .A1(n5275), .A2(n5274), .ZN(n9725) );
  INV_X1 U5415 ( .A(n9604), .ZN(n9838) );
  NAND2_X1 U5416 ( .A1(n7789), .A2(n7788), .ZN(n9324) );
  OR2_X1 U5417 ( .A1(n9636), .A2(n6776), .ZN(n7789) );
  INV_X1 U5418 ( .A(n9892), .ZN(n9699) );
  NAND2_X1 U5419 ( .A1(n6681), .A2(n10205), .ZN(n9376) );
  AND2_X1 U5420 ( .A1(n6665), .A2(n6388), .ZN(n10005) );
  NAND2_X1 U5421 ( .A1(n9504), .A2(n4654), .ZN(n4653) );
  INV_X1 U5422 ( .A(n4655), .ZN(n4654) );
  OAI21_X1 U5423 ( .B1(n9505), .B2(n10152), .A(n10121), .ZN(n4655) );
  NOR2_X1 U5424 ( .A1(n5368), .A2(n9778), .ZN(n9510) );
  INV_X1 U5425 ( .A(n9967), .ZN(n9622) );
  AND4_X1 U5426 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n9911)
         );
  NAND2_X1 U5427 ( .A1(n5241), .A2(n5240), .ZN(n9804) );
  NAND2_X1 U5428 ( .A1(n5222), .A2(n5221), .ZN(n9200) );
  INV_X1 U5429 ( .A(n7483), .ZN(n10199) );
  NAND2_X1 U5430 ( .A1(n6659), .A2(n4811), .ZN(n7017) );
  AND2_X1 U5431 ( .A1(n6973), .A2(n7281), .ZN(n4811) );
  INV_X1 U5432 ( .A(n9833), .ZN(n9935) );
  INV_X1 U5433 ( .A(n8059), .ZN(n6936) );
  XNOR2_X1 U5434 ( .A(n5350), .B(n5349), .ZN(n10014) );
  OAI21_X1 U5435 ( .B1(n5346), .B2(n5345), .A(n5344), .ZN(n5350) );
  NAND2_X1 U5436 ( .A1(n4451), .A2(n4704), .ZN(n4703) );
  INV_X1 U5437 ( .A(n5786), .ZN(n4704) );
  AND2_X1 U5438 ( .A1(n4706), .A2(n5534), .ZN(n4705) );
  NAND2_X1 U5439 ( .A1(n7455), .A2(n5720), .ZN(n4706) );
  OR2_X1 U5440 ( .A1(n5739), .A2(n5720), .ZN(n4707) );
  INV_X1 U5441 ( .A(n7860), .ZN(n4834) );
  INV_X1 U5442 ( .A(n4835), .ZN(n4838) );
  OR2_X1 U5443 ( .A1(n7861), .A2(n7860), .ZN(n4839) );
  AOI21_X1 U5444 ( .B1(n5572), .B2(n5844), .A(n4701), .ZN(n4700) );
  NAND2_X1 U5445 ( .A1(n9790), .A2(n5740), .ZN(n4701) );
  NOR2_X1 U5446 ( .A1(n5846), .A2(n5720), .ZN(n4699) );
  NAND2_X1 U5447 ( .A1(n4528), .A2(n4527), .ZN(n7879) );
  NAND2_X1 U5448 ( .A1(n7876), .A2(n4530), .ZN(n4527) );
  NAND2_X1 U5449 ( .A1(n4531), .A2(n4529), .ZN(n4528) );
  INV_X1 U5450 ( .A(n5606), .ZN(n4702) );
  NAND2_X1 U5451 ( .A1(n4861), .A2(n4860), .ZN(n4859) );
  NOR2_X1 U5452 ( .A1(n7913), .A2(n8675), .ZN(n4860) );
  NAND2_X1 U5453 ( .A1(n5639), .A2(n5814), .ZN(n5632) );
  NAND2_X1 U5454 ( .A1(n8601), .A2(n7924), .ZN(n4532) );
  NAND2_X1 U5455 ( .A1(n4725), .A2(n5648), .ZN(n4724) );
  AND2_X1 U5456 ( .A1(n4696), .A2(n4695), .ZN(n5802) );
  AND2_X1 U5457 ( .A1(n9771), .A2(n9790), .ZN(n4695) );
  NAND2_X1 U5458 ( .A1(n5568), .A2(n4697), .ZN(n4696) );
  INV_X1 U5459 ( .A(n5740), .ZN(n4697) );
  INV_X1 U5460 ( .A(n7953), .ZN(n4850) );
  INV_X1 U5461 ( .A(n4848), .ZN(n4847) );
  AOI21_X1 U5462 ( .B1(n4851), .B2(n7947), .A(n4476), .ZN(n4848) );
  OR2_X1 U5463 ( .A1(n9591), .A2(n9590), .ZN(n8132) );
  OAI22_X1 U5464 ( .A1(n4470), .A2(n6845), .B1(n4715), .B2(n5784), .ZN(n4710)
         );
  OR2_X1 U5465 ( .A1(n5693), .A2(n5692), .ZN(n4716) );
  AND2_X1 U5466 ( .A1(n5766), .A2(n5767), .ZN(n5826) );
  INV_X1 U5467 ( .A(n4894), .ZN(n4893) );
  OAI21_X1 U5468 ( .B1(n5315), .B2(n4895), .A(n5320), .ZN(n4894) );
  INV_X1 U5469 ( .A(n5107), .ZN(n4895) );
  INV_X1 U5470 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4828) );
  NOR2_X1 U5471 ( .A1(n4927), .A2(n5084), .ZN(n4926) );
  NOR2_X1 U5472 ( .A1(n5253), .A2(SI_14_), .ZN(n4933) );
  NAND2_X1 U5473 ( .A1(n5245), .A2(n4934), .ZN(n4932) );
  AND2_X1 U5474 ( .A1(n5069), .A2(n4935), .ZN(n4934) );
  NAND2_X1 U5475 ( .A1(n5253), .A2(SI_14_), .ZN(n4935) );
  INV_X1 U5476 ( .A(n5208), .ZN(n4617) );
  NAND2_X1 U5477 ( .A1(n8035), .A2(n4855), .ZN(n8036) );
  NOR2_X1 U5478 ( .A1(n7994), .A2(n7962), .ZN(n4633) );
  NAND2_X1 U5479 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5480 ( .A1(n4879), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4878) );
  INV_X1 U5481 ( .A(n6715), .ZN(n4872) );
  AOI21_X1 U5482 ( .B1(n6716), .B2(n6715), .A(n4876), .ZN(n4871) );
  NOR2_X1 U5483 ( .A1(n6821), .A2(n6820), .ZN(n4876) );
  NAND2_X1 U5484 ( .A1(n7364), .A2(n7365), .ZN(n7515) );
  NAND2_X1 U5485 ( .A1(n8424), .A2(n4523), .ZN(n8461) );
  INV_X1 U5486 ( .A(n4786), .ZN(n4781) );
  NAND2_X1 U5487 ( .A1(n7222), .A2(n7877), .ZN(n4732) );
  OAI21_X1 U5488 ( .B1(n6344), .B2(P2_D_REG_0__SCAN_IN), .A(n6451), .ZN(n6737)
         );
  NAND2_X1 U5489 ( .A1(n4982), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5922) );
  OR2_X1 U5490 ( .A1(n6344), .A2(n6357), .ZN(n6372) );
  OR2_X1 U5491 ( .A1(n7963), .A2(n7964), .ZN(n7994) );
  INV_X1 U5492 ( .A(n7960), .ZN(n4742) );
  NOR2_X1 U5493 ( .A1(n4447), .A2(n8533), .ZN(n4804) );
  NAND2_X1 U5494 ( .A1(n6212), .A2(n7996), .ZN(n7955) );
  NAND2_X1 U5495 ( .A1(n4468), .A2(n4772), .ZN(n4771) );
  NOR2_X1 U5496 ( .A1(n4774), .A2(n4776), .ZN(n4772) );
  INV_X1 U5497 ( .A(n6298), .ZN(n4776) );
  NAND2_X1 U5498 ( .A1(n4770), .A2(n6304), .ZN(n4769) );
  INV_X1 U5499 ( .A(n4774), .ZN(n4770) );
  INV_X1 U5500 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4768) );
  NOR2_X1 U5501 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4858) );
  INV_X1 U5502 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5503 ( .A1(n4823), .A2(n7826), .ZN(n7696) );
  INV_X1 U5504 ( .A(n6924), .ZN(n4823) );
  INV_X1 U5505 ( .A(n4554), .ZN(n4553) );
  AOI21_X1 U5506 ( .B1(n4552), .B2(n4554), .A(n4504), .ZN(n4551) );
  INV_X1 U5507 ( .A(n4555), .ZN(n4552) );
  NAND2_X1 U5508 ( .A1(n9263), .A2(n4555), .ZN(n4550) );
  OR2_X1 U5509 ( .A1(n7736), .A2(n7738), .ZN(n4538) );
  AND2_X1 U5510 ( .A1(n7736), .A2(n7738), .ZN(n4540) );
  OAI211_X1 U5511 ( .C1(n4716), .C2(n4712), .A(n4711), .B(n4709), .ZN(n5713)
         );
  OAI21_X1 U5512 ( .B1(n4714), .B2(n4710), .A(n4713), .ZN(n4709) );
  NAND2_X1 U5513 ( .A1(n4713), .A2(n5720), .ZN(n4712) );
  OR2_X1 U5514 ( .A1(n5693), .A2(n4471), .ZN(n4711) );
  NOR2_X1 U5515 ( .A1(n5713), .A2(n9941), .ZN(n5716) );
  NOR4_X1 U5516 ( .A1(n5863), .A2(n5869), .A3(n5762), .A4(n5761), .ZN(n5871)
         );
  INV_X1 U5517 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4937) );
  OR2_X1 U5518 ( .A1(n9622), .A2(n9631), .ZN(n5647) );
  NAND2_X1 U5519 ( .A1(n9676), .A2(n9675), .ZN(n4955) );
  INV_X1 U5520 ( .A(n5613), .ZN(n5619) );
  NAND2_X1 U5521 ( .A1(n4936), .A2(n4463), .ZN(n5839) );
  NAND2_X1 U5522 ( .A1(n7267), .A2(n5790), .ZN(n4936) );
  OR2_X1 U5523 ( .A1(n9563), .A2(n9576), .ZN(n5729) );
  NAND2_X1 U5524 ( .A1(n4449), .A2(n4666), .ZN(n4665) );
  INV_X1 U5525 ( .A(n8129), .ZN(n4666) );
  INV_X1 U5526 ( .A(n4449), .ZN(n4667) );
  OR2_X1 U5527 ( .A1(n9619), .A2(n9838), .ZN(n9598) );
  AND2_X1 U5528 ( .A1(n9625), .A2(n8133), .ZN(n9589) );
  OR2_X1 U5529 ( .A1(n9650), .A2(n9664), .ZN(n5775) );
  NAND2_X1 U5530 ( .A1(n9722), .A2(n4443), .ZN(n4676) );
  NOR2_X1 U5531 ( .A1(n6974), .A2(n6936), .ZN(n6986) );
  NAND2_X1 U5532 ( .A1(n4897), .A2(n4896), .ZN(n5336) );
  AOI21_X1 U5533 ( .B1(n4899), .B2(n4901), .A(n4522), .ZN(n4896) );
  AND2_X1 U5534 ( .A1(n5116), .A2(n5115), .ZN(n5323) );
  AOI21_X1 U5535 ( .B1(n4907), .B2(n4432), .A(n4505), .ZN(n4905) );
  NOR2_X1 U5536 ( .A1(n4906), .A2(n4628), .ZN(n4627) );
  INV_X1 U5537 ( .A(n5089), .ZN(n4628) );
  INV_X1 U5538 ( .A(n4907), .ZN(n4906) );
  OR2_X1 U5539 ( .A1(n5090), .A2(n5296), .ZN(n4904) );
  NAND2_X1 U5540 ( .A1(n4506), .A2(n5080), .ZN(n4928) );
  INV_X1 U5541 ( .A(n5075), .ZN(n4929) );
  NAND2_X1 U5542 ( .A1(n4495), .A2(n5080), .ZN(n4927) );
  NAND2_X1 U5543 ( .A1(n5065), .A2(SI_13_), .ZN(n5069) );
  INV_X1 U5544 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5010) );
  XNOR2_X1 U5545 ( .A(n4421), .B(n6746), .ZN(n6747) );
  NAND2_X1 U5546 ( .A1(n4978), .A2(n6762), .ZN(n6914) );
  AND2_X1 U5547 ( .A1(n6690), .A2(n6602), .ZN(n7845) );
  NAND2_X1 U5548 ( .A1(n8230), .A2(n4980), .ZN(n8295) );
  OR2_X1 U5549 ( .A1(n8081), .A2(n8591), .ZN(n5000) );
  OR2_X1 U5550 ( .A1(n6743), .A2(n8367), .ZN(n6744) );
  NAND2_X1 U5551 ( .A1(n4975), .A2(n4462), .ZN(n4974) );
  NAND2_X1 U5552 ( .A1(n7006), .A2(n4976), .ZN(n4975) );
  INV_X1 U5553 ( .A(n6913), .ZN(n4976) );
  AND2_X1 U5554 ( .A1(n6762), .A2(n7006), .ZN(n4977) );
  INV_X1 U5555 ( .A(n8074), .ZN(n4970) );
  NAND2_X1 U5556 ( .A1(n4972), .A2(n4973), .ZN(n4971) );
  INV_X1 U5557 ( .A(n8215), .ZN(n4972) );
  NAND2_X1 U5558 ( .A1(n4982), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4984) );
  OAI21_X1 U5559 ( .B1(n6572), .B2(n6323), .A(n5905), .ZN(n5906) );
  NAND2_X1 U5560 ( .A1(n4877), .A2(n6525), .ZN(n6527) );
  INV_X1 U5561 ( .A(n4878), .ZN(n4877) );
  NOR2_X1 U5562 ( .A1(n6519), .A2(n6520), .ZN(n6541) );
  NAND2_X1 U5563 ( .A1(n6546), .A2(n4875), .ZN(n6547) );
  NAND2_X1 U5564 ( .A1(n4870), .A2(n6715), .ZN(n6819) );
  NAND2_X1 U5565 ( .A1(n4873), .A2(n4875), .ZN(n4870) );
  AND2_X1 U5566 ( .A1(n4869), .A2(n4868), .ZN(n7173) );
  NAND2_X1 U5567 ( .A1(n7250), .A2(n7251), .ZN(n7253) );
  NAND2_X1 U5568 ( .A1(n7253), .A2(n7252), .ZN(n7364) );
  OR2_X1 U5569 ( .A1(n7239), .A2(n7238), .ZN(n7351) );
  XNOR2_X1 U5570 ( .A(n7515), .B(n7509), .ZN(n7366) );
  AND2_X1 U5571 ( .A1(n7351), .A2(n7350), .ZN(n7508) );
  NAND2_X1 U5572 ( .A1(n8372), .A2(n8373), .ZN(n8399) );
  NOR2_X1 U5573 ( .A1(n8421), .A2(n4882), .ZN(n8453) );
  AND2_X1 U5574 ( .A1(n8422), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4882) );
  XNOR2_X1 U5575 ( .A(n8461), .B(n8452), .ZN(n8426) );
  NAND2_X1 U5576 ( .A1(n8426), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8465) );
  AND2_X1 U5577 ( .A1(n7684), .A2(n6326), .ZN(n7976) );
  NAND2_X1 U5578 ( .A1(n6227), .A2(n6226), .ZN(n6238) );
  INV_X1 U5579 ( .A(n6228), .ZN(n6227) );
  NAND2_X1 U5580 ( .A1(n6195), .A2(n6194), .ZN(n6216) );
  NAND2_X1 U5581 ( .A1(n6182), .A2(n6181), .ZN(n6204) );
  INV_X1 U5582 ( .A(n6183), .ZN(n6182) );
  OR2_X1 U5583 ( .A1(n6175), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6183) );
  AND2_X1 U5584 ( .A1(n7943), .A2(n7933), .ZN(n8595) );
  NAND2_X1 U5585 ( .A1(n6141), .A2(n6140), .ZN(n6155) );
  INV_X1 U5586 ( .A(n6142), .ZN(n6141) );
  OR2_X1 U5587 ( .A1(n6125), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U5588 ( .A1(n6113), .A2(n6112), .ZN(n6125) );
  INV_X1 U5589 ( .A(n6114), .ZN(n6113) );
  NAND2_X1 U5590 ( .A1(n6095), .A2(n8340), .ZN(n6114) );
  INV_X1 U5591 ( .A(n6096), .ZN(n6095) );
  NAND2_X1 U5592 ( .A1(n6062), .A2(n6061), .ZN(n6073) );
  NAND2_X1 U5593 ( .A1(n7499), .A2(n7500), .ZN(n4733) );
  INV_X1 U5594 ( .A(n6037), .ZN(n6036) );
  NAND2_X1 U5595 ( .A1(n4790), .A2(n6290), .ZN(n7441) );
  NAND2_X1 U5596 ( .A1(n4791), .A2(n4793), .ZN(n4790) );
  INV_X1 U5597 ( .A(n7303), .ZN(n4791) );
  AND4_X1 U5598 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n7403)
         );
  NAND2_X1 U5599 ( .A1(n6012), .A2(n6011), .ZN(n6024) );
  INV_X1 U5600 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6011) );
  INV_X1 U5601 ( .A(n6013), .ZN(n6012) );
  AND4_X1 U5602 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n7336)
         );
  NOR2_X1 U5603 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n5969) );
  AND4_X1 U5604 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n7060)
         );
  NOR2_X1 U5605 ( .A1(n5927), .A2(n5928), .ZN(n4730) );
  NAND2_X1 U5606 ( .A1(n8001), .A2(n7846), .ZN(n6687) );
  INV_X1 U5607 ( .A(n7994), .ZN(n8515) );
  AOI21_X1 U5608 ( .B1(n8567), .B2(n7949), .A(n6190), .ZN(n8557) );
  AND2_X1 U5609 ( .A1(n7950), .A2(n7949), .ZN(n8568) );
  NAND2_X1 U5610 ( .A1(n7924), .A2(n7929), .ZN(n8635) );
  NAND2_X1 U5611 ( .A1(n6299), .A2(n6298), .ZN(n8646) );
  OR2_X1 U5612 ( .A1(n8646), .A2(n8645), .ZN(n8649) );
  NAND2_X1 U5613 ( .A1(n4857), .A2(n4855), .ZN(n8764) );
  AND2_X1 U5614 ( .A1(n6587), .A2(n6456), .ZN(n6594) );
  XNOR2_X1 U5615 ( .A(n6278), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8034) );
  AND2_X1 U5616 ( .A1(n4428), .A2(n4482), .ZN(n4596) );
  NAND2_X1 U5617 ( .A1(n6044), .A2(n6046), .ZN(n6070) );
  OR2_X1 U5618 ( .A1(n7737), .A2(n7736), .ZN(n4824) );
  AND2_X1 U5619 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5502) );
  OR2_X1 U5620 ( .A1(n5521), .A2(n5520), .ZN(n5537) );
  INV_X1 U5621 ( .A(n4542), .ZN(n4541) );
  OAI21_X1 U5622 ( .B1(n4821), .B2(n7294), .A(n7690), .ZN(n4542) );
  NAND2_X1 U5623 ( .A1(n4822), .A2(n7312), .ZN(n4821) );
  OR2_X1 U5624 ( .A1(n5573), .A2(n9317), .ZN(n5580) );
  NOR2_X1 U5625 ( .A1(n5451), .A2(n9240), .ZN(n5444) );
  INV_X1 U5626 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5509) );
  AND2_X1 U5627 ( .A1(n5593), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5595) );
  INV_X1 U5628 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U5629 ( .A1(n6633), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5630 ( .A1(n10056), .A2(n6614), .ZN(n10065) );
  NOR2_X1 U5631 ( .A1(n10023), .A2(n4517), .ZN(n10112) );
  NOR2_X1 U5632 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  NOR2_X1 U5633 ( .A1(n10140), .A2(n4650), .ZN(n9466) );
  AND2_X1 U5634 ( .A1(n10148), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5635 ( .A1(n9598), .A2(n4607), .ZN(n9542) );
  NAND2_X1 U5636 ( .A1(n9542), .A2(n8144), .ZN(n9543) );
  NAND2_X1 U5637 ( .A1(n5647), .A2(n8154), .ZN(n9613) );
  NOR3_X1 U5638 ( .A1(n9665), .A2(n9650), .A3(n9867), .ZN(n5001) );
  NOR3_X1 U5639 ( .A1(n9665), .A2(n9650), .A3(n4601), .ZN(n9634) );
  AND2_X1 U5640 ( .A1(n5310), .A2(n5309), .ZN(n9636) );
  NAND2_X1 U5641 ( .A1(n4955), .A2(n5857), .ZN(n8148) );
  AND2_X1 U5642 ( .A1(n9762), .A2(n4514), .ZN(n9677) );
  NAND2_X1 U5643 ( .A1(n9762), .A2(n9905), .ZN(n9742) );
  NAND2_X1 U5644 ( .A1(n7589), .A2(n4434), .ZN(n9776) );
  NAND2_X1 U5645 ( .A1(n7589), .A2(n4605), .ZN(n9801) );
  AND2_X1 U5646 ( .A1(n5735), .A2(n5849), .ZN(n9774) );
  OR2_X1 U5647 ( .A1(n5561), .A2(n5560), .ZN(n5573) );
  NAND2_X1 U5648 ( .A1(n4670), .A2(n4669), .ZN(n9798) );
  AOI21_X1 U5649 ( .B1(n4671), .B2(n4673), .A(n4435), .ZN(n4669) );
  NAND2_X1 U5650 ( .A1(n7584), .A2(n7583), .ZN(n7609) );
  NOR2_X1 U5651 ( .A1(n5009), .A2(n4416), .ZN(n7588) );
  AOI21_X1 U5652 ( .B1(n7479), .B2(n4662), .A(n4472), .ZN(n4661) );
  INV_X1 U5653 ( .A(n7382), .ZN(n4662) );
  NAND2_X1 U5654 ( .A1(n5174), .A2(n4598), .ZN(n7478) );
  NOR2_X1 U5655 ( .A1(n10210), .A2(n7381), .ZN(n4598) );
  INV_X1 U5656 ( .A(n7270), .ZN(n5174) );
  NAND2_X1 U5657 ( .A1(n5174), .A2(n7275), .ZN(n7271) );
  NAND2_X1 U5658 ( .A1(n5136), .A2(n5135), .ZN(n8188) );
  INV_X1 U5659 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U5660 ( .A1(n9560), .A2(n8158), .ZN(n9547) );
  NAND2_X1 U5661 ( .A1(n5729), .A2(n8158), .ZN(n9557) );
  AND2_X1 U5662 ( .A1(n8156), .A2(n5730), .ZN(n9575) );
  AND2_X1 U5663 ( .A1(n5775), .A2(n5776), .ZN(n9648) );
  AND2_X1 U5664 ( .A1(n5816), .A2(n5857), .ZN(n9675) );
  AND4_X1 U5665 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n9912)
         );
  AND4_X1 U5666 ( .A1(n5585), .A2(n5584), .A3(n5583), .A4(n5582), .ZN(n10276)
         );
  AND2_X1 U5667 ( .A1(n4943), .A2(n4940), .ZN(n5468) );
  NAND2_X1 U5668 ( .A1(n5167), .A2(n4941), .ZN(n4940) );
  NAND2_X1 U5669 ( .A1(n4478), .A2(n4942), .ZN(n4941) );
  NOR2_X1 U5670 ( .A1(n5412), .A2(n6952), .ZN(n5420) );
  AND2_X1 U5671 ( .A1(n5381), .A2(n6842), .ZN(n10234) );
  NAND2_X1 U5672 ( .A1(n5395), .A2(n5394), .ZN(n10004) );
  AND2_X1 U5673 ( .A1(n4690), .A2(n5131), .ZN(n4689) );
  AND2_X1 U5674 ( .A1(n4958), .A2(n4691), .ZN(n4690) );
  NOR2_X1 U5675 ( .A1(n5132), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4957) );
  INV_X1 U5676 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5385) );
  INV_X1 U5677 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U5678 ( .A1(n4930), .A2(n5075), .ZN(n5277) );
  NAND2_X1 U5679 ( .A1(n4612), .A2(n4609), .ZN(n5243) );
  NOR2_X1 U5680 ( .A1(n4465), .A2(n4610), .ZN(n4609) );
  NOR2_X1 U5681 ( .A1(n4618), .A2(n4611), .ZN(n4610) );
  AND2_X1 U5682 ( .A1(n5232), .A2(n5239), .ZN(n6644) );
  NAND2_X1 U5683 ( .A1(n5218), .A2(n5059), .ZN(n5224) );
  NAND2_X1 U5684 ( .A1(n4717), .A2(n4720), .ZN(n5191) );
  AOI21_X1 U5685 ( .B1(n5185), .B2(n4722), .A(n4721), .ZN(n4720) );
  INV_X1 U5686 ( .A(n5044), .ZN(n4721) );
  AND2_X1 U5687 ( .A1(n5048), .A2(n5047), .ZN(n5190) );
  INV_X1 U5688 ( .A(n5025), .ZN(n5027) );
  NAND2_X1 U5689 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  NAND2_X1 U5690 ( .A1(n4988), .A2(n5007), .ZN(n8205) );
  AND3_X1 U5691 ( .A1(n6170), .A2(n6169), .A3(n6168), .ZN(n8579) );
  NAND2_X1 U5692 ( .A1(n6174), .A2(n6173), .ZN(n8251) );
  NAND2_X1 U5693 ( .A1(n6914), .A2(n6913), .ZN(n7007) );
  NAND2_X1 U5694 ( .A1(n4581), .A2(n4585), .ZN(n8275) );
  NAND2_X1 U5695 ( .A1(n8262), .A2(n4586), .ZN(n4581) );
  NAND2_X1 U5696 ( .A1(n6164), .A2(n6163), .ZN(n8596) );
  AND2_X1 U5697 ( .A1(n4962), .A2(n4966), .ZN(n4961) );
  AOI21_X1 U5698 ( .B1(n4577), .B2(n4579), .A(n4479), .ZN(n4576) );
  NAND2_X1 U5699 ( .A1(n4992), .A2(n8087), .ZN(n8304) );
  OAI21_X1 U5700 ( .B1(n8230), .B2(n4579), .A(n4577), .ZN(n4992) );
  NOR2_X1 U5701 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  INV_X1 U5702 ( .A(n8335), .ZN(n8344) );
  INV_X1 U5703 ( .A(n8342), .ZN(n8331) );
  NAND2_X1 U5704 ( .A1(n4585), .A2(n4587), .ZN(n4580) );
  INV_X1 U5705 ( .A(n4583), .ZN(n4582) );
  NAND2_X1 U5706 ( .A1(n6599), .A2(n6598), .ZN(n8332) );
  NAND2_X1 U5707 ( .A1(n4593), .A2(n4592), .ZN(n7149) );
  AND2_X1 U5708 ( .A1(n4593), .A2(n4594), .ZN(n7009) );
  INV_X1 U5709 ( .A(n4974), .ZN(n4594) );
  AND2_X1 U5710 ( .A1(n4971), .A2(n4445), .ZN(n8347) );
  NAND2_X1 U5711 ( .A1(n4971), .A2(n8074), .ZN(n8349) );
  AND2_X1 U5712 ( .A1(n6581), .A2(n6580), .ZN(n8348) );
  NAND2_X1 U5713 ( .A1(n6574), .A2(n8683), .ZN(n8353) );
  NAND2_X1 U5714 ( .A1(n6244), .A2(n6243), .ZN(n8526) );
  AND4_X1 U5715 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n7442)
         );
  INV_X1 U5716 ( .A(n7403), .ZN(n8361) );
  OR2_X1 U5717 ( .A1(n7679), .A2(n5932), .ZN(n5933) );
  OR2_X1 U5718 ( .A1(n6323), .A2(n6462), .ZN(n5934) );
  NAND2_X1 U5719 ( .A1(n4879), .A2(n6525), .ZN(n6498) );
  XNOR2_X1 U5720 ( .A(n4561), .B(n6554), .ZN(n6711) );
  OAI22_X1 U5721 ( .A1(n6711), .A2(n6710), .B1(n6709), .B2(n4560), .ZN(n6712)
         );
  INV_X1 U5722 ( .A(n4561), .ZN(n4560) );
  NAND2_X1 U5723 ( .A1(n4564), .A2(n4562), .ZN(n7031) );
  NAND2_X1 U5724 ( .A1(n4563), .A2(n4566), .ZN(n4562) );
  INV_X1 U5725 ( .A(n6862), .ZN(n4566) );
  AND2_X1 U5726 ( .A1(n4565), .A2(n4569), .ZN(n6861) );
  NAND2_X1 U5727 ( .A1(n6860), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4565) );
  XNOR2_X1 U5728 ( .A(n4866), .B(n7249), .ZN(n7193) );
  NOR2_X1 U5729 ( .A1(n7503), .A2(n7193), .ZN(n7234) );
  XNOR2_X1 U5730 ( .A(n7509), .B(n7508), .ZN(n7352) );
  XNOR2_X1 U5731 ( .A(n8399), .B(n8393), .ZN(n8374) );
  INV_X1 U5732 ( .A(n8457), .ZN(n8451) );
  AOI21_X1 U5733 ( .B1(n8465), .B2(n8463), .A(n8464), .ZN(n8479) );
  AND2_X1 U5734 ( .A1(n6438), .A2(n8489), .ZN(n8499) );
  NAND2_X1 U5735 ( .A1(n6259), .A2(n6258), .ZN(n7675) );
  NOR2_X1 U5736 ( .A1(n8623), .A2(n4739), .ZN(n4738) );
  INV_X1 U5737 ( .A(n7929), .ZN(n4739) );
  NAND2_X1 U5738 ( .A1(n8629), .A2(n7929), .ZN(n8624) );
  NAND2_X1 U5739 ( .A1(n6138), .A2(n6137), .ZN(n8737) );
  NAND2_X1 U5740 ( .A1(n4782), .A2(n4785), .ZN(n7501) );
  INV_X1 U5741 ( .A(n4784), .ZN(n4785) );
  NAND2_X1 U5742 ( .A1(n4810), .A2(n6285), .ZN(n7398) );
  NAND2_X1 U5743 ( .A1(n6565), .A2(n6594), .ZN(n8683) );
  OR2_X1 U5744 ( .A1(n5952), .A2(n5024), .ZN(n4993) );
  INV_X1 U5745 ( .A(n4995), .ZN(n4994) );
  NAND2_X1 U5747 ( .A1(n7970), .A2(n7969), .ZN(n8703) );
  INV_X1 U5748 ( .A(n8772), .ZN(n7564) );
  NAND2_X1 U5749 ( .A1(n6247), .A2(n6246), .ZN(n8779) );
  NAND2_X1 U5750 ( .A1(n6237), .A2(n6236), .ZN(n8785) );
  NAND2_X1 U5751 ( .A1(n6225), .A2(n6224), .ZN(n8791) );
  OAI21_X1 U5752 ( .B1(n8567), .B2(n4747), .A(n4743), .ZN(n8523) );
  NAND2_X1 U5753 ( .A1(n6215), .A2(n6214), .ZN(n8797) );
  NAND2_X1 U5754 ( .A1(n4801), .A2(n4806), .ZN(n8534) );
  NAND2_X1 U5755 ( .A1(n4809), .A2(n4447), .ZN(n4801) );
  NAND2_X1 U5756 ( .A1(n4748), .A2(n4429), .ZN(n8532) );
  NAND2_X1 U5757 ( .A1(n8567), .A2(n4750), .ZN(n4748) );
  NAND2_X1 U5758 ( .A1(n4808), .A2(n5002), .ZN(n8544) );
  NAND2_X1 U5759 ( .A1(n4809), .A2(n4446), .ZN(n4808) );
  NAND2_X1 U5760 ( .A1(n6203), .A2(n6202), .ZN(n8809) );
  NAND2_X1 U5761 ( .A1(n6180), .A2(n6179), .ZN(n8815) );
  NAND2_X1 U5762 ( .A1(n6154), .A2(n6153), .ZN(n8829) );
  NAND2_X1 U5763 ( .A1(n6111), .A2(n6110), .ZN(n8842) );
  OAI21_X1 U5764 ( .B1(n6079), .B2(n4758), .A(n4755), .ZN(n8644) );
  NAND2_X1 U5765 ( .A1(n6094), .A2(n6093), .ZN(n8848) );
  NAND2_X1 U5766 ( .A1(n4760), .A2(n7843), .ZN(n8656) );
  NAND2_X1 U5767 ( .A1(n6079), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5768 ( .A1(n6083), .A2(n6082), .ZN(n8855) );
  NAND2_X1 U5769 ( .A1(n6079), .A2(n7911), .ZN(n8674) );
  NAND2_X1 U5770 ( .A1(n6072), .A2(n6071), .ZN(n8861) );
  INV_X1 U5771 ( .A(n8835), .ZN(n8862) );
  AND2_X1 U5772 ( .A1(n6368), .A2(n6367), .ZN(n10341) );
  NOR2_X1 U5773 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4989) );
  NAND2_X1 U5774 ( .A1(n6339), .A2(n6341), .ZN(n8879) );
  NAND2_X1 U5775 ( .A1(n6332), .A2(n5911), .ZN(n6340) );
  XNOR2_X1 U5776 ( .A(n6337), .B(n6336), .ZN(n7649) );
  NAND2_X1 U5777 ( .A1(n6334), .A2(n6335), .ZN(n7651) );
  XNOR2_X1 U5778 ( .A(n4595), .B(n4727), .ZN(n8485) );
  NAND2_X1 U5779 ( .A1(n6152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4595) );
  NOR2_X1 U5780 ( .A1(n5950), .A2(n5887), .ZN(n6031) );
  XNOR2_X1 U5781 ( .A(n5960), .B(n5959), .ZN(n6542) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U5783 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4884) );
  NAND2_X1 U5784 ( .A1(n6106), .A2(n5884), .ZN(n4883) );
  NAND2_X1 U5785 ( .A1(n7313), .A2(n7312), .ZN(n7692) );
  NAND2_X1 U5786 ( .A1(n4824), .A2(n7739), .ZN(n9181) );
  NAND2_X1 U5787 ( .A1(n9188), .A2(n9189), .ZN(n4544) );
  AND2_X1 U5788 ( .A1(n5295), .A2(n5294), .ZN(n9874) );
  NOR2_X1 U5789 ( .A1(n8194), .A2(n4820), .ZN(n4819) );
  INV_X1 U5790 ( .A(n7816), .ZN(n4820) );
  INV_X1 U5791 ( .A(n9804), .ZN(n10269) );
  AND4_X1 U5792 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(n9842)
         );
  AND2_X1 U5793 ( .A1(n4556), .A2(n4444), .ZN(n9271) );
  NAND2_X1 U5794 ( .A1(n9263), .A2(n9264), .ZN(n4556) );
  AND2_X1 U5795 ( .A1(n4816), .A2(n7797), .ZN(n4815) );
  AND2_X1 U5796 ( .A1(n6784), .A2(n6783), .ZN(n9357) );
  AND2_X1 U5797 ( .A1(n7125), .A2(n7122), .ZN(n7123) );
  XNOR2_X1 U5798 ( .A(n9188), .B(n9189), .ZN(n9325) );
  INV_X1 U5799 ( .A(n4545), .ZN(n9323) );
  AND4_X1 U5800 ( .A1(n5567), .A2(n5566), .A3(n5565), .A4(n5564), .ZN(n10274)
         );
  INV_X1 U5801 ( .A(n9359), .ZN(n9372) );
  AND2_X1 U5802 ( .A1(n6784), .A2(n6671), .ZN(n9352) );
  INV_X1 U5803 ( .A(n9361), .ZN(n9374) );
  AND4_X1 U5804 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n9528)
         );
  INV_X1 U5805 ( .A(n9664), .ZN(n9384) );
  NAND4_X1 U5806 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n9930)
         );
  NAND4_X1 U5807 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n9393)
         );
  NAND4_X1 U5808 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n9395)
         );
  OR2_X1 U5809 ( .A1(n5711), .A2(n6477), .ZN(n5466) );
  OR2_X1 U5810 ( .A1(n5490), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U5811 ( .A1(n9397), .A2(n9407), .ZN(n9396) );
  INV_X1 U5812 ( .A(n4649), .ZN(n10086) );
  INV_X1 U5813 ( .A(n4647), .ZN(n10096) );
  INV_X1 U5814 ( .A(n4645), .ZN(n10095) );
  NOR2_X1 U5815 ( .A1(n10110), .A2(n4642), .ZN(n6615) );
  AND2_X1 U5816 ( .A1(n6644), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4642) );
  NAND2_X1 U5817 ( .A1(n6615), .A2(n6616), .ZN(n9462) );
  NOR2_X1 U5818 ( .A1(n10129), .A2(n4651), .ZN(n10142) );
  AND2_X1 U5819 ( .A1(n10134), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4651) );
  NOR2_X1 U5820 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  XNOR2_X1 U5821 ( .A(n9466), .B(n9465), .ZN(n10158) );
  OR2_X1 U5822 ( .A1(n9482), .A2(n9483), .ZN(n9502) );
  OR2_X1 U5823 ( .A1(n6648), .A2(n6617), .ZN(n10156) );
  OR2_X1 U5824 ( .A1(n6648), .A2(n9408), .ZN(n10121) );
  NAND2_X1 U5825 ( .A1(n4909), .A2(n5343), .ZN(n9520) );
  NAND2_X1 U5826 ( .A1(n9516), .A2(n9932), .ZN(n9808) );
  XNOR2_X1 U5827 ( .A(n9515), .B(n9941), .ZN(n9516) );
  NAND2_X1 U5828 ( .A1(n4688), .A2(n8145), .ZN(n9533) );
  NAND2_X1 U5829 ( .A1(n4688), .A2(n4686), .ZN(n9812) );
  AND2_X1 U5830 ( .A1(n5318), .A2(n5317), .ZN(n9604) );
  AND4_X1 U5831 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n9841)
         );
  AND2_X1 U5832 ( .A1(n9647), .A2(n8151), .ZN(n9630) );
  INV_X1 U5833 ( .A(n9636), .ZN(n9854) );
  NAND2_X1 U5834 ( .A1(n4950), .A2(n5854), .ZN(n9711) );
  NOR2_X1 U5835 ( .A1(n9719), .A2(n4683), .ZN(n9706) );
  NAND2_X1 U5836 ( .A1(n5259), .A2(n5258), .ZN(n9914) );
  NAND2_X1 U5837 ( .A1(n9769), .A2(n5849), .ZN(n9754) );
  NAND2_X1 U5838 ( .A1(n7578), .A2(n5844), .ZN(n7617) );
  NAND2_X1 U5839 ( .A1(n6004), .A2(n5352), .ZN(n5207) );
  NAND2_X1 U5840 ( .A1(n7476), .A2(n7479), .ZN(n7475) );
  NAND2_X1 U5841 ( .A1(n7383), .A2(n7382), .ZN(n7476) );
  INV_X1 U5842 ( .A(n10191), .ZN(n10213) );
  NAND4_X1 U5843 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .ZN(n9391)
         );
  INV_X1 U5844 ( .A(n10236), .ZN(n8056) );
  NAND2_X1 U5845 ( .A1(n10005), .A2(n6680), .ZN(n10205) );
  INV_X1 U5846 ( .A(n10198), .ZN(n10211) );
  OR2_X1 U5847 ( .A1(n5711), .A2(n5456), .ZN(n5460) );
  OR2_X1 U5848 ( .A1(n5698), .A2(n6972), .ZN(n5461) );
  AND2_X1 U5849 ( .A1(n8188), .A2(n9833), .ZN(n8169) );
  AND2_X1 U5850 ( .A1(n10296), .A2(n10280), .ZN(n9833) );
  INV_X1 U5851 ( .A(n9520), .ZN(n9941) );
  AND2_X1 U5852 ( .A1(n9808), .A2(n9807), .ZN(n9939) );
  AND2_X1 U5853 ( .A1(n8188), .A2(n9955), .ZN(n8189) );
  XNOR2_X1 U5854 ( .A(n8147), .B(n8162), .ZN(n8186) );
  INV_X1 U5855 ( .A(n4686), .ZN(n4685) );
  OR2_X1 U5856 ( .A1(n5143), .A2(n10019), .ZN(n5329) );
  NAND2_X1 U5857 ( .A1(n8875), .A2(n5352), .ZN(n5330) );
  NAND2_X1 U5858 ( .A1(n5322), .A2(n5321), .ZN(n9956) );
  NAND2_X1 U5859 ( .A1(n7647), .A2(n5352), .ZN(n5322) );
  AND2_X1 U5860 ( .A1(n5314), .A2(n5313), .ZN(n9967) );
  OR2_X1 U5861 ( .A1(n5143), .A2(n7494), .ZN(n5313) );
  AND2_X1 U5862 ( .A1(n4679), .A2(n4682), .ZN(n9688) );
  NAND2_X1 U5863 ( .A1(n4680), .A2(n4443), .ZN(n4679) );
  INV_X1 U5864 ( .A(n9200), .ZN(n7607) );
  AND3_X1 U5865 ( .A1(n5201), .A2(n5200), .A3(n5199), .ZN(n7547) );
  AND2_X1 U5866 ( .A1(n5189), .A2(n4483), .ZN(n4547) );
  NAND2_X1 U5867 ( .A1(n4549), .A2(n5352), .ZN(n4548) );
  AND2_X1 U5868 ( .A1(n10289), .A2(n10280), .ZN(n9955) );
  AND3_X1 U5869 ( .A1(n5163), .A2(n5162), .A3(n5161), .ZN(n7103) );
  AND3_X1 U5870 ( .A1(n5153), .A2(n5152), .A3(n5151), .ZN(n8059) );
  NAND2_X1 U5871 ( .A1(n10008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5375) );
  XNOR2_X1 U5872 ( .A(n5134), .B(n4691), .ZN(n10021) );
  NAND2_X1 U5873 ( .A1(n5392), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U5874 ( .A(n5312), .B(n5311), .ZN(n7495) );
  NAND2_X1 U5875 ( .A1(n5357), .A2(n5356), .ZN(n5365) );
  INV_X1 U5876 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U5877 ( .A1(n4916), .A2(n4915), .ZN(n5237) );
  NAND2_X1 U5878 ( .A1(n4916), .A2(n4917), .ZN(n5236) );
  NAND2_X1 U5879 ( .A1(n4620), .A2(n4450), .ZN(n5216) );
  INV_X1 U5880 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U5881 ( .A1(n5186), .A2(n5185), .ZN(n5188) );
  NAND2_X1 U5882 ( .A1(n5180), .A2(n5039), .ZN(n5186) );
  NAND2_X1 U5883 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4641) );
  AOI21_X1 U5884 ( .B1(n10138), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9509), .ZN(
        n4656) );
  NAND2_X1 U5885 ( .A1(n4653), .A2(n6973), .ZN(n4652) );
  NAND2_X1 U5886 ( .A1(n9508), .A2(n5722), .ZN(n4657) );
  OAI21_X1 U5887 ( .B1(n9514), .B2(n9935), .A(n5416), .ZN(n5417) );
  OAI21_X1 U5888 ( .B1(n9514), .B2(n10000), .A(n5423), .ZN(n5424) );
  AND2_X1 U5889 ( .A1(n4574), .A2(n4765), .ZN(n6044) );
  AND2_X1 U5890 ( .A1(n5306), .A2(n5305), .ZN(n7781) );
  OR2_X1 U5891 ( .A1(n8815), .A2(n8578), .ZN(n7950) );
  NOR2_X1 U5892 ( .A1(n7872), .A2(n7873), .ZN(n4427) );
  INV_X1 U5893 ( .A(n5706), .ZN(n4713) );
  NAND2_X1 U5894 ( .A1(n5925), .A2(n5884), .ZN(n5937) );
  AND3_X1 U5895 ( .A1(n4467), .A2(n4825), .A3(n4938), .ZN(n5363) );
  NAND2_X1 U5896 ( .A1(n6044), .A2(n4455), .ZN(n6269) );
  AND2_X1 U5897 ( .A1(n6046), .A2(n4597), .ZN(n4428) );
  AND2_X1 U5898 ( .A1(n6213), .A2(n4749), .ZN(n4429) );
  INV_X1 U5899 ( .A(n7871), .ZN(n4832) );
  AND2_X1 U5900 ( .A1(n8139), .A2(n4665), .ZN(n4430) );
  OR2_X1 U5901 ( .A1(n8699), .A2(n8355), .ZN(n4431) );
  NAND2_X1 U5902 ( .A1(n6192), .A2(n6191), .ZN(n8803) );
  NOR2_X1 U5903 ( .A1(n5090), .A2(n5296), .ZN(n4432) );
  AND2_X1 U5904 ( .A1(n4475), .A2(n4858), .ZN(n4433) );
  AND2_X1 U5905 ( .A1(n4605), .A2(n4604), .ZN(n4434) );
  AND2_X1 U5906 ( .A1(n8118), .A2(n9794), .ZN(n4435) );
  NOR2_X1 U5907 ( .A1(n8791), .A2(n8258), .ZN(n4436) );
  INV_X1 U5908 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5894) );
  AND2_X1 U5909 ( .A1(n7151), .A2(n7148), .ZN(n4437) );
  OR2_X1 U5910 ( .A1(n8737), .A2(n8234), .ZN(n8601) );
  AND2_X1 U5911 ( .A1(n5354), .A2(n5130), .ZN(n4438) );
  AND2_X1 U5912 ( .A1(n4603), .A2(n4602), .ZN(n4439) );
  AND2_X1 U5913 ( .A1(n5850), .A2(n5849), .ZN(n4440) );
  AND2_X1 U5914 ( .A1(n6286), .A2(n6285), .ZN(n4441) );
  AND2_X1 U5915 ( .A1(n7629), .A2(n8359), .ZN(n7597) );
  AND2_X1 U5916 ( .A1(n4596), .A2(n6108), .ZN(n4442) );
  AND2_X1 U5917 ( .A1(n4681), .A2(n8124), .ZN(n4443) );
  INV_X1 U5918 ( .A(n7046), .ZN(n4536) );
  INV_X1 U5919 ( .A(n7781), .ZN(n9650) );
  NAND2_X1 U5920 ( .A1(n9762), .A2(n4603), .ZN(n5008) );
  NAND2_X1 U5921 ( .A1(n8160), .A2(n5728), .ZN(n9546) );
  INV_X1 U5922 ( .A(n8128), .ZN(n4668) );
  INV_X1 U5923 ( .A(n5720), .ZN(n6845) );
  NAND2_X1 U5924 ( .A1(n7754), .A2(n7753), .ZN(n4444) );
  INV_X1 U5925 ( .A(n6289), .ZN(n4793) );
  NAND2_X1 U5926 ( .A1(n4874), .A2(n6546), .ZN(n4873) );
  NAND2_X2 U5927 ( .A1(n5167), .A2(n6392), .ZN(n5143) );
  NAND2_X2 U5928 ( .A1(n6385), .A2(n5928), .ZN(n5952) );
  NAND2_X1 U5929 ( .A1(n4936), .A2(n5495), .ZN(n5786) );
  NAND2_X1 U5930 ( .A1(n6385), .A2(n6392), .ZN(n5953) );
  NOR2_X1 U5931 ( .A1(n5194), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5196) );
  XNOR2_X1 U5932 ( .A(n5913), .B(n5912), .ZN(n6318) );
  NOR2_X1 U5933 ( .A1(n8350), .A2(n4970), .ZN(n4445) );
  INV_X1 U5934 ( .A(n7653), .ZN(n4966) );
  NAND2_X1 U5935 ( .A1(n6271), .A2(n5894), .ZN(n6275) );
  NAND2_X1 U5936 ( .A1(n9647), .A2(n4947), .ZN(n9607) );
  OR2_X1 U5937 ( .A1(n8809), .A2(n8570), .ZN(n4446) );
  AND2_X1 U5938 ( .A1(n5003), .A2(n4446), .ZN(n4447) );
  NOR3_X1 U5939 ( .A1(n9598), .A2(n4607), .A3(n4466), .ZN(n4606) );
  AND2_X1 U5940 ( .A1(n8155), .A2(n5778), .ZN(n4448) );
  AND2_X1 U5941 ( .A1(n8131), .A2(n4668), .ZN(n4449) );
  INV_X1 U5942 ( .A(n4747), .ZN(n4746) );
  NAND2_X1 U5943 ( .A1(n4429), .A2(n7958), .ZN(n4747) );
  NAND2_X1 U5944 ( .A1(n5914), .A2(n4989), .ZN(n5902) );
  OR2_X1 U5945 ( .A1(n5054), .A2(SI_9_), .ZN(n4450) );
  AND4_X1 U5946 ( .A1(n5531), .A2(n6845), .A3(n5837), .A4(n5794), .ZN(n4451)
         );
  NAND2_X1 U5947 ( .A1(n4664), .A2(n4663), .ZN(n9572) );
  NAND2_X1 U5948 ( .A1(n8295), .A2(n8083), .ZN(n8246) );
  AND2_X1 U5949 ( .A1(n7790), .A2(n4817), .ZN(n4452) );
  AND2_X1 U5950 ( .A1(n5128), .A2(n4937), .ZN(n4453) );
  NAND2_X1 U5951 ( .A1(n5330), .A2(n5329), .ZN(n9946) );
  INV_X1 U5952 ( .A(n7925), .ZN(n4754) );
  AOI21_X1 U5953 ( .B1(n6330), .B2(n8690), .A(n6329), .ZN(n7668) );
  NAND2_X1 U5954 ( .A1(n8230), .A2(n5000), .ZN(n8294) );
  AND2_X1 U5955 ( .A1(n4645), .A2(n4644), .ZN(n4454) );
  AND2_X1 U5956 ( .A1(n5893), .A2(n4991), .ZN(n4455) );
  OR2_X1 U5957 ( .A1(n7550), .A2(n9930), .ZN(n4456) );
  NAND2_X1 U5958 ( .A1(n6044), .A2(n5893), .ZN(n6267) );
  OR2_X1 U5959 ( .A1(n7323), .A2(n6776), .ZN(n4457) );
  NOR2_X1 U5960 ( .A1(n5569), .A2(n6845), .ZN(n4458) );
  AND2_X1 U5961 ( .A1(n6542), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U5962 ( .A1(n4639), .A2(n4850), .ZN(n4460) );
  AND2_X1 U5963 ( .A1(n9607), .A2(n8153), .ZN(n4461) );
  NAND2_X1 U5964 ( .A1(n7005), .A2(n7011), .ZN(n4462) );
  AND2_X1 U5965 ( .A1(n5837), .A2(n5495), .ZN(n4463) );
  AND2_X1 U5966 ( .A1(n4702), .A2(n6845), .ZN(n4464) );
  INV_X1 U5967 ( .A(n7323), .ZN(n9389) );
  AND4_X1 U5968 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n7323)
         );
  INV_X1 U5969 ( .A(n7296), .ZN(n9390) );
  AND4_X1 U5970 ( .A1(n5507), .A2(n5506), .A3(n5505), .A4(n5504), .ZN(n7296)
         );
  OAI21_X1 U5971 ( .B1(n4919), .B2(n4914), .A(n5064), .ZN(n4913) );
  OR2_X1 U5972 ( .A1(n4913), .A2(n4615), .ZN(n4465) );
  INV_X1 U5973 ( .A(n6304), .ZN(n4777) );
  OR2_X1 U5974 ( .A1(n9814), .A2(n9946), .ZN(n4466) );
  OR2_X1 U5975 ( .A1(n6997), .A2(n6890), .ZN(n7863) );
  OR2_X1 U5976 ( .A1(n8797), .A2(n6223), .ZN(n7958) );
  AND2_X1 U5977 ( .A1(n4438), .A2(n5131), .ZN(n4467) );
  NAND2_X1 U5978 ( .A1(n6885), .A2(n5940), .ZN(n8003) );
  INV_X1 U5979 ( .A(n4918), .ZN(n4917) );
  NOR2_X1 U5980 ( .A1(n5060), .A2(SI_11_), .ZN(n4918) );
  INV_X1 U5981 ( .A(n6602), .ZN(n5917) );
  NOR2_X1 U5982 ( .A1(n8645), .A2(n6302), .ZN(n4468) );
  AND2_X1 U5983 ( .A1(n5828), .A2(n5766), .ZN(n8162) );
  INV_X1 U5984 ( .A(n8162), .ZN(n4714) );
  NAND2_X1 U5985 ( .A1(n5803), .A2(n5736), .ZN(n4469) );
  AND2_X1 U5986 ( .A1(n7958), .A2(n7957), .ZN(n8533) );
  INV_X1 U5987 ( .A(n8533), .ZN(n4805) );
  AND3_X1 U5988 ( .A1(n5893), .A2(n4766), .A3(n4765), .ZN(n6271) );
  NAND2_X1 U5989 ( .A1(n7985), .A2(n7971), .ZN(n8029) );
  INV_X1 U5990 ( .A(n8029), .ZN(n4632) );
  INV_X1 U5991 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5410) );
  INV_X1 U5992 ( .A(n4915), .ZN(n4914) );
  NOR2_X1 U5993 ( .A1(n5235), .A2(n4918), .ZN(n4915) );
  NAND2_X1 U5994 ( .A1(n5694), .A2(n5727), .ZN(n4470) );
  OR3_X1 U5995 ( .A1(n5706), .A2(n5824), .A3(n4715), .ZN(n4471) );
  AND2_X1 U5997 ( .A1(n7323), .A2(n10199), .ZN(n4472) );
  AND2_X1 U5998 ( .A1(n4747), .A2(n4742), .ZN(n4473) );
  OR2_X1 U5999 ( .A1(n4966), .A2(n4963), .ZN(n4474) );
  AND2_X1 U6000 ( .A1(n5897), .A2(n5896), .ZN(n4475) );
  AND2_X1 U6001 ( .A1(n4638), .A2(n4637), .ZN(n4476) );
  NAND2_X1 U6002 ( .A1(n8767), .A2(n6998), .ZN(n5930) );
  AND2_X1 U6003 ( .A1(n7992), .A2(n7991), .ZN(n4477) );
  OR2_X1 U6004 ( .A1(n4436), .A2(n7960), .ZN(n8524) );
  OR2_X1 U6005 ( .A1(n6393), .A2(n6392), .ZN(n4478) );
  NAND2_X1 U6006 ( .A1(n8088), .A2(n8087), .ZN(n4479) );
  OR2_X1 U6007 ( .A1(n5005), .A2(n4807), .ZN(n4480) );
  OR2_X1 U6008 ( .A1(n7470), .A2(n7623), .ZN(n4792) );
  AND2_X1 U6009 ( .A1(n4743), .A2(n4742), .ZN(n4481) );
  AND3_X1 U6010 ( .A1(n6104), .A2(n6103), .A3(n6102), .ZN(n4482) );
  OR2_X1 U6011 ( .A1(n6429), .A2(n10105), .ZN(n4483) );
  AND2_X1 U6012 ( .A1(n6201), .A2(n6200), .ZN(n8285) );
  AND2_X1 U6013 ( .A1(n6069), .A2(n7900), .ZN(n4484) );
  AND2_X1 U6014 ( .A1(n4947), .A2(n8154), .ZN(n4485) );
  AND2_X1 U6015 ( .A1(n6030), .A2(n7885), .ZN(n4486) );
  AND2_X1 U6016 ( .A1(n5356), .A2(n4813), .ZN(n4487) );
  AND2_X1 U6017 ( .A1(n5911), .A2(n4979), .ZN(n4488) );
  AND2_X1 U6018 ( .A1(n9540), .A2(n4948), .ZN(n4489) );
  AND2_X1 U6019 ( .A1(n4805), .A2(n4806), .ZN(n4490) );
  OR2_X1 U6020 ( .A1(n7597), .A2(n4966), .ZN(n4491) );
  OR2_X1 U6021 ( .A1(n8076), .A2(n8672), .ZN(n4492) );
  INV_X1 U6022 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6023 ( .A1(n7859), .A2(n7863), .ZN(n4835) );
  INV_X1 U6024 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4597) );
  OAI21_X1 U6025 ( .B1(n7293), .B2(n4821), .A(n4541), .ZN(n9226) );
  AND3_X1 U6026 ( .A1(n4938), .A2(n5196), .A3(n4453), .ZN(n5272) );
  OR2_X1 U6027 ( .A1(n9665), .A2(n9867), .ZN(n4493) );
  NAND2_X1 U6028 ( .A1(n7737), .A2(n7736), .ZN(n7739) );
  XNOR2_X1 U6029 ( .A(n5339), .B(SI_29_), .ZN(n8192) );
  AND2_X1 U6030 ( .A1(n9762), .A2(n4439), .ZN(n4494) );
  AND3_X1 U6031 ( .A1(n5173), .A2(n5172), .A3(n5171), .ZN(n7275) );
  INV_X1 U6032 ( .A(n8273), .ZN(n4587) );
  NAND2_X1 U6033 ( .A1(n9365), .A2(n7746), .ZN(n9263) );
  INV_X1 U6034 ( .A(n7973), .ZN(n7977) );
  INV_X1 U6035 ( .A(n7977), .ZN(n4530) );
  OAI22_X1 U6036 ( .A1(n8262), .A2(n4580), .B1(n8273), .B2(n4582), .ZN(n8322)
         );
  NAND2_X1 U6037 ( .A1(n7609), .A2(n7608), .ZN(n8121) );
  OAI21_X1 U6038 ( .B1(n8667), .B2(n6296), .A(n6295), .ZN(n8657) );
  AOI22_X1 U6039 ( .A1(n10014), .A2(n7968), .B1(n7677), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U6040 ( .A1(n5301), .A2(n5300), .ZN(n9867) );
  AND2_X1 U6041 ( .A1(n4571), .A2(n4570), .ZN(n8072) );
  INV_X1 U6042 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4886) );
  OR2_X1 U6043 ( .A1(n5074), .A2(SI_16_), .ZN(n4495) );
  XNOR2_X1 U6044 ( .A(n4641), .B(n8881), .ZN(n6620) );
  NAND2_X1 U6045 ( .A1(n5281), .A2(n5280), .ZN(n9888) );
  INV_X1 U6046 ( .A(n9888), .ZN(n4602) );
  INV_X1 U6047 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4691) );
  AND2_X1 U6048 ( .A1(n9273), .A2(n7759), .ZN(n4496) );
  AND3_X1 U6049 ( .A1(n4824), .A2(n7739), .A3(n7738), .ZN(n4497) );
  NAND2_X1 U6050 ( .A1(n5196), .A2(n4938), .ZN(n4498) );
  OR2_X1 U6051 ( .A1(n6382), .A2(n8835), .ZN(n4499) );
  AND4_X1 U6052 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9527)
         );
  NAND2_X1 U6053 ( .A1(n4732), .A2(n7885), .ZN(n7301) );
  NAND2_X1 U6054 ( .A1(n5196), .A2(n5127), .ZN(n5255) );
  INV_X1 U6055 ( .A(n9794), .ZN(n8119) );
  AND4_X1 U6056 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n9794)
         );
  OR2_X1 U6057 ( .A1(n6382), .A2(n8742), .ZN(n4500) );
  AND2_X1 U6058 ( .A1(n5265), .A2(n5264), .ZN(n9905) );
  INV_X1 U6059 ( .A(n9905), .ZN(n9747) );
  INV_X1 U6060 ( .A(n9294), .ZN(n9388) );
  AND4_X1 U6061 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n9294)
         );
  INV_X1 U6062 ( .A(n9232), .ZN(n9928) );
  AND4_X1 U6063 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5539), .ZN(n9232)
         );
  INV_X1 U6064 ( .A(n10254), .ZN(n9387) );
  AND4_X1 U6065 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n10254)
         );
  OR3_X1 U6066 ( .A1(n7914), .A2(n8686), .A3(n7973), .ZN(n4501) );
  AND2_X1 U6067 ( .A1(n9604), .A2(n9842), .ZN(n4502) );
  AND2_X1 U6068 ( .A1(n8079), .A2(n8234), .ZN(n4503) );
  OR2_X1 U6069 ( .A1(n7769), .A2(n7768), .ZN(n4504) );
  AND2_X1 U6070 ( .A1(n5091), .A2(SI_21_), .ZN(n4505) );
  INV_X1 U6071 ( .A(n4585), .ZN(n4584) );
  NAND2_X1 U6072 ( .A1(n8263), .A2(n8659), .ZN(n4585) );
  NAND2_X1 U6073 ( .A1(n5334), .A2(n5333), .ZN(n9814) );
  INV_X1 U6074 ( .A(n9722), .ZN(n4677) );
  AND2_X1 U6075 ( .A1(n5732), .A2(n5854), .ZN(n9722) );
  NAND2_X1 U6076 ( .A1(n5286), .A2(n5285), .ZN(n9701) );
  OR2_X1 U6077 ( .A1(n5276), .A2(n4929), .ZN(n4506) );
  OR2_X1 U6078 ( .A1(n4557), .A2(n4496), .ZN(n4507) );
  AND2_X1 U6079 ( .A1(n6044), .A2(n4596), .ZN(n4508) );
  OR2_X1 U6080 ( .A1(n5091), .A2(SI_21_), .ZN(n4509) );
  NOR2_X1 U6081 ( .A1(n7628), .A2(n7597), .ZN(n4510) );
  NOR2_X1 U6082 ( .A1(n4933), .A2(n9032), .ZN(n4511) );
  AND2_X1 U6083 ( .A1(n9687), .A2(n4682), .ZN(n4512) );
  AND2_X1 U6084 ( .A1(n5326), .A2(n5325), .ZN(n9824) );
  INV_X1 U6085 ( .A(n9824), .ZN(n9563) );
  OR2_X1 U6086 ( .A1(n4625), .A2(n5287), .ZN(n4513) );
  AND2_X1 U6087 ( .A1(n9882), .A2(n4439), .ZN(n4514) );
  AND2_X1 U6088 ( .A1(n9814), .A2(n8146), .ZN(n4515) );
  NOR2_X1 U6089 ( .A1(n6277), .A2(n6276), .ZN(n8043) );
  INV_X1 U6090 ( .A(n8043), .ZN(n4857) );
  NAND2_X1 U6091 ( .A1(n4978), .A2(n4977), .ZN(n4593) );
  NAND2_X1 U6092 ( .A1(n8043), .A2(n8034), .ZN(n7973) );
  OAI22_X1 U6093 ( .A1(n4591), .A2(n4590), .B1(n4437), .B2(n4589), .ZN(n7411)
         );
  NOR2_X1 U6094 ( .A1(n6781), .A2(n6782), .ZN(n6929) );
  OR2_X1 U6095 ( .A1(n9931), .A2(n10184), .ZN(n5009) );
  AND2_X1 U6096 ( .A1(n7589), .A2(n8118), .ZN(n4516) );
  AND2_X1 U6097 ( .A1(n7588), .A2(n7607), .ZN(n7589) );
  AND2_X1 U6098 ( .A1(n6642), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4517) );
  AND2_X1 U6099 ( .A1(n5414), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4518) );
  AND2_X1 U6100 ( .A1(n10287), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U6101 ( .A1(n7293), .A2(n7294), .ZN(n7313) );
  NAND2_X1 U6102 ( .A1(n4733), .A2(n7900), .ZN(n7556) );
  OR2_X1 U6103 ( .A1(n7412), .A2(n7623), .ZN(n4520) );
  INV_X1 U6104 ( .A(n4788), .ZN(n4787) );
  NOR2_X1 U6105 ( .A1(n6291), .A2(n4789), .ZN(n4788) );
  AND2_X1 U6106 ( .A1(n7149), .A2(n4437), .ZN(n4521) );
  INV_X1 U6107 ( .A(n8216), .ZN(n4973) );
  AND2_X1 U6108 ( .A1(n5124), .A2(n5123), .ZN(n4522) );
  INV_X1 U6109 ( .A(n4444), .ZN(n4557) );
  NAND2_X1 U6110 ( .A1(n5251), .A2(n5250), .ZN(n10279) );
  INV_X1 U6111 ( .A(n10279), .ZN(n4604) );
  NAND2_X1 U6112 ( .A1(n4983), .A2(n4986), .ZN(n6690) );
  OR2_X1 U6113 ( .A1(n8425), .A2(n8745), .ZN(n4523) );
  INV_X1 U6114 ( .A(n4873), .ZN(n6717) );
  INV_X1 U6115 ( .A(n8034), .ZN(n4855) );
  INV_X1 U6116 ( .A(n6517), .ZN(n4880) );
  XOR2_X1 U6117 ( .A(n10050), .B(P1_REG2_REG_8__SCAN_IN), .Z(n4524) );
  AND2_X1 U6118 ( .A1(n8034), .A2(n8038), .ZN(n4525) );
  INV_X1 U6119 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6120 ( .A1(n4724), .A2(n4448), .ZN(n5654) );
  NAND2_X1 U6121 ( .A1(n4698), .A2(n4693), .ZN(n5602) );
  NAND2_X1 U6122 ( .A1(n5570), .A2(n5802), .ZN(n4694) );
  NAND2_X1 U6123 ( .A1(n5155), .A2(n5154), .ZN(n5157) );
  NAND2_X1 U6124 ( .A1(n5209), .A2(n5208), .ZN(n4620) );
  INV_X1 U6125 ( .A(n4965), .ZN(n4964) );
  NAND2_X1 U6126 ( .A1(n4831), .A2(n8037), .ZN(n4830) );
  NAND2_X1 U6127 ( .A1(n4859), .A2(n4501), .ZN(n7921) );
  NAND2_X1 U6128 ( .A1(n4863), .A2(n4862), .ZN(n4861) );
  AOI21_X1 U6129 ( .B1(n7926), .B2(n7925), .A(n4532), .ZN(n7927) );
  NAND2_X1 U6130 ( .A1(n4841), .A2(n4635), .ZN(n4634) );
  XNOR2_X1 U6131 ( .A(n8453), .B(n8452), .ZN(n8423) );
  OAI21_X1 U6132 ( .B1(n4873), .B2(n4872), .A(n4871), .ZN(n6822) );
  NOR2_X1 U6133 ( .A1(n8661), .A2(n8370), .ZN(n8394) );
  NOR2_X1 U6134 ( .A1(n7173), .A2(n7172), .ZN(n7191) );
  NAND2_X1 U6135 ( .A1(n4608), .A2(n5052), .ZN(n5209) );
  AOI21_X1 U6136 ( .B1(n8187), .B2(n10296), .A(n4533), .ZN(n8170) );
  AOI21_X1 U6137 ( .B1(n8187), .B2(n10289), .A(n4534), .ZN(n8190) );
  NAND2_X1 U6138 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  AOI21_X2 U6139 ( .B1(n8457), .B2(n8456), .A(n8455), .ZN(n8476) );
  INV_X1 U6140 ( .A(n6496), .ZN(n4881) );
  NOR2_X1 U6141 ( .A1(n7510), .A2(n7511), .ZN(n7514) );
  INV_X1 U6142 ( .A(n7169), .ZN(n4869) );
  NAND2_X1 U6143 ( .A1(n4537), .A2(n7746), .ZN(n9368) );
  OR2_X1 U6144 ( .A1(n7737), .A2(n4540), .ZN(n4539) );
  OAI21_X2 U6145 ( .B1(n9263), .B2(n4553), .A(n4551), .ZN(n4558) );
  AOI21_X2 U6146 ( .B1(n4558), .B2(n7779), .A(n9304), .ZN(n9237) );
  NAND2_X1 U6147 ( .A1(n6860), .A2(n4567), .ZN(n4564) );
  NOR2_X1 U6148 ( .A1(n7031), .A2(n4568), .ZN(n7163) );
  NAND2_X1 U6149 ( .A1(n6858), .A2(n6859), .ZN(n4569) );
  INV_X1 U6150 ( .A(n6750), .ZN(n6752) );
  NAND2_X1 U6151 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  INV_X1 U6152 ( .A(n4572), .ZN(n7630) );
  AOI22_X1 U6153 ( .A1(n4961), .A2(n7597), .B1(n4964), .B2(n4491), .ZN(n4570)
         );
  OAI21_X1 U6154 ( .B1(n4961), .B2(n4964), .A(n4572), .ZN(n4571) );
  NAND2_X1 U6155 ( .A1(n8230), .A2(n4577), .ZN(n4575) );
  NAND2_X1 U6156 ( .A1(n4575), .A2(n4576), .ZN(n8223) );
  INV_X1 U6157 ( .A(n4593), .ZN(n4591) );
  NAND2_X1 U6158 ( .A1(n6044), .A2(n4442), .ZN(n6134) );
  NAND3_X1 U6159 ( .A1(n7781), .A2(n9967), .A3(n4600), .ZN(n4599) );
  AND3_X1 U6160 ( .A1(n4825), .A2(n4438), .A3(n4938), .ZN(n5360) );
  NAND4_X1 U6161 ( .A1(n4467), .A2(n4825), .A3(n4958), .A4(n4938), .ZN(n5392)
         );
  INV_X1 U6162 ( .A(n4606), .ZN(n8168) );
  NAND2_X1 U6163 ( .A1(n5204), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U6164 ( .A1(n4621), .A2(n4623), .ZN(n5312) );
  NAND3_X1 U6165 ( .A1(n7949), .A2(n7973), .A3(n8550), .ZN(n4637) );
  MUX2_X1 U6166 ( .A(n5456), .B(P1_REG2_REG_1__SCAN_IN), .S(n6620), .Z(n9397)
         );
  NAND3_X1 U6167 ( .A1(n4657), .A2(n4656), .A3(n4652), .ZN(P1_U3262) );
  OAI21_X1 U6168 ( .B1(n7383), .B2(n4659), .A(n4661), .ZN(n7385) );
  NAND3_X1 U6169 ( .A1(n4660), .A2(n4658), .A3(n7384), .ZN(n7457) );
  NAND2_X1 U6170 ( .A1(n4661), .A2(n4659), .ZN(n4658) );
  INV_X1 U6171 ( .A(n7479), .ZN(n4659) );
  NAND2_X1 U6172 ( .A1(n7383), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U6173 ( .A1(n9660), .A2(n4430), .ZN(n4664) );
  AOI21_X1 U6174 ( .B1(n9660), .B2(n8129), .A(n8128), .ZN(n9643) );
  NAND2_X1 U6175 ( .A1(n7584), .A2(n4671), .ZN(n4670) );
  INV_X1 U6176 ( .A(n9720), .ZN(n4678) );
  NAND2_X1 U6177 ( .A1(n4674), .A2(n4675), .ZN(n9686) );
  NAND2_X1 U6178 ( .A1(n9720), .A2(n4443), .ZN(n4674) );
  AND2_X1 U6179 ( .A1(n9725), .A2(n9901), .ZN(n4683) );
  NAND2_X1 U6180 ( .A1(n9541), .A2(n9546), .ZN(n4688) );
  OAI21_X1 U6181 ( .B1(n9541), .B2(n4685), .A(n4684), .ZN(n8147) );
  AOI21_X1 U6182 ( .B1(n4686), .B2(n8159), .A(n4515), .ZN(n4684) );
  NAND2_X1 U6183 ( .A1(n5360), .A2(n4689), .ZN(n4692) );
  INV_X1 U6184 ( .A(n4692), .ZN(n5373) );
  NAND4_X1 U6185 ( .A1(n4707), .A2(n4705), .A3(n5535), .A4(n4703), .ZN(n5545)
         );
  MUX2_X1 U6186 ( .A(n9074), .B(n9007), .S(n6392), .Z(n5113) );
  MUX2_X1 U6187 ( .A(n10016), .B(n6245), .S(n6392), .Z(n5124) );
  NAND2_X1 U6188 ( .A1(n5012), .A2(n4708), .ZN(n5015) );
  NAND2_X1 U6189 ( .A1(n6392), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U6190 ( .A1(n5178), .A2(n5177), .ZN(n5180) );
  NAND2_X1 U6191 ( .A1(n5178), .A2(n4718), .ZN(n4717) );
  NAND3_X1 U6192 ( .A1(n5646), .A2(n4726), .A3(n9629), .ZN(n4725) );
  INV_X1 U6193 ( .A(n6004), .ZN(n6408) );
  XNOR2_X1 U6194 ( .A(n5204), .B(n5205), .ZN(n6004) );
  NAND4_X1 U6195 ( .A1(n6103), .A2(n4597), .A3(n5890), .A4(n4727), .ZN(n5891)
         );
  OAI211_X2 U6196 ( .C1(n5952), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n4729), .B(
        n4728), .ZN(n6741) );
  NAND2_X1 U6197 ( .A1(n6385), .A2(n4730), .ZN(n4728) );
  NAND2_X1 U6198 ( .A1(n4731), .A2(n6458), .ZN(n4729) );
  INV_X2 U6199 ( .A(n6385), .ZN(n4731) );
  INV_X2 U6200 ( .A(n8001), .ZN(n6280) );
  AND2_X2 U6201 ( .A1(n5930), .A2(n7848), .ZN(n8001) );
  NAND2_X1 U6202 ( .A1(n4732), .A2(n4486), .ZN(n7439) );
  NAND2_X1 U6203 ( .A1(n4733), .A2(n4484), .ZN(n8761) );
  INV_X1 U6204 ( .A(n7993), .ZN(n4735) );
  NAND2_X1 U6205 ( .A1(n4481), .A2(n8567), .ZN(n4740) );
  NAND2_X1 U6206 ( .A1(n4752), .A2(n4753), .ZN(n6120) );
  NAND2_X1 U6207 ( .A1(n6079), .A2(n4755), .ZN(n4752) );
  INV_X1 U6208 ( .A(n5950), .ZN(n4765) );
  NAND4_X1 U6209 ( .A1(n5893), .A2(n4764), .A3(n4858), .A4(n4763), .ZN(n4778)
         );
  NAND3_X1 U6210 ( .A1(n4991), .A2(n5888), .A3(n4768), .ZN(n4767) );
  OAI21_X2 U6211 ( .B1(n6299), .B2(n4775), .A(n4773), .ZN(n8603) );
  AOI21_X2 U6212 ( .B1(n8603), .B2(n6307), .A(n6306), .ZN(n8588) );
  NAND2_X1 U6213 ( .A1(n4792), .A2(n4787), .ZN(n4780) );
  NAND2_X1 U6214 ( .A1(n4788), .A2(n6289), .ZN(n4786) );
  NAND2_X1 U6215 ( .A1(n4796), .A2(n6688), .ZN(n4794) );
  NAND3_X1 U6216 ( .A1(n6281), .A2(n4795), .A3(n4794), .ZN(n6794) );
  NAND2_X1 U6217 ( .A1(n8003), .A2(n6885), .ZN(n4795) );
  NOR2_X1 U6218 ( .A1(n4799), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U6219 ( .A1(n4798), .A2(n7847), .ZN(n6884) );
  NAND2_X1 U6220 ( .A1(n6688), .A2(n6999), .ZN(n4798) );
  INV_X1 U6221 ( .A(n6999), .ZN(n4799) );
  INV_X1 U6222 ( .A(n8559), .ZN(n4809) );
  NAND2_X1 U6223 ( .A1(n4800), .A2(n4802), .ZN(n8525) );
  NAND2_X1 U6224 ( .A1(n8559), .A2(n4490), .ZN(n4800) );
  NAND2_X1 U6225 ( .A1(n4810), .A2(n4441), .ZN(n7214) );
  OAI21_X2 U6226 ( .B1(n8684), .B2(n7904), .A(n7902), .ZN(n8667) );
  NAND2_X1 U6227 ( .A1(n5357), .A2(n4487), .ZN(n5367) );
  NAND2_X1 U6228 ( .A1(n4814), .A2(n4815), .ZN(n9280) );
  NAND2_X1 U6229 ( .A1(n9237), .A2(n4452), .ZN(n4814) );
  NAND2_X1 U6230 ( .A1(n9237), .A2(n9238), .ZN(n9236) );
  NAND2_X1 U6231 ( .A1(n9353), .A2(n4819), .ZN(n8196) );
  NAND2_X1 U6232 ( .A1(n9353), .A2(n7816), .ZN(n8195) );
  NAND2_X4 U6233 ( .A1(n6660), .A2(n6661), .ZN(n7826) );
  INV_X2 U6234 ( .A(n6924), .ZN(n7798) );
  NOR2_X2 U6235 ( .A1(n5194), .A2(n4826), .ZN(n4825) );
  XNOR2_X1 U6236 ( .A(n4829), .B(n8485), .ZN(n8046) );
  OAI21_X1 U6237 ( .B1(n7982), .B2(n4830), .A(n8039), .ZN(n4829) );
  NAND2_X1 U6238 ( .A1(n7984), .A2(n7983), .ZN(n4831) );
  NAND2_X1 U6239 ( .A1(n4837), .A2(n4836), .ZN(n7865) );
  NAND3_X1 U6240 ( .A1(n7861), .A2(n7868), .A3(n4838), .ZN(n4837) );
  NAND2_X1 U6241 ( .A1(n4839), .A2(n7859), .ZN(n7870) );
  INV_X1 U6242 ( .A(n7948), .ZN(n4840) );
  INV_X1 U6243 ( .A(n7946), .ZN(n4853) );
  NAND3_X1 U6244 ( .A1(n4865), .A2(n4864), .A3(n6069), .ZN(n4863) );
  NAND3_X1 U6245 ( .A1(n7896), .A2(n7898), .A3(n4530), .ZN(n4864) );
  NAND3_X1 U6246 ( .A1(n7901), .A2(n7977), .A3(n7900), .ZN(n4865) );
  NOR2_X4 U6247 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5925) );
  INV_X1 U6248 ( .A(n4866), .ZN(n7232) );
  NAND2_X1 U6249 ( .A1(n7170), .A2(n7171), .ZN(n4868) );
  INV_X1 U6250 ( .A(n6716), .ZN(n4875) );
  AND2_X1 U6251 ( .A1(n6714), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4874) );
  NAND2_X1 U6252 ( .A1(n4878), .A2(n6525), .ZN(n6523) );
  OR2_X2 U6253 ( .A1(n8423), .A2(n9059), .ZN(n8457) );
  OAI211_X1 U6254 ( .C1(n4425), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4885), .ZN(n5014) );
  NAND2_X1 U6255 ( .A1(n4425), .A2(n4886), .ZN(n4885) );
  AND2_X4 U6256 ( .A1(n4887), .A2(n4888), .ZN(n6392) );
  NAND2_X2 U6257 ( .A1(n6909), .A2(n5011), .ZN(n4887) );
  NAND2_X1 U6258 ( .A1(n6908), .A2(n5010), .ZN(n4888) );
  NAND2_X1 U6259 ( .A1(n5316), .A2(n4893), .ZN(n4891) );
  NAND2_X1 U6260 ( .A1(n5327), .A2(n4899), .ZN(n4897) );
  NAND2_X1 U6261 ( .A1(n5327), .A2(n5328), .ZN(n4898) );
  NAND2_X1 U6262 ( .A1(n5299), .A2(n4904), .ZN(n4903) );
  NAND2_X1 U6263 ( .A1(n8114), .A2(n5352), .ZN(n4909) );
  NAND2_X1 U6264 ( .A1(n5073), .A2(n5072), .ZN(n5266) );
  NAND3_X1 U6265 ( .A1(n5073), .A2(n5072), .A3(n4922), .ZN(n4921) );
  NAND3_X1 U6266 ( .A1(n5073), .A2(n5072), .A3(n4926), .ZN(n4925) );
  NAND3_X1 U6267 ( .A1(n5073), .A2(n5072), .A3(n4495), .ZN(n4930) );
  NAND2_X1 U6268 ( .A1(n4932), .A2(n4511), .ZN(n5071) );
  NAND3_X1 U6269 ( .A1(n5196), .A2(n4938), .A3(n5128), .ZN(n5269) );
  NAND2_X1 U6270 ( .A1(n5167), .A2(n5928), .ZN(n5148) );
  NAND3_X1 U6271 ( .A1(n5381), .A2(n10021), .A3(n9401), .ZN(n4943) );
  NAND2_X1 U6272 ( .A1(n4944), .A2(n8154), .ZN(n4945) );
  INV_X1 U6273 ( .A(n8153), .ZN(n4944) );
  NAND2_X1 U6274 ( .A1(n9647), .A2(n4485), .ZN(n4946) );
  NAND2_X1 U6275 ( .A1(n4946), .A2(n4945), .ZN(n9595) );
  NAND2_X1 U6276 ( .A1(n4950), .A2(n4949), .ZN(n9689) );
  NAND2_X1 U6277 ( .A1(n7578), .A2(n4951), .ZN(n7618) );
  NAND3_X1 U6278 ( .A1(n5149), .A2(n5168), .A3(n4952), .ZN(n5183) );
  NAND4_X1 U6279 ( .A1(n5149), .A2(n5168), .A3(n5125), .A4(n4952), .ZN(n5194)
         );
  INV_X1 U6280 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6281 ( .A1(n9560), .A2(n4956), .ZN(n9550) );
  AND2_X1 U6282 ( .A1(n5363), .A2(n4957), .ZN(n5390) );
  NAND2_X1 U6283 ( .A1(n5363), .A2(n5410), .ZN(n5383) );
  NAND2_X1 U6284 ( .A1(n6332), .A2(n4488), .ZN(n6339) );
  NAND3_X1 U6285 ( .A1(n4983), .A2(n4986), .A3(n5917), .ZN(n6742) );
  AND2_X1 U6286 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  INV_X1 U6287 ( .A(n5906), .ZN(n4985) );
  NAND2_X1 U6288 ( .A1(n6139), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6289 ( .A1(n8330), .A2(n8258), .ZN(n4988) );
  NAND2_X1 U6290 ( .A1(n8207), .A2(n8105), .ZN(n8108) );
  NAND2_X1 U6291 ( .A1(n5914), .A2(n5898), .ZN(n5900) );
  NAND2_X1 U6292 ( .A1(n5925), .A2(n4990), .ZN(n5950) );
  NAND2_X2 U6293 ( .A1(n5907), .A2(n5908), .ZN(n6127) );
  NAND3_X1 U6294 ( .A1(n5907), .A2(n5908), .A3(P2_REG3_REG_2__SCAN_IN), .ZN(
        n5935) );
  NAND3_X1 U6295 ( .A1(n5907), .A2(n5908), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n5919) );
  XNOR2_X1 U6296 ( .A(n6758), .B(n6997), .ZN(n6754) );
  OAI22_X1 U6297 ( .A1(n5953), .A2(n6404), .B1(n6517), .B2(n6385), .ZN(n4995)
         );
  NOR2_X2 U6298 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6908) );
  INV_X1 U6299 ( .A(n9946), .ZN(n8144) );
  INV_X1 U6300 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5011) );
  AND2_X1 U6301 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U6302 ( .A1(n7741), .A2(n7742), .ZN(n7746) );
  XNOR2_X1 U6303 ( .A(n5331), .B(n5332), .ZN(n8871) );
  OAI21_X1 U6304 ( .B1(n6746), .B2(n5917), .A(n6742), .ZN(n8239) );
  AND2_X1 U6305 ( .A1(n7439), .A2(n7302), .ZN(n7305) );
  XNOR2_X1 U6306 ( .A(n5324), .B(n5323), .ZN(n8116) );
  NAND2_X1 U6307 ( .A1(n5324), .A2(n5323), .ZN(n5117) );
  XOR2_X1 U6308 ( .A(n9546), .B(n9541), .Z(n9948) );
  NAND2_X1 U6309 ( .A1(n5726), .A2(n5725), .ZN(n5877) );
  NAND2_X1 U6310 ( .A1(n5900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U6311 ( .A1(n9686), .A2(n8125), .ZN(n9674) );
  MUX2_X2 U6312 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n6380), .S(n8772), .Z(n6381)
         );
  MUX2_X2 U6313 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n6380), .S(n10338), .Z(n6369) );
  XNOR2_X1 U6314 ( .A(n9556), .B(n9557), .ZN(n9952) );
  NAND2_X2 U6315 ( .A1(n6280), .A2(n6689), .ZN(n6688) );
  NAND2_X1 U6316 ( .A1(n5393), .A2(n5392), .ZN(n8117) );
  OR2_X1 U6317 ( .A1(n5390), .A2(n5228), .ZN(n5391) );
  OAI21_X2 U6318 ( .B1(n7059), .B2(n7058), .A(n7056), .ZN(n7085) );
  INV_X1 U6319 ( .A(n8262), .ZN(n8265) );
  OR2_X1 U6320 ( .A1(n6777), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U6321 ( .A1(n5468), .A2(n8056), .ZN(n6974) );
  INV_X1 U6322 ( .A(n5468), .ZN(n5469) );
  XNOR2_X1 U6323 ( .A(n6741), .B(n6746), .ZN(n6743) );
  INV_X1 U6324 ( .A(n6754), .ZN(n6751) );
  OAI22_X1 U6325 ( .A1(n8525), .A2(n6311), .B1(n8258), .B2(n6310), .ZN(n8516)
         );
  NOR2_X1 U6326 ( .A1(n8150), .A2(n9645), .ZN(n4996) );
  AND2_X1 U6327 ( .A1(n10269), .A2(n10274), .ZN(n4997) );
  AND2_X1 U6328 ( .A1(n7290), .A2(n7289), .ZN(n4998) );
  NOR2_X1 U6329 ( .A1(n9528), .A2(n10275), .ZN(n4999) );
  INV_X1 U6330 ( .A(n6318), .ZN(n6414) );
  AND2_X1 U6331 ( .A1(n8214), .A2(n8336), .ZN(n5004) );
  AND2_X2 U6332 ( .A1(n5420), .A2(n6956), .ZN(n10289) );
  AND4_X1 U6333 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n9713)
         );
  INV_X1 U6334 ( .A(n8037), .ZN(n8038) );
  AND2_X1 U6335 ( .A1(n8803), .A2(n8561), .ZN(n5005) );
  INV_X1 U6336 ( .A(n9548), .ZN(n8146) );
  NAND2_X1 U6337 ( .A1(n6957), .A2(n10205), .ZN(n10208) );
  INV_X1 U6338 ( .A(n10208), .ZN(n10220) );
  INV_X1 U6339 ( .A(n10208), .ZN(n9728) );
  INV_X2 U6340 ( .A(n5929), .ZN(n6998) );
  INV_X1 U6341 ( .A(n7275), .ZN(n10210) );
  AND2_X1 U6342 ( .A1(n5861), .A2(n9380), .ZN(n5006) );
  INV_X1 U6343 ( .A(n9932), .ZN(n9778) );
  AND2_X1 U6344 ( .A1(n10235), .A2(n7281), .ZN(n9932) );
  AND2_X2 U6345 ( .A1(n5420), .A2(n6670), .ZN(n10296) );
  INV_X1 U6346 ( .A(n7999), .ZN(n6030) );
  MUX2_X1 U6347 ( .A(n7928), .B(n7927), .S(n7973), .Z(n7939) );
  NAND2_X1 U6348 ( .A1(n8154), .A2(n5441), .ZN(n5772) );
  INV_X1 U6349 ( .A(n5772), .ZN(n5779) );
  INV_X1 U6350 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U6351 ( .A1(n8034), .A2(n8037), .ZN(n6735) );
  INV_X1 U6352 ( .A(n8699), .ZN(n7991) );
  NAND2_X1 U6353 ( .A1(n5833), .A2(n5864), .ZN(n5865) );
  INV_X1 U6354 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5888) );
  NOR2_X1 U6355 ( .A1(n9213), .A2(n9346), .ZN(n7768) );
  INV_X1 U6356 ( .A(n7783), .ZN(n7784) );
  INV_X1 U6357 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5989) );
  INV_X1 U6358 ( .A(n6204), .ZN(n6193) );
  INV_X1 U6359 ( .A(n6063), .ZN(n6062) );
  AND2_X1 U6360 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND2_X1 U6361 ( .A1(n7782), .A2(n7784), .ZN(n7785) );
  INV_X1 U6362 ( .A(n9546), .ZN(n8159) );
  INV_X1 U6363 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5131) );
  INV_X1 U6364 ( .A(n5267), .ZN(n5074) );
  INV_X1 U6365 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6366 ( .A1(n5928), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6367 ( .A1(n5990), .A2(n5989), .ZN(n6013) );
  OR2_X1 U6368 ( .A1(n5953), .A2(n6394), .ZN(n5938) );
  OR2_X1 U6369 ( .A1(n8073), .A2(n8686), .ZN(n8074) );
  INV_X1 U6370 ( .A(n4423), .ZN(n6263) );
  OR2_X1 U6371 ( .A1(n6216), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6228) );
  OR2_X1 U6372 ( .A1(n6084), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U6373 ( .A1(n6036), .A2(n6035), .ZN(n6051) );
  INV_X1 U6374 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U6375 ( .B1(n7087), .B2(n7872), .A(n7864), .ZN(n7395) );
  INV_X1 U6376 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6150) );
  INV_X1 U6377 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6106) );
  NOR2_X1 U6378 ( .A1(n5580), .A2(n5579), .ZN(n5593) );
  AND2_X1 U6379 ( .A1(n5552), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5554) );
  AOI22_X1 U6380 ( .A1(n5469), .A2(n7696), .B1(n6777), .B2(n4419), .ZN(n6778)
         );
  INV_X1 U6381 ( .A(n7131), .ZN(n7132) );
  NOR2_X1 U6382 ( .A1(n5537), .A2(n5536), .ZN(n5552) );
  NOR2_X1 U6383 ( .A1(n9515), .A2(n9520), .ZN(n5353) );
  NAND2_X1 U6384 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  OR2_X1 U6385 ( .A1(n5143), .A2(n7636), .ZN(n5317) );
  INV_X1 U6386 ( .A(n9644), .ZN(n9646) );
  INV_X1 U6387 ( .A(n9756), .ZN(n5850) );
  INV_X1 U6388 ( .A(n5282), .ZN(n5084) );
  NAND2_X1 U6389 ( .A1(n5061), .A2(SI_12_), .ZN(n5064) );
  INV_X1 U6390 ( .A(n8093), .ZN(n8283) );
  NAND2_X1 U6391 ( .A1(n5969), .A2(n5968), .ZN(n5976) );
  OR2_X1 U6392 ( .A1(P2_U3150), .A2(n6416), .ZN(n8441) );
  OR2_X1 U6393 ( .A1(n6238), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6250) );
  INV_X1 U6394 ( .A(n8623), .ZN(n6149) );
  INV_X1 U6395 ( .A(n8357), .ZN(n8672) );
  AND2_X1 U6396 ( .A1(n6375), .A2(n6346), .ZN(n6371) );
  INV_X1 U6397 ( .A(n8016), .ZN(n8695) );
  NAND2_X1 U6398 ( .A1(n6731), .A2(n7977), .ZN(n8671) );
  INV_X1 U6399 ( .A(n8690), .ZN(n8668) );
  NOR2_X1 U6400 ( .A1(n5626), .A2(n9221), .ZN(n5625) );
  OR2_X1 U6401 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  NAND2_X1 U6402 ( .A1(n7130), .A2(n7132), .ZN(n7133) );
  XNOR2_X1 U6403 ( .A(n7121), .B(n7798), .ZN(n7130) );
  NAND2_X1 U6404 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  INV_X1 U6405 ( .A(n9357), .ZN(n9370) );
  NOR2_X1 U6406 ( .A1(n6675), .A2(n6952), .ZN(n6784) );
  OR2_X1 U6407 ( .A1(n6648), .A2(n6647), .ZN(n10152) );
  XNOR2_X1 U6408 ( .A(n5353), .B(n9514), .ZN(n5368) );
  NAND2_X1 U6409 ( .A1(n6958), .A2(n6959), .ZN(n6960) );
  OR2_X1 U6410 ( .A1(n10004), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6411 ( .A1(n5143), .A2(n8047), .ZN(n5321) );
  NAND2_X1 U6412 ( .A1(n9701), .A2(n9871), .ZN(n8125) );
  INV_X1 U6413 ( .A(n10280), .ZN(n10268) );
  AND2_X1 U6414 ( .A1(n6427), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6388) );
  AND2_X1 U6415 ( .A1(n5107), .A2(n5106), .ZN(n5315) );
  AND2_X1 U6416 ( .A1(n5069), .A2(n5068), .ZN(n5242) );
  XNOR2_X1 U6417 ( .A(n5053), .B(SI_9_), .ZN(n5208) );
  AND2_X1 U6418 ( .A1(n5039), .A2(n5038), .ZN(n5177) );
  INV_X1 U6419 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  OR2_X1 U6420 ( .A1(n5976), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5991) );
  OR2_X1 U6421 ( .A1(n7669), .A2(n6127), .ZN(n7684) );
  AND4_X1 U6422 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n7599)
         );
  INV_X1 U6423 ( .A(n8486), .ZN(n8450) );
  INV_X1 U6424 ( .A(n8666), .ZN(n8696) );
  INV_X1 U6425 ( .A(n8683), .ZN(n10311) );
  INV_X1 U6426 ( .A(n8742), .ZN(n8755) );
  AND2_X1 U6427 ( .A1(n7998), .A2(n7997), .ZN(n8604) );
  INV_X1 U6428 ( .A(n6941), .ZN(n8760) );
  OR2_X1 U6429 ( .A1(n6582), .A2(n6366), .ZN(n6367) );
  INV_X1 U6430 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5959) );
  XNOR2_X1 U6431 ( .A(n7130), .B(n7131), .ZN(n7125) );
  NAND2_X1 U6432 ( .A1(n7094), .A2(n7492), .ZN(n9361) );
  INV_X1 U6433 ( .A(n7492), .ZN(n5878) );
  AND4_X1 U6434 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n9548)
         );
  AND4_X1 U6435 ( .A1(n5631), .A2(n5630), .A3(n5629), .A4(n5628), .ZN(n9662)
         );
  INV_X1 U6436 ( .A(n10121), .ZN(n10171) );
  AND2_X1 U6437 ( .A1(n9408), .A2(n6842), .ZN(n9929) );
  INV_X1 U6438 ( .A(n10296), .ZN(n5414) );
  AOI22_X1 U6439 ( .A1(n9757), .A2(n9756), .B1(n8122), .B2(n10276), .ZN(n9735)
         );
  NAND2_X1 U6440 ( .A1(n6834), .A2(n6833), .ZN(n9927) );
  INV_X1 U6441 ( .A(n6670), .ZN(n6956) );
  AND2_X1 U6442 ( .A1(n5198), .A2(n5197), .ZN(n10045) );
  INV_X1 U6443 ( .A(n8785), .ZN(n8214) );
  INV_X1 U6444 ( .A(n8332), .ZN(n8346) );
  NAND2_X1 U6445 ( .A1(n6256), .A2(n6255), .ZN(n8517) );
  INV_X1 U6446 ( .A(n8285), .ZN(n8561) );
  OR2_X1 U6447 ( .A1(n6587), .A2(n6387), .ZN(n8368) );
  OR2_X1 U6448 ( .A1(n8368), .A2(n8040), .ZN(n8494) );
  OR2_X1 U6449 ( .A1(n6433), .A2(n8489), .ZN(n8501) );
  INV_X1 U6450 ( .A(n7305), .ZN(n7487) );
  AND2_X1 U6451 ( .A1(n6570), .A2(n8683), .ZN(n10310) );
  NAND2_X1 U6452 ( .A1(n8678), .A2(n6792), .ZN(n8666) );
  XOR2_X1 U6453 ( .A(n8505), .B(n8506), .Z(n8782) );
  OR2_X1 U6454 ( .A1(n10341), .A2(n8764), .ZN(n8835) );
  OR2_X1 U6455 ( .A1(n8741), .A2(n8740), .ZN(n8833) );
  INV_X2 U6456 ( .A(n10341), .ZN(n10338) );
  AND2_X1 U6457 ( .A1(n6594), .A2(n6344), .ZN(n6450) );
  AND2_X1 U6458 ( .A1(n6586), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6456) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9083) );
  AND2_X1 U6460 ( .A1(n6430), .A2(n6480), .ZN(n10138) );
  INV_X1 U6461 ( .A(n9701), .ZN(n9882) );
  INV_X1 U6462 ( .A(n9352), .ZN(n9378) );
  INV_X1 U6463 ( .A(n9841), .ZN(n9857) );
  INV_X1 U6464 ( .A(n9912), .ZN(n9893) );
  INV_X1 U6465 ( .A(n10138), .ZN(n10180) );
  OR2_X1 U6466 ( .A1(n10220), .A2(n6971), .ZN(n10198) );
  INV_X1 U6467 ( .A(n10216), .ZN(n9753) );
  INV_X1 U6468 ( .A(n9816), .ZN(n9909) );
  INV_X1 U6469 ( .A(n9943), .ZN(n9996) );
  INV_X1 U6470 ( .A(n9955), .ZN(n10000) );
  INV_X1 U6471 ( .A(n10289), .ZN(n10287) );
  INV_X1 U6472 ( .A(n10231), .ZN(n10232) );
  AND2_X1 U6473 ( .A1(n10005), .A2(n10004), .ZN(n10231) );
  INV_X1 U6474 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10349) );
  XNOR2_X1 U6475 ( .A(n5015), .B(n5014), .ZN(n5137) );
  NAND2_X1 U6476 ( .A1(n5137), .A2(SI_1_), .ZN(n5141) );
  INV_X1 U6477 ( .A(n5014), .ZN(n5016) );
  NAND2_X1 U6478 ( .A1(n5016), .A2(n5015), .ZN(n5017) );
  NAND2_X1 U6479 ( .A1(n5141), .A2(n5017), .ZN(n5145) );
  MUX2_X1 U6480 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6392), .Z(n5020) );
  INV_X1 U6481 ( .A(n5020), .ZN(n5019) );
  INV_X1 U6482 ( .A(SI_2_), .ZN(n5018) );
  NAND2_X1 U6483 ( .A1(n5019), .A2(n5018), .ZN(n5021) );
  NAND2_X1 U6484 ( .A1(n5020), .A2(SI_2_), .ZN(n5022) );
  AND2_X2 U6485 ( .A1(n5021), .A2(n5022), .ZN(n5144) );
  NAND2_X1 U6486 ( .A1(n5145), .A2(n5144), .ZN(n5147) );
  NAND2_X1 U6487 ( .A1(n5147), .A2(n5022), .ZN(n5155) );
  NAND2_X1 U6488 ( .A1(n5025), .A2(SI_3_), .ZN(n5029) );
  INV_X1 U6489 ( .A(SI_3_), .ZN(n5026) );
  NAND2_X1 U6490 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  NAND2_X1 U6491 ( .A1(n5157), .A2(n5029), .ZN(n5166) );
  MUX2_X1 U6492 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5928), .Z(n5030) );
  NAND2_X1 U6493 ( .A1(n5030), .A2(SI_4_), .ZN(n5034) );
  INV_X1 U6494 ( .A(n5030), .ZN(n5032) );
  INV_X1 U6495 ( .A(SI_4_), .ZN(n5031) );
  NAND2_X1 U6496 ( .A1(n5032), .A2(n5031), .ZN(n5033) );
  NAND2_X1 U6497 ( .A1(n5166), .A2(n5165), .ZN(n5035) );
  NAND2_X1 U6498 ( .A1(n5035), .A2(n5034), .ZN(n5178) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5928), .Z(n5036) );
  NAND2_X1 U6500 ( .A1(n5036), .A2(SI_5_), .ZN(n5039) );
  INV_X1 U6501 ( .A(n5036), .ZN(n5037) );
  INV_X1 U6502 ( .A(SI_5_), .ZN(n9149) );
  NAND2_X1 U6503 ( .A1(n5037), .A2(n9149), .ZN(n5038) );
  MUX2_X1 U6504 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5928), .Z(n5040) );
  NAND2_X1 U6505 ( .A1(n5040), .A2(SI_6_), .ZN(n5044) );
  INV_X1 U6506 ( .A(n5040), .ZN(n5042) );
  INV_X1 U6507 ( .A(SI_6_), .ZN(n5041) );
  NAND2_X1 U6508 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5928), .Z(n5045) );
  NAND2_X1 U6510 ( .A1(n5045), .A2(SI_7_), .ZN(n5048) );
  INV_X1 U6511 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6512 ( .A1(n5046), .A2(n9071), .ZN(n5047) );
  NAND2_X1 U6513 ( .A1(n5191), .A2(n5190), .ZN(n5193) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5928), .Z(n5049) );
  INV_X1 U6515 ( .A(n5049), .ZN(n5051) );
  INV_X1 U6516 ( .A(SI_8_), .ZN(n5050) );
  NAND2_X1 U6517 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  MUX2_X1 U6518 ( .A(n9083), .B(n6411), .S(n5928), .Z(n5053) );
  INV_X1 U6519 ( .A(n5053), .ZN(n5054) );
  MUX2_X1 U6520 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5928), .Z(n5055) );
  NAND2_X1 U6521 ( .A1(n5055), .A2(SI_10_), .ZN(n5059) );
  INV_X1 U6522 ( .A(n5055), .ZN(n5057) );
  INV_X1 U6523 ( .A(SI_10_), .ZN(n5056) );
  NAND2_X1 U6524 ( .A1(n5057), .A2(n5056), .ZN(n5058) );
  MUX2_X1 U6525 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5928), .Z(n5060) );
  MUX2_X1 U6526 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5928), .Z(n5061) );
  INV_X1 U6527 ( .A(n5061), .ZN(n5062) );
  INV_X1 U6528 ( .A(SI_12_), .ZN(n8984) );
  NAND2_X1 U6529 ( .A1(n5062), .A2(n8984), .ZN(n5063) );
  MUX2_X1 U6530 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5928), .Z(n5065) );
  INV_X1 U6531 ( .A(n5065), .ZN(n5067) );
  INV_X1 U6532 ( .A(SI_13_), .ZN(n5066) );
  NAND2_X1 U6533 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  MUX2_X1 U6534 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5928), .Z(n5253) );
  MUX2_X1 U6535 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5928), .Z(n5260) );
  INV_X1 U6536 ( .A(n5260), .ZN(n5070) );
  NAND2_X1 U6537 ( .A1(n5071), .A2(n5070), .ZN(n5073) );
  INV_X1 U6538 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6727) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U6540 ( .A(n6727), .B(n6728), .S(n5928), .Z(n5267) );
  NAND2_X1 U6541 ( .A1(n5074), .A2(SI_16_), .ZN(n5075) );
  INV_X1 U6542 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6857) );
  MUX2_X1 U6543 ( .A(n6857), .B(n8974), .S(n5928), .Z(n5077) );
  INV_X1 U6544 ( .A(SI_17_), .ZN(n5076) );
  NAND2_X1 U6545 ( .A1(n5077), .A2(n5076), .ZN(n5080) );
  INV_X1 U6546 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6547 ( .A1(n5078), .A2(SI_17_), .ZN(n5079) );
  NAND2_X1 U6548 ( .A1(n5080), .A2(n5079), .ZN(n5276) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7068) );
  INV_X1 U6550 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7030) );
  MUX2_X1 U6551 ( .A(n7068), .B(n7030), .S(n5928), .Z(n5081) );
  XNOR2_X1 U6552 ( .A(n5081), .B(SI_18_), .ZN(n5282) );
  INV_X1 U6553 ( .A(n5081), .ZN(n5082) );
  NAND2_X1 U6554 ( .A1(n5082), .A2(SI_18_), .ZN(n5083) );
  INV_X1 U6555 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7160) );
  INV_X1 U6556 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7161) );
  MUX2_X1 U6557 ( .A(n7160), .B(n7161), .S(n5928), .Z(n5086) );
  INV_X1 U6558 ( .A(SI_19_), .ZN(n5085) );
  NAND2_X1 U6559 ( .A1(n5086), .A2(n5085), .ZN(n5089) );
  INV_X1 U6560 ( .A(n5086), .ZN(n5087) );
  NAND2_X1 U6561 ( .A1(n5087), .A2(SI_19_), .ZN(n5088) );
  NAND2_X1 U6562 ( .A1(n5089), .A2(n5088), .ZN(n5287) );
  INV_X1 U6563 ( .A(SI_20_), .ZN(n5296) );
  MUX2_X1 U6564 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5928), .Z(n5297) );
  INV_X1 U6565 ( .A(n5297), .ZN(n5090) );
  INV_X1 U6566 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7327) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7333) );
  MUX2_X1 U6568 ( .A(n7327), .B(n7333), .S(n5928), .Z(n5302) );
  INV_X1 U6569 ( .A(n5302), .ZN(n5091) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7540) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7537) );
  MUX2_X1 U6572 ( .A(n7540), .B(n7537), .S(n5928), .Z(n5093) );
  INV_X1 U6573 ( .A(SI_22_), .ZN(n5092) );
  NAND2_X1 U6574 ( .A1(n5093), .A2(n5092), .ZN(n5096) );
  INV_X1 U6575 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6576 ( .A1(n5094), .A2(SI_22_), .ZN(n5095) );
  NAND2_X1 U6577 ( .A1(n5096), .A2(n5095), .ZN(n5307) );
  INV_X1 U6578 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7498) );
  INV_X1 U6579 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7494) );
  MUX2_X1 U6580 ( .A(n7498), .B(n7494), .S(n5928), .Z(n5098) );
  INV_X1 U6581 ( .A(SI_23_), .ZN(n5097) );
  NAND2_X1 U6582 ( .A1(n5098), .A2(n5097), .ZN(n5101) );
  INV_X1 U6583 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6584 ( .A1(n5099), .A2(SI_23_), .ZN(n5100) );
  NAND2_X1 U6585 ( .A1(n5312), .A2(n5311), .ZN(n5102) );
  NAND2_X1 U6586 ( .A1(n5102), .A2(n5101), .ZN(n5316) );
  INV_X1 U6587 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7650) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7636) );
  MUX2_X1 U6589 ( .A(n7650), .B(n7636), .S(n5928), .Z(n5104) );
  INV_X1 U6590 ( .A(SI_24_), .ZN(n5103) );
  NAND2_X1 U6591 ( .A1(n5104), .A2(n5103), .ZN(n5107) );
  INV_X1 U6592 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6593 ( .A1(n5105), .A2(SI_24_), .ZN(n5106) );
  INV_X1 U6594 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7648) );
  INV_X1 U6595 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8047) );
  MUX2_X1 U6596 ( .A(n7648), .B(n8047), .S(n5928), .Z(n5108) );
  INV_X1 U6597 ( .A(SI_25_), .ZN(n9046) );
  NAND2_X1 U6598 ( .A1(n5108), .A2(n9046), .ZN(n5111) );
  INV_X1 U6599 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6600 ( .A1(n5109), .A2(SI_25_), .ZN(n5110) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9007) );
  INV_X1 U6602 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9074) );
  INV_X1 U6603 ( .A(SI_26_), .ZN(n5112) );
  NAND2_X1 U6604 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  INV_X1 U6605 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6606 ( .A1(n5114), .A2(SI_26_), .ZN(n5115) );
  INV_X1 U6607 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6235) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10019) );
  MUX2_X1 U6609 ( .A(n6235), .B(n10019), .S(n5928), .Z(n5119) );
  INV_X1 U6610 ( .A(SI_27_), .ZN(n5118) );
  NAND2_X1 U6611 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U6612 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6613 ( .A1(n5120), .A2(SI_27_), .ZN(n5121) );
  INV_X1 U6614 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6245) );
  INV_X1 U6615 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10016) );
  XNOR2_X1 U6616 ( .A(n5124), .B(SI_28_), .ZN(n5332) );
  INV_X1 U6617 ( .A(SI_28_), .ZN(n5123) );
  INV_X1 U6618 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8193) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8868) );
  MUX2_X1 U6620 ( .A(n8193), .B(n8868), .S(n6392), .Z(n5335) );
  NOR2_X1 U6621 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5354) );
  NOR2_X1 U6622 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5130) );
  NAND2_X1 U6623 ( .A1(n5387), .A2(n5385), .ZN(n5132) );
  INV_X1 U6624 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6625 ( .A1(n8192), .A2(n5352), .ZN(n5136) );
  OR2_X1 U6626 ( .A1(n5143), .A2(n8193), .ZN(n5135) );
  INV_X1 U6627 ( .A(n5137), .ZN(n5139) );
  INV_X1 U6628 ( .A(SI_1_), .ZN(n5138) );
  NAND2_X1 U6629 ( .A1(n5139), .A2(n5138), .ZN(n5140) );
  AND2_X1 U6630 ( .A1(n5141), .A2(n5140), .ZN(n5927) );
  INV_X1 U6631 ( .A(n5927), .ZN(n6393) );
  INV_X1 U6632 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9038) );
  INV_X1 U6633 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U6634 ( .A1(n5928), .A2(SI_0_), .ZN(n5142) );
  XNOR2_X1 U6635 ( .A(n5142), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U6636 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10022), .S(n5167), .Z(n10236)
         );
  INV_X1 U6637 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6395) );
  OR2_X1 U6638 ( .A1(n5143), .A2(n6395), .ZN(n5153) );
  OR2_X1 U6639 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  NAND2_X1 U6640 ( .A1(n5147), .A2(n5146), .ZN(n6394) );
  OR2_X1 U6641 ( .A1(n5148), .A2(n6394), .ZN(n5152) );
  OR2_X1 U6642 ( .A1(n5149), .A2(n5228), .ZN(n5170) );
  INV_X1 U6643 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6644 ( .A1(n5170), .A2(n5150), .ZN(n5158) );
  OAI21_X1 U6645 ( .B1(n5170), .B2(n5150), .A(n5158), .ZN(n9414) );
  OR2_X1 U6646 ( .A1(n6429), .A2(n9414), .ZN(n5151) );
  INV_X1 U6647 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6405) );
  OR2_X1 U6648 ( .A1(n5143), .A2(n6405), .ZN(n5163) );
  OR2_X1 U6649 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6650 ( .A1(n5157), .A2(n5156), .ZN(n6404) );
  OR2_X1 U6651 ( .A1(n5148), .A2(n6404), .ZN(n5162) );
  NAND2_X1 U6652 ( .A1(n5158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5160) );
  INV_X1 U6653 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6654 ( .A(n5160), .B(n5159), .ZN(n9425) );
  OR2_X1 U6655 ( .A1(n6429), .A2(n9425), .ZN(n5161) );
  NAND2_X1 U6656 ( .A1(n6986), .A2(n7103), .ZN(n7270) );
  INV_X1 U6657 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5164) );
  OR2_X1 U6658 ( .A1(n5143), .A2(n5164), .ZN(n5173) );
  XNOR2_X1 U6659 ( .A(n5166), .B(n5165), .ZN(n6396) );
  OR2_X1 U6660 ( .A1(n5148), .A2(n6396), .ZN(n5172) );
  OR2_X1 U6661 ( .A1(n5168), .A2(n5228), .ZN(n5169) );
  NAND2_X1 U6662 ( .A1(n5170), .A2(n5169), .ZN(n5175) );
  XNOR2_X1 U6663 ( .A(n5175), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9442) );
  OR2_X1 U6664 ( .A1(n6429), .A2(n9442), .ZN(n5171) );
  OAI21_X1 U6665 ( .B1(n5175), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5176) );
  XNOR2_X1 U6666 ( .A(n5176), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10091) );
  INV_X1 U6667 ( .A(n10091), .ZN(n6398) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6400) );
  OR2_X1 U6669 ( .A1(n5143), .A2(n6400), .ZN(n5182) );
  OR2_X1 U6670 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6671 ( .A1(n5180), .A2(n5179), .ZN(n6399) );
  OR2_X1 U6672 ( .A1(n5148), .A2(n6399), .ZN(n5181) );
  NAND2_X1 U6673 ( .A1(n5183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6674 ( .A(n5184), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6633) );
  INV_X1 U6675 ( .A(n6633), .ZN(n10105) );
  OR2_X1 U6676 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6677 ( .A1(n5188), .A2(n5187), .ZN(n6403) );
  INV_X1 U6678 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6402) );
  OR2_X1 U6679 ( .A1(n5143), .A2(n6402), .ZN(n5189) );
  OR2_X1 U6680 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6681 ( .A1(n5193), .A2(n5192), .ZN(n6407) );
  OR2_X1 U6682 ( .A1(n5148), .A2(n6407), .ZN(n5201) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6406) );
  OR2_X1 U6684 ( .A1(n5143), .A2(n6406), .ZN(n5200) );
  NAND2_X1 U6685 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5195) );
  MUX2_X1 U6686 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5195), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n5198) );
  INV_X1 U6687 ( .A(n5196), .ZN(n5197) );
  INV_X1 U6688 ( .A(n10045), .ZN(n6613) );
  OR2_X1 U6689 ( .A1(n6429), .A2(n6613), .ZN(n5199) );
  NAND2_X1 U6690 ( .A1(n7477), .A2(n7547), .ZN(n9931) );
  OR2_X1 U6691 ( .A1(n5196), .A2(n5228), .ZN(n5203) );
  INV_X1 U6692 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6693 ( .A1(n5203), .A2(n5202), .ZN(n5210) );
  OAI21_X1 U6694 ( .B1(n5203), .B2(n5202), .A(n5210), .ZN(n10050) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9131) );
  OR2_X1 U6696 ( .A1(n5143), .A2(n9131), .ZN(n5206) );
  XNOR2_X1 U6697 ( .A(n5209), .B(n5208), .ZN(n6409) );
  NAND2_X1 U6698 ( .A1(n6409), .A2(n5352), .ZN(n5213) );
  NAND2_X1 U6699 ( .A1(n5210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U6700 ( .A(n5211), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U6701 ( .A1(n5292), .A2(n6640), .ZN(n5212) );
  INV_X1 U6702 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6703 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6704 ( .A1(n5218), .A2(n5217), .ZN(n9172) );
  OR2_X1 U6705 ( .A1(n9172), .A2(n5148), .ZN(n5222) );
  AND2_X1 U6706 ( .A1(n5196), .A2(n5219), .ZN(n5226) );
  OR2_X1 U6707 ( .A1(n5226), .A2(n5228), .ZN(n5220) );
  XNOR2_X1 U6708 ( .A(n5220), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U6709 ( .A1(n5293), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5292), .B2(
        n6642), .ZN(n5221) );
  XNOR2_X1 U6710 ( .A(n5224), .B(n5223), .ZN(n6424) );
  NAND2_X1 U6711 ( .A1(n6424), .A2(n5352), .ZN(n5234) );
  AND2_X1 U6712 ( .A1(n5226), .A2(n5225), .ZN(n5231) );
  NOR2_X1 U6713 ( .A1(n5231), .A2(n5228), .ZN(n5227) );
  MUX2_X1 U6714 ( .A(n5228), .B(n5227), .S(P1_IR_REG_11__SCAN_IN), .Z(n5229)
         );
  INV_X1 U6715 ( .A(n5229), .ZN(n5232) );
  NAND2_X1 U6716 ( .A1(n5231), .A2(n5230), .ZN(n5239) );
  AOI22_X1 U6717 ( .A1(n5293), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5292), .B2(
        n6644), .ZN(n5233) );
  NAND2_X1 U6718 ( .A1(n5236), .A2(n5235), .ZN(n5238) );
  NAND2_X1 U6719 ( .A1(n5238), .A2(n5237), .ZN(n6432) );
  OR2_X1 U6720 ( .A1(n6432), .A2(n5148), .ZN(n5241) );
  NAND2_X1 U6721 ( .A1(n5239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6722 ( .A(n5247), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U6723 ( .A1(n5293), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5292), .B2(
        n9463), .ZN(n5240) );
  OR2_X1 U6724 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  NAND2_X1 U6725 ( .A1(n5245), .A2(n5244), .ZN(n6486) );
  OR2_X1 U6726 ( .A1(n6486), .A2(n5148), .ZN(n5251) );
  INV_X1 U6727 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6728 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  NAND2_X1 U6729 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6730 ( .A(n5249), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U6731 ( .A1(n5293), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5292), .B2(
        n10134), .ZN(n5250) );
  XNOR2_X1 U6732 ( .A(n5253), .B(SI_14_), .ZN(n5254) );
  XNOR2_X1 U6733 ( .A(n5252), .B(n5254), .ZN(n6533) );
  NAND2_X1 U6734 ( .A1(n6533), .A2(n5352), .ZN(n5259) );
  NAND2_X1 U6735 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  MUX2_X1 U6736 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5256), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5257) );
  AND2_X1 U6737 ( .A1(n5257), .A2(n4498), .ZN(n10148) );
  AOI22_X1 U6738 ( .A1(n5293), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5292), .B2(
        n10148), .ZN(n5258) );
  XNOR2_X1 U6739 ( .A(n5260), .B(SI_15_), .ZN(n5261) );
  XNOR2_X1 U6740 ( .A(n5262), .B(n5261), .ZN(n6657) );
  NAND2_X1 U6741 ( .A1(n6657), .A2(n5352), .ZN(n5265) );
  NAND2_X1 U6742 ( .A1(n4498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6743 ( .A(n5263), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U6744 ( .A1(n5293), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5292), .B2(
        n10161), .ZN(n5264) );
  XNOR2_X1 U6745 ( .A(n5267), .B(SI_16_), .ZN(n5268) );
  XNOR2_X1 U6746 ( .A(n5266), .B(n5268), .ZN(n6726) );
  NAND2_X1 U6747 ( .A1(n6726), .A2(n5352), .ZN(n5275) );
  NAND2_X1 U6748 ( .A1(n5269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5270) );
  MUX2_X1 U6749 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5270), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5271) );
  INV_X1 U6750 ( .A(n5271), .ZN(n5273) );
  NOR2_X1 U6751 ( .A1(n5273), .A2(n5272), .ZN(n9485) );
  AOI22_X1 U6752 ( .A1(n5293), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5292), .B2(
        n9485), .ZN(n5274) );
  XNOR2_X1 U6753 ( .A(n5277), .B(n5276), .ZN(n6855) );
  NAND2_X1 U6754 ( .A1(n6855), .A2(n5352), .ZN(n5281) );
  INV_X1 U6755 ( .A(n5272), .ZN(n5278) );
  NAND2_X1 U6756 ( .A1(n5278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5279) );
  XNOR2_X1 U6757 ( .A(n5279), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U6758 ( .A1(n5293), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5292), .B2(
        n10172), .ZN(n5280) );
  XNOR2_X1 U6759 ( .A(n5283), .B(n5282), .ZN(n7029) );
  NAND2_X1 U6760 ( .A1(n7029), .A2(n5352), .ZN(n5286) );
  NAND2_X1 U6761 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5357) );
  XNOR2_X1 U6762 ( .A(n5357), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U6763 ( .A1(n5293), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5292), .B2(
        n9476), .ZN(n5285) );
  XNOR2_X1 U6764 ( .A(n5288), .B(n5287), .ZN(n7159) );
  NAND2_X1 U6765 ( .A1(n7159), .A2(n5352), .ZN(n5295) );
  INV_X1 U6766 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6767 ( .A1(n5357), .A2(n5289), .ZN(n5290) );
  NAND2_X1 U6768 ( .A1(n5290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X2 U6769 ( .A(n5291), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6973) );
  AOI22_X1 U6770 ( .A1(n5293), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6973), .B2(
        n5292), .ZN(n5294) );
  NAND2_X1 U6771 ( .A1(n9677), .A2(n9874), .ZN(n9665) );
  XNOR2_X1 U6772 ( .A(n5297), .B(n5296), .ZN(n5298) );
  XNOR2_X1 U6773 ( .A(n5299), .B(n5298), .ZN(n7263) );
  NAND2_X1 U6774 ( .A1(n7263), .A2(n5352), .ZN(n5301) );
  INV_X1 U6775 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7279) );
  OR2_X1 U6776 ( .A1(n5143), .A2(n7279), .ZN(n5300) );
  XNOR2_X1 U6777 ( .A(n5302), .B(SI_21_), .ZN(n5303) );
  XNOR2_X1 U6778 ( .A(n5304), .B(n5303), .ZN(n6172) );
  NAND2_X1 U6779 ( .A1(n6172), .A2(n5352), .ZN(n5306) );
  OR2_X1 U6780 ( .A1(n5143), .A2(n7333), .ZN(n5305) );
  XNOR2_X1 U6781 ( .A(n5308), .B(n5307), .ZN(n7536) );
  NAND2_X1 U6782 ( .A1(n7536), .A2(n5352), .ZN(n5310) );
  OR2_X1 U6783 ( .A1(n5143), .A2(n7537), .ZN(n5309) );
  NAND2_X1 U6784 ( .A1(n7495), .A2(n5352), .ZN(n5314) );
  XNOR2_X1 U6785 ( .A(n5316), .B(n5315), .ZN(n7635) );
  NAND2_X1 U6786 ( .A1(n7635), .A2(n5352), .ZN(n5318) );
  NAND2_X1 U6787 ( .A1(n8116), .A2(n5352), .ZN(n5326) );
  OR2_X1 U6788 ( .A1(n5143), .A2(n9074), .ZN(n5325) );
  NAND2_X1 U6789 ( .A1(n8871), .A2(n5352), .ZN(n5334) );
  OR2_X1 U6790 ( .A1(n5143), .A2(n10016), .ZN(n5333) );
  INV_X1 U6791 ( .A(SI_29_), .ZN(n5338) );
  INV_X1 U6792 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8172) );
  INV_X1 U6793 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8115) );
  MUX2_X1 U6794 ( .A(n8172), .B(n8115), .S(n6392), .Z(n5340) );
  INV_X1 U6795 ( .A(SI_30_), .ZN(n9009) );
  NAND2_X1 U6796 ( .A1(n5340), .A2(n9009), .ZN(n5344) );
  INV_X1 U6797 ( .A(n5340), .ZN(n5341) );
  NAND2_X1 U6798 ( .A1(n5341), .A2(SI_30_), .ZN(n5342) );
  NAND2_X1 U6799 ( .A1(n5344), .A2(n5342), .ZN(n5345) );
  OR2_X1 U6800 ( .A1(n5143), .A2(n8172), .ZN(n5343) );
  INV_X1 U6801 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10010) );
  INV_X1 U6802 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5347) );
  MUX2_X1 U6803 ( .A(n10010), .B(n5347), .S(n6392), .Z(n5348) );
  XNOR2_X1 U6804 ( .A(n5348), .B(SI_31_), .ZN(n5349) );
  NOR2_X1 U6805 ( .A1(n5143), .A2(n10010), .ZN(n5351) );
  INV_X1 U6806 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6807 ( .A1(n5355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5356) );
  INV_X1 U6808 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5358) );
  INV_X1 U6809 ( .A(n5360), .ZN(n5361) );
  NAND2_X1 U6810 ( .A1(n5361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5362) );
  MUX2_X1 U6811 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5362), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n5364) );
  INV_X1 U6812 ( .A(n5363), .ZN(n5409) );
  NAND2_X1 U6813 ( .A1(n5365), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6814 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5369) );
  NAND2_X1 U6815 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  XNOR2_X2 U6816 ( .A(n5371), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5377) );
  NOR2_X1 U6817 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5372) );
  NAND2_X1 U6818 ( .A1(n5373), .A2(n5372), .ZN(n10008) );
  XNOR2_X2 U6819 ( .A(n5375), .B(n5374), .ZN(n5376) );
  NAND2_X4 U6820 ( .A1(n5377), .A2(n5428), .ZN(n5711) );
  INV_X1 U6821 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6822 ( .A1(n5708), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5379) );
  NAND2_X4 U6823 ( .A1(n5429), .A2(n5376), .ZN(n5490) );
  INV_X1 U6824 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5415) );
  OR2_X1 U6825 ( .A1(n5490), .A2(n5415), .ZN(n5378) );
  OAI211_X1 U6826 ( .C1(n5711), .C2(n5380), .A(n5379), .B(n5378), .ZN(n9380)
         );
  INV_X1 U6827 ( .A(n5381), .ZN(n9408) );
  INV_X1 U6828 ( .A(n7538), .ZN(n6832) );
  INV_X1 U6829 ( .A(n10021), .ZN(n6647) );
  NAND2_X1 U6830 ( .A1(n6647), .A2(P1_B_REG_SCAN_IN), .ZN(n5382) );
  AND2_X1 U6831 ( .A1(n10234), .A2(n5382), .ZN(n8164) );
  AND2_X1 U6832 ( .A1(n9380), .A2(n8164), .ZN(n9511) );
  NOR2_X1 U6833 ( .A1(n9510), .A2(n9511), .ZN(n5421) );
  NAND2_X1 U6834 ( .A1(n5383), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6835 ( .A1(n5388), .A2(n5387), .ZN(n5384) );
  NAND2_X1 U6836 ( .A1(n5384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6837 ( .A1(n8049), .A2(P1_B_REG_SCAN_IN), .ZN(n5389) );
  XNOR2_X1 U6838 ( .A(n5388), .B(n5387), .ZN(n7637) );
  MUX2_X1 U6839 ( .A(P1_B_REG_SCAN_IN), .B(n5389), .S(n7637), .Z(n5395) );
  MUX2_X1 U6840 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5391), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5393) );
  INV_X1 U6841 ( .A(n8117), .ZN(n5394) );
  OR2_X1 U6842 ( .A1(n10004), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6843 ( .A1(n8117), .A2(n8049), .ZN(n10006) );
  NAND2_X1 U6844 ( .A1(n5396), .A2(n10006), .ZN(n6669) );
  NAND2_X1 U6845 ( .A1(n5722), .A2(n7281), .ZN(n5880) );
  NAND2_X1 U6846 ( .A1(n6842), .A2(n5880), .ZN(n6953) );
  NAND2_X1 U6847 ( .A1(n9932), .A2(n6973), .ZN(n6679) );
  NAND3_X1 U6848 ( .A1(n6669), .A2(n6953), .A3(n6679), .ZN(n5412) );
  NOR4_X1 U6849 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5405) );
  NOR4_X1 U6850 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5404) );
  INV_X1 U6851 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10223) );
  INV_X1 U6852 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10226) );
  INV_X1 U6853 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10222) );
  INV_X1 U6854 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10230) );
  NAND4_X1 U6855 ( .A1(n10223), .A2(n10226), .A3(n10222), .A4(n10230), .ZN(
        n5402) );
  NOR4_X1 U6856 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5400) );
  NOR4_X1 U6857 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5399) );
  NOR4_X1 U6858 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5398) );
  NOR4_X1 U6859 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5397) );
  NAND4_X1 U6860 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n5401)
         );
  NOR4_X1 U6861 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        n5402), .A4(n5401), .ZN(n5403) );
  AND3_X1 U6862 ( .A1(n5405), .A2(n5404), .A3(n5403), .ZN(n5406) );
  NAND2_X1 U6863 ( .A1(n5409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U6864 ( .A(n5411), .B(n5410), .ZN(n6427) );
  NAND2_X1 U6865 ( .A1(n8117), .A2(n7637), .ZN(n10007) );
  OR2_X1 U6866 ( .A1(n5421), .A2(n5414), .ZN(n5419) );
  OR2_X1 U6867 ( .A1(n10296), .A2(n5415), .ZN(n5416) );
  INV_X1 U6868 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6869 ( .A1(n5419), .A2(n5418), .ZN(P1_U3553) );
  OR2_X1 U6870 ( .A1(n5421), .A2(n10287), .ZN(n5426) );
  INV_X1 U6871 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5422) );
  OR2_X1 U6872 ( .A1(n10289), .A2(n5422), .ZN(n5423) );
  INV_X1 U6873 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6874 ( .A1(n5426), .A2(n5425), .ZN(P1_U3521) );
  INV_X1 U6875 ( .A(n9514), .ZN(n5714) );
  INV_X1 U6876 ( .A(n9380), .ZN(n5427) );
  INV_X1 U6877 ( .A(n5869), .ZN(n5721) );
  NAND2_X1 U6878 ( .A1(n7538), .A2(n6973), .ZN(n5720) );
  NAND2_X1 U6879 ( .A1(n5695), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5435) );
  INV_X1 U6880 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9965) );
  OR2_X1 U6881 ( .A1(n5697), .A2(n9965), .ZN(n5434) );
  NAND2_X4 U6882 ( .A1(n5429), .A2(n5428), .ZN(n5698) );
  NAND2_X1 U6883 ( .A1(n5502), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5510) );
  NOR2_X1 U6884 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  NAND2_X1 U6885 ( .A1(n5511), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5521) );
  INV_X1 U6886 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5520) );
  INV_X1 U6887 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6888 ( .A1(n5554), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5561) );
  INV_X1 U6889 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5560) );
  INV_X1 U6890 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9317) );
  INV_X1 U6891 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6892 ( .A1(n5595), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5587) );
  INV_X1 U6893 ( .A(n5587), .ZN(n5614) );
  NAND2_X1 U6894 ( .A1(n5614), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6895 ( .A1(n5619), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5626) );
  INV_X1 U6896 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U6897 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n5625), .ZN(n5451) );
  INV_X1 U6898 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U6899 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5444), .ZN(n5436) );
  INV_X1 U6900 ( .A(n5436), .ZN(n5430) );
  NAND2_X1 U6901 ( .A1(n5430), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5665) );
  INV_X1 U6902 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U6903 ( .A1(n5436), .A2(n9194), .ZN(n5431) );
  NAND2_X1 U6904 ( .A1(n5665), .A2(n5431), .ZN(n9615) );
  OR2_X1 U6905 ( .A1(n5698), .A2(n9615), .ZN(n5433) );
  INV_X1 U6906 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9849) );
  OR2_X1 U6907 ( .A1(n5490), .A2(n9849), .ZN(n5432) );
  NAND2_X1 U6908 ( .A1(n9622), .A2(n9631), .ZN(n8154) );
  NAND2_X1 U6909 ( .A1(n5708), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5440) );
  INV_X1 U6910 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9638) );
  OR2_X1 U6911 ( .A1(n5711), .A2(n9638), .ZN(n5439) );
  OAI21_X1 U6912 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5444), .A(n5436), .ZN(
        n9637) );
  OR2_X1 U6913 ( .A1(n5698), .A2(n9637), .ZN(n5438) );
  INV_X1 U6914 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9855) );
  OR2_X1 U6915 ( .A1(n5490), .A2(n9855), .ZN(n5437) );
  OR2_X1 U6916 ( .A1(n9636), .A2(n9857), .ZN(n5441) );
  NAND2_X1 U6917 ( .A1(n5772), .A2(n5647), .ZN(n5443) );
  NOR2_X1 U6918 ( .A1(n9854), .A2(n9841), .ZN(n8152) );
  INV_X1 U6919 ( .A(n8152), .ZN(n9608) );
  NAND2_X1 U6920 ( .A1(n5647), .A2(n9608), .ZN(n5442) );
  NAND2_X1 U6921 ( .A1(n5442), .A2(n8154), .ZN(n5768) );
  MUX2_X1 U6922 ( .A(n5443), .B(n5768), .S(n6845), .Z(n5648) );
  NAND2_X1 U6923 ( .A1(n5695), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5450) );
  INV_X1 U6924 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9973) );
  OR2_X1 U6925 ( .A1(n5697), .A2(n9973), .ZN(n5449) );
  INV_X1 U6926 ( .A(n5451), .ZN(n5446) );
  INV_X1 U6927 ( .A(n5444), .ZN(n5445) );
  OAI21_X1 U6928 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n5446), .A(n5445), .ZN(
        n9651) );
  OR2_X1 U6929 ( .A1(n5698), .A2(n9651), .ZN(n5448) );
  INV_X1 U6930 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9862) );
  OR2_X1 U6931 ( .A1(n5490), .A2(n9862), .ZN(n5447) );
  NAND2_X1 U6932 ( .A1(n5695), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5455) );
  INV_X1 U6933 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9977) );
  OR2_X1 U6934 ( .A1(n5697), .A2(n9977), .ZN(n5454) );
  OAI21_X1 U6935 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5625), .A(n5451), .ZN(
        n9668) );
  OR2_X1 U6936 ( .A1(n5698), .A2(n9668), .ZN(n5453) );
  INV_X1 U6937 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9868) );
  OR2_X1 U6938 ( .A1(n5490), .A2(n9868), .ZN(n5452) );
  NAND4_X1 U6939 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n9870)
         );
  INV_X1 U6940 ( .A(n9870), .ZN(n9654) );
  OR2_X1 U6941 ( .A1(n9867), .A2(n9654), .ZN(n5731) );
  NAND2_X1 U6942 ( .A1(n5775), .A2(n5731), .ZN(n5819) );
  INV_X1 U6943 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6972) );
  INV_X1 U6944 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6945 ( .A1(n5479), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5459) );
  INV_X1 U6946 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5457) );
  INV_X1 U6947 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5462) );
  OR2_X1 U6948 ( .A1(n5698), .A2(n5462), .ZN(n5467) );
  INV_X1 U6949 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6477) );
  INV_X1 U6950 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6951 ( .A1(n5479), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6952 ( .A1(n6962), .A2(n6837), .ZN(n6964) );
  NAND2_X1 U6953 ( .A1(n5479), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5476) );
  INV_X1 U6954 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6939) );
  OR2_X1 U6955 ( .A1(n5698), .A2(n6939), .ZN(n5475) );
  INV_X1 U6956 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5471) );
  OR2_X1 U6957 ( .A1(n5490), .A2(n5471), .ZN(n5474) );
  INV_X1 U6958 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5472) );
  OR2_X1 U6959 ( .A1(n5711), .A2(n5472), .ZN(n5473) );
  OAI21_X1 U6960 ( .B1(n6836), .B2(n7102), .A(n6936), .ZN(n5478) );
  NAND2_X1 U6961 ( .A1(n6836), .A2(n7102), .ZN(n5477) );
  NAND2_X1 U6962 ( .A1(n5478), .A2(n5477), .ZN(n6979) );
  NAND2_X1 U6963 ( .A1(n5479), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6964 ( .A1(n5698), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5482) );
  OR2_X1 U6965 ( .A1(n5490), .A2(n6624), .ZN(n5481) );
  INV_X1 U6966 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6607) );
  OR2_X1 U6967 ( .A1(n5711), .A2(n6607), .ZN(n5480) );
  NAND4_X1 U6968 ( .A1(n5483), .A2(n5482), .A3(n5481), .A4(n5480), .ZN(n9392)
         );
  XNOR2_X1 U6969 ( .A(n9392), .B(n7103), .ZN(n6983) );
  INV_X1 U6970 ( .A(n6983), .ZN(n6980) );
  NAND2_X1 U6971 ( .A1(n6979), .A2(n6980), .ZN(n5485) );
  INV_X1 U6972 ( .A(n9392), .ZN(n8060) );
  INV_X1 U6973 ( .A(n7103), .ZN(n6989) );
  NAND2_X1 U6974 ( .A1(n8060), .A2(n6989), .ZN(n5484) );
  NAND2_X1 U6975 ( .A1(n5485), .A2(n5484), .ZN(n7267) );
  NAND2_X1 U6976 ( .A1(n5708), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5494) );
  INV_X1 U6977 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10207) );
  OR2_X1 U6978 ( .A1(n5711), .A2(n10207), .ZN(n5493) );
  INV_X1 U6979 ( .A(n5502), .ZN(n5488) );
  INV_X1 U6980 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6981 ( .A1(n7020), .A2(n5486), .ZN(n5487) );
  NAND2_X1 U6982 ( .A1(n5488), .A2(n5487), .ZN(n10206) );
  OR2_X1 U6983 ( .A1(n5698), .A2(n10206), .ZN(n5492) );
  INV_X1 U6984 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5489) );
  OR2_X1 U6985 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U6986 ( .A1(n9391), .A2(n7275), .ZN(n5790) );
  INV_X1 U6987 ( .A(n9391), .ZN(n7141) );
  NAND2_X1 U6988 ( .A1(n7141), .A2(n10210), .ZN(n5495) );
  NAND2_X1 U6989 ( .A1(n5708), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5501) );
  OR2_X1 U6990 ( .A1(n5511), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6991 ( .A1(n5521), .A2(n5496), .ZN(n7386) );
  OR2_X1 U6992 ( .A1(n5698), .A2(n7386), .ZN(n5500) );
  INV_X1 U6993 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6634) );
  OR2_X1 U6994 ( .A1(n5490), .A2(n6634), .ZN(n5499) );
  INV_X1 U6995 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5497) );
  OR2_X1 U6996 ( .A1(n5711), .A2(n5497), .ZN(n5498) );
  XNOR2_X1 U6997 ( .A(n9930), .B(n7547), .ZN(n7384) );
  INV_X1 U6998 ( .A(n7384), .ZN(n5531) );
  NAND2_X1 U6999 ( .A1(n5708), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5507) );
  INV_X1 U7000 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7080) );
  OR2_X1 U7001 ( .A1(n5711), .A2(n7080), .ZN(n5506) );
  OAI21_X1 U7002 ( .B1(n5502), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5510), .ZN(
        n7139) );
  OR2_X1 U7003 ( .A1(n5698), .A2(n7139), .ZN(n5505) );
  INV_X1 U7004 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5503) );
  OR2_X1 U7005 ( .A1(n5490), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U7006 ( .A1(n7296), .A2(n7381), .ZN(n5837) );
  NAND2_X1 U7007 ( .A1(n5708), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5517) );
  INV_X1 U7008 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5508) );
  OR2_X1 U7009 ( .A1(n5711), .A2(n5508), .ZN(n5516) );
  AND2_X1 U7010 ( .A1(n5510), .A2(n5509), .ZN(n5512) );
  OR2_X1 U7011 ( .A1(n5512), .A2(n5511), .ZN(n10193) );
  OR2_X1 U7012 ( .A1(n5698), .A2(n10193), .ZN(n5515) );
  INV_X1 U7013 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5513) );
  OR2_X1 U7014 ( .A1(n5490), .A2(n5513), .ZN(n5514) );
  NAND2_X1 U7015 ( .A1(n7323), .A2(n7483), .ZN(n5794) );
  NAND2_X1 U7016 ( .A1(n9389), .A2(n10199), .ZN(n7376) );
  INV_X1 U7017 ( .A(n7381), .ZN(n10248) );
  NAND2_X1 U7018 ( .A1(n9390), .A2(n10248), .ZN(n5792) );
  NAND3_X1 U7019 ( .A1(n7376), .A2(n5792), .A3(n5720), .ZN(n5518) );
  NOR2_X1 U7020 ( .A1(n7384), .A2(n5518), .ZN(n5519) );
  NAND2_X1 U7021 ( .A1(n5786), .A2(n5519), .ZN(n5535) );
  NAND2_X1 U7022 ( .A1(n5708), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5526) );
  INV_X1 U7023 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6637) );
  OR2_X1 U7024 ( .A1(n5490), .A2(n6637), .ZN(n5525) );
  NAND2_X1 U7025 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U7026 ( .A1(n5537), .A2(n5522), .ZN(n10181) );
  OR2_X1 U7027 ( .A1(n5698), .A2(n10181), .ZN(n5524) );
  INV_X1 U7028 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10182) );
  OR2_X1 U7029 ( .A1(n5711), .A2(n10182), .ZN(n5523) );
  NAND2_X1 U7030 ( .A1(n9388), .A2(n4418), .ZN(n7458) );
  NAND2_X1 U7031 ( .A1(n9930), .A2(n7547), .ZN(n5527) );
  AOI21_X1 U7032 ( .B1(n7376), .B2(n5792), .A(n5720), .ZN(n5528) );
  NAND2_X1 U7033 ( .A1(n5528), .A2(n5794), .ZN(n5530) );
  NAND4_X1 U7034 ( .A1(n7376), .A2(n7296), .A3(n5720), .A4(n7381), .ZN(n5529)
         );
  OAI211_X1 U7035 ( .C1(n6845), .C2(n5794), .A(n5530), .B(n5529), .ZN(n5532)
         );
  NAND2_X1 U7036 ( .A1(n5532), .A2(n5531), .ZN(n5534) );
  NAND2_X1 U7037 ( .A1(n9294), .A2(n10184), .ZN(n7459) );
  INV_X1 U7038 ( .A(n9930), .ZN(n5533) );
  INV_X1 U7039 ( .A(n7547), .ZN(n7550) );
  NAND2_X1 U7040 ( .A1(n5533), .A2(n7550), .ZN(n9922) );
  NAND2_X1 U7041 ( .A1(n7459), .A2(n9922), .ZN(n7455) );
  NAND2_X1 U7042 ( .A1(n5708), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5542) );
  OR2_X1 U7043 ( .A1(n5490), .A2(n7571), .ZN(n5541) );
  AND2_X1 U7044 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  OR2_X1 U7045 ( .A1(n5538), .A2(n5552), .ZN(n9297) );
  OR2_X1 U7046 ( .A1(n5698), .A2(n9297), .ZN(n5540) );
  INV_X1 U7047 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7464) );
  OR2_X1 U7048 ( .A1(n5711), .A2(n7464), .ZN(n5539) );
  AND2_X1 U7049 ( .A1(n7453), .A2(n7458), .ZN(n5745) );
  NAND2_X1 U7050 ( .A1(n9232), .A2(n4416), .ZN(n7454) );
  AND2_X1 U7051 ( .A1(n7454), .A2(n7459), .ZN(n5543) );
  MUX2_X1 U7052 ( .A(n5745), .B(n5543), .S(n6845), .Z(n5544) );
  NAND2_X1 U7053 ( .A1(n5545), .A2(n5544), .ZN(n5571) );
  INV_X2 U7054 ( .A(n8118), .ZN(n10257) );
  NAND2_X1 U7055 ( .A1(n5708), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5550) );
  INV_X1 U7056 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7612) );
  OR2_X1 U7057 ( .A1(n5711), .A2(n7612), .ZN(n5549) );
  OR2_X1 U7058 ( .A1(n5554), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7059 ( .A1(n5561), .A2(n5546), .ZN(n9339) );
  OR2_X1 U7060 ( .A1(n5698), .A2(n9339), .ZN(n5548) );
  INV_X1 U7061 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6643) );
  OR2_X1 U7062 ( .A1(n5490), .A2(n6643), .ZN(n5547) );
  NAND2_X1 U7063 ( .A1(n10257), .A2(n9794), .ZN(n5736) );
  NAND2_X1 U7064 ( .A1(n5708), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5559) );
  INV_X1 U7065 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5551) );
  OR2_X1 U7066 ( .A1(n5490), .A2(n5551), .ZN(n5558) );
  NOR2_X1 U7067 ( .A1(n5552), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5553) );
  OR2_X1 U7068 ( .A1(n5554), .A2(n5553), .ZN(n7585) );
  OR2_X1 U7069 ( .A1(n5698), .A2(n7585), .ZN(n5557) );
  INV_X1 U7070 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7071 ( .A1(n5711), .A2(n5555), .ZN(n5556) );
  NAND2_X1 U7072 ( .A1(n9200), .A2(n10254), .ZN(n5844) );
  AND2_X1 U7073 ( .A1(n5736), .A2(n5844), .ZN(n5568) );
  NAND3_X1 U7074 ( .A1(n5571), .A2(n5568), .A3(n7454), .ZN(n5570) );
  NAND2_X1 U7075 ( .A1(n5708), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5567) );
  INV_X1 U7076 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9800) );
  OR2_X1 U7077 ( .A1(n5711), .A2(n9800), .ZN(n5566) );
  NAND2_X1 U7078 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  NAND2_X1 U7079 ( .A1(n5573), .A2(n5562), .ZN(n9799) );
  OR2_X1 U7080 ( .A1(n5698), .A2(n9799), .ZN(n5565) );
  INV_X1 U7081 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5563) );
  OR2_X1 U7082 ( .A1(n5490), .A2(n5563), .ZN(n5564) );
  INV_X1 U7083 ( .A(n5568), .ZN(n5800) );
  OR2_X1 U7084 ( .A1(n10254), .A2(n9200), .ZN(n5740) );
  NAND2_X1 U7085 ( .A1(n9804), .A2(n10274), .ZN(n5803) );
  INV_X1 U7086 ( .A(n5803), .ZN(n5569) );
  NAND2_X1 U7087 ( .A1(n5571), .A2(n7453), .ZN(n5572) );
  INV_X1 U7088 ( .A(n9771), .ZN(n5846) );
  NAND2_X1 U7089 ( .A1(n5708), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5578) );
  INV_X1 U7090 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9455) );
  OR2_X1 U7091 ( .A1(n5490), .A2(n9455), .ZN(n5577) );
  NAND2_X1 U7092 ( .A1(n5573), .A2(n9317), .ZN(n5574) );
  NAND2_X1 U7093 ( .A1(n5580), .A2(n5574), .ZN(n9780) );
  OR2_X1 U7094 ( .A1(n5698), .A2(n9780), .ZN(n5576) );
  INV_X1 U7095 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9781) );
  OR2_X1 U7096 ( .A1(n5711), .A2(n9781), .ZN(n5575) );
  NAND2_X1 U7097 ( .A1(n10279), .A2(n9911), .ZN(n5849) );
  NAND2_X1 U7098 ( .A1(n5708), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5585) );
  INV_X1 U7099 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9759) );
  OR2_X1 U7100 ( .A1(n5711), .A2(n9759), .ZN(n5584) );
  AND2_X1 U7101 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  OR2_X1 U7102 ( .A1(n5581), .A2(n5593), .ZN(n9758) );
  OR2_X1 U7103 ( .A1(n5698), .A2(n9758), .ZN(n5583) );
  INV_X1 U7104 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9094) );
  OR2_X1 U7105 ( .A1(n5490), .A2(n9094), .ZN(n5582) );
  OR2_X1 U7106 ( .A1(n10279), .A2(n9911), .ZN(n5735) );
  AND2_X1 U7107 ( .A1(n5851), .A2(n5735), .ZN(n5809) );
  INV_X1 U7108 ( .A(n5809), .ZN(n5586) );
  AOI21_X1 U7109 ( .B1(n5602), .B2(n5849), .A(n5586), .ZN(n5600) );
  NAND2_X1 U7110 ( .A1(n9914), .A2(n10276), .ZN(n5734) );
  INV_X1 U7111 ( .A(n5734), .ZN(n5603) );
  NAND2_X1 U7112 ( .A1(n5695), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5592) );
  INV_X1 U7113 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9990) );
  OR2_X1 U7114 ( .A1(n5697), .A2(n9990), .ZN(n5591) );
  OR2_X1 U7115 ( .A1(n5595), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7116 ( .A1(n5588), .A2(n5587), .ZN(n9726) );
  OR2_X1 U7117 ( .A1(n5698), .A2(n9726), .ZN(n5590) );
  INV_X1 U7118 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9899) );
  OR2_X1 U7119 ( .A1(n5490), .A2(n9899), .ZN(n5589) );
  OR2_X1 U7120 ( .A1(n9725), .A2(n9712), .ZN(n5732) );
  NAND2_X1 U7121 ( .A1(n5708), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5599) );
  INV_X1 U7122 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9744) );
  OR2_X1 U7123 ( .A1(n5711), .A2(n9744), .ZN(n5598) );
  NOR2_X1 U7124 ( .A1(n5593), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5594) );
  OR2_X1 U7125 ( .A1(n5595), .A2(n5594), .ZN(n9743) );
  OR2_X1 U7126 ( .A1(n5698), .A2(n9743), .ZN(n5597) );
  INV_X1 U7127 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10154) );
  OR2_X1 U7128 ( .A1(n5490), .A2(n10154), .ZN(n5596) );
  OR2_X1 U7129 ( .A1(n9747), .A2(n9912), .ZN(n5733) );
  AND2_X1 U7130 ( .A1(n5732), .A2(n5733), .ZN(n5785) );
  OAI21_X1 U7131 ( .B1(n5600), .B2(n5603), .A(n5785), .ZN(n5607) );
  INV_X1 U7132 ( .A(n5849), .ZN(n5601) );
  OAI21_X1 U7133 ( .B1(n5602), .B2(n5601), .A(n5809), .ZN(n5605) );
  NAND2_X1 U7134 ( .A1(n9725), .A2(n9712), .ZN(n5854) );
  NAND2_X1 U7135 ( .A1(n9747), .A2(n9912), .ZN(n5853) );
  NAND2_X1 U7136 ( .A1(n5854), .A2(n5853), .ZN(n5608) );
  NOR2_X1 U7137 ( .A1(n5608), .A2(n5603), .ZN(n5806) );
  INV_X1 U7138 ( .A(n5732), .ZN(n5604) );
  AOI21_X1 U7139 ( .B1(n5605), .B2(n5806), .A(n5604), .ZN(n5606) );
  AOI22_X1 U7140 ( .A1(n5608), .A2(n5732), .B1(n6845), .B2(n9905), .ZN(n5610)
         );
  AOI21_X1 U7141 ( .B1(n5854), .B2(n9893), .A(n5720), .ZN(n5609) );
  OR2_X1 U7142 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  NAND2_X1 U7143 ( .A1(n5708), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5618) );
  INV_X1 U7144 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5612) );
  OR2_X1 U7145 ( .A1(n5711), .A2(n5612), .ZN(n5617) );
  OAI21_X1 U7146 ( .B1(P1_REG3_REG_17__SCAN_IN), .B2(n5614), .A(n5613), .ZN(
        n9707) );
  OR2_X1 U7147 ( .A1(n5698), .A2(n9707), .ZN(n5616) );
  INV_X1 U7148 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9486) );
  OR2_X1 U7149 ( .A1(n5490), .A2(n9486), .ZN(n5615) );
  NAND4_X1 U7150 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n9892)
         );
  OR2_X1 U7151 ( .A1(n9888), .A2(n9699), .ZN(n9690) );
  NAND2_X1 U7152 ( .A1(n9888), .A2(n9699), .ZN(n5624) );
  NAND2_X1 U7153 ( .A1(n9690), .A2(n5624), .ZN(n9710) );
  INV_X1 U7154 ( .A(n9710), .ZN(n9705) );
  NAND2_X1 U7155 ( .A1(n5708), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5623) );
  INV_X1 U7156 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9696) );
  OR2_X1 U7157 ( .A1(n5711), .A2(n9696), .ZN(n5622) );
  OAI21_X1 U7158 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(n5619), .A(n5626), .ZN(
        n9695) );
  OR2_X1 U7159 ( .A1(n5698), .A2(n9695), .ZN(n5621) );
  INV_X1 U7160 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9885) );
  OR2_X1 U7161 ( .A1(n5490), .A2(n9885), .ZN(n5620) );
  NAND2_X1 U7162 ( .A1(n9701), .A2(n9713), .ZN(n5856) );
  AND2_X1 U7163 ( .A1(n5856), .A2(n5624), .ZN(n5814) );
  INV_X1 U7164 ( .A(n9874), .ZN(n9682) );
  NAND2_X1 U7165 ( .A1(n5695), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5631) );
  AOI21_X1 U7166 ( .B1(n5626), .B2(n9221), .A(n5625), .ZN(n9678) );
  INV_X1 U7167 ( .A(n9678), .ZN(n5627) );
  OR2_X1 U7168 ( .A1(n5698), .A2(n5627), .ZN(n5630) );
  INV_X1 U7169 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9877) );
  OR2_X1 U7170 ( .A1(n5490), .A2(n9877), .ZN(n5629) );
  INV_X1 U7171 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9981) );
  OR2_X1 U7172 ( .A1(n5697), .A2(n9981), .ZN(n5628) );
  OR2_X1 U7173 ( .A1(n9682), .A2(n9662), .ZN(n5816) );
  OR2_X1 U7174 ( .A1(n9701), .A2(n9713), .ZN(n5815) );
  NAND4_X1 U7175 ( .A1(n5632), .A2(n5816), .A3(n5720), .A4(n5815), .ZN(n5645)
         );
  NAND2_X1 U7176 ( .A1(n9867), .A2(n9654), .ZN(n5773) );
  NAND2_X1 U7177 ( .A1(n5776), .A2(n5773), .ZN(n5640) );
  NAND2_X1 U7178 ( .A1(n9682), .A2(n9662), .ZN(n5857) );
  INV_X1 U7179 ( .A(n5857), .ZN(n5633) );
  OR3_X1 U7180 ( .A1(n5640), .A2(n6845), .A3(n5633), .ZN(n5637) );
  NAND3_X1 U7181 ( .A1(n5819), .A2(n5720), .A3(n5776), .ZN(n5636) );
  NAND3_X1 U7182 ( .A1(n5640), .A2(n6845), .A3(n5775), .ZN(n5635) );
  NAND4_X1 U7183 ( .A1(n5775), .A2(n6845), .A3(n5731), .A4(n5816), .ZN(n5634)
         );
  NAND4_X1 U7184 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n5644)
         );
  AND2_X1 U7185 ( .A1(n5815), .A2(n9690), .ZN(n5810) );
  NAND3_X1 U7186 ( .A1(n5857), .A2(n6845), .A3(n5856), .ZN(n5638) );
  AOI21_X1 U7187 ( .B1(n5639), .B2(n5810), .A(n5638), .ZN(n5642) );
  INV_X1 U7188 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7189 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  OAI211_X1 U7190 ( .C1(n5819), .C2(n5645), .A(n5644), .B(n5643), .ZN(n5646)
         );
  XNOR2_X1 U7191 ( .A(n9854), .B(n9857), .ZN(n9629) );
  INV_X1 U7192 ( .A(n9629), .ZN(n9627) );
  NAND2_X1 U7193 ( .A1(n5695), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5652) );
  INV_X1 U7194 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9961) );
  OR2_X1 U7195 ( .A1(n5697), .A2(n9961), .ZN(n5651) );
  INV_X1 U7196 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9282) );
  XNOR2_X1 U7197 ( .A(n5665), .B(n9282), .ZN(n9600) );
  OR2_X1 U7198 ( .A1(n5698), .A2(n9600), .ZN(n5650) );
  INV_X1 U7199 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9839) );
  OR2_X1 U7200 ( .A1(n5490), .A2(n9839), .ZN(n5649) );
  NAND2_X1 U7201 ( .A1(n9838), .A2(n9842), .ZN(n5778) );
  MUX2_X1 U7202 ( .A(n5778), .B(n8155), .S(n6845), .Z(n5653) );
  NAND2_X1 U7203 ( .A1(n5654), .A2(n5653), .ZN(n5674) );
  INV_X1 U7204 ( .A(n5674), .ZN(n5673) );
  NAND2_X1 U7205 ( .A1(n5695), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5663) );
  INV_X1 U7206 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9950) );
  OR2_X1 U7207 ( .A1(n5697), .A2(n9950), .ZN(n5662) );
  INV_X1 U7208 ( .A(n5665), .ZN(n5656) );
  AND2_X1 U7209 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5655) );
  NAND2_X1 U7210 ( .A1(n5656), .A2(n5655), .ZN(n5666) );
  INV_X1 U7211 ( .A(n5666), .ZN(n5657) );
  NAND2_X1 U7212 ( .A1(n5657), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5685) );
  INV_X1 U7213 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7214 ( .A1(n5666), .A2(n5658), .ZN(n5659) );
  NAND2_X1 U7215 ( .A1(n5685), .A2(n5659), .ZN(n9356) );
  OR2_X1 U7216 ( .A1(n5698), .A2(n9356), .ZN(n5661) );
  INV_X1 U7217 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9828) );
  OR2_X1 U7218 ( .A1(n5490), .A2(n9828), .ZN(n5660) );
  NAND2_X1 U7219 ( .A1(n5695), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5671) );
  INV_X1 U7220 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9953) );
  OR2_X1 U7221 ( .A1(n5697), .A2(n9953), .ZN(n5670) );
  INV_X1 U7222 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5664) );
  OAI21_X1 U7223 ( .B1(n5665), .B2(n9282), .A(n5664), .ZN(n5667) );
  NAND2_X1 U7224 ( .A1(n5667), .A2(n5666), .ZN(n9257) );
  OR2_X1 U7225 ( .A1(n5698), .A2(n9257), .ZN(n5669) );
  INV_X1 U7226 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9832) );
  OR2_X1 U7227 ( .A1(n5490), .A2(n9832), .ZN(n5668) );
  NAND4_X1 U7228 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n9821)
         );
  INV_X1 U7229 ( .A(n9821), .ZN(n9566) );
  NAND2_X1 U7230 ( .A1(n5729), .A2(n8156), .ZN(n5771) );
  NAND2_X1 U7231 ( .A1(n9956), .A2(n9566), .ZN(n5730) );
  INV_X1 U7232 ( .A(n5730), .ZN(n5672) );
  NAND2_X1 U7233 ( .A1(n5729), .A2(n5672), .ZN(n5780) );
  OAI211_X1 U7234 ( .C1(n5673), .C2(n5771), .A(n8158), .B(n5780), .ZN(n5679)
         );
  INV_X1 U7235 ( .A(n5771), .ZN(n5677) );
  NAND2_X1 U7236 ( .A1(n5674), .A2(n5730), .ZN(n5676) );
  INV_X1 U7237 ( .A(n8158), .ZN(n5675) );
  AOI21_X1 U7238 ( .B1(n5677), .B2(n5676), .A(n5675), .ZN(n5678) );
  MUX2_X1 U7239 ( .A(n5679), .B(n5678), .S(n6845), .Z(n5693) );
  NAND2_X1 U7240 ( .A1(n5695), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5684) );
  INV_X1 U7241 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9146) );
  OR2_X1 U7242 ( .A1(n5697), .A2(n9146), .ZN(n5683) );
  INV_X1 U7243 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U7244 ( .A(n5685), .B(n8199), .ZN(n8198) );
  OR2_X1 U7245 ( .A1(n5698), .A2(n8198), .ZN(n5682) );
  INV_X1 U7246 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5680) );
  OR2_X1 U7247 ( .A1(n5490), .A2(n5680), .ZN(n5681) );
  INV_X1 U7248 ( .A(n8160), .ZN(n5824) );
  NAND2_X1 U7249 ( .A1(n5695), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5691) );
  INV_X1 U7250 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9069) );
  OR2_X1 U7251 ( .A1(n5697), .A2(n9069), .ZN(n5690) );
  INV_X1 U7252 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9000) );
  OAI21_X1 U7253 ( .B1(n5685), .B2(n8199), .A(n9000), .ZN(n5686) );
  OR3_X1 U7254 ( .A1(n5685), .A2(n9000), .A3(n8199), .ZN(n8176) );
  NAND2_X1 U7255 ( .A1(n5686), .A2(n8176), .ZN(n7833) );
  OR2_X1 U7256 ( .A1(n5698), .A2(n7833), .ZN(n5689) );
  INV_X1 U7257 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5687) );
  OR2_X1 U7258 ( .A1(n5490), .A2(n5687), .ZN(n5688) );
  NAND2_X1 U7259 ( .A1(n9814), .A2(n9548), .ZN(n5727) );
  NAND2_X1 U7260 ( .A1(n9946), .A2(n9527), .ZN(n5728) );
  AND2_X1 U7261 ( .A1(n5727), .A2(n5728), .ZN(n5784) );
  INV_X1 U7262 ( .A(n5784), .ZN(n5692) );
  NAND2_X1 U7263 ( .A1(n8161), .A2(n8160), .ZN(n5694) );
  NAND2_X1 U7264 ( .A1(n5695), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5703) );
  INV_X1 U7265 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5696) );
  OR2_X1 U7266 ( .A1(n5697), .A2(n5696), .ZN(n5702) );
  OR2_X1 U7267 ( .A1(n5698), .A2(n8176), .ZN(n5701) );
  INV_X1 U7268 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5699) );
  OR2_X1 U7269 ( .A1(n5490), .A2(n5699), .ZN(n5700) );
  NAND2_X1 U7270 ( .A1(n8188), .A2(n9528), .ZN(n5766) );
  INV_X1 U7271 ( .A(n5766), .ZN(n5705) );
  INV_X1 U7272 ( .A(n5828), .ZN(n5704) );
  MUX2_X1 U7273 ( .A(n5705), .B(n5704), .S(n6845), .Z(n5706) );
  INV_X1 U7274 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9517) );
  INV_X1 U7275 ( .A(n5490), .ZN(n5707) );
  NAND2_X1 U7276 ( .A1(n5707), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7277 ( .A1(n5708), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U7278 ( .C1(n5711), .C2(n9517), .A(n5710), .B(n5709), .ZN(n9381)
         );
  AOI22_X1 U7279 ( .A1(n9520), .A2(n5720), .B1(n9380), .B2(n9381), .ZN(n5712)
         );
  AND2_X1 U7280 ( .A1(n9514), .A2(n9380), .ZN(n5863) );
  INV_X1 U7281 ( .A(n5863), .ZN(n5833) );
  OAI211_X1 U7282 ( .C1(n5716), .C2(n5713), .A(n5712), .B(n5833), .ZN(n5719)
         );
  OAI211_X1 U7283 ( .C1(n9520), .C2(n5720), .A(n5714), .B(n9381), .ZN(n5715)
         );
  OAI21_X1 U7284 ( .B1(n5716), .B2(n5715), .A(n5721), .ZN(n5717) );
  INV_X1 U7285 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7286 ( .A1(n5719), .A2(n5718), .ZN(n5765) );
  OAI21_X1 U7287 ( .B1(n5721), .B2(n5720), .A(n5765), .ZN(n5726) );
  NOR3_X1 U7288 ( .A1(n7335), .A2(n6832), .A3(n7281), .ZN(n5723) );
  INV_X1 U7289 ( .A(n5724), .ZN(n5725) );
  AOI211_X1 U7290 ( .C1(n6659), .C2(n6845), .A(n7281), .B(n5722), .ZN(n5764)
         );
  NAND2_X1 U7291 ( .A1(n5731), .A2(n5773), .ZN(n9661) );
  NAND2_X1 U7292 ( .A1(n5815), .A2(n5856), .ZN(n9687) );
  INV_X1 U7293 ( .A(n9687), .ZN(n9692) );
  NAND2_X1 U7294 ( .A1(n5733), .A2(n5853), .ZN(n9737) );
  INV_X1 U7295 ( .A(n9737), .ZN(n5751) );
  NAND2_X1 U7296 ( .A1(n5851), .A2(n5734), .ZN(n9756) );
  NAND2_X1 U7297 ( .A1(n9790), .A2(n5736), .ZN(n7616) );
  INV_X1 U7298 ( .A(n7616), .ZN(n7610) );
  NAND2_X1 U7299 ( .A1(n9771), .A2(n5803), .ZN(n9797) );
  INV_X1 U7300 ( .A(n9797), .ZN(n9792) );
  AND2_X1 U7301 ( .A1(n8056), .A2(n9395), .ZN(n5788) );
  OR2_X1 U7302 ( .A1(n5788), .A2(n6962), .ZN(n10237) );
  NAND2_X1 U7303 ( .A1(n5794), .A2(n7376), .ZN(n7479) );
  NOR2_X1 U7304 ( .A1(n10237), .A2(n7479), .ZN(n5738) );
  NAND2_X1 U7305 ( .A1(n5837), .A2(n5792), .ZN(n7076) );
  NOR2_X1 U7306 ( .A1(n7076), .A2(n6659), .ZN(n5737) );
  XNOR2_X1 U7307 ( .A(n9393), .B(n8059), .ZN(n6839) );
  INV_X1 U7308 ( .A(n6839), .ZN(n6835) );
  AND4_X1 U7309 ( .A1(n5738), .A2(n5737), .A3(n6837), .A4(n6835), .ZN(n5744)
         );
  NAND2_X1 U7310 ( .A1(n5739), .A2(n7453), .ZN(n5797) );
  INV_X1 U7311 ( .A(n5797), .ZN(n5743) );
  NAND2_X1 U7312 ( .A1(n5740), .A2(n5844), .ZN(n7583) );
  INV_X1 U7313 ( .A(n7583), .ZN(n5742) );
  NOR2_X1 U7314 ( .A1(n6983), .A2(n7268), .ZN(n5741) );
  NAND4_X1 U7315 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n5747)
         );
  NAND2_X1 U7316 ( .A1(n7455), .A2(n5745), .ZN(n5746) );
  NAND2_X1 U7317 ( .A1(n5746), .A2(n7454), .ZN(n5798) );
  NOR2_X1 U7318 ( .A1(n5747), .A2(n5798), .ZN(n5748) );
  NAND4_X1 U7319 ( .A1(n9774), .A2(n7610), .A3(n9792), .A4(n5748), .ZN(n5749)
         );
  NOR2_X1 U7320 ( .A1(n9756), .A2(n5749), .ZN(n5750) );
  NAND3_X1 U7321 ( .A1(n9722), .A2(n5751), .A3(n5750), .ZN(n5752) );
  NOR2_X1 U7322 ( .A1(n9710), .A2(n5752), .ZN(n5753) );
  NAND3_X1 U7323 ( .A1(n9675), .A2(n9692), .A3(n5753), .ZN(n5754) );
  NOR2_X1 U7324 ( .A1(n9661), .A2(n5754), .ZN(n5755) );
  NAND2_X1 U7325 ( .A1(n9648), .A2(n5755), .ZN(n5756) );
  NOR2_X1 U7326 ( .A1(n9613), .A2(n5756), .ZN(n5757) );
  NAND4_X1 U7327 ( .A1(n9575), .A2(n4448), .A3(n5757), .A4(n9629), .ZN(n5758)
         );
  NOR2_X1 U7328 ( .A1(n9557), .A2(n5758), .ZN(n5759) );
  NAND4_X1 U7329 ( .A1(n8162), .A2(n9532), .A3(n8159), .A4(n5759), .ZN(n5762)
         );
  INV_X1 U7330 ( .A(n9381), .ZN(n5760) );
  NOR2_X1 U7331 ( .A1(n9520), .A2(n5760), .ZN(n5861) );
  INV_X1 U7332 ( .A(n5861), .ZN(n5831) );
  NAND2_X1 U7333 ( .A1(n5831), .A2(n5767), .ZN(n5761) );
  INV_X1 U7334 ( .A(n5871), .ZN(n5763) );
  OAI211_X1 U7335 ( .C1(n5765), .C2(n7335), .A(n5764), .B(n5763), .ZN(n5876)
         );
  NAND2_X1 U7336 ( .A1(n6973), .A2(n7281), .ZN(n5836) );
  NAND2_X1 U7337 ( .A1(n5768), .A2(n8155), .ZN(n5769) );
  AND2_X1 U7338 ( .A1(n5769), .A2(n5778), .ZN(n5770) );
  OR2_X1 U7339 ( .A1(n5771), .A2(n5770), .ZN(n5820) );
  INV_X1 U7340 ( .A(n5773), .ZN(n5774) );
  NAND2_X1 U7341 ( .A1(n5775), .A2(n5774), .ZN(n5777) );
  AND3_X1 U7342 ( .A1(n5779), .A2(n5778), .A3(n8151), .ZN(n5781) );
  OAI21_X1 U7343 ( .B1(n5820), .B2(n5781), .A(n5780), .ZN(n5782) );
  NAND2_X1 U7344 ( .A1(n5782), .A2(n8160), .ZN(n5783) );
  AND2_X1 U7345 ( .A1(n5784), .A2(n5783), .ZN(n5825) );
  NAND3_X1 U7346 ( .A1(n5826), .A2(n5825), .A3(n8158), .ZN(n5858) );
  INV_X1 U7347 ( .A(n5785), .ZN(n5813) );
  OAI22_X1 U7348 ( .A1(n7102), .A2(n6936), .B1(n8060), .B2(n6989), .ZN(n5787)
         );
  AOI211_X1 U7349 ( .C1(n5468), .C2(n6777), .A(n7335), .B(n5787), .ZN(n5791)
         );
  INV_X1 U7350 ( .A(n5788), .ZN(n5789) );
  AND3_X1 U7351 ( .A1(n5791), .A2(n5790), .A3(n5789), .ZN(n5793) );
  OAI21_X1 U7352 ( .B1(n5839), .B2(n5793), .A(n5792), .ZN(n5795) );
  INV_X1 U7353 ( .A(n5794), .ZN(n7377) );
  NOR2_X1 U7354 ( .A1(n5798), .A2(n7377), .ZN(n5840) );
  NAND2_X1 U7355 ( .A1(n5795), .A2(n5840), .ZN(n5801) );
  INV_X1 U7356 ( .A(n7376), .ZN(n5796) );
  NOR2_X1 U7357 ( .A1(n5797), .A2(n5796), .ZN(n5799) );
  OR2_X1 U7358 ( .A1(n5799), .A2(n5798), .ZN(n5841) );
  AOI21_X1 U7359 ( .B1(n5801), .B2(n5841), .A(n5800), .ZN(n5805) );
  INV_X1 U7360 ( .A(n5802), .ZN(n5804) );
  OAI211_X1 U7361 ( .C1(n5805), .C2(n5804), .A(n5849), .B(n5803), .ZN(n5808)
         );
  INV_X1 U7362 ( .A(n5806), .ZN(n5807) );
  AOI21_X1 U7363 ( .B1(n5809), .B2(n5808), .A(n5807), .ZN(n5812) );
  INV_X1 U7364 ( .A(n5810), .ZN(n5811) );
  AOI211_X1 U7365 ( .C1(n5854), .C2(n5813), .A(n5812), .B(n5811), .ZN(n5818)
         );
  INV_X1 U7366 ( .A(n5814), .ZN(n5817) );
  OAI211_X1 U7367 ( .C1(n5818), .C2(n5817), .A(n5816), .B(n5815), .ZN(n5822)
         );
  NOR2_X1 U7368 ( .A1(n5820), .A2(n5819), .ZN(n5859) );
  INV_X1 U7369 ( .A(n5859), .ZN(n5821) );
  AOI21_X1 U7370 ( .B1(n5857), .B2(n5822), .A(n5821), .ZN(n5832) );
  INV_X1 U7371 ( .A(n8161), .ZN(n5823) );
  AOI21_X1 U7372 ( .B1(n5825), .B2(n5824), .A(n5823), .ZN(n5829) );
  INV_X1 U7373 ( .A(n5826), .ZN(n5827) );
  AOI21_X1 U7374 ( .B1(n5829), .B2(n5828), .A(n5827), .ZN(n5862) );
  INV_X1 U7375 ( .A(n5862), .ZN(n5830) );
  OAI211_X1 U7376 ( .C1(n5858), .C2(n5832), .A(n5831), .B(n5830), .ZN(n5834)
         );
  AOI21_X1 U7377 ( .B1(n5834), .B2(n5833), .A(n5869), .ZN(n5835) );
  MUX2_X1 U7378 ( .A(n5836), .B(n5880), .S(n5835), .Z(n5874) );
  NAND2_X1 U7379 ( .A1(n7076), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U7380 ( .A1(n5839), .A2(n5838), .ZN(n7375) );
  NAND2_X1 U7381 ( .A1(n7375), .A2(n5840), .ZN(n5842) );
  NAND2_X1 U7382 ( .A1(n5842), .A2(n5841), .ZN(n7580) );
  INV_X1 U7383 ( .A(n7580), .ZN(n5843) );
  NAND2_X1 U7384 ( .A1(n7618), .A2(n9790), .ZN(n5845) );
  NAND2_X1 U7385 ( .A1(n5845), .A2(n9792), .ZN(n9770) );
  INV_X1 U7386 ( .A(n9774), .ZN(n5847) );
  NOR2_X1 U7387 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  INV_X1 U7388 ( .A(n5851), .ZN(n9738) );
  NOR2_X1 U7389 ( .A1(n9737), .A2(n9738), .ZN(n5852) );
  NAND2_X1 U7390 ( .A1(n9736), .A2(n5852), .ZN(n9740) );
  AND2_X1 U7391 ( .A1(n9692), .A2(n9690), .ZN(n5855) );
  NAND2_X1 U7392 ( .A1(n9689), .A2(n5855), .ZN(n9691) );
  AOI21_X1 U7393 ( .B1(n5859), .B2(n8148), .A(n5858), .ZN(n5860) );
  INV_X1 U7394 ( .A(n5860), .ZN(n5867) );
  NOR2_X1 U7395 ( .A1(n5862), .A2(n5006), .ZN(n5866) );
  NAND2_X1 U7396 ( .A1(n9514), .A2(n9520), .ZN(n5864) );
  AOI21_X1 U7397 ( .B1(n5867), .B2(n5866), .A(n5865), .ZN(n5870) );
  INV_X1 U7398 ( .A(n6842), .ZN(n5868) );
  NOR3_X1 U7399 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n5872) );
  OAI211_X1 U7400 ( .C1(n5872), .C2(n5871), .A(n6673), .B(n5722), .ZN(n5873)
         );
  NAND3_X1 U7401 ( .A1(n5877), .A2(n5876), .A3(n5875), .ZN(n5879) );
  OR2_X1 U7402 ( .A1(n6427), .A2(P1_U3086), .ZN(n7492) );
  NAND2_X1 U7403 ( .A1(n5879), .A2(n5878), .ZN(n5883) );
  NAND4_X1 U7404 ( .A1(n9929), .A2(n10005), .A3(n6844), .A4(n6647), .ZN(n5881)
         );
  OAI211_X1 U7405 ( .C1(n6832), .C2(n7492), .A(n5881), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5882) );
  NAND2_X1 U7406 ( .A1(n5883), .A2(n5882), .ZN(P1_U3242) );
  INV_X1 U7407 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6572) );
  INV_X1 U7408 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5884) );
  NOR2_X1 U7409 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5886) );
  NOR2_X1 U7410 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5889) );
  NAND4_X1 U7411 ( .A1(n5889), .A2(n6104), .A3(n6046), .A4(n6150), .ZN(n5892)
         );
  NOR2_X2 U7412 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  INV_X1 U7413 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5895) );
  INV_X1 U7414 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7415 ( .A1(n6333), .A2(n6336), .ZN(n5910) );
  INV_X1 U7416 ( .A(n5910), .ZN(n5897) );
  NOR2_X1 U7417 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5896) );
  INV_X1 U7418 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5898) );
  INV_X1 U7419 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7664) );
  XNOR2_X2 U7420 ( .A(n5899), .B(n7664), .ZN(n5904) );
  NAND2_X4 U7421 ( .A1(n5907), .A2(n8869), .ZN(n6323) );
  NAND2_X1 U7422 ( .A1(n5943), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5905) );
  INV_X2 U7423 ( .A(n8869), .ZN(n5908) );
  NAND2_X4 U7424 ( .A1(n5904), .A2(n5908), .ZN(n7679) );
  INV_X1 U7425 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6439) );
  INV_X1 U7426 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U7427 ( .A1(n6392), .A2(SI_0_), .ZN(n5909) );
  XNOR2_X1 U7428 ( .A(n5909), .B(n4886), .ZN(n9179) );
  NAND2_X1 U7429 ( .A1(n5910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  INV_X1 U7430 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5912) );
  INV_X1 U7431 ( .A(n5914), .ZN(n5915) );
  NAND2_X1 U7432 ( .A1(n5915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X2 U7433 ( .A(n5916), .B(n5898), .ZN(n6417) );
  MUX2_X1 U7434 ( .A(n6440), .B(n9179), .S(n6385), .Z(n6602) );
  INV_X1 U7435 ( .A(n6742), .ZN(n7846) );
  INV_X1 U7436 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6697) );
  OR2_X1 U7437 ( .A1(n6323), .A2(n6697), .ZN(n5923) );
  NAND2_X1 U7438 ( .A1(n4422), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5920) );
  INV_X1 U7439 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5918) );
  AND2_X1 U7440 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  NAND3_X1 U7441 ( .A1(n5923), .A2(n5922), .A3(n5921), .ZN(n5929) );
  NAND2_X1 U7442 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5924) );
  MUX2_X1 U7443 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5924), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5926) );
  INV_X1 U7444 ( .A(n5925), .ZN(n6441) );
  NAND2_X1 U7445 ( .A1(n5926), .A2(n6441), .ZN(n6458) );
  INV_X1 U7446 ( .A(n6458), .ZN(n6447) );
  NAND2_X1 U7447 ( .A1(n6741), .A2(n5929), .ZN(n7848) );
  NAND2_X1 U7448 ( .A1(n6687), .A2(n5930), .ZN(n6995) );
  NAND2_X1 U7449 ( .A1(n4423), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5936) );
  INV_X1 U7450 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5931) );
  INV_X1 U7451 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6462) );
  INV_X1 U7452 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5932) );
  NAND4_X2 U7453 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n8366)
         );
  INV_X1 U7454 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6390) );
  OR2_X1 U7455 ( .A1(n5952), .A2(n6390), .ZN(n5939) );
  OAI211_X1 U7456 ( .C1(n6385), .C2(n4417), .A(n5939), .B(n5938), .ZN(n5941)
         );
  OR2_X2 U7457 ( .A1(n8366), .A2(n4421), .ZN(n6885) );
  NAND2_X1 U7458 ( .A1(n8366), .A2(n4421), .ZN(n5940) );
  NAND2_X1 U7459 ( .A1(n6995), .A2(n8003), .ZN(n5942) );
  INV_X1 U7460 ( .A(n8366), .ZN(n7856) );
  NAND2_X1 U7461 ( .A1(n7856), .A2(n4421), .ZN(n7855) );
  NAND2_X1 U7462 ( .A1(n5942), .A2(n7855), .ZN(n6883) );
  NAND2_X1 U7463 ( .A1(n4423), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5948) );
  INV_X1 U7464 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7465 ( .A1(n7679), .A2(n5944), .ZN(n5947) );
  INV_X1 U7466 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6889) );
  OR2_X1 U7467 ( .A1(n6323), .A2(n6889), .ZN(n5946) );
  OR2_X1 U7468 ( .A1(n6127), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7469 ( .A1(n5937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  MUX2_X1 U7470 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5949), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5951) );
  NAND2_X1 U7471 ( .A1(n5951), .A2(n5950), .ZN(n6517) );
  NAND2_X1 U7472 ( .A1(n6997), .A2(n6890), .ZN(n7866) );
  NAND2_X1 U7473 ( .A1(n7863), .A2(n7866), .ZN(n6281) );
  INV_X1 U7474 ( .A(n6281), .ZN(n8002) );
  NAND2_X1 U7475 ( .A1(n6883), .A2(n8002), .ZN(n6882) );
  NAND2_X1 U7476 ( .A1(n6882), .A2(n7866), .ZN(n6790) );
  NAND2_X1 U7477 ( .A1(n4423), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5958) );
  INV_X1 U7478 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7479 ( .A1(n7679), .A2(n5954), .ZN(n5957) );
  XNOR2_X1 U7480 ( .A(n5968), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n6766) );
  OR2_X1 U7481 ( .A1(n6127), .A2(n6766), .ZN(n5956) );
  INV_X1 U7482 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6800) );
  OR2_X1 U7483 ( .A1(n6323), .A2(n6800), .ZN(n5955) );
  NAND2_X1 U7484 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5960) );
  OR2_X1 U7485 ( .A1(n5953), .A2(n6396), .ZN(n5962) );
  INV_X1 U7486 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6391) );
  OR2_X1 U7487 ( .A1(n5952), .A2(n6391), .ZN(n5961) );
  OAI211_X1 U7488 ( .C1(n6385), .C2(n6542), .A(n5962), .B(n5961), .ZN(n6802)
         );
  OR2_X1 U7489 ( .A1(n7060), .A2(n6802), .ZN(n7867) );
  NAND2_X1 U7490 ( .A1(n7060), .A2(n6802), .ZN(n7862) );
  NAND2_X1 U7491 ( .A1(n7867), .A2(n7862), .ZN(n8005) );
  INV_X1 U7492 ( .A(n8005), .ZN(n7859) );
  NAND2_X1 U7493 ( .A1(n6790), .A2(n7859), .ZN(n5963) );
  NAND2_X1 U7494 ( .A1(n5963), .A2(n7862), .ZN(n7055) );
  OR2_X1 U7495 ( .A1(n5950), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7496 ( .A1(n5982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5964) );
  INV_X1 U7497 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7498 ( .A(n5964), .B(n5983), .ZN(n6554) );
  OR2_X1 U7499 ( .A1(n5953), .A2(n6399), .ZN(n5966) );
  INV_X1 U7500 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6397) );
  OR2_X1 U7501 ( .A1(n5952), .A2(n6397), .ZN(n5965) );
  OAI211_X1 U7502 ( .C1(n6385), .C2(n6554), .A(n5966), .B(n5965), .ZN(n7112)
         );
  INV_X1 U7503 ( .A(n7112), .ZN(n7064) );
  NAND2_X1 U7504 ( .A1(n4982), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5974) );
  INV_X1 U7505 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5967) );
  OR2_X1 U7506 ( .A1(n6263), .A2(n5967), .ZN(n5973) );
  OAI21_X1 U7507 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5970) );
  AND2_X1 U7508 ( .A1(n5976), .A2(n5970), .ZN(n6915) );
  OR2_X1 U7509 ( .A1(n6127), .A2(n6915), .ZN(n5972) );
  INV_X1 U7510 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7110) );
  OR2_X1 U7511 ( .A1(n6323), .A2(n7110), .ZN(n5971) );
  NAND4_X1 U7512 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n8364)
         );
  NAND2_X1 U7513 ( .A1(n7064), .A2(n8364), .ZN(n7868) );
  NAND2_X1 U7514 ( .A1(n7055), .A2(n7868), .ZN(n5975) );
  INV_X1 U7515 ( .A(n8364), .ZN(n7011) );
  NAND2_X1 U7516 ( .A1(n7011), .A2(n7112), .ZN(n7871) );
  NAND2_X1 U7517 ( .A1(n5975), .A2(n7871), .ZN(n7087) );
  NAND2_X1 U7518 ( .A1(n4423), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5981) );
  INV_X1 U7519 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6708) );
  OR2_X1 U7520 ( .A1(n7679), .A2(n6708), .ZN(n5980) );
  NAND2_X1 U7521 ( .A1(n5976), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5977) );
  AND2_X1 U7522 ( .A1(n5991), .A2(n5977), .ZN(n7088) );
  OR2_X1 U7523 ( .A1(n6127), .A2(n7088), .ZN(n5979) );
  INV_X1 U7524 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6820) );
  OR2_X1 U7525 ( .A1(n6323), .A2(n6820), .ZN(n5978) );
  NAND4_X1 U7526 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n8363)
         );
  INV_X1 U7527 ( .A(n8363), .ZN(n7399) );
  INV_X1 U7528 ( .A(n5982), .ZN(n5984) );
  NAND2_X1 U7529 ( .A1(n5984), .A2(n5983), .ZN(n5997) );
  NAND2_X1 U7530 ( .A1(n5997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7531 ( .A(n5985), .B(n5998), .ZN(n6721) );
  OR2_X1 U7532 ( .A1(n5953), .A2(n6403), .ZN(n5987) );
  INV_X1 U7533 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6401) );
  OR2_X1 U7534 ( .A1(n5952), .A2(n6401), .ZN(n5986) );
  OAI211_X1 U7535 ( .C1(n6385), .C2(n6721), .A(n5987), .B(n5986), .ZN(n7014)
         );
  AND2_X1 U7536 ( .A1(n7399), .A2(n7014), .ZN(n7872) );
  INV_X1 U7537 ( .A(n7014), .ZN(n7228) );
  NAND2_X1 U7538 ( .A1(n7228), .A2(n8363), .ZN(n7864) );
  NAND2_X1 U7539 ( .A1(n4982), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5996) );
  INV_X1 U7540 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7541 ( .A1(n6263), .A2(n5988), .ZN(n5995) );
  NAND2_X1 U7542 ( .A1(n5991), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5992) );
  AND2_X1 U7543 ( .A1(n6013), .A2(n5992), .ZN(n7155) );
  OR2_X1 U7544 ( .A1(n6127), .A2(n7155), .ZN(n5994) );
  OR2_X1 U7545 ( .A1(n6323), .A2(n6824), .ZN(n5993) );
  INV_X1 U7546 ( .A(n5997), .ZN(n5999) );
  NAND2_X1 U7547 ( .A1(n5999), .A2(n5998), .ZN(n6005) );
  NAND2_X1 U7548 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6000) );
  INV_X1 U7549 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U7550 ( .A(n6000), .B(n6006), .ZN(n6859) );
  OR2_X1 U7551 ( .A1(n6407), .A2(n5953), .ZN(n6003) );
  INV_X1 U7552 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7553 ( .A1(n5952), .A2(n6001), .ZN(n6002) );
  OAI211_X1 U7554 ( .C1(n6385), .C2(n6859), .A(n6003), .B(n6002), .ZN(n10306)
         );
  OR2_X1 U7555 ( .A1(n7336), .A2(n10306), .ZN(n7223) );
  NAND2_X1 U7556 ( .A1(n7336), .A2(n10306), .ZN(n7884) );
  NAND2_X1 U7557 ( .A1(n7395), .A2(n8007), .ZN(n7222) );
  NAND2_X1 U7558 ( .A1(n6004), .A2(n7968), .ZN(n6010) );
  INV_X1 U7559 ( .A(n6005), .ZN(n6007) );
  NAND2_X1 U7560 ( .A1(n6007), .A2(n6006), .ZN(n6019) );
  NAND2_X1 U7561 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7562 ( .A(n6008), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U7563 ( .A1(n7677), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4731), .B2(
        n7046), .ZN(n6009) );
  NAND2_X1 U7564 ( .A1(n6010), .A2(n6009), .ZN(n7340) );
  NAND2_X1 U7565 ( .A1(n4423), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6018) );
  INV_X1 U7566 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6863) );
  OR2_X1 U7567 ( .A1(n7679), .A2(n6863), .ZN(n6017) );
  NAND2_X1 U7568 ( .A1(n6013), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6014) );
  AND2_X1 U7569 ( .A1(n6024), .A2(n6014), .ZN(n7341) );
  OR2_X1 U7570 ( .A1(n6127), .A2(n7341), .ZN(n6016) );
  INV_X1 U7571 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7220) );
  OR2_X1 U7572 ( .A1(n6323), .A2(n7220), .ZN(n6015) );
  OR2_X1 U7573 ( .A1(n7340), .A2(n7403), .ZN(n7880) );
  AND2_X1 U7574 ( .A1(n7880), .A2(n7223), .ZN(n7877) );
  NAND2_X1 U7575 ( .A1(n7340), .A2(n7403), .ZN(n7885) );
  NAND2_X1 U7576 ( .A1(n6409), .A2(n7968), .ZN(n6022) );
  OAI21_X1 U7577 ( .B1(n6019), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6020) );
  XNOR2_X1 U7578 ( .A(n6020), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7164) );
  AOI22_X1 U7579 ( .A1(n7677), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4731), .B2(
        n7164), .ZN(n6021) );
  NAND2_X1 U7580 ( .A1(n6022), .A2(n6021), .ZN(n7490) );
  NAND2_X1 U7581 ( .A1(n4982), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6029) );
  INV_X1 U7582 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6023) );
  OR2_X1 U7583 ( .A1(n6263), .A2(n6023), .ZN(n6028) );
  NAND2_X1 U7584 ( .A1(n6024), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6025) );
  AND2_X1 U7585 ( .A1(n6037), .A2(n6025), .ZN(n7430) );
  OR2_X1 U7586 ( .A1(n6127), .A2(n7430), .ZN(n6027) );
  INV_X1 U7587 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7033) );
  OR2_X1 U7588 ( .A1(n6323), .A2(n7033), .ZN(n6026) );
  NAND2_X1 U7589 ( .A1(n7490), .A2(n7442), .ZN(n7886) );
  NAND2_X1 U7590 ( .A1(n7881), .A2(n7886), .ZN(n7999) );
  OR2_X1 U7591 ( .A1(n9172), .A2(n5953), .ZN(n6034) );
  OR2_X1 U7592 ( .A1(n6031), .A2(n6106), .ZN(n6032) );
  XNOR2_X1 U7593 ( .A(n6032), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9174) );
  AOI22_X1 U7594 ( .A1(n7677), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4731), .B2(
        n9174), .ZN(n6033) );
  NAND2_X1 U7595 ( .A1(n6034), .A2(n6033), .ZN(n7450) );
  NAND2_X1 U7596 ( .A1(n4423), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6042) );
  INV_X1 U7597 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7178) );
  OR2_X1 U7598 ( .A1(n7679), .A2(n7178), .ZN(n6041) );
  INV_X1 U7599 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7600 ( .A1(n6037), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6038) );
  AND2_X1 U7601 ( .A1(n6051), .A2(n6038), .ZN(n7447) );
  OR2_X1 U7602 ( .A1(n6127), .A2(n7447), .ZN(n6040) );
  INV_X1 U7603 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7448) );
  OR2_X1 U7604 ( .A1(n6323), .A2(n7448), .ZN(n6039) );
  OR2_X1 U7605 ( .A1(n7450), .A2(n7623), .ZN(n7897) );
  AND2_X1 U7606 ( .A1(n7897), .A2(n7881), .ZN(n7891) );
  NAND2_X1 U7607 ( .A1(n7439), .A2(n7891), .ZN(n6043) );
  NAND2_X1 U7608 ( .A1(n7450), .A2(n7623), .ZN(n7895) );
  NAND2_X1 U7609 ( .A1(n6043), .A2(n7895), .ZN(n7499) );
  NAND2_X1 U7610 ( .A1(n6424), .A2(n7968), .ZN(n6050) );
  NOR2_X1 U7611 ( .A1(n6044), .A2(n6106), .ZN(n6045) );
  MUX2_X1 U7612 ( .A(n6106), .B(n6045), .S(P2_IR_REG_11__SCAN_IN), .Z(n6048)
         );
  INV_X1 U7613 ( .A(n6070), .ZN(n6047) );
  OR2_X1 U7614 ( .A1(n6048), .A2(n6047), .ZN(n7249) );
  INV_X1 U7615 ( .A(n7249), .ZN(n7233) );
  AOI22_X1 U7616 ( .A1(n7677), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4731), .B2(
        n7233), .ZN(n6049) );
  NAND2_X1 U7617 ( .A1(n4423), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6056) );
  INV_X1 U7618 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7503) );
  OR2_X1 U7619 ( .A1(n6323), .A2(n7503), .ZN(n6055) );
  NAND2_X1 U7620 ( .A1(n6051), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6052) );
  AND2_X1 U7621 ( .A1(n6063), .A2(n6052), .ZN(n7627) );
  OR2_X1 U7622 ( .A1(n6127), .A2(n7627), .ZN(n6054) );
  INV_X1 U7623 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7195) );
  OR2_X1 U7624 ( .A1(n7679), .A2(n7195), .ZN(n6053) );
  NAND2_X1 U7625 ( .A1(n7633), .A2(n7599), .ZN(n7900) );
  INV_X1 U7626 ( .A(n8014), .ZN(n7500) );
  OR2_X1 U7627 ( .A1(n6432), .A2(n5953), .ZN(n6059) );
  NAND2_X1 U7628 ( .A1(n6070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6057) );
  XNOR2_X1 U7629 ( .A(n6057), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7254) );
  AOI22_X1 U7630 ( .A1(n7677), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4731), .B2(
        n7254), .ZN(n6058) );
  NAND2_X1 U7631 ( .A1(n4982), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6068) );
  INV_X1 U7632 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7633 ( .A1(n6263), .A2(n6060), .ZN(n6067) );
  INV_X1 U7634 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7635 ( .A1(n6063), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6064) );
  AND2_X1 U7636 ( .A1(n6073), .A2(n6064), .ZN(n7603) );
  OR2_X1 U7637 ( .A1(n6127), .A2(n7603), .ZN(n6066) );
  INV_X1 U7638 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8966) );
  OR2_X1 U7639 ( .A1(n6323), .A2(n8966), .ZN(n6065) );
  NAND4_X1 U7640 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n8688)
         );
  INV_X1 U7641 ( .A(n8688), .ZN(n7657) );
  XNOR2_X1 U7642 ( .A(n7906), .B(n7657), .ZN(n7557) );
  INV_X1 U7643 ( .A(n7557), .ZN(n6069) );
  OR2_X1 U7644 ( .A1(n7906), .A2(n7657), .ZN(n7905) );
  NAND2_X1 U7645 ( .A1(n8761), .A2(n7905), .ZN(n8694) );
  OR2_X1 U7646 ( .A1(n6486), .A2(n5953), .ZN(n6072) );
  NAND2_X1 U7647 ( .A1(n6105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6080) );
  XNOR2_X1 U7648 ( .A(n6080), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7509) );
  AOI22_X1 U7649 ( .A1(n7677), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4731), .B2(
        n7509), .ZN(n6071) );
  NAND2_X1 U7650 ( .A1(n4423), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6078) );
  INV_X1 U7651 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8754) );
  OR2_X1 U7652 ( .A1(n7679), .A2(n8754), .ZN(n6077) );
  NAND2_X1 U7653 ( .A1(n6073), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6074) );
  AND2_X1 U7654 ( .A1(n6084), .A2(n6074), .ZN(n8682) );
  OR2_X1 U7655 ( .A1(n6127), .A2(n8682), .ZN(n6076) );
  INV_X1 U7656 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7354) );
  OR2_X1 U7657 ( .A1(n6323), .A2(n7354), .ZN(n6075) );
  NAND4_X1 U7658 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n8358)
         );
  INV_X1 U7659 ( .A(n8358), .ZN(n8670) );
  NAND2_X1 U7660 ( .A1(n8861), .A2(n8670), .ZN(n7910) );
  NAND2_X1 U7661 ( .A1(n8694), .A2(n7910), .ZN(n6079) );
  OR2_X1 U7662 ( .A1(n8861), .A2(n8670), .ZN(n7911) );
  NAND2_X1 U7663 ( .A1(n6533), .A2(n7968), .ZN(n6083) );
  NAND2_X1 U7664 ( .A1(n6080), .A2(n6103), .ZN(n6081) );
  NAND2_X1 U7665 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7666 ( .A(n6090), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7522) );
  AOI22_X1 U7667 ( .A1(n7677), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4731), .B2(
        n7522), .ZN(n6082) );
  NAND2_X1 U7668 ( .A1(n4423), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6089) );
  INV_X1 U7669 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9020) );
  OR2_X1 U7670 ( .A1(n7679), .A2(n9020), .ZN(n6088) );
  NAND2_X1 U7671 ( .A1(n6084), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6085) );
  AND2_X1 U7672 ( .A1(n6096), .A2(n6085), .ZN(n8676) );
  OR2_X1 U7673 ( .A1(n6127), .A2(n8676), .ZN(n6087) );
  INV_X1 U7674 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8677) );
  OR2_X1 U7675 ( .A1(n6323), .A2(n8677), .ZN(n6086) );
  NAND4_X1 U7676 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n8686)
         );
  INV_X1 U7677 ( .A(n8686), .ZN(n8341) );
  NOR2_X1 U7678 ( .A1(n8855), .A2(n8341), .ZN(n7915) );
  NAND2_X1 U7679 ( .A1(n8855), .A2(n8341), .ZN(n7843) );
  NAND2_X1 U7680 ( .A1(n6657), .A2(n7968), .ZN(n6094) );
  NAND2_X1 U7681 ( .A1(n6090), .A2(n6104), .ZN(n6091) );
  NAND2_X1 U7682 ( .A1(n6091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6092) );
  XNOR2_X1 U7683 ( .A(n6092), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8393) );
  AOI22_X1 U7684 ( .A1(n7677), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4731), .B2(
        n8393), .ZN(n6093) );
  NAND2_X1 U7685 ( .A1(n4423), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6101) );
  INV_X1 U7686 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9107) );
  OR2_X1 U7687 ( .A1(n7679), .A2(n9107), .ZN(n6100) );
  INV_X1 U7688 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U7689 ( .A1(n6096), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6097) );
  AND2_X1 U7690 ( .A1(n6114), .A2(n6097), .ZN(n8662) );
  OR2_X1 U7691 ( .A1(n6127), .A2(n8662), .ZN(n6099) );
  INV_X1 U7692 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8661) );
  OR2_X1 U7693 ( .A1(n6323), .A2(n8661), .ZN(n6098) );
  NAND4_X1 U7694 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n8357)
         );
  NAND2_X1 U7695 ( .A1(n8848), .A2(n8672), .ZN(n6297) );
  INV_X1 U7696 ( .A(n6297), .ZN(n7919) );
  NAND2_X1 U7697 ( .A1(n6726), .A2(n7968), .ZN(n6111) );
  INV_X1 U7698 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7699 ( .A1(n4508), .A2(n6106), .ZN(n6107) );
  INV_X1 U7700 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6108) );
  MUX2_X1 U7701 ( .A(n6107), .B(P2_IR_REG_31__SCAN_IN), .S(n6108), .Z(n6109)
         );
  NAND2_X1 U7702 ( .A1(n6109), .A2(n6134), .ZN(n8422) );
  INV_X1 U7703 ( .A(n8422), .ZN(n8425) );
  AOI22_X1 U7704 ( .A1(n7677), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4731), .B2(
        n8425), .ZN(n6110) );
  NAND2_X1 U7705 ( .A1(n4423), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6119) );
  INV_X1 U7706 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8745) );
  OR2_X1 U7707 ( .A1(n7679), .A2(n8745), .ZN(n6118) );
  INV_X1 U7708 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7709 ( .A1(n6114), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6115) );
  AND2_X1 U7710 ( .A1(n6125), .A2(n6115), .ZN(n8652) );
  OR2_X1 U7711 ( .A1(n6127), .A2(n8652), .ZN(n6117) );
  INV_X1 U7712 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8651) );
  OR2_X1 U7713 ( .A1(n6323), .A2(n8651), .ZN(n6116) );
  NAND4_X1 U7714 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n8659)
         );
  INV_X1 U7715 ( .A(n8659), .ZN(n8276) );
  NAND2_X1 U7716 ( .A1(n8842), .A2(n8276), .ZN(n7925) );
  NAND2_X1 U7717 ( .A1(n6120), .A2(n7923), .ZN(n8628) );
  INV_X1 U7718 ( .A(n8628), .ZN(n6133) );
  NAND2_X1 U7719 ( .A1(n6855), .A2(n7968), .ZN(n6123) );
  NAND2_X1 U7720 ( .A1(n6134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7721 ( .A(n6121), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8452) );
  AOI22_X1 U7722 ( .A1(n7677), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4731), .B2(
        n8452), .ZN(n6122) );
  NAND2_X1 U7723 ( .A1(n4423), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6131) );
  INV_X1 U7724 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7725 ( .A1(n7679), .A2(n6124), .ZN(n6130) );
  NAND2_X1 U7726 ( .A1(n6125), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6126) );
  AND2_X1 U7727 ( .A1(n6142), .A2(n6126), .ZN(n8632) );
  OR2_X1 U7728 ( .A1(n6127), .A2(n8632), .ZN(n6129) );
  INV_X1 U7729 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9059) );
  OR2_X1 U7730 ( .A1(n6323), .A2(n9059), .ZN(n6128) );
  OR2_X1 U7731 ( .A1(n8631), .A2(n8647), .ZN(n7924) );
  NAND2_X1 U7732 ( .A1(n8631), .A2(n8647), .ZN(n7929) );
  INV_X1 U7733 ( .A(n8635), .ZN(n6132) );
  NAND2_X1 U7734 ( .A1(n7029), .A2(n7968), .ZN(n6138) );
  INV_X1 U7735 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7736 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7737 ( .A(n6151), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8467) );
  AOI22_X1 U7738 ( .A1(n7677), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4731), .B2(
        n8467), .ZN(n6137) );
  INV_X1 U7739 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7740 ( .A1(n6142), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7741 ( .A1(n6155), .A2(n6143), .ZN(n8619) );
  NAND2_X1 U7742 ( .A1(n6139), .A2(n8619), .ZN(n6148) );
  INV_X1 U7743 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8462) );
  OR2_X1 U7744 ( .A1(n7679), .A2(n8462), .ZN(n6147) );
  INV_X1 U7745 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6144) );
  OR2_X1 U7746 ( .A1(n6263), .A2(n6144), .ZN(n6146) );
  INV_X1 U7747 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8621) );
  OR2_X1 U7748 ( .A1(n6323), .A2(n8621), .ZN(n6145) );
  NAND4_X1 U7749 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n8637)
         );
  INV_X1 U7750 ( .A(n8637), .ZN(n8234) );
  NAND2_X1 U7751 ( .A1(n8737), .A2(n8234), .ZN(n7937) );
  NAND2_X1 U7752 ( .A1(n8601), .A2(n7937), .ZN(n8623) );
  NAND2_X1 U7753 ( .A1(n7159), .A2(n7968), .ZN(n6154) );
  NAND2_X1 U7754 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  INV_X1 U7755 ( .A(n8485), .ZN(n6363) );
  AOI22_X1 U7756 ( .A1(n7677), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6363), .B2(
        n4731), .ZN(n6153) );
  NAND2_X1 U7757 ( .A1(n6155), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7758 ( .A1(n6166), .A2(n6156), .ZN(n8608) );
  NAND2_X1 U7759 ( .A1(n6139), .A2(n8608), .ZN(n6160) );
  NAND2_X1 U7760 ( .A1(n6260), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6159) );
  INV_X1 U7761 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8732) );
  OR2_X1 U7762 ( .A1(n7679), .A2(n8732), .ZN(n6158) );
  INV_X1 U7763 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9134) );
  OR2_X1 U7764 ( .A1(n6263), .A2(n9134), .ZN(n6157) );
  NAND4_X1 U7765 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8615)
         );
  INV_X1 U7766 ( .A(n8615), .ZN(n8591) );
  OR2_X1 U7767 ( .A1(n8829), .A2(n8591), .ZN(n7998) );
  AND2_X1 U7768 ( .A1(n7998), .A2(n8601), .ZN(n7930) );
  NAND2_X1 U7769 ( .A1(n8736), .A2(n7930), .ZN(n6161) );
  NAND2_X1 U7770 ( .A1(n8829), .A2(n8591), .ZN(n7997) );
  NAND2_X1 U7771 ( .A1(n6161), .A2(n7997), .ZN(n8594) );
  NAND2_X1 U7772 ( .A1(n7263), .A2(n7968), .ZN(n6164) );
  INV_X1 U7773 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6162) );
  OR2_X1 U7774 ( .A1(n5952), .A2(n6162), .ZN(n6163) );
  AOI22_X1 U7775 ( .A1(n4982), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n4423), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6170) );
  INV_X1 U7776 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U7777 ( .A1(n6166), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7778 ( .A1(n6175), .A2(n6167), .ZN(n8597) );
  NAND2_X1 U7779 ( .A1(n8597), .A2(n6139), .ZN(n6169) );
  NAND2_X1 U7780 ( .A1(n6260), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7781 ( .A1(n8594), .A2(n7943), .ZN(n6171) );
  NAND2_X1 U7782 ( .A1(n8596), .A2(n8579), .ZN(n7933) );
  NAND2_X1 U7783 ( .A1(n6171), .A2(n7933), .ZN(n8581) );
  NAND2_X1 U7784 ( .A1(n6172), .A2(n7968), .ZN(n6174) );
  OR2_X1 U7785 ( .A1(n5952), .A2(n7327), .ZN(n6173) );
  INV_X1 U7786 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U7787 ( .A1(n6175), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7788 ( .A1(n6183), .A2(n6176), .ZN(n8580) );
  NAND2_X1 U7789 ( .A1(n8580), .A2(n6139), .ZN(n6178) );
  AOI22_X1 U7790 ( .A1(n4982), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n4423), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7791 ( .C1(n6323), .C2(n8584), .A(n6178), .B(n6177), .ZN(n8589)
         );
  INV_X1 U7792 ( .A(n8589), .ZN(n8085) );
  NAND2_X1 U7793 ( .A1(n8251), .A2(n8085), .ZN(n7944) );
  INV_X1 U7794 ( .A(n7944), .ZN(n7934) );
  OAI21_X2 U7795 ( .B1(n8581), .B2(n7934), .A(n7945), .ZN(n8567) );
  NAND2_X1 U7796 ( .A1(n7536), .A2(n7968), .ZN(n6180) );
  OR2_X1 U7797 ( .A1(n5952), .A2(n7540), .ZN(n6179) );
  INV_X1 U7798 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7799 ( .A1(n6183), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7800 ( .A1(n6204), .A2(n6184), .ZN(n8573) );
  NAND2_X1 U7801 ( .A1(n8573), .A2(n6139), .ZN(n6189) );
  INV_X1 U7802 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U7803 ( .A1(n4982), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7804 ( .A1(n4423), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6185) );
  OAI211_X1 U7805 ( .C1(n8572), .C2(n6323), .A(n6186), .B(n6185), .ZN(n6187)
         );
  INV_X1 U7806 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7807 ( .A1(n6189), .A2(n6188), .ZN(n8560) );
  INV_X1 U7808 ( .A(n8560), .ZN(n8578) );
  NAND2_X1 U7809 ( .A1(n8815), .A2(n8578), .ZN(n7949) );
  INV_X1 U7810 ( .A(n7950), .ZN(n6190) );
  NAND2_X1 U7811 ( .A1(n7635), .A2(n7968), .ZN(n6192) );
  OR2_X1 U7812 ( .A1(n5952), .A2(n7650), .ZN(n6191) );
  INV_X1 U7813 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9010) );
  INV_X1 U7814 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6194) );
  INV_X1 U7815 ( .A(n6195), .ZN(n6206) );
  NAND2_X1 U7816 ( .A1(n6206), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7817 ( .A1(n6216), .A2(n6196), .ZN(n8548) );
  NAND2_X1 U7818 ( .A1(n8548), .A2(n6139), .ZN(n6201) );
  NAND2_X1 U7819 ( .A1(n4423), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7820 ( .A1(n4982), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7821 ( .C1(n9001), .C2(n6323), .A(n6198), .B(n6197), .ZN(n6199)
         );
  INV_X1 U7822 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7823 ( .A1(n8803), .A2(n8285), .ZN(n7995) );
  NAND2_X1 U7824 ( .A1(n7495), .A2(n7968), .ZN(n6203) );
  OR2_X1 U7825 ( .A1(n5952), .A2(n7498), .ZN(n6202) );
  NAND2_X1 U7826 ( .A1(n6204), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7827 ( .A1(n6206), .A2(n6205), .ZN(n8564) );
  NAND2_X1 U7828 ( .A1(n8564), .A2(n6139), .ZN(n6211) );
  INV_X1 U7829 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U7830 ( .A1(n4423), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7831 ( .A1(n4982), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6207) );
  OAI211_X1 U7832 ( .C1(n8563), .C2(n6323), .A(n6208), .B(n6207), .ZN(n6209)
         );
  INV_X1 U7833 ( .A(n6209), .ZN(n6210) );
  NAND2_X1 U7834 ( .A1(n7995), .A2(n8550), .ZN(n7951) );
  OR2_X1 U7835 ( .A1(n8809), .A2(n8307), .ZN(n8552) );
  OR2_X1 U7836 ( .A1(n7951), .A2(n8552), .ZN(n6212) );
  INV_X1 U7837 ( .A(n7955), .ZN(n6213) );
  NAND2_X1 U7838 ( .A1(n7647), .A2(n7968), .ZN(n6215) );
  OR2_X1 U7839 ( .A1(n5952), .A2(n7648), .ZN(n6214) );
  NAND2_X1 U7840 ( .A1(n6216), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7841 ( .A1(n6228), .A2(n6217), .ZN(n8537) );
  NAND2_X1 U7842 ( .A1(n8537), .A2(n6139), .ZN(n6222) );
  INV_X1 U7843 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U7844 ( .A1(n4423), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6219) );
  INV_X1 U7845 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9016) );
  OR2_X1 U7846 ( .A1(n7679), .A2(n9016), .ZN(n6218) );
  OAI211_X1 U7847 ( .C1(n8952), .C2(n6323), .A(n6219), .B(n6218), .ZN(n6220)
         );
  INV_X1 U7848 ( .A(n6220), .ZN(n6221) );
  INV_X1 U7849 ( .A(n8545), .ZN(n6223) );
  NAND2_X1 U7850 ( .A1(n8797), .A2(n6223), .ZN(n7957) );
  NAND2_X1 U7851 ( .A1(n8116), .A2(n7968), .ZN(n6225) );
  OR2_X1 U7852 ( .A1(n5952), .A2(n9007), .ZN(n6224) );
  INV_X1 U7853 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7854 ( .A1(n6228), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7855 ( .A1(n6238), .A2(n6229), .ZN(n8529) );
  NAND2_X1 U7856 ( .A1(n8529), .A2(n6139), .ZN(n6234) );
  INV_X1 U7857 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U7858 ( .A1(n4982), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7859 ( .A1(n4423), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6230) );
  OAI211_X1 U7860 ( .C1(n8528), .C2(n6323), .A(n6231), .B(n6230), .ZN(n6232)
         );
  INV_X1 U7861 ( .A(n6232), .ZN(n6233) );
  NAND2_X1 U7862 ( .A1(n8875), .A2(n7968), .ZN(n6237) );
  OR2_X1 U7863 ( .A1(n5952), .A2(n6235), .ZN(n6236) );
  NAND2_X1 U7864 ( .A1(n6238), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7865 ( .A1(n6250), .A2(n6239), .ZN(n8520) );
  NAND2_X1 U7866 ( .A1(n8520), .A2(n6139), .ZN(n6244) );
  INV_X1 U7867 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U7868 ( .A1(n4423), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7869 ( .A1(n6260), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6240) );
  OAI211_X1 U7870 ( .C1(n8708), .C2(n7679), .A(n6241), .B(n6240), .ZN(n6242)
         );
  INV_X1 U7871 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7872 ( .A1(n8785), .A2(n8336), .ZN(n7961) );
  NAND2_X1 U7873 ( .A1(n8871), .A2(n7968), .ZN(n6247) );
  OR2_X1 U7874 ( .A1(n5952), .A2(n6245), .ZN(n6246) );
  INV_X1 U7875 ( .A(n8779), .ZN(n7981) );
  INV_X1 U7876 ( .A(n6250), .ZN(n6249) );
  INV_X1 U7877 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7878 ( .A1(n6249), .A2(n6248), .ZN(n7669) );
  NAND2_X1 U7879 ( .A1(n6250), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7880 ( .A1(n7669), .A2(n6251), .ZN(n8511) );
  NAND2_X1 U7881 ( .A1(n8511), .A2(n6139), .ZN(n6256) );
  INV_X1 U7882 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U7883 ( .A1(n6260), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7884 ( .A1(n5943), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6252) );
  OAI211_X1 U7885 ( .C1(n7679), .C2(n9003), .A(n6253), .B(n6252), .ZN(n6254)
         );
  INV_X1 U7886 ( .A(n6254), .ZN(n6255) );
  NOR2_X1 U7887 ( .A1(n7981), .A2(n8517), .ZN(n6257) );
  INV_X1 U7888 ( .A(n8517), .ZN(n6328) );
  NAND2_X1 U7889 ( .A1(n8192), .A2(n7968), .ZN(n6259) );
  OR2_X1 U7890 ( .A1(n5952), .A2(n8868), .ZN(n6258) );
  INV_X1 U7891 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U7892 ( .A1(n4982), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7893 ( .A1(n6260), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6261) );
  OAI211_X1 U7894 ( .C1(n6263), .C2(n8988), .A(n6262), .B(n6261), .ZN(n6264)
         );
  INV_X1 U7895 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U7896 ( .A1(n7684), .A2(n6265), .ZN(n8508) );
  INV_X1 U7897 ( .A(n8508), .ZN(n6266) );
  NAND2_X1 U7898 ( .A1(n7675), .A2(n6266), .ZN(n7971) );
  XNOR2_X1 U7899 ( .A(n7990), .B(n4632), .ZN(n7672) );
  NAND2_X1 U7900 ( .A1(n6267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6268) );
  MUX2_X1 U7901 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6268), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6270) );
  NAND2_X1 U7902 ( .A1(n6270), .A2(n6269), .ZN(n8037) );
  INV_X1 U7903 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U7904 ( .A1(n6272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6273) );
  MUX2_X1 U7905 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6273), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n6274) );
  INV_X1 U7906 ( .A(n6274), .ZN(n6277) );
  INV_X1 U7907 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U7908 ( .A1(n6269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6278) );
  OR2_X1 U7909 ( .A1(n6739), .A2(n7973), .ZN(n6595) );
  NAND2_X1 U7910 ( .A1(n6595), .A2(n8764), .ZN(n6566) );
  NAND2_X1 U7911 ( .A1(n8485), .A2(n8043), .ZN(n6373) );
  AND2_X1 U7912 ( .A1(n6739), .A2(n6373), .ZN(n6279) );
  OR2_X1 U7913 ( .A1(n6566), .A2(n6279), .ZN(n7446) );
  NAND2_X1 U7914 ( .A1(n6363), .A2(n8037), .ZN(n10312) );
  OR2_X1 U7915 ( .A1(n10312), .A2(n8043), .ZN(n7486) );
  AND2_X1 U7916 ( .A1(n7446), .A2(n7486), .ZN(n6941) );
  OR2_X1 U7917 ( .A1(n7672), .A2(n6941), .ZN(n6331) );
  NAND2_X1 U7918 ( .A1(n5917), .A2(n6690), .ZN(n6689) );
  NAND2_X1 U7919 ( .A1(n6998), .A2(n6741), .ZN(n6999) );
  INV_X1 U7920 ( .A(n8003), .ZN(n7847) );
  INV_X1 U7921 ( .A(n6890), .ZN(n6947) );
  NAND2_X1 U7922 ( .A1(n6997), .A2(n6947), .ZN(n6795) );
  NAND2_X1 U7923 ( .A1(n6794), .A2(n6795), .ZN(n6282) );
  NAND2_X1 U7924 ( .A1(n6282), .A2(n8005), .ZN(n6793) );
  INV_X1 U7925 ( .A(n6802), .ZN(n6943) );
  NAND2_X1 U7926 ( .A1(n7060), .A2(n6943), .ZN(n6283) );
  NAND2_X1 U7927 ( .A1(n6793), .A2(n6283), .ZN(n7059) );
  NOR2_X1 U7928 ( .A1(n8364), .A2(n7112), .ZN(n7058) );
  NAND2_X1 U7929 ( .A1(n8364), .A2(n7112), .ZN(n7056) );
  OR2_X1 U7930 ( .A1(n8363), .A2(n7014), .ZN(n6284) );
  NAND2_X1 U7931 ( .A1(n8363), .A2(n7014), .ZN(n6285) );
  NAND2_X1 U7932 ( .A1(n7880), .A2(n7885), .ZN(n8009) );
  INV_X1 U7933 ( .A(n10306), .ZN(n7396) );
  NAND2_X1 U7934 ( .A1(n7396), .A2(n7336), .ZN(n7215) );
  AND2_X1 U7935 ( .A1(n8009), .A2(n7215), .ZN(n6287) );
  NAND2_X1 U7936 ( .A1(n7214), .A2(n6287), .ZN(n7213) );
  NAND2_X1 U7937 ( .A1(n7340), .A2(n8361), .ZN(n6288) );
  NAND2_X1 U7938 ( .A1(n7213), .A2(n6288), .ZN(n7303) );
  AND2_X1 U7939 ( .A1(n7490), .A2(n7425), .ZN(n6289) );
  OR2_X1 U7940 ( .A1(n7490), .A2(n7425), .ZN(n6290) );
  INV_X1 U7941 ( .A(n7623), .ZN(n8360) );
  NOR2_X1 U7942 ( .A1(n7450), .A2(n8360), .ZN(n6291) );
  INV_X1 U7943 ( .A(n7450), .ZN(n7470) );
  INV_X1 U7944 ( .A(n7599), .ZN(n8359) );
  NAND2_X1 U7945 ( .A1(n7633), .A2(n8359), .ZN(n6292) );
  AND2_X1 U7946 ( .A1(n7906), .A2(n8688), .ZN(n6294) );
  NOR2_X1 U7947 ( .A1(n8861), .A2(n8358), .ZN(n7904) );
  NAND2_X1 U7948 ( .A1(n8861), .A2(n8358), .ZN(n7902) );
  AND2_X1 U7949 ( .A1(n8855), .A2(n8686), .ZN(n6296) );
  OR2_X1 U7950 ( .A1(n8855), .A2(n8686), .ZN(n6295) );
  NAND2_X1 U7951 ( .A1(n7916), .A2(n6297), .ZN(n8658) );
  NAND2_X1 U7952 ( .A1(n8657), .A2(n8658), .ZN(n6299) );
  OR2_X1 U7953 ( .A1(n8848), .A2(n8357), .ZN(n6298) );
  INV_X1 U7954 ( .A(n8647), .ZN(n8616) );
  NAND2_X1 U7955 ( .A1(n8631), .A2(n8616), .ZN(n8612) );
  INV_X1 U7956 ( .A(n8612), .ZN(n6300) );
  NOR2_X1 U7957 ( .A1(n6300), .A2(n8635), .ZN(n6302) );
  NAND2_X1 U7958 ( .A1(n8842), .A2(n8659), .ZN(n8611) );
  AND2_X1 U7959 ( .A1(n8611), .A2(n8612), .ZN(n6301) );
  OR2_X1 U7960 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  OR2_X1 U7961 ( .A1(n8737), .A2(n8637), .ZN(n6305) );
  AND2_X1 U7962 ( .A1(n8737), .A2(n8637), .ZN(n6304) );
  NAND2_X1 U7963 ( .A1(n8829), .A2(n8615), .ZN(n6307) );
  NOR2_X1 U7964 ( .A1(n8829), .A2(n8615), .ZN(n6306) );
  INV_X1 U7965 ( .A(n8579), .ZN(n8605) );
  NAND2_X1 U7966 ( .A1(n7945), .A2(n7944), .ZN(n8582) );
  INV_X1 U7967 ( .A(n8251), .ZN(n8820) );
  AOI22_X1 U7968 ( .A1(n8576), .A2(n8582), .B1(n8085), .B2(n8820), .ZN(n8569)
         );
  OAI21_X1 U7969 ( .B1(n8569), .B2(n8568), .A(n6308), .ZN(n8559) );
  INV_X1 U7970 ( .A(n8809), .ZN(n6309) );
  NOR2_X1 U7971 ( .A1(n8791), .A2(n8535), .ZN(n6311) );
  INV_X1 U7972 ( .A(n8791), .ZN(n6310) );
  INV_X1 U7973 ( .A(n8516), .ZN(n6313) );
  AOI21_X2 U7974 ( .B1(n6313), .B2(n6312), .A(n5004), .ZN(n8507) );
  NAND2_X1 U7975 ( .A1(n7981), .A2(n6328), .ZN(n6314) );
  AOI22_X1 U7976 ( .A1(n8507), .A2(n6314), .B1(n8779), .B2(n8517), .ZN(n6315)
         );
  XNOR2_X1 U7977 ( .A(n6315), .B(n8029), .ZN(n6330) );
  OR2_X1 U7978 ( .A1(n8485), .A2(n4857), .ZN(n6317) );
  NAND2_X1 U7979 ( .A1(n8034), .A2(n8038), .ZN(n6316) );
  INV_X1 U7980 ( .A(n6417), .ZN(n8040) );
  NAND2_X1 U7981 ( .A1(n6414), .A2(n8040), .ZN(n6319) );
  AND2_X1 U7982 ( .A1(n6385), .A2(n6319), .ZN(n6731) );
  INV_X1 U7983 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7984 ( .A1(n4423), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6322) );
  INV_X1 U7985 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6320) );
  OR2_X1 U7986 ( .A1(n7679), .A2(n6320), .ZN(n6321) );
  OAI211_X1 U7987 ( .C1(n6324), .C2(n6323), .A(n6322), .B(n6321), .ZN(n6325)
         );
  INV_X1 U7988 ( .A(n6325), .ZN(n6326) );
  NAND2_X1 U7989 ( .A1(n6385), .A2(P2_B_REG_SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7990 ( .A1(n8685), .A2(n6327), .ZN(n7685) );
  OAI22_X1 U7991 ( .A1(n6328), .A2(n8671), .B1(n7976), .B2(n7685), .ZN(n6329)
         );
  NAND2_X1 U7992 ( .A1(n6331), .A2(n7668), .ZN(n6380) );
  OR2_X1 U7993 ( .A1(n6332), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7994 ( .A1(n6332), .A2(n6333), .ZN(n6335) );
  XNOR2_X1 U7995 ( .A(n7651), .B(P2_B_REG_SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7996 ( .A1(n6335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7997 ( .A1(n6338), .A2(n7649), .ZN(n6343) );
  NAND2_X1 U7998 ( .A1(n6340), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7999 ( .A1(n8879), .A2(n7651), .ZN(n6451) );
  INV_X1 U8000 ( .A(n6737), .ZN(n6375) );
  OR2_X1 U8001 ( .A1(n6344), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8002 ( .A1(n7649), .A2(n8879), .ZN(n6454) );
  NAND2_X1 U8003 ( .A1(n6345), .A2(n6454), .ZN(n6560) );
  INV_X1 U8004 ( .A(n6560), .ZN(n6346) );
  NOR2_X1 U8005 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .ZN(
        n6350) );
  NOR4_X1 U8006 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6349) );
  NOR4_X1 U8007 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6348) );
  NOR4_X1 U8008 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6347) );
  NAND4_X1 U8009 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n6356)
         );
  NOR4_X1 U8010 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6354) );
  NOR4_X1 U8011 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6353) );
  NOR4_X1 U8012 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6352) );
  NOR4_X1 U8013 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6351) );
  NAND4_X1 U8014 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6355)
         );
  NOR2_X1 U8015 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  NAND2_X1 U8016 ( .A1(n6371), .A2(n6372), .ZN(n6584) );
  INV_X1 U8017 ( .A(n6584), .ZN(n6361) );
  NOR2_X1 U8018 ( .A1(n8879), .A2(n7651), .ZN(n6359) );
  INV_X1 U8019 ( .A(n7649), .ZN(n6358) );
  NAND2_X1 U8020 ( .A1(n6359), .A2(n6358), .ZN(n6587) );
  NAND2_X1 U8021 ( .A1(n6275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6360) );
  XNOR2_X1 U8022 ( .A(n6360), .B(n5895), .ZN(n6586) );
  NOR3_X1 U8023 ( .A1(n4857), .A2(n8034), .A3(n8037), .ZN(n6362) );
  NAND2_X1 U8024 ( .A1(n6363), .A2(n6362), .ZN(n6578) );
  NAND2_X1 U8025 ( .A1(n6595), .A2(n6578), .ZN(n6364) );
  NAND2_X1 U8026 ( .A1(n6577), .A2(n6364), .ZN(n6368) );
  AND3_X1 U8027 ( .A1(n6737), .A2(n6560), .A3(n6372), .ZN(n6585) );
  NAND2_X1 U8028 ( .A1(n6585), .A2(n6594), .ZN(n6582) );
  NAND2_X1 U8029 ( .A1(n10312), .A2(n8766), .ZN(n8547) );
  NOR2_X1 U8030 ( .A1(n7977), .A2(n8766), .ZN(n6365) );
  NAND2_X1 U8031 ( .A1(n6578), .A2(n6365), .ZN(n6575) );
  NAND2_X1 U8032 ( .A1(n8547), .A2(n6575), .ZN(n6583) );
  INV_X1 U8033 ( .A(n6583), .ZN(n6366) );
  INV_X1 U8034 ( .A(n6369), .ZN(n6370) );
  INV_X1 U8035 ( .A(n7675), .ZN(n6382) );
  NAND2_X1 U8036 ( .A1(n6370), .A2(n4499), .ZN(P2_U3456) );
  INV_X1 U8037 ( .A(n6371), .ZN(n6379) );
  NAND2_X1 U8038 ( .A1(n6739), .A2(n7977), .ZN(n6588) );
  NAND3_X1 U8039 ( .A1(n6594), .A2(n6372), .A3(n6588), .ZN(n6559) );
  NOR2_X1 U8040 ( .A1(n7486), .A2(n8034), .ZN(n6565) );
  NOR2_X1 U8041 ( .A1(n6559), .A2(n6565), .ZN(n6378) );
  INV_X1 U8042 ( .A(n6373), .ZN(n6374) );
  AOI21_X1 U8043 ( .B1(n6374), .B2(n8038), .A(n7977), .ZN(n6377) );
  NAND2_X1 U8044 ( .A1(n6375), .A2(n6377), .ZN(n6376) );
  OAI21_X1 U8045 ( .B1(n6377), .B2(n6560), .A(n6376), .ZN(n6563) );
  AND3_X2 U8046 ( .A1(n6379), .A2(n6378), .A3(n6563), .ZN(n8772) );
  INV_X1 U8047 ( .A(n6381), .ZN(n6383) );
  NAND2_X1 U8048 ( .A1(n8772), .A2(n8766), .ZN(n8742) );
  NAND2_X1 U8049 ( .A1(n6383), .A2(n4500), .ZN(P2_U3488) );
  NAND2_X1 U8050 ( .A1(n6587), .A2(n7973), .ZN(n6384) );
  NAND2_X1 U8051 ( .A1(n6384), .A2(n6586), .ZN(n6418) );
  NAND2_X1 U8052 ( .A1(n6418), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U8053 ( .A1(n6386), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8054 ( .A(n6456), .ZN(n6387) );
  INV_X2 U8055 ( .A(n8368), .ZN(P2_U3893) );
  INV_X1 U8056 ( .A(n6388), .ZN(n6389) );
  OR2_X1 U8057 ( .A1(n6665), .A2(n6389), .ZN(n9394) );
  XNOR2_X1 U8058 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8059 ( .A1(n4425), .A2(P2_U3151), .ZN(n9175) );
  NOR2_X1 U8060 ( .A1(n4424), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9173) );
  INV_X2 U8061 ( .A(n9173), .ZN(n8878) );
  OAI222_X1 U8062 ( .A1(n8874), .A2(n6393), .B1(n6458), .B2(P2_U3151), .C1(
        n5013), .C2(n8878), .ZN(P2_U3294) );
  OAI222_X1 U8063 ( .A1(n8878), .A2(n5024), .B1(n6517), .B2(P2_U3151), .C1(
        n8874), .C2(n6404), .ZN(P2_U3292) );
  OAI222_X1 U8064 ( .A1(n8878), .A2(n6390), .B1(n4417), .B2(P2_U3151), .C1(
        n8874), .C2(n6394), .ZN(P2_U3293) );
  OAI222_X1 U8065 ( .A1(n8878), .A2(n6391), .B1(n8874), .B2(n6396), .C1(
        P2_U3151), .C2(n6542), .ZN(P2_U3291) );
  NAND2_X1 U8066 ( .A1(n4425), .A2(P1_U3086), .ZN(n10009) );
  NOR2_X1 U8067 ( .A1(n6392), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10013) );
  OAI222_X1 U8068 ( .A1(n10009), .A2(n9038), .B1(n8174), .B2(n6393), .C1(
        P1_U3086), .C2(n6620), .ZN(P1_U3354) );
  OAI222_X1 U8069 ( .A1(n10009), .A2(n6395), .B1(n8174), .B2(n6394), .C1(
        P1_U3086), .C2(n9414), .ZN(P1_U3353) );
  OAI222_X1 U8070 ( .A1(P1_U3086), .A2(n9442), .B1(n8174), .B2(n6396), .C1(
        n10009), .C2(n5164), .ZN(P1_U3351) );
  OAI222_X1 U8071 ( .A1(n8874), .A2(n6399), .B1(n6554), .B2(P2_U3151), .C1(
        n6397), .C2(n8878), .ZN(P2_U3290) );
  OAI222_X1 U8072 ( .A1(n10009), .A2(n6400), .B1(n8174), .B2(n6399), .C1(
        P1_U3086), .C2(n6398), .ZN(P1_U3350) );
  OAI222_X1 U8073 ( .A1(n8874), .A2(n6403), .B1(n6721), .B2(P2_U3151), .C1(
        n6401), .C2(n8878), .ZN(P2_U3289) );
  OAI222_X1 U8074 ( .A1(P1_U3086), .A2(n10105), .B1(n8174), .B2(n6403), .C1(
        n6402), .C2(n10009), .ZN(P1_U3349) );
  INV_X1 U8075 ( .A(n10009), .ZN(n6483) );
  INV_X1 U8076 ( .A(n6483), .ZN(n10018) );
  OAI222_X1 U8077 ( .A1(n10018), .A2(n6405), .B1(n8174), .B2(n6404), .C1(
        P1_U3086), .C2(n9425), .ZN(P1_U3352) );
  OAI222_X1 U8078 ( .A1(n8874), .A2(n6407), .B1(n8878), .B2(n6001), .C1(
        P2_U3151), .C2(n6859), .ZN(P2_U3288) );
  OAI222_X1 U8079 ( .A1(P1_U3086), .A2(n6613), .B1(n8174), .B2(n6407), .C1(
        n6406), .C2(n10009), .ZN(P1_U3348) );
  INV_X1 U8080 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9126) );
  OAI222_X1 U8081 ( .A1(n8878), .A2(n9126), .B1(n8874), .B2(n6408), .C1(
        P2_U3151), .C2(n4536), .ZN(P2_U3287) );
  OAI222_X1 U8082 ( .A1(n10050), .A2(P1_U3086), .B1(n8174), .B2(n6408), .C1(
        n9131), .C2(n10009), .ZN(P1_U3347) );
  INV_X1 U8083 ( .A(n6409), .ZN(n6410) );
  INV_X1 U8084 ( .A(n7164), .ZN(n7171) );
  OAI222_X1 U8085 ( .A1(n8874), .A2(n6410), .B1(n7171), .B2(P2_U3151), .C1(
        n9083), .C2(n8878), .ZN(P2_U3286) );
  INV_X1 U8086 ( .A(n6640), .ZN(n10074) );
  OAI222_X1 U8087 ( .A1(P1_U3086), .A2(n10074), .B1(n8174), .B2(n6410), .C1(
        n6411), .C2(n10009), .ZN(P1_U3346) );
  INV_X1 U8088 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9120) );
  NOR2_X1 U8089 ( .A1(n6450), .A2(n9120), .ZN(P2_U3252) );
  INV_X1 U8090 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9017) );
  NOR2_X1 U8091 ( .A1(n6450), .A2(n9017), .ZN(P2_U3250) );
  INV_X1 U8092 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9138) );
  NOR2_X1 U8093 ( .A1(n6450), .A2(n9138), .ZN(P2_U3235) );
  INV_X1 U8094 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U8095 ( .A1(n6450), .A2(n8964), .ZN(P2_U3261) );
  INV_X1 U8096 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9006) );
  NOR2_X1 U8097 ( .A1(n6450), .A2(n9006), .ZN(P2_U3249) );
  INV_X1 U8098 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9135) );
  NOR2_X1 U8099 ( .A1(n6450), .A2(n9135), .ZN(P2_U3240) );
  INV_X1 U8100 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n8954) );
  NOR2_X1 U8101 ( .A1(n6450), .A2(n8954), .ZN(P2_U3238) );
  INV_X1 U8102 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9004) );
  NOR2_X1 U8103 ( .A1(n6450), .A2(n9004), .ZN(P2_U3260) );
  INV_X1 U8104 ( .A(n6642), .ZN(n10033) );
  INV_X1 U8105 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9137) );
  OAI222_X1 U8106 ( .A1(P1_U3086), .A2(n10033), .B1(n8174), .B2(n9172), .C1(
        n9137), .C2(n10009), .ZN(P1_U3345) );
  MUX2_X1 U8107 ( .A(n6411), .B(n7442), .S(P2_U3893), .Z(n6412) );
  INV_X1 U8108 ( .A(n6412), .ZN(P2_U3500) );
  INV_X1 U8109 ( .A(n7060), .ZN(n6916) );
  NAND2_X1 U8110 ( .A1(n6916), .A2(P2_U3893), .ZN(n6413) );
  OAI21_X1 U8111 ( .B1(P2_U3893), .B2(n5164), .A(n6413), .ZN(P2_U3495) );
  NOR2_X1 U8112 ( .A1(n8489), .A2(P2_U3151), .ZN(n8876) );
  NAND2_X1 U8113 ( .A1(n8876), .A2(n6418), .ZN(n6415) );
  MUX2_X1 U8114 ( .A(n8368), .B(n6415), .S(n6417), .Z(n8486) );
  INV_X1 U8115 ( .A(n6586), .ZN(n7496) );
  NOR2_X1 U8116 ( .A1(n6587), .A2(n7496), .ZN(n6416) );
  INV_X1 U8117 ( .A(n8441), .ZN(n8482) );
  AOI22_X1 U8118 ( .A1(n8482), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6422) );
  NOR2_X1 U8119 ( .A1(n6417), .A2(P2_U3151), .ZN(n8872) );
  AND2_X1 U8120 ( .A1(n6418), .A2(n8872), .ZN(n6438) );
  INV_X1 U8121 ( .A(n8494), .ZN(n8382) );
  MUX2_X1 U8122 ( .A(n6572), .B(n6439), .S(n8489), .Z(n6419) );
  NAND2_X1 U8123 ( .A1(n6419), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6460) );
  OAI21_X1 U8124 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6419), .A(n6460), .ZN(n6420) );
  OAI21_X1 U8125 ( .B1(n6438), .B2(n8382), .A(n6420), .ZN(n6421) );
  OAI211_X1 U8126 ( .C1(n8486), .C2(n6440), .A(n6422), .B(n6421), .ZN(P2_U3182) );
  INV_X1 U8127 ( .A(n6450), .ZN(n6423) );
  AND2_X1 U8128 ( .A1(n6423), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8129 ( .A1(n6423), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8130 ( .A1(n6423), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8131 ( .A1(n6423), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8132 ( .A1(n6423), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8133 ( .A1(n6423), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8134 ( .A1(n6423), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  INV_X1 U8135 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9092) );
  INV_X1 U8136 ( .A(n6424), .ZN(n6426) );
  OAI222_X1 U8137 ( .A1(n8878), .A2(n9092), .B1(n8874), .B2(n6426), .C1(
        P2_U3151), .C2(n7249), .ZN(P2_U3284) );
  INV_X1 U8138 ( .A(n6644), .ZN(n10120) );
  INV_X1 U8139 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6425) );
  OAI222_X1 U8140 ( .A1(n10120), .A2(P1_U3086), .B1(n8174), .B2(n6426), .C1(
        n6425), .C2(n10009), .ZN(P1_U3344) );
  NAND2_X1 U8141 ( .A1(n6842), .A2(n6427), .ZN(n6428) );
  AND2_X1 U8142 ( .A1(n6429), .A2(n6428), .ZN(n6479) );
  INV_X1 U8143 ( .A(n6479), .ZN(n6430) );
  INV_X1 U8144 ( .A(n10005), .ZN(n6677) );
  NAND2_X1 U8145 ( .A1(n6677), .A2(n7492), .ZN(n6480) );
  NOR2_X1 U8146 ( .A1(n10138), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8147 ( .A(n7254), .ZN(n7363) );
  INV_X1 U8148 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6431) );
  OAI222_X1 U8149 ( .A1(n8874), .A2(n6432), .B1(n7363), .B2(P2_U3151), .C1(
        n6431), .C2(n8878), .ZN(P2_U3283) );
  INV_X1 U8150 ( .A(n9463), .ZN(n6652) );
  INV_X1 U8151 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9063) );
  OAI222_X1 U8152 ( .A1(P1_U3086), .A2(n6652), .B1(n8174), .B2(n6432), .C1(
        n9063), .C2(n10018), .ZN(P1_U3343) );
  MUX2_X1 U8153 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6318), .Z(n6459) );
  XNOR2_X1 U8154 ( .A(n6459), .B(n6447), .ZN(n6461) );
  XNOR2_X1 U8155 ( .A(n6461), .B(n6460), .ZN(n6449) );
  INV_X1 U8156 ( .A(n6438), .ZN(n6433) );
  AND2_X1 U8157 ( .A1(n6440), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8158 ( .A1(n5925), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6463) );
  OAI21_X1 U8159 ( .B1(n6458), .B2(n6434), .A(n6463), .ZN(n6436) );
  INV_X1 U8160 ( .A(n6464), .ZN(n6435) );
  AOI21_X1 U8161 ( .B1(n6697), .B2(n6436), .A(n6435), .ZN(n6437) );
  OAI22_X1 U8162 ( .A1(n8501), .A2(n6437), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5918), .ZN(n6446) );
  INV_X1 U8163 ( .A(n8499), .ZN(n7053) );
  OAI21_X1 U8164 ( .B1(n6441), .B2(n6439), .A(n6458), .ZN(n6443) );
  NAND3_X1 U8165 ( .A1(n6441), .A2(P2_REG1_REG_0__SCAN_IN), .A3(n6440), .ZN(
        n6442) );
  NAND2_X1 U8166 ( .A1(n6443), .A2(n6442), .ZN(n6469) );
  XOR2_X1 U8167 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6469), .Z(n6444) );
  INV_X1 U8168 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10346) );
  OAI22_X1 U8169 ( .A1(n7053), .A2(n6444), .B1(n10346), .B2(n8441), .ZN(n6445)
         );
  AOI211_X1 U8170 ( .C1(n6447), .C2(n8450), .A(n6446), .B(n6445), .ZN(n6448)
         );
  OAI21_X1 U8171 ( .B1(n8494), .B2(n6449), .A(n6448), .ZN(P2_U3183) );
  AND2_X1 U8172 ( .A1(n6423), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8173 ( .A1(n6423), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8174 ( .A1(n6423), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8175 ( .A1(n6423), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8176 ( .A1(n6423), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8177 ( .A1(n6423), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8178 ( .A1(n6423), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8179 ( .A1(n6423), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8180 ( .A1(n6423), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8181 ( .A1(n6423), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8182 ( .A1(n6423), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8183 ( .A1(n6423), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8184 ( .A1(n6423), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8185 ( .A1(n6423), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8186 ( .A1(n6423), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8187 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6453) );
  INV_X1 U8188 ( .A(n6451), .ZN(n6452) );
  AOI22_X1 U8189 ( .A1(n6423), .A2(n6453), .B1(n6456), .B2(n6452), .ZN(
        P2_U3376) );
  INV_X1 U8190 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6457) );
  INV_X1 U8191 ( .A(n6454), .ZN(n6455) );
  AOI22_X1 U8192 ( .A1(n6423), .A2(n6457), .B1(n6456), .B2(n6455), .ZN(
        P2_U3377) );
  AOI22_X1 U8193 ( .A1(n6461), .A2(n6460), .B1(n6459), .B2(n6458), .ZN(n6491)
         );
  MUX2_X1 U8194 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8489), .Z(n6487) );
  XNOR2_X1 U8195 ( .A(n6487), .B(n4417), .ZN(n6490) );
  XNOR2_X1 U8196 ( .A(n6491), .B(n6490), .ZN(n6476) );
  INV_X1 U8197 ( .A(n4417), .ZN(n6489) );
  INV_X1 U8198 ( .A(n8501), .ZN(n8458) );
  XNOR2_X1 U8199 ( .A(n4417), .B(n6462), .ZN(n6466) );
  NAND2_X1 U8200 ( .A1(n6466), .A2(n6465), .ZN(n6495) );
  OAI21_X1 U8201 ( .B1(n6466), .B2(n6465), .A(n6495), .ZN(n6467) );
  NAND2_X1 U8202 ( .A1(n8458), .A2(n6467), .ZN(n6468) );
  OAI21_X1 U8203 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5931), .A(n6468), .ZN(n6474) );
  MUX2_X1 U8204 ( .A(n5932), .B(P2_REG1_REG_2__SCAN_IN), .S(n4417), .Z(n6471)
         );
  AOI22_X1 U8205 ( .A1(n6469), .A2(P2_REG1_REG_1__SCAN_IN), .B1(n5925), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U8206 ( .A1(n6471), .A2(n6470), .ZN(n6500) );
  AOI21_X1 U8207 ( .B1(n6471), .B2(n6470), .A(n6500), .ZN(n6472) );
  INV_X1 U8208 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9155) );
  OAI22_X1 U8209 ( .A1(n7053), .A2(n6472), .B1(n9155), .B2(n8441), .ZN(n6473)
         );
  AOI211_X1 U8210 ( .C1(n6489), .C2(n8450), .A(n6474), .B(n6473), .ZN(n6475)
         );
  OAI21_X1 U8211 ( .B1(n8494), .B2(n6476), .A(n6475), .ZN(P2_U3184) );
  AOI21_X1 U8212 ( .B1(n6647), .B2(n6477), .A(n5381), .ZN(n9411) );
  OAI21_X1 U8213 ( .B1(n6647), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9411), .ZN(
        n6478) );
  XOR2_X1 U8214 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6478), .Z(n6482) );
  NAND2_X1 U8215 ( .A1(n6480), .A2(n6479), .ZN(n6648) );
  AOI22_X1 U8216 ( .A1(n10138), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6481) );
  OAI21_X1 U8217 ( .B1(n6482), .B2(n6648), .A(n6481), .ZN(P1_U3243) );
  AOI22_X1 U8218 ( .A1(n10134), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6483), .ZN(n6484) );
  OAI21_X1 U8219 ( .B1(n6486), .B2(n8174), .A(n6484), .ZN(P1_U3342) );
  INV_X1 U8220 ( .A(n7509), .ZN(n7516) );
  INV_X1 U8221 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6485) );
  OAI222_X1 U8222 ( .A1(n8874), .A2(n6486), .B1(n7516), .B2(P2_U3151), .C1(
        n6485), .C2(n8878), .ZN(P2_U3282) );
  MUX2_X1 U8223 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8489), .Z(n6509) );
  XNOR2_X1 U8224 ( .A(n6509), .B(n6517), .ZN(n6493) );
  INV_X1 U8225 ( .A(n6487), .ZN(n6488) );
  OAI22_X1 U8226 ( .A1(n6491), .A2(n6490), .B1(n6489), .B2(n6488), .ZN(n6492)
         );
  NOR2_X1 U8227 ( .A1(n6492), .A2(n6493), .ZN(n6512) );
  AOI21_X1 U8228 ( .B1(n6493), .B2(n6492), .A(n6512), .ZN(n6506) );
  NAND2_X1 U8229 ( .A1(n4417), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8230 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  INV_X1 U8231 ( .A(n6527), .ZN(n6497) );
  AOI21_X1 U8232 ( .B1(n6889), .B2(n6498), .A(n6497), .ZN(n6499) );
  NAND2_X1 U8233 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6733) );
  OAI21_X1 U8234 ( .B1(n8501), .B2(n6499), .A(n6733), .ZN(n6504) );
  AOI21_X1 U8235 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n4417), .A(n6500), .ZN(
        n6515) );
  XNOR2_X1 U8236 ( .A(n6515), .B(n6517), .ZN(n6518) );
  XOR2_X1 U8237 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6518), .Z(n6502) );
  INV_X1 U8238 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9132) );
  OAI22_X1 U8239 ( .A1(n7053), .A2(n6502), .B1(n9132), .B2(n8441), .ZN(n6503)
         );
  AOI211_X1 U8240 ( .C1(n4880), .C2(n8450), .A(n6504), .B(n6503), .ZN(n6505)
         );
  OAI21_X1 U8241 ( .B1(n6506), .B2(n8494), .A(n6505), .ZN(P2_U3185) );
  NAND2_X1 U8242 ( .A1(n9930), .A2(P1_U3973), .ZN(n6507) );
  OAI21_X1 U8243 ( .B1(P1_U3973), .B2(n6001), .A(n6507), .ZN(P1_U3561) );
  NAND2_X1 U8244 ( .A1(n9870), .A2(P1_U3973), .ZN(n6508) );
  OAI21_X1 U8245 ( .B1(n6162), .B2(P1_U3973), .A(n6508), .ZN(P1_U3574) );
  NOR2_X1 U8246 ( .A1(n6509), .A2(n6517), .ZN(n6511) );
  MUX2_X1 U8247 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8489), .Z(n6540) );
  XNOR2_X1 U8248 ( .A(n6540), .B(n6542), .ZN(n6510) );
  NOR3_X1 U8249 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(n6539) );
  INV_X1 U8250 ( .A(n6539), .ZN(n6514) );
  OAI21_X1 U8251 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6513) );
  NAND3_X1 U8252 ( .A1(n6514), .A2(n8382), .A3(n6513), .ZN(n6532) );
  MUX2_X1 U8253 ( .A(n5954), .B(P2_REG1_REG_4__SCAN_IN), .S(n6542), .Z(n6520)
         );
  INV_X1 U8254 ( .A(n6515), .ZN(n6516) );
  AOI22_X1 U8255 ( .A1(n6518), .A2(P2_REG1_REG_3__SCAN_IN), .B1(n6517), .B2(
        n6516), .ZN(n6519) );
  AOI21_X1 U8256 ( .B1(n6520), .B2(n6519), .A(n6541), .ZN(n6522) );
  INV_X1 U8257 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6521) );
  OAI22_X1 U8258 ( .A1(n7053), .A2(n6522), .B1(n6521), .B2(n8441), .ZN(n6530)
         );
  AND2_X1 U8259 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6767) );
  XNOR2_X1 U8260 ( .A(n6542), .B(n6800), .ZN(n6524) );
  NAND2_X1 U8261 ( .A1(n6523), .A2(n6524), .ZN(n6544) );
  INV_X1 U8262 ( .A(n6524), .ZN(n6526) );
  NAND3_X1 U8263 ( .A1(n6527), .A2(n6526), .A3(n6525), .ZN(n6528) );
  AOI21_X1 U8264 ( .B1(n6544), .B2(n6528), .A(n8501), .ZN(n6529) );
  NOR3_X1 U8265 ( .A1(n6530), .A2(n6767), .A3(n6529), .ZN(n6531) );
  OAI211_X1 U8266 ( .C1(n8486), .C2(n6542), .A(n6532), .B(n6531), .ZN(P2_U3186) );
  INV_X1 U8267 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9073) );
  INV_X1 U8268 ( .A(n6533), .ZN(n6535) );
  INV_X1 U8269 ( .A(n7522), .ZN(n8371) );
  OAI222_X1 U8270 ( .A1(n8878), .A2(n9073), .B1(n8874), .B2(n6535), .C1(
        P2_U3151), .C2(n8371), .ZN(P2_U3281) );
  INV_X1 U8271 ( .A(n10148), .ZN(n9464) );
  INV_X1 U8272 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6534) );
  OAI222_X1 U8273 ( .A1(n9464), .A2(P1_U3086), .B1(n8174), .B2(n6535), .C1(
        n6534), .C2(n10018), .ZN(P1_U3341) );
  NOR2_X1 U8274 ( .A1(n6998), .A2(n8673), .ZN(n6569) );
  INV_X1 U8275 ( .A(n7845), .ZN(n6536) );
  NAND2_X1 U8276 ( .A1(n6742), .A2(n6536), .ZN(n8004) );
  INV_X1 U8277 ( .A(n8004), .ZN(n6567) );
  AOI21_X1 U8278 ( .B1(n6941), .B2(n8668), .A(n6567), .ZN(n6537) );
  AOI211_X1 U8279 ( .C1(n8766), .C2(n5917), .A(n6569), .B(n6537), .ZN(n10321)
         );
  NAND2_X1 U8280 ( .A1(n7564), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6538) );
  OAI21_X1 U8281 ( .B1(n10321), .B2(n7564), .A(n6538), .ZN(P2_U3459) );
  AOI21_X1 U8282 ( .B1(n6540), .B2(n6542), .A(n6539), .ZN(n6704) );
  MUX2_X1 U8283 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8489), .Z(n6701) );
  XNOR2_X1 U8284 ( .A(n6701), .B(n6554), .ZN(n6703) );
  XNOR2_X1 U8285 ( .A(n6704), .B(n6703), .ZN(n6558) );
  INV_X1 U8286 ( .A(n6554), .ZN(n6709) );
  XOR2_X1 U8287 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6711), .Z(n6556) );
  NAND2_X1 U8288 ( .A1(n6542), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8289 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U8290 ( .A1(n6545), .A2(n6554), .ZN(n6714) );
  OR2_X1 U8291 ( .A1(n6545), .A2(n6554), .ZN(n6546) );
  NAND2_X1 U8292 ( .A1(n6547), .A2(n7110), .ZN(n6548) );
  NAND2_X1 U8293 ( .A1(n4873), .A2(n6548), .ZN(n6550) );
  NAND2_X1 U8294 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6917) );
  INV_X1 U8295 ( .A(n6917), .ZN(n6549) );
  AOI21_X1 U8296 ( .B1(n8458), .B2(n6550), .A(n6549), .ZN(n6553) );
  INV_X1 U8297 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6551) );
  OR2_X1 U8298 ( .A1(n8441), .A2(n6551), .ZN(n6552) );
  OAI211_X1 U8299 ( .C1(n8486), .C2(n6554), .A(n6553), .B(n6552), .ZN(n6555)
         );
  AOI21_X1 U8300 ( .B1(n6556), .B2(n8499), .A(n6555), .ZN(n6557) );
  OAI21_X1 U8301 ( .B1(n6558), .B2(n8494), .A(n6557), .ZN(P2_U3187) );
  INV_X1 U8302 ( .A(n6559), .ZN(n6562) );
  NAND2_X1 U8303 ( .A1(n6737), .A2(n6560), .ZN(n6561) );
  NAND2_X1 U8304 ( .A1(n6562), .A2(n6561), .ZN(n6564) );
  OR2_X1 U8305 ( .A1(n6564), .A2(n6563), .ZN(n6570) );
  NOR2_X2 U8306 ( .A1(n6570), .A2(n8547), .ZN(n10307) );
  INV_X1 U8307 ( .A(n10307), .ZN(n8633) );
  NOR2_X1 U8308 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  AOI211_X1 U8309 ( .C1(n10311), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6569), .B(
        n6568), .ZN(n6571) );
  INV_X2 U8310 ( .A(n10310), .ZN(n8678) );
  MUX2_X1 U8311 ( .A(n6572), .B(n6571), .S(n8678), .Z(n6573) );
  OAI21_X1 U8312 ( .B1(n8633), .B2(n6602), .A(n6573), .ZN(P2_U3233) );
  NAND2_X1 U8313 ( .A1(n6577), .A2(n8766), .ZN(n6574) );
  INV_X1 U8314 ( .A(n8353), .ZN(n8311) );
  INV_X1 U8315 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U8316 ( .A1(n6577), .A2(n6576), .ZN(n6581) );
  INV_X1 U8317 ( .A(n6582), .ZN(n6579) );
  INV_X1 U8318 ( .A(n6578), .ZN(n6590) );
  NAND2_X1 U8319 ( .A1(n6579), .A2(n6590), .ZN(n6580) );
  INV_X1 U8320 ( .A(n8348), .ZN(n8315) );
  OR2_X1 U8321 ( .A1(n6582), .A2(n6595), .ZN(n6730) );
  OR2_X1 U8322 ( .A1(n6730), .A2(n6731), .ZN(n8335) );
  INV_X1 U8323 ( .A(n6998), .ZN(n8367) );
  AOI22_X1 U8324 ( .A1(n8315), .A2(n8004), .B1(n8344), .B2(n8367), .ZN(n6601)
         );
  NAND2_X1 U8325 ( .A1(n6584), .A2(n6583), .ZN(n6592) );
  INV_X1 U8326 ( .A(n6585), .ZN(n6597) );
  NAND3_X1 U8327 ( .A1(n6588), .A2(n6587), .A3(n6586), .ZN(n6589) );
  AOI21_X1 U8328 ( .B1(n6597), .B2(n6590), .A(n6589), .ZN(n6591) );
  NAND2_X1 U8329 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  NAND2_X1 U8330 ( .A1(n6593), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6599) );
  INV_X1 U8331 ( .A(n6594), .ZN(n6596) );
  NOR2_X1 U8332 ( .A1(n6596), .A2(n6595), .ZN(n8041) );
  NAND2_X1 U8333 ( .A1(n6597), .A2(n8041), .ZN(n6598) );
  OR2_X1 U8334 ( .A1(n8332), .A2(P2_U3151), .ZN(n8317) );
  NAND2_X1 U8335 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n8317), .ZN(n6600) );
  OAI211_X1 U8336 ( .C1(n8311), .C2(n6602), .A(n6601), .B(n6600), .ZN(P2_U3172) );
  AOI22_X1 U8337 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9463), .B1(n6652), .B2(
        n9800), .ZN(n6616) );
  NAND2_X1 U8338 ( .A1(n6642), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6603) );
  OAI21_X1 U8339 ( .B1(n6642), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6603), .ZN(
        n10025) );
  NOR2_X1 U8340 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6640), .ZN(n6604) );
  AOI21_X1 U8341 ( .B1(n6640), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6604), .ZN(
        n10066) );
  MUX2_X1 U8342 ( .A(n5472), .B(P1_REG2_REG_2__SCAN_IN), .S(n9414), .Z(n9421)
         );
  AND2_X1 U8343 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9407) );
  INV_X1 U8344 ( .A(n6620), .ZN(n9401) );
  NAND2_X1 U8345 ( .A1(n9401), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8346 ( .A1(n9396), .A2(n6605), .ZN(n9420) );
  NAND2_X1 U8347 ( .A1(n9421), .A2(n9420), .ZN(n9419) );
  INV_X1 U8348 ( .A(n9414), .ZN(n6622) );
  NAND2_X1 U8349 ( .A1(n6622), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8350 ( .A1(n9419), .A2(n6606), .ZN(n9434) );
  MUX2_X1 U8351 ( .A(n6607), .B(P1_REG2_REG_3__SCAN_IN), .S(n9425), .Z(n9435)
         );
  NAND2_X1 U8352 ( .A1(n9434), .A2(n9435), .ZN(n9433) );
  OR2_X1 U8353 ( .A1(n9425), .A2(n6607), .ZN(n6608) );
  NAND2_X1 U8354 ( .A1(n9433), .A2(n6608), .ZN(n9445) );
  XNOR2_X1 U8355 ( .A(n9442), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U8356 ( .A1(n9445), .A2(n9446), .ZN(n9444) );
  INV_X1 U8357 ( .A(n9442), .ZN(n6626) );
  NAND2_X1 U8358 ( .A1(n6626), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U8359 ( .A1(n9444), .A2(n6609), .ZN(n10084) );
  OR2_X1 U8360 ( .A1(n10091), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8361 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10091), .ZN(n6610) );
  AND2_X1 U8362 ( .A1(n6611), .A2(n6610), .ZN(n10085) );
  NAND2_X1 U8363 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6633), .ZN(n6612) );
  OAI21_X1 U8364 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6633), .A(n6612), .ZN(
        n10097) );
  AOI22_X1 U8365 ( .A1(n10045), .A2(n5497), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6613), .ZN(n10042) );
  NOR2_X1 U8366 ( .A1(n4454), .A2(n10042), .ZN(n10041) );
  NOR2_X1 U8367 ( .A1(n10050), .A2(n10182), .ZN(n6614) );
  NAND2_X1 U8368 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  OAI21_X1 U8369 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6640), .A(n10064), .ZN(
        n10024) );
  NOR2_X1 U8370 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  AOI22_X1 U8371 ( .A1(n6644), .A2(n7612), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n10120), .ZN(n10111) );
  OAI21_X1 U8372 ( .B1(n6616), .B2(n6615), .A(n9462), .ZN(n6654) );
  OR2_X1 U8373 ( .A1(n5381), .A2(n10021), .ZN(n6617) );
  OR2_X1 U8374 ( .A1(n6642), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8375 ( .A1(n6642), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8376 ( .A1(n6619), .A2(n6618), .ZN(n10028) );
  XNOR2_X1 U8377 ( .A(n10050), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U8378 ( .A1(n10045), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U8379 ( .A(n5471), .B(P1_REG1_REG_2__SCAN_IN), .S(n9414), .Z(n9418)
         );
  MUX2_X1 U8380 ( .A(n5457), .B(P1_REG1_REG_1__SCAN_IN), .S(n6620), .Z(n9400)
         );
  AND2_X1 U8381 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9399) );
  NAND2_X1 U8382 ( .A1(n9400), .A2(n9399), .ZN(n9398) );
  NAND2_X1 U8383 ( .A1(n9401), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U8384 ( .A1(n9398), .A2(n6621), .ZN(n9417) );
  NAND2_X1 U8385 ( .A1(n9418), .A2(n9417), .ZN(n9416) );
  NAND2_X1 U8386 ( .A1(n6622), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8387 ( .A1(n9416), .A2(n6623), .ZN(n9431) );
  INV_X1 U8388 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6624) );
  MUX2_X1 U8389 ( .A(n6624), .B(P1_REG1_REG_3__SCAN_IN), .S(n9425), .Z(n9432)
         );
  NAND2_X1 U8390 ( .A1(n9431), .A2(n9432), .ZN(n9430) );
  OR2_X1 U8391 ( .A1(n9425), .A2(n6624), .ZN(n6625) );
  NAND2_X1 U8392 ( .A1(n9430), .A2(n6625), .ZN(n9448) );
  XNOR2_X1 U8393 ( .A(n9442), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U8394 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
  NAND2_X1 U8395 ( .A1(n6626), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8396 ( .A1(n9447), .A2(n6627), .ZN(n10079) );
  OR2_X1 U8397 ( .A1(n10091), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U8398 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10091), .ZN(n6628) );
  AND2_X1 U8399 ( .A1(n6629), .A2(n6628), .ZN(n10080) );
  AND2_X1 U8400 ( .A1(n10079), .A2(n10080), .ZN(n10081) );
  AND2_X1 U8401 ( .A1(n10091), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U8402 ( .A1(n10081), .A2(n6630), .ZN(n10101) );
  OR2_X1 U8403 ( .A1(n6633), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8404 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6633), .ZN(n6631) );
  NAND2_X1 U8405 ( .A1(n6632), .A2(n6631), .ZN(n10100) );
  NOR2_X1 U8406 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  AOI21_X1 U8407 ( .B1(n6633), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10099), .ZN(
        n10040) );
  MUX2_X1 U8408 ( .A(n6634), .B(P1_REG1_REG_7__SCAN_IN), .S(n10045), .Z(n10039) );
  NOR2_X1 U8409 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  INV_X1 U8410 ( .A(n10038), .ZN(n6635) );
  NAND2_X1 U8411 ( .A1(n6636), .A2(n6635), .ZN(n10051) );
  AND2_X1 U8412 ( .A1(n10052), .A2(n10051), .ZN(n10053) );
  NOR2_X1 U8413 ( .A1(n10050), .A2(n6637), .ZN(n6638) );
  NOR2_X1 U8414 ( .A1(n10053), .A2(n6638), .ZN(n10069) );
  NOR2_X1 U8415 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6640), .ZN(n6639) );
  AOI21_X1 U8416 ( .B1(n6640), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6639), .ZN(
        n10070) );
  NAND2_X1 U8417 ( .A1(n10069), .A2(n10070), .ZN(n10068) );
  OR2_X1 U8418 ( .A1(n6640), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8419 ( .A1(n10068), .A2(n6641), .ZN(n10029) );
  NOR2_X1 U8420 ( .A1(n10028), .A2(n10029), .ZN(n10027) );
  AOI21_X1 U8421 ( .B1(n6642), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10027), .ZN(
        n10115) );
  MUX2_X1 U8422 ( .A(n6643), .B(P1_REG1_REG_11__SCAN_IN), .S(n6644), .Z(n10116) );
  NOR2_X1 U8423 ( .A1(n10115), .A2(n10116), .ZN(n10114) );
  AOI21_X1 U8424 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6644), .A(n10114), .ZN(
        n6646) );
  AOI22_X1 U8425 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9463), .B1(n6652), .B2(
        n5563), .ZN(n6645) );
  NAND2_X1 U8426 ( .A1(n6646), .A2(n6645), .ZN(n9454) );
  OAI21_X1 U8427 ( .B1(n6646), .B2(n6645), .A(n9454), .ZN(n6649) );
  INV_X1 U8428 ( .A(n10152), .ZN(n10174) );
  NAND2_X1 U8429 ( .A1(n6649), .A2(n10174), .ZN(n6651) );
  AND2_X1 U8430 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9249) );
  AOI21_X1 U8431 ( .B1(n10138), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9249), .ZN(
        n6650) );
  OAI211_X1 U8432 ( .C1(n10121), .C2(n6652), .A(n6651), .B(n6650), .ZN(n6653)
         );
  AOI21_X1 U8433 ( .B1(n6654), .B2(n10175), .A(n6653), .ZN(n6655) );
  INV_X1 U8434 ( .A(n6655), .ZN(P1_U3255) );
  NAND2_X1 U8435 ( .A1(n9394), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6656) );
  OAI21_X1 U8436 ( .B1(n9528), .B2(n9394), .A(n6656), .ZN(P1_U3583) );
  INV_X1 U8437 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9147) );
  INV_X1 U8438 ( .A(n6657), .ZN(n6658) );
  INV_X1 U8439 ( .A(n8393), .ZN(n8400) );
  OAI222_X1 U8440 ( .A1(n8878), .A2(n9147), .B1(n8874), .B2(n6658), .C1(
        P2_U3151), .C2(n8400), .ZN(P2_U3280) );
  INV_X1 U8441 ( .A(n10161), .ZN(n9465) );
  INV_X1 U8442 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9111) );
  OAI222_X1 U8443 ( .A1(n9465), .A2(P1_U3086), .B1(n8174), .B2(n6658), .C1(
        n9111), .C2(n10018), .ZN(P1_U3340) );
  INV_X1 U8444 ( .A(n6665), .ZN(n7092) );
  INV_X1 U8445 ( .A(n9395), .ZN(n6785) );
  NAND2_X1 U8446 ( .A1(n6844), .A2(n7538), .ZN(n6661) );
  NOR2_X1 U8447 ( .A1(n6973), .A2(n7538), .ZN(n6843) );
  INV_X1 U8448 ( .A(n6843), .ZN(n6662) );
  NAND2_X1 U8449 ( .A1(n9395), .A2(n7807), .ZN(n6668) );
  NAND2_X1 U8450 ( .A1(n10236), .A2(n7808), .ZN(n6667) );
  NAND2_X1 U8451 ( .A1(n7092), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6666) );
  AND3_X1 U8452 ( .A1(n6668), .A2(n6667), .A3(n6666), .ZN(n6774) );
  XNOR2_X1 U8453 ( .A(n6775), .B(n6774), .ZN(n9406) );
  INV_X1 U8454 ( .A(n6669), .ZN(n6954) );
  NAND2_X1 U8455 ( .A1(n6954), .A2(n6670), .ZN(n6675) );
  NOR2_X1 U8456 ( .A1(n10280), .A2(n6842), .ZN(n6671) );
  INV_X1 U8457 ( .A(n6672), .ZN(n6674) );
  NAND2_X1 U8458 ( .A1(n10235), .A2(n6673), .ZN(n6971) );
  INV_X1 U8459 ( .A(n6971), .ZN(n6678) );
  OAI22_X1 U8460 ( .A1(n6675), .A2(n6674), .B1(n6678), .B2(n10268), .ZN(n6676)
         );
  NAND2_X1 U8461 ( .A1(n6676), .A2(n6953), .ZN(n7093) );
  NOR2_X1 U8462 ( .A1(n7093), .A2(n6677), .ZN(n6940) );
  INV_X1 U8463 ( .A(n6940), .ZN(n6684) );
  NAND2_X1 U8464 ( .A1(n6784), .A2(n6678), .ZN(n6681) );
  INV_X1 U8465 ( .A(n6679), .ZN(n6680) );
  INV_X1 U8466 ( .A(n9376), .ZN(n9364) );
  INV_X1 U8467 ( .A(n6777), .ZN(n6934) );
  AND2_X1 U8468 ( .A1(n10234), .A2(n6844), .ZN(n6682) );
  NAND2_X1 U8469 ( .A1(n6784), .A2(n6682), .ZN(n9359) );
  OAI22_X1 U8470 ( .A1(n9364), .A2(n8056), .B1(n6934), .B2(n9359), .ZN(n6683)
         );
  AOI21_X1 U8471 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6684), .A(n6683), .ZN(
        n6685) );
  OAI21_X1 U8472 ( .B1(n9406), .B2(n9378), .A(n6685), .ZN(P1_U3232) );
  NAND2_X1 U8473 ( .A1(n6280), .A2(n6742), .ZN(n6686) );
  NAND2_X1 U8474 ( .A1(n6687), .A2(n6686), .ZN(n8769) );
  INV_X1 U8475 ( .A(n8769), .ZN(n6700) );
  OR2_X1 U8476 ( .A1(n10312), .A2(n4855), .ZN(n6791) );
  OR2_X1 U8477 ( .A1(n10320), .A2(n6791), .ZN(n10314) );
  OAI21_X1 U8478 ( .B1(n6689), .B2(n6280), .A(n6688), .ZN(n6694) );
  NAND2_X1 U8479 ( .A1(n6690), .A2(n8687), .ZN(n6692) );
  NAND2_X1 U8480 ( .A1(n8366), .A2(n8685), .ZN(n6691) );
  NAND2_X1 U8481 ( .A1(n6692), .A2(n6691), .ZN(n6693) );
  AOI21_X1 U8482 ( .B1(n6694), .B2(n8690), .A(n6693), .ZN(n6696) );
  INV_X1 U8483 ( .A(n7446), .ZN(n10299) );
  NAND2_X1 U8484 ( .A1(n8769), .A2(n10299), .ZN(n6695) );
  AND2_X1 U8485 ( .A1(n6696), .A2(n6695), .ZN(n8771) );
  MUX2_X1 U8486 ( .A(n8771), .B(n6697), .S(n10320), .Z(n6699) );
  AOI22_X1 U8487 ( .A1(n10307), .A2(n8767), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10311), .ZN(n6698) );
  OAI211_X1 U8488 ( .C1(n6700), .C2(n10314), .A(n6699), .B(n6698), .ZN(
        P2_U3232) );
  INV_X1 U8489 ( .A(n6701), .ZN(n6702) );
  OAI22_X1 U8490 ( .A1(n6704), .A2(n6703), .B1(n6709), .B2(n6702), .ZN(n6707)
         );
  MUX2_X1 U8491 ( .A(n6820), .B(n6708), .S(n8489), .Z(n6705) );
  INV_X1 U8492 ( .A(n6721), .ZN(n6821) );
  NAND2_X1 U8493 ( .A1(n6705), .A2(n6821), .ZN(n6807) );
  OAI21_X1 U8494 ( .B1(n6705), .B2(n6821), .A(n6807), .ZN(n6706) );
  NOR2_X1 U8495 ( .A1(n6707), .A2(n6706), .ZN(n6814) );
  AOI21_X1 U8496 ( .B1(n6707), .B2(n6706), .A(n6814), .ZN(n6725) );
  MUX2_X1 U8497 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6708), .S(n6721), .Z(n6713)
         );
  INV_X1 U8498 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8499 ( .A1(n6712), .A2(n6713), .ZN(n6806) );
  OAI21_X1 U8500 ( .B1(n6713), .B2(n6712), .A(n6806), .ZN(n6723) );
  INV_X1 U8501 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9036) );
  NOR2_X1 U8502 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9036), .ZN(n7013) );
  MUX2_X1 U8503 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6820), .S(n6721), .Z(n6715)
         );
  INV_X1 U8504 ( .A(n6714), .ZN(n6716) );
  OR3_X1 U8505 ( .A1(n6717), .A2(n6715), .A3(n6716), .ZN(n6718) );
  AOI21_X1 U8506 ( .B1(n6718), .B2(n6819), .A(n8501), .ZN(n6719) );
  AOI211_X1 U8507 ( .C1(n8482), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7013), .B(
        n6719), .ZN(n6720) );
  OAI21_X1 U8508 ( .B1(n6721), .B2(n8486), .A(n6720), .ZN(n6722) );
  AOI21_X1 U8509 ( .B1(n8499), .B2(n6723), .A(n6722), .ZN(n6724) );
  OAI21_X1 U8510 ( .B1(n6725), .B2(n8494), .A(n6724), .ZN(P2_U3188) );
  INV_X1 U8511 ( .A(n6726), .ZN(n6729) );
  OAI222_X1 U8512 ( .A1(n8874), .A2(n6729), .B1(n8422), .B2(P2_U3151), .C1(
        n6727), .C2(n8878), .ZN(P2_U3279) );
  INV_X1 U8513 ( .A(n9485), .ZN(n9468) );
  OAI222_X1 U8514 ( .A1(P1_U3086), .A2(n9468), .B1(n8174), .B2(n6729), .C1(
        n6728), .C2(n10018), .ZN(P1_U3339) );
  INV_X1 U8515 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8976) );
  INV_X1 U8516 ( .A(n6730), .ZN(n6732) );
  NAND2_X1 U8517 ( .A1(n6732), .A2(n6731), .ZN(n8342) );
  AOI22_X1 U8518 ( .A1(n8331), .A2(n8366), .B1(n8344), .B2(n6916), .ZN(n6734)
         );
  OAI211_X1 U8519 ( .C1(n6947), .C2(n8311), .A(n6734), .B(n6733), .ZN(n6756)
         );
  OAI21_X1 U8520 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6738) );
  INV_X1 U8521 ( .A(n6738), .ZN(n6740) );
  XNOR2_X1 U8522 ( .A(n6743), .B(n6998), .ZN(n8240) );
  NAND2_X1 U8523 ( .A1(n8240), .A2(n8239), .ZN(n6745) );
  NAND2_X1 U8524 ( .A1(n6745), .A2(n6744), .ZN(n8313) );
  XNOR2_X1 U8525 ( .A(n8366), .B(n6747), .ZN(n8314) );
  NAND2_X1 U8526 ( .A1(n8313), .A2(n8314), .ZN(n6749) );
  NAND2_X1 U8527 ( .A1(n6747), .A2(n7856), .ZN(n6748) );
  NAND2_X1 U8528 ( .A1(n6752), .A2(n6751), .ZN(n6761) );
  INV_X1 U8529 ( .A(n6761), .ZN(n6753) );
  AOI211_X1 U8530 ( .C1(n6754), .C2(n6750), .A(n8348), .B(n6753), .ZN(n6755)
         );
  AOI211_X1 U8531 ( .C1(n8976), .C2(n8332), .A(n6756), .B(n6755), .ZN(n6757)
         );
  INV_X1 U8532 ( .A(n6757), .ZN(P2_U3158) );
  XNOR2_X1 U8533 ( .A(n6746), .B(n6802), .ZN(n6912) );
  XNOR2_X1 U8534 ( .A(n6912), .B(n7060), .ZN(n6765) );
  INV_X1 U8535 ( .A(n6758), .ZN(n6759) );
  INV_X1 U8536 ( .A(n6997), .ZN(n8365) );
  NAND2_X1 U8537 ( .A1(n6759), .A2(n8365), .ZN(n6760) );
  NAND2_X1 U8538 ( .A1(n6761), .A2(n6760), .ZN(n6764) );
  INV_X1 U8539 ( .A(n6914), .ZN(n6763) );
  AOI21_X1 U8540 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(n6772) );
  INV_X1 U8541 ( .A(n6766), .ZN(n6801) );
  AOI22_X1 U8542 ( .A1(n8331), .A2(n8365), .B1(n8344), .B2(n8364), .ZN(n6769)
         );
  INV_X1 U8543 ( .A(n6767), .ZN(n6768) );
  OAI211_X1 U8544 ( .C1(n6943), .C2(n8311), .A(n6769), .B(n6768), .ZN(n6770)
         );
  AOI21_X1 U8545 ( .B1(n6801), .B2(n8332), .A(n6770), .ZN(n6771) );
  OAI21_X1 U8546 ( .B1(n6772), .B2(n8348), .A(n6771), .ZN(P2_U3170) );
  OAI22_X1 U8547 ( .A1(n6775), .A2(n6774), .B1(n7798), .B2(n6773), .ZN(n6782)
         );
  XNOR2_X1 U8548 ( .A(n6778), .B(n7798), .ZN(n6780) );
  AOI22_X1 U8549 ( .A1(n5469), .A2(n7808), .B1(n6777), .B2(n7807), .ZN(n6779)
         );
  NAND2_X1 U8550 ( .A1(n6780), .A2(n6779), .ZN(n6922) );
  OAI21_X1 U8551 ( .B1(n6780), .B2(n6779), .A(n6922), .ZN(n6781) );
  AOI21_X1 U8552 ( .B1(n6782), .B2(n6781), .A(n6929), .ZN(n6789) );
  NOR2_X1 U8553 ( .A1(n6940), .A2(n6972), .ZN(n6787) );
  AND2_X1 U8554 ( .A1(n9929), .A2(n6844), .ZN(n6783) );
  OAI22_X1 U8555 ( .A1(n9370), .A2(n6785), .B1(n7102), .B2(n9359), .ZN(n6786)
         );
  AOI211_X1 U8556 ( .C1(n5469), .C2(n9376), .A(n6787), .B(n6786), .ZN(n6788)
         );
  OAI21_X1 U8557 ( .B1(n6789), .B2(n9378), .A(n6788), .ZN(P1_U3222) );
  XNOR2_X1 U8558 ( .A(n6790), .B(n7859), .ZN(n6945) );
  INV_X1 U8559 ( .A(n6945), .ZN(n6805) );
  NAND2_X1 U8560 ( .A1(n7446), .A2(n6791), .ZN(n6792) );
  NAND3_X1 U8561 ( .A1(n6794), .A2(n7859), .A3(n6795), .ZN(n6796) );
  NAND2_X1 U8562 ( .A1(n6793), .A2(n6796), .ZN(n6799) );
  NAND2_X1 U8563 ( .A1(n8364), .A2(n8685), .ZN(n6797) );
  OAI21_X1 U8564 ( .B1(n6997), .B2(n8671), .A(n6797), .ZN(n6798) );
  AOI21_X1 U8565 ( .B1(n6799), .B2(n8690), .A(n6798), .ZN(n6942) );
  MUX2_X1 U8566 ( .A(n6800), .B(n6942), .S(n8678), .Z(n6804) );
  AOI22_X1 U8567 ( .A1(n10307), .A2(n6802), .B1(n10311), .B2(n6801), .ZN(n6803) );
  OAI211_X1 U8568 ( .C1(n6805), .C2(n8666), .A(n6804), .B(n6803), .ZN(P2_U3229) );
  OAI21_X1 U8569 ( .B1(n6821), .B2(n6708), .A(n6806), .ZN(n6858) );
  INV_X1 U8570 ( .A(n6859), .ZN(n6828) );
  INV_X1 U8571 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6808) );
  XNOR2_X1 U8572 ( .A(n6860), .B(n6808), .ZN(n6831) );
  INV_X1 U8573 ( .A(n6807), .ZN(n6813) );
  MUX2_X1 U8574 ( .A(n6824), .B(n6808), .S(n8489), .Z(n6809) );
  NAND2_X1 U8575 ( .A1(n6809), .A2(n6828), .ZN(n6868) );
  INV_X1 U8576 ( .A(n6809), .ZN(n6810) );
  NAND2_X1 U8577 ( .A1(n6810), .A2(n6859), .ZN(n6811) );
  AND2_X1 U8578 ( .A1(n6868), .A2(n6811), .ZN(n6812) );
  OAI21_X1 U8579 ( .B1(n6814), .B2(n6813), .A(n6812), .ZN(n6869) );
  INV_X1 U8580 ( .A(n6869), .ZN(n6816) );
  NOR3_X1 U8581 ( .A1(n6814), .A2(n6813), .A3(n6812), .ZN(n6815) );
  OAI21_X1 U8582 ( .B1(n6816), .B2(n6815), .A(n8382), .ZN(n6830) );
  INV_X1 U8583 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6818) );
  AND2_X1 U8584 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7154) );
  INV_X1 U8585 ( .A(n7154), .ZN(n6817) );
  OAI21_X1 U8586 ( .B1(n8441), .B2(n6818), .A(n6817), .ZN(n6827) );
  INV_X1 U8587 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8588 ( .A1(n6822), .A2(n6859), .ZN(n6872) );
  OAI21_X1 U8589 ( .B1(n6822), .B2(n6859), .A(n6872), .ZN(n6823) );
  AOI21_X1 U8590 ( .B1(n6824), .B2(n6823), .A(n6875), .ZN(n6825) );
  NOR2_X1 U8591 ( .A1(n6825), .A2(n8501), .ZN(n6826) );
  AOI211_X1 U8592 ( .C1(n8450), .C2(n6828), .A(n6827), .B(n6826), .ZN(n6829)
         );
  OAI211_X1 U8593 ( .C1(n6831), .C2(n7053), .A(n6830), .B(n6829), .ZN(P2_U3189) );
  OR2_X1 U8594 ( .A1(n7335), .A2(n7281), .ZN(n6834) );
  NAND2_X1 U8595 ( .A1(n6832), .A2(n6973), .ZN(n6833) );
  XNOR2_X1 U8596 ( .A(n6836), .B(n6835), .ZN(n8066) );
  INV_X1 U8597 ( .A(n6837), .ZN(n6958) );
  NAND2_X1 U8598 ( .A1(n9395), .A2(n10236), .ZN(n6959) );
  NAND2_X1 U8599 ( .A1(n6934), .A2(n5468), .ZN(n6838) );
  NAND2_X1 U8600 ( .A1(n6960), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8601 ( .A1(n6840), .A2(n6839), .ZN(n6982) );
  OAI21_X1 U8602 ( .B1(n6840), .B2(n6839), .A(n6982), .ZN(n6841) );
  INV_X1 U8603 ( .A(n6841), .ZN(n8069) );
  NAND2_X1 U8604 ( .A1(n6842), .A2(n6844), .ZN(n8051) );
  INV_X1 U8605 ( .A(n10235), .ZN(n8050) );
  OAI211_X1 U8606 ( .C1(n6844), .C2(n6843), .A(n8051), .B(n8050), .ZN(n7018)
         );
  NAND2_X1 U8607 ( .A1(n6845), .A2(n7281), .ZN(n10260) );
  NAND2_X1 U8608 ( .A1(n7018), .A2(n10260), .ZN(n10285) );
  INV_X1 U8609 ( .A(n10285), .ZN(n10233) );
  AOI22_X1 U8610 ( .A1(n9929), .A2(n6777), .B1(n9392), .B2(n10234), .ZN(n6848)
         );
  INV_X1 U8611 ( .A(n6974), .ZN(n6847) );
  INV_X1 U8612 ( .A(n6986), .ZN(n6846) );
  OAI211_X1 U8613 ( .C1(n8059), .C2(n6847), .A(n6846), .B(n9932), .ZN(n8062)
         );
  OAI211_X1 U8614 ( .C1(n8069), .C2(n10233), .A(n6848), .B(n8062), .ZN(n6849)
         );
  AOI21_X1 U8615 ( .B1(n9927), .B2(n8066), .A(n6849), .ZN(n6854) );
  INV_X1 U8616 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6850) );
  OAI22_X1 U8617 ( .A1(n10000), .A2(n8059), .B1(n10289), .B2(n6850), .ZN(n6851) );
  INV_X1 U8618 ( .A(n6851), .ZN(n6852) );
  OAI21_X1 U8619 ( .B1(n6854), .B2(n10287), .A(n6852), .ZN(P1_U3459) );
  AOI22_X1 U8620 ( .A1(n9833), .A2(n6936), .B1(n5414), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6853) );
  OAI21_X1 U8621 ( .B1(n6854), .B2(n5414), .A(n6853), .ZN(P1_U3524) );
  INV_X1 U8622 ( .A(n10172), .ZN(n9487) );
  INV_X1 U8623 ( .A(n6855), .ZN(n6856) );
  OAI222_X1 U8624 ( .A1(n9487), .A2(P1_U3086), .B1(n8174), .B2(n6856), .C1(
        n8974), .C2(n10018), .ZN(P1_U3338) );
  INV_X1 U8625 ( .A(n8452), .ZN(n8460) );
  OAI222_X1 U8626 ( .A1(n8878), .A2(n6857), .B1(n8874), .B2(n6856), .C1(
        P2_U3151), .C2(n8460), .ZN(P2_U3278) );
  MUX2_X1 U8627 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6863), .S(n7046), .Z(n6862)
         );
  AOI21_X1 U8628 ( .B1(n6862), .B2(n6861), .A(n7031), .ZN(n6881) );
  MUX2_X1 U8629 ( .A(n7220), .B(n6863), .S(n8489), .Z(n6864) );
  NAND2_X1 U8630 ( .A1(n6864), .A2(n7046), .ZN(n7032) );
  INV_X1 U8631 ( .A(n6864), .ZN(n6865) );
  NAND2_X1 U8632 ( .A1(n6865), .A2(n4536), .ZN(n6866) );
  NAND2_X1 U8633 ( .A1(n7032), .A2(n6866), .ZN(n6867) );
  AOI21_X1 U8634 ( .B1(n6869), .B2(n6868), .A(n6867), .ZN(n7039) );
  AND3_X1 U8635 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n6870) );
  OAI21_X1 U8636 ( .B1(n7039), .B2(n6870), .A(n8382), .ZN(n6880) );
  INV_X1 U8637 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8972) );
  AND2_X1 U8638 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7339) );
  INV_X1 U8639 ( .A(n7339), .ZN(n6871) );
  OAI21_X1 U8640 ( .B1(n8441), .B2(n8972), .A(n6871), .ZN(n6878) );
  INV_X1 U8641 ( .A(n6872), .ZN(n6873) );
  MUX2_X1 U8642 ( .A(n7220), .B(P2_REG2_REG_8__SCAN_IN), .S(n7046), .Z(n6874)
         );
  OR3_X1 U8643 ( .A1(n6875), .A2(n6874), .A3(n6873), .ZN(n6876) );
  AOI21_X1 U8644 ( .B1(n7045), .B2(n6876), .A(n8501), .ZN(n6877) );
  AOI211_X1 U8645 ( .C1(n8450), .C2(n7046), .A(n6878), .B(n6877), .ZN(n6879)
         );
  OAI211_X1 U8646 ( .C1(n6881), .C2(n7053), .A(n6880), .B(n6879), .ZN(P2_U3190) );
  OAI21_X1 U8647 ( .B1(n6883), .B2(n8002), .A(n6882), .ZN(n6950) );
  INV_X1 U8648 ( .A(n6950), .ZN(n6893) );
  NAND3_X1 U8649 ( .A1(n6884), .A2(n8002), .A3(n6885), .ZN(n6886) );
  AND2_X1 U8650 ( .A1(n6794), .A2(n6886), .ZN(n6887) );
  OAI222_X1 U8651 ( .A1(n8673), .A2(n7060), .B1(n8671), .B2(n7856), .C1(n8668), 
        .C2(n6887), .ZN(n6948) );
  INV_X1 U8652 ( .A(n6948), .ZN(n6888) );
  MUX2_X1 U8653 ( .A(n6889), .B(n6888), .S(n8678), .Z(n6892) );
  AOI22_X1 U8654 ( .A1(n10307), .A2(n6890), .B1(n8976), .B2(n10311), .ZN(n6891) );
  OAI211_X1 U8655 ( .C1(n6893), .C2(n8666), .A(n6892), .B(n6891), .ZN(P2_U3230) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10351) );
  INV_X1 U8657 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10179) );
  INV_X1 U8658 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9148) );
  AOI22_X1 U8659 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10179), .B2(n9148), .ZN(n10356) );
  NOR2_X1 U8660 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6894) );
  AOI21_X1 U8661 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6894), .ZN(n10359) );
  INV_X1 U8662 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10165) );
  INV_X1 U8663 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U8664 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n10165), .B2(n6895), .ZN(n10362) );
  NOR2_X1 U8665 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6896) );
  AOI21_X1 U8666 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6896), .ZN(n10365) );
  NOR2_X1 U8667 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6897) );
  AOI21_X1 U8668 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6897), .ZN(n10368) );
  NOR2_X1 U8669 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6898) );
  AOI21_X1 U8670 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6898), .ZN(n10371) );
  NOR2_X1 U8671 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6899) );
  AOI21_X1 U8672 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6899), .ZN(n10374) );
  INV_X1 U8673 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10037) );
  INV_X1 U8674 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7174) );
  AOI22_X1 U8675 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .B1(n10037), .B2(n7174), .ZN(n10377) );
  INV_X1 U8676 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10078) );
  INV_X1 U8677 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7044) );
  AOI22_X1 U8678 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(n10078), .B2(n7044), .ZN(n10386) );
  NOR2_X1 U8679 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6900) );
  AOI21_X1 U8680 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6900), .ZN(n10392) );
  NOR2_X1 U8681 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6901) );
  AOI21_X1 U8682 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6901), .ZN(n10389) );
  NOR2_X1 U8683 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6902) );
  AOI21_X1 U8684 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6902), .ZN(n10380) );
  NOR2_X1 U8685 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6903) );
  AOI21_X1 U8686 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6903), .ZN(n10383) );
  INV_X1 U8687 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10348) );
  NOR2_X1 U8688 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  NOR2_X1 U8689 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10347), .ZN(n10343) );
  INV_X1 U8690 ( .A(n10343), .ZN(n10344) );
  NAND3_X1 U8691 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U8692 ( .A1(n10346), .A2(n10345), .ZN(n10342) );
  NAND2_X1 U8693 ( .A1(n10344), .A2(n10342), .ZN(n10395) );
  NAND2_X1 U8694 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6904) );
  OAI21_X1 U8695 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6904), .ZN(n10394) );
  NOR2_X1 U8696 ( .A1(n10395), .A2(n10394), .ZN(n10393) );
  AOI21_X1 U8697 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10393), .ZN(n10398) );
  NAND2_X1 U8698 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6905) );
  OAI21_X1 U8699 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6905), .ZN(n10397) );
  NOR2_X1 U8700 ( .A1(n10398), .A2(n10397), .ZN(n10396) );
  AOI21_X1 U8701 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10396), .ZN(n10401) );
  NOR2_X1 U8702 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6906) );
  AOI21_X1 U8703 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6906), .ZN(n10400) );
  NAND2_X1 U8704 ( .A1(n10401), .A2(n10400), .ZN(n10399) );
  OAI21_X1 U8705 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10399), .ZN(n10382) );
  NAND2_X1 U8706 ( .A1(n10383), .A2(n10382), .ZN(n10381) );
  OAI21_X1 U8707 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10381), .ZN(n10379) );
  NAND2_X1 U8708 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  OAI21_X1 U8709 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10378), .ZN(n10388) );
  NAND2_X1 U8710 ( .A1(n10389), .A2(n10388), .ZN(n10387) );
  OAI21_X1 U8711 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10387), .ZN(n10391) );
  NAND2_X1 U8712 ( .A1(n10392), .A2(n10391), .ZN(n10390) );
  OAI21_X1 U8713 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10390), .ZN(n10385) );
  NAND2_X1 U8714 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  OAI21_X1 U8715 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10384), .ZN(n10376) );
  NAND2_X1 U8716 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  OAI21_X1 U8717 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10375), .ZN(n10373) );
  NAND2_X1 U8718 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  OAI21_X1 U8719 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10372), .ZN(n10370) );
  NAND2_X1 U8720 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  OAI21_X1 U8721 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10369), .ZN(n10367) );
  NAND2_X1 U8722 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  OAI21_X1 U8723 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10366), .ZN(n10364) );
  NAND2_X1 U8724 ( .A1(n10365), .A2(n10364), .ZN(n10363) );
  OAI21_X1 U8725 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10363), .ZN(n10361) );
  NAND2_X1 U8726 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OAI21_X1 U8727 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10360), .ZN(n10358) );
  NAND2_X1 U8728 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  OAI21_X1 U8729 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10357), .ZN(n10355) );
  NAND2_X1 U8730 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  OAI21_X1 U8731 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10354), .ZN(n10352) );
  NOR2_X1 U8732 ( .A1(n10351), .A2(n10352), .ZN(n6907) );
  NAND2_X1 U8733 ( .A1(n10351), .A2(n10352), .ZN(n10350) );
  OAI21_X1 U8734 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6907), .A(n10350), .ZN(
        n6911) );
  NOR2_X1 U8735 ( .A1(n6908), .A2(n6909), .ZN(n6910) );
  XNOR2_X1 U8736 ( .A(n6911), .B(n6910), .ZN(ADD_1068_U4) );
  NAND2_X1 U8737 ( .A1(n6912), .A2(n7060), .ZN(n6913) );
  XNOR2_X1 U8738 ( .A(n6746), .B(n7112), .ZN(n7005) );
  XNOR2_X1 U8739 ( .A(n7005), .B(n8364), .ZN(n7006) );
  XOR2_X1 U8740 ( .A(n7007), .B(n7006), .Z(n6921) );
  INV_X1 U8741 ( .A(n6915), .ZN(n7111) );
  AOI22_X1 U8742 ( .A1(n8331), .A2(n6916), .B1(n8344), .B2(n8363), .ZN(n6918)
         );
  OAI211_X1 U8743 ( .C1(n7064), .C2(n8311), .A(n6918), .B(n6917), .ZN(n6919)
         );
  AOI21_X1 U8744 ( .B1(n7111), .B2(n8332), .A(n6919), .ZN(n6920) );
  OAI21_X1 U8745 ( .B1(n6921), .B2(n8348), .A(n6920), .ZN(P2_U3167) );
  INV_X1 U8746 ( .A(n6922), .ZN(n6931) );
  NAND2_X1 U8747 ( .A1(n9393), .A2(n7808), .ZN(n6923) );
  OAI21_X1 U8748 ( .B1(n8059), .B2(n7812), .A(n6923), .ZN(n6925) );
  XNOR2_X1 U8749 ( .A(n6925), .B(n6924), .ZN(n6927) );
  AOI22_X1 U8750 ( .A1(n6936), .A2(n7808), .B1(n9393), .B2(n7807), .ZN(n6926)
         );
  NAND2_X1 U8751 ( .A1(n6927), .A2(n6926), .ZN(n7097) );
  OR2_X1 U8752 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  AND2_X1 U8753 ( .A1(n7097), .A2(n6928), .ZN(n6930) );
  INV_X1 U8754 ( .A(n7098), .ZN(n6933) );
  NOR3_X1 U8755 ( .A1(n6929), .A2(n6931), .A3(n6930), .ZN(n6932) );
  OAI21_X1 U8756 ( .B1(n6933), .B2(n6932), .A(n9352), .ZN(n6938) );
  OAI22_X1 U8757 ( .A1(n9370), .A2(n6934), .B1(n8060), .B2(n9359), .ZN(n6935)
         );
  AOI21_X1 U8758 ( .B1(n6936), .B2(n9376), .A(n6935), .ZN(n6937) );
  OAI211_X1 U8759 ( .C1(n6940), .C2(n6939), .A(n6938), .B(n6937), .ZN(P1_U3237) );
  OAI21_X1 U8760 ( .B1(n6943), .B2(n8764), .A(n6942), .ZN(n6944) );
  AOI21_X1 U8761 ( .B1(n6945), .B2(n8760), .A(n6944), .ZN(n10329) );
  OR2_X1 U8762 ( .A1(n8772), .A2(n5954), .ZN(n6946) );
  OAI21_X1 U8763 ( .B1(n10329), .B2(n7564), .A(n6946), .ZN(P2_U3463) );
  NOR2_X1 U8764 ( .A1(n6947), .A2(n8764), .ZN(n6949) );
  AOI211_X1 U8765 ( .C1(n8760), .C2(n6950), .A(n6949), .B(n6948), .ZN(n10327)
         );
  OR2_X1 U8766 ( .A1(n10327), .A2(n7564), .ZN(n6951) );
  OAI21_X1 U8767 ( .B1(n8772), .B2(n5944), .A(n6951), .ZN(P2_U3462) );
  INV_X1 U8768 ( .A(n6952), .ZN(n6955) );
  NAND4_X1 U8769 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6957)
         );
  INV_X1 U8770 ( .A(n7017), .ZN(n6970) );
  OR2_X1 U8771 ( .A1(n6958), .A2(n6959), .ZN(n6961) );
  NAND2_X1 U8772 ( .A1(n6961), .A2(n6960), .ZN(n10241) );
  INV_X1 U8773 ( .A(n7018), .ZN(n10264) );
  NAND2_X1 U8774 ( .A1(n10241), .A2(n10264), .ZN(n6969) );
  AOI22_X1 U8775 ( .A1(n9929), .A2(n9395), .B1(n9393), .B2(n10234), .ZN(n6968)
         );
  INV_X1 U8776 ( .A(n6962), .ZN(n6963) );
  NAND2_X1 U8777 ( .A1(n6963), .A2(n6958), .ZN(n6965) );
  NAND2_X1 U8778 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  NAND2_X1 U8779 ( .A1(n6966), .A2(n9927), .ZN(n6967) );
  NAND3_X1 U8780 ( .A1(n6969), .A2(n6968), .A3(n6967), .ZN(n10245) );
  AOI21_X1 U8781 ( .B1(n6970), .B2(n10241), .A(n10245), .ZN(n6978) );
  OAI22_X1 U8782 ( .A1(n10208), .A2(n5456), .B1(n6972), .B2(n10205), .ZN(n6976) );
  NOR2_X2 U8783 ( .A1(n9728), .A2(n6973), .ZN(n10191) );
  OAI211_X1 U8784 ( .C1(n8056), .C2(n5468), .A(n9932), .B(n6974), .ZN(n10242)
         );
  NOR2_X1 U8785 ( .A1(n10213), .A2(n10242), .ZN(n6975) );
  AOI211_X1 U8786 ( .C1(n10211), .C2(n5469), .A(n6976), .B(n6975), .ZN(n6977)
         );
  OAI21_X1 U8787 ( .B1(n10220), .B2(n6978), .A(n6977), .ZN(P1_U3292) );
  XNOR2_X1 U8788 ( .A(n6979), .B(n6980), .ZN(n7025) );
  NAND2_X1 U8789 ( .A1(n7102), .A2(n8059), .ZN(n6981) );
  NAND2_X1 U8790 ( .A1(n6982), .A2(n6981), .ZN(n6984) );
  NAND2_X1 U8791 ( .A1(n6984), .A2(n6983), .ZN(n7074) );
  OAI21_X1 U8792 ( .B1(n6984), .B2(n6983), .A(n7074), .ZN(n6985) );
  INV_X1 U8793 ( .A(n6985), .ZN(n7028) );
  AOI22_X1 U8794 ( .A1(n9929), .A2(n9393), .B1(n9391), .B2(n10234), .ZN(n6987)
         );
  OAI211_X1 U8795 ( .C1(n6986), .C2(n7103), .A(n7270), .B(n9932), .ZN(n7022)
         );
  OAI211_X1 U8796 ( .C1(n7028), .C2(n10233), .A(n6987), .B(n7022), .ZN(n6988)
         );
  AOI21_X1 U8797 ( .B1(n9927), .B2(n7025), .A(n6988), .ZN(n6994) );
  AOI22_X1 U8798 ( .A1(n9833), .A2(n6989), .B1(n5414), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6990) );
  OAI21_X1 U8799 ( .B1(n6994), .B2(n5414), .A(n6990), .ZN(P1_U3525) );
  INV_X1 U8800 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6991) );
  OAI22_X1 U8801 ( .A1(n10000), .A2(n7103), .B1(n10289), .B2(n6991), .ZN(n6992) );
  INV_X1 U8802 ( .A(n6992), .ZN(n6993) );
  OAI21_X1 U8803 ( .B1(n6994), .B2(n10287), .A(n6993), .ZN(P1_U3462) );
  INV_X1 U8804 ( .A(n7486), .ZN(n8768) );
  XNOR2_X1 U8805 ( .A(n6995), .B(n8003), .ZN(n10316) );
  INV_X1 U8806 ( .A(n4421), .ZN(n6996) );
  NOR2_X1 U8807 ( .A1(n6996), .A2(n8764), .ZN(n10313) );
  OAI22_X1 U8808 ( .A1(n6998), .A2(n8671), .B1(n6997), .B2(n8673), .ZN(n7002)
         );
  NAND3_X1 U8809 ( .A1(n6688), .A2(n8003), .A3(n6999), .ZN(n7000) );
  AOI21_X1 U8810 ( .B1(n6884), .B2(n7000), .A(n8668), .ZN(n7001) );
  AOI211_X1 U8811 ( .C1(n10299), .C2(n10316), .A(n7002), .B(n7001), .ZN(n10319) );
  INV_X1 U8812 ( .A(n10319), .ZN(n7003) );
  AOI211_X1 U8813 ( .C1(n8768), .C2(n10316), .A(n10313), .B(n7003), .ZN(n10325) );
  OR2_X1 U8814 ( .A1(n10325), .A2(n7564), .ZN(n7004) );
  OAI21_X1 U8815 ( .B1(n8772), .B2(n5932), .A(n7004), .ZN(P2_U3461) );
  XNOR2_X1 U8816 ( .A(n6746), .B(n7014), .ZN(n7146) );
  XNOR2_X1 U8817 ( .A(n7146), .B(n8363), .ZN(n7008) );
  OAI211_X1 U8818 ( .C1(n7009), .C2(n7008), .A(n7149), .B(n8315), .ZN(n7016)
         );
  INV_X1 U8819 ( .A(n7336), .ZN(n8362) );
  NAND2_X1 U8820 ( .A1(n8344), .A2(n8362), .ZN(n7010) );
  OAI21_X1 U8821 ( .B1(n7011), .B2(n8342), .A(n7010), .ZN(n7012) );
  AOI211_X1 U8822 ( .C1(n7014), .C2(n8353), .A(n7013), .B(n7012), .ZN(n7015)
         );
  OAI211_X1 U8823 ( .C1(n7088), .C2(n8346), .A(n7016), .B(n7015), .ZN(P2_U3179) );
  AND2_X1 U8824 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  NOR2_X2 U8825 ( .A1(n10220), .A2(n7019), .ZN(n10216) );
  NOR2_X2 U8826 ( .A1(n9728), .A2(n10275), .ZN(n9784) );
  INV_X1 U8827 ( .A(n10205), .ZN(n10194) );
  INV_X1 U8828 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U8829 ( .A1(n9728), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10194), .B2(
        n7020), .ZN(n7021) );
  OAI21_X1 U8830 ( .B1(n10198), .B2(n7103), .A(n7021), .ZN(n7024) );
  OR2_X1 U8831 ( .A1(n10220), .A2(n10273), .ZN(n9779) );
  OAI22_X1 U8832 ( .A1(n7022), .A2(n10213), .B1(n7102), .B2(n9779), .ZN(n7023)
         );
  AOI211_X1 U8833 ( .C1(n9784), .C2(n9391), .A(n7024), .B(n7023), .ZN(n7027)
         );
  NOR2_X1 U8834 ( .A1(n9728), .A2(n10283), .ZN(n9751) );
  NAND2_X1 U8835 ( .A1(n7025), .A2(n9751), .ZN(n7026) );
  OAI211_X1 U8836 ( .C1(n7028), .C2(n9753), .A(n7027), .B(n7026), .ZN(P1_U3290) );
  INV_X1 U8837 ( .A(n7029), .ZN(n7067) );
  INV_X1 U8838 ( .A(n9476), .ZN(n9494) );
  OAI222_X1 U8839 ( .A1(n10009), .A2(n7030), .B1(n8174), .B2(n7067), .C1(
        P1_U3086), .C2(n9494), .ZN(P1_U3337) );
  XNOR2_X1 U8840 ( .A(n7163), .B(n7164), .ZN(n7166) );
  XNOR2_X1 U8841 ( .A(n7166), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7054) );
  INV_X1 U8842 ( .A(n7032), .ZN(n7038) );
  INV_X1 U8843 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7165) );
  MUX2_X1 U8844 ( .A(n7033), .B(n7165), .S(n8489), .Z(n7034) );
  NAND2_X1 U8845 ( .A1(n7034), .A2(n7164), .ZN(n7183) );
  INV_X1 U8846 ( .A(n7034), .ZN(n7035) );
  NAND2_X1 U8847 ( .A1(n7035), .A2(n7171), .ZN(n7036) );
  AND2_X1 U8848 ( .A1(n7183), .A2(n7036), .ZN(n7037) );
  OAI21_X1 U8849 ( .B1(n7039), .B2(n7038), .A(n7037), .ZN(n7184) );
  INV_X1 U8850 ( .A(n7184), .ZN(n7041) );
  NOR3_X1 U8851 ( .A1(n7039), .A2(n7038), .A3(n7037), .ZN(n7040) );
  OAI21_X1 U8852 ( .B1(n7041), .B2(n7040), .A(n8382), .ZN(n7052) );
  INV_X1 U8853 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7042) );
  NOR2_X1 U8854 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7042), .ZN(n7429) );
  INV_X1 U8855 ( .A(n7429), .ZN(n7043) );
  OAI21_X1 U8856 ( .B1(n8441), .B2(n7044), .A(n7043), .ZN(n7050) );
  XNOR2_X1 U8857 ( .A(n7170), .B(n7171), .ZN(n7047) );
  NOR2_X1 U8858 ( .A1(n7047), .A2(n7033), .ZN(n7169) );
  AOI21_X1 U8859 ( .B1(n7033), .B2(n7047), .A(n7169), .ZN(n7048) );
  NOR2_X1 U8860 ( .A1(n7048), .A2(n8501), .ZN(n7049) );
  AOI211_X1 U8861 ( .C1(n8450), .C2(n7164), .A(n7050), .B(n7049), .ZN(n7051)
         );
  OAI211_X1 U8862 ( .C1(n7054), .C2(n7053), .A(n7052), .B(n7051), .ZN(P2_U3191) );
  INV_X1 U8863 ( .A(n7056), .ZN(n7057) );
  OR2_X1 U8864 ( .A1(n7058), .A2(n7057), .ZN(n8000) );
  XOR2_X1 U8865 ( .A(n7055), .B(n8000), .Z(n7115) );
  XOR2_X1 U8866 ( .A(n8000), .B(n7059), .Z(n7062) );
  OAI22_X1 U8867 ( .A1(n7399), .A2(n8673), .B1(n7060), .B2(n8671), .ZN(n7061)
         );
  AOI21_X1 U8868 ( .B1(n7062), .B2(n8690), .A(n7061), .ZN(n7063) );
  OAI21_X1 U8869 ( .B1(n7115), .B2(n7446), .A(n7063), .ZN(n7108) );
  OAI22_X1 U8870 ( .A1(n7115), .A2(n7486), .B1(n7064), .B2(n8764), .ZN(n7065)
         );
  NOR2_X1 U8871 ( .A1(n7108), .A2(n7065), .ZN(n10331) );
  NAND2_X1 U8872 ( .A1(n7564), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7066) );
  OAI21_X1 U8873 ( .B1(n10331), .B2(n7564), .A(n7066), .ZN(P2_U3464) );
  INV_X1 U8874 ( .A(n8467), .ZN(n8480) );
  OAI222_X1 U8875 ( .A1(n8878), .A2(n7068), .B1(n8480), .B2(P2_U3151), .C1(
        n8874), .C2(n7067), .ZN(P2_U3277) );
  INV_X1 U8876 ( .A(n7076), .ZN(n7069) );
  XNOR2_X1 U8877 ( .A(n5786), .B(n7069), .ZN(n7072) );
  NAND2_X1 U8878 ( .A1(n9391), .A2(n9929), .ZN(n7070) );
  OAI21_X1 U8879 ( .B1(n7323), .B2(n10275), .A(n7070), .ZN(n7071) );
  AOI21_X1 U8880 ( .B1(n7072), .B2(n9927), .A(n7071), .ZN(n10252) );
  NAND2_X1 U8881 ( .A1(n8060), .A2(n7103), .ZN(n7073) );
  NAND2_X1 U8882 ( .A1(n7074), .A2(n7073), .ZN(n7264) );
  NAND2_X1 U8883 ( .A1(n7264), .A2(n7268), .ZN(n7266) );
  NAND2_X1 U8884 ( .A1(n7141), .A2(n7275), .ZN(n7075) );
  NAND2_X1 U8885 ( .A1(n7266), .A2(n7075), .ZN(n7077) );
  NAND2_X1 U8886 ( .A1(n7077), .A2(n7076), .ZN(n7383) );
  OR2_X1 U8887 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  NAND2_X1 U8888 ( .A1(n7383), .A2(n7078), .ZN(n10250) );
  AOI21_X1 U8889 ( .B1(n7271), .B2(n7381), .A(n9778), .ZN(n7079) );
  NAND2_X1 U8890 ( .A1(n7079), .A2(n7478), .ZN(n10247) );
  OAI22_X1 U8891 ( .A1(n10208), .A2(n7080), .B1(n7139), .B2(n10205), .ZN(n7081) );
  AOI21_X1 U8892 ( .B1(n10211), .B2(n7381), .A(n7081), .ZN(n7082) );
  OAI21_X1 U8893 ( .B1(n10247), .B2(n10213), .A(n7082), .ZN(n7083) );
  AOI21_X1 U8894 ( .B1(n10250), .B2(n10216), .A(n7083), .ZN(n7084) );
  OAI21_X1 U8895 ( .B1(n10252), .B2(n10220), .A(n7084), .ZN(P1_U3288) );
  INV_X1 U8896 ( .A(n7864), .ZN(n7873) );
  XNOR2_X1 U8897 ( .A(n7085), .B(n4427), .ZN(n7086) );
  AOI222_X1 U8898 ( .A1(n8690), .A2(n7086), .B1(n8362), .B2(n8685), .C1(n8364), 
        .C2(n8687), .ZN(n7227) );
  XNOR2_X1 U8899 ( .A(n7087), .B(n4427), .ZN(n7230) );
  NOR2_X1 U8900 ( .A1(n8633), .A2(n7228), .ZN(n7090) );
  OAI22_X1 U8901 ( .A1(n8678), .A2(n6820), .B1(n7088), .B2(n8683), .ZN(n7089)
         );
  AOI211_X1 U8902 ( .C1(n7230), .C2(n8696), .A(n7090), .B(n7089), .ZN(n7091)
         );
  OAI21_X1 U8903 ( .B1(n7227), .B2(n10310), .A(n7091), .ZN(P2_U3227) );
  OAI21_X1 U8904 ( .B1(n7093), .B2(n7092), .A(P1_STATE_REG_SCAN_IN), .ZN(n7094) );
  OAI22_X1 U8905 ( .A1(n8060), .A2(n7826), .B1(n7103), .B2(n6776), .ZN(n7117)
         );
  NAND2_X1 U8906 ( .A1(n9392), .A2(n7808), .ZN(n7095) );
  OAI21_X1 U8907 ( .B1(n7103), .B2(n7812), .A(n7095), .ZN(n7096) );
  XNOR2_X1 U8908 ( .A(n7096), .B(n7798), .ZN(n7116) );
  XOR2_X1 U8909 ( .A(n7117), .B(n7116), .Z(n7100) );
  NAND2_X1 U8910 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  NAND2_X1 U8911 ( .A1(n7099), .A2(n7100), .ZN(n7124) );
  OAI21_X1 U8912 ( .B1(n7100), .B2(n7099), .A(n7124), .ZN(n7101) );
  NAND2_X1 U8913 ( .A1(n7101), .A2(n9352), .ZN(n7107) );
  NAND2_X1 U8914 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9426) );
  INV_X1 U8915 ( .A(n9426), .ZN(n7105) );
  OAI22_X1 U8916 ( .A1(n7103), .A2(n9364), .B1(n9370), .B2(n7102), .ZN(n7104)
         );
  AOI211_X1 U8917 ( .C1(n9372), .C2(n9391), .A(n7105), .B(n7104), .ZN(n7106)
         );
  OAI211_X1 U8918 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9374), .A(n7107), .B(
        n7106), .ZN(P1_U3218) );
  INV_X1 U8919 ( .A(n7108), .ZN(n7109) );
  MUX2_X1 U8920 ( .A(n7110), .B(n7109), .S(n8678), .Z(n7114) );
  AOI22_X1 U8921 ( .A1(n10307), .A2(n7112), .B1(n10311), .B2(n7111), .ZN(n7113) );
  OAI211_X1 U8922 ( .C1(n7115), .C2(n10314), .A(n7114), .B(n7113), .ZN(
        P2_U3228) );
  INV_X1 U8923 ( .A(n7116), .ZN(n7119) );
  INV_X1 U8924 ( .A(n7117), .ZN(n7118) );
  NAND2_X1 U8925 ( .A1(n7119), .A2(n7118), .ZN(n7122) );
  AND2_X1 U8926 ( .A1(n7124), .A2(n7122), .ZN(n7126) );
  NAND2_X1 U8927 ( .A1(n9391), .A2(n7808), .ZN(n7120) );
  OAI21_X1 U8928 ( .B1(n7275), .B2(n7812), .A(n7120), .ZN(n7121) );
  AOI22_X1 U8929 ( .A1(n10210), .A2(n7808), .B1(n9391), .B2(n7807), .ZN(n7131)
         );
  NAND2_X1 U8930 ( .A1(n7124), .A2(n7123), .ZN(n7134) );
  OAI211_X1 U8931 ( .C1(n7126), .C2(n7125), .A(n9352), .B(n7134), .ZN(n7129)
         );
  AND2_X1 U8932 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9439) );
  OAI22_X1 U8933 ( .A1(n9364), .A2(n7275), .B1(n7296), .B2(n9359), .ZN(n7127)
         );
  AOI211_X1 U8934 ( .C1(n9357), .C2(n9392), .A(n9439), .B(n7127), .ZN(n7128)
         );
  OAI211_X1 U8935 ( .C1(n9374), .C2(n10206), .A(n7129), .B(n7128), .ZN(
        P1_U3230) );
  NAND2_X1 U8936 ( .A1(n7134), .A2(n7133), .ZN(n7292) );
  OAI22_X1 U8937 ( .A1(n7296), .A2(n6776), .B1(n10248), .B2(n7812), .ZN(n7135)
         );
  XNOR2_X1 U8938 ( .A(n7135), .B(n6924), .ZN(n7288) );
  OR2_X1 U8939 ( .A1(n7296), .A2(n7826), .ZN(n7137) );
  NAND2_X1 U8940 ( .A1(n7381), .A2(n7808), .ZN(n7136) );
  AND2_X1 U8941 ( .A1(n7137), .A2(n7136), .ZN(n7287) );
  INV_X1 U8942 ( .A(n7287), .ZN(n7289) );
  XNOR2_X1 U8943 ( .A(n7288), .B(n7289), .ZN(n7138) );
  XNOR2_X1 U8944 ( .A(n7292), .B(n7138), .ZN(n7145) );
  INV_X1 U8945 ( .A(n7139), .ZN(n7143) );
  AOI22_X1 U8946 ( .A1(n9372), .A2(n9389), .B1(n9376), .B2(n7381), .ZN(n7140)
         );
  NAND2_X1 U8947 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10092) );
  OAI211_X1 U8948 ( .C1(n7141), .C2(n9370), .A(n7140), .B(n10092), .ZN(n7142)
         );
  AOI21_X1 U8949 ( .B1(n7143), .B2(n9361), .A(n7142), .ZN(n7144) );
  OAI21_X1 U8950 ( .B1(n7145), .B2(n9378), .A(n7144), .ZN(P1_U3227) );
  XNOR2_X1 U8951 ( .A(n6746), .B(n10306), .ZN(n7337) );
  XNOR2_X1 U8952 ( .A(n7337), .B(n7336), .ZN(n7152) );
  INV_X1 U8953 ( .A(n7146), .ZN(n7147) );
  NAND2_X1 U8954 ( .A1(n7147), .A2(n8363), .ZN(n7148) );
  INV_X1 U8955 ( .A(n7152), .ZN(n7151) );
  AOI21_X1 U8956 ( .B1(n7152), .B2(n7150), .A(n4521), .ZN(n7158) );
  NOR2_X1 U8957 ( .A1(n8342), .A2(n7399), .ZN(n7153) );
  AOI211_X1 U8958 ( .C1(n8344), .C2(n8361), .A(n7154), .B(n7153), .ZN(n7157)
         );
  INV_X1 U8959 ( .A(n7155), .ZN(n10300) );
  AOI22_X1 U8960 ( .A1(n8353), .A2(n10306), .B1(n8332), .B2(n10300), .ZN(n7156) );
  OAI211_X1 U8961 ( .C1(n7158), .C2(n8348), .A(n7157), .B(n7156), .ZN(P2_U3153) );
  INV_X1 U8962 ( .A(n7159), .ZN(n7162) );
  OAI222_X1 U8963 ( .A1(n8878), .A2(n7160), .B1(n8874), .B2(n7162), .C1(n8485), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8964 ( .A1(n5722), .A2(P1_U3086), .B1(n8174), .B2(n7162), .C1(
        n7161), .C2(n10018), .ZN(P1_U3336) );
  OAI22_X1 U8965 ( .A1(n7166), .A2(n7165), .B1(n7164), .B2(n7163), .ZN(n7168)
         );
  INV_X1 U8966 ( .A(n9174), .ZN(n7192) );
  AOI22_X1 U8967 ( .A1(n9174), .A2(n7178), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7192), .ZN(n7167) );
  NAND2_X1 U8968 ( .A1(n7167), .A2(n7168), .ZN(n7204) );
  OAI21_X1 U8969 ( .B1(n7168), .B2(n7167), .A(n7204), .ZN(n7189) );
  AOI22_X1 U8970 ( .A1(n9174), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7448), .B2(
        n7192), .ZN(n7172) );
  AOI21_X1 U8971 ( .B1(n7173), .B2(n7172), .A(n7191), .ZN(n7177) );
  AND2_X1 U8972 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7414) );
  NOR2_X1 U8973 ( .A1(n8441), .A2(n7174), .ZN(n7175) );
  AOI211_X1 U8974 ( .C1(n8450), .C2(n9174), .A(n7414), .B(n7175), .ZN(n7176)
         );
  OAI21_X1 U8975 ( .B1(n7177), .B2(n8501), .A(n7176), .ZN(n7188) );
  MUX2_X1 U8976 ( .A(n7448), .B(n7178), .S(n8489), .Z(n7179) );
  NAND2_X1 U8977 ( .A1(n7179), .A2(n9174), .ZN(n7194) );
  INV_X1 U8978 ( .A(n7179), .ZN(n7180) );
  NAND2_X1 U8979 ( .A1(n7180), .A2(n7192), .ZN(n7181) );
  NAND2_X1 U8980 ( .A1(n7194), .A2(n7181), .ZN(n7182) );
  AOI21_X1 U8981 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7201) );
  INV_X1 U8982 ( .A(n7201), .ZN(n7186) );
  NAND3_X1 U8983 ( .A1(n7184), .A2(n7183), .A3(n7182), .ZN(n7185) );
  AOI21_X1 U8984 ( .B1(n7186), .B2(n7185), .A(n8494), .ZN(n7187) );
  AOI211_X1 U8985 ( .C1(n8499), .C2(n7189), .A(n7188), .B(n7187), .ZN(n7190)
         );
  INV_X1 U8986 ( .A(n7190), .ZN(P2_U3192) );
  AOI21_X1 U8987 ( .B1(n7503), .B2(n7193), .A(n7234), .ZN(n7212) );
  INV_X1 U8988 ( .A(n7194), .ZN(n7200) );
  MUX2_X1 U8989 ( .A(n7503), .B(n7195), .S(n8489), .Z(n7196) );
  NAND2_X1 U8990 ( .A1(n7196), .A2(n7233), .ZN(n7245) );
  INV_X1 U8991 ( .A(n7196), .ZN(n7197) );
  NAND2_X1 U8992 ( .A1(n7197), .A2(n7249), .ZN(n7198) );
  AND2_X1 U8993 ( .A1(n7245), .A2(n7198), .ZN(n7199) );
  OAI21_X1 U8994 ( .B1(n7201), .B2(n7200), .A(n7199), .ZN(n7246) );
  INV_X1 U8995 ( .A(n7246), .ZN(n7203) );
  NOR3_X1 U8996 ( .A1(n7201), .A2(n7200), .A3(n7199), .ZN(n7202) );
  OAI21_X1 U8997 ( .B1(n7203), .B2(n7202), .A(n8382), .ZN(n7211) );
  OAI21_X1 U8998 ( .B1(n9174), .B2(n7178), .A(n7204), .ZN(n7248) );
  XNOR2_X1 U8999 ( .A(n7248), .B(n7233), .ZN(n7205) );
  NAND2_X1 U9000 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7205), .ZN(n7250) );
  OAI21_X1 U9001 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7205), .A(n7250), .ZN(
        n7209) );
  INV_X1 U9002 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7206) );
  NOR2_X1 U9003 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7206), .ZN(n7625) );
  AOI21_X1 U9004 ( .B1(n8482), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7625), .ZN(
        n7207) );
  OAI21_X1 U9005 ( .B1(n7249), .B2(n8486), .A(n7207), .ZN(n7208) );
  AOI21_X1 U9006 ( .B1(n7209), .B2(n8499), .A(n7208), .ZN(n7210) );
  OAI211_X1 U9007 ( .C1(n7212), .C2(n8501), .A(n7211), .B(n7210), .ZN(P2_U3193) );
  INV_X1 U9008 ( .A(n7213), .ZN(n7217) );
  AOI21_X1 U9009 ( .B1(n7214), .B2(n7215), .A(n8009), .ZN(n7216) );
  NOR3_X1 U9010 ( .A1(n7217), .A2(n7216), .A3(n8668), .ZN(n7219) );
  OAI22_X1 U9011 ( .A1(n7336), .A2(n8671), .B1(n7442), .B2(n8673), .ZN(n7218)
         );
  NOR2_X1 U9012 ( .A1(n7219), .A2(n7218), .ZN(n7328) );
  OAI22_X1 U9013 ( .A1(n8678), .A2(n7220), .B1(n7341), .B2(n8683), .ZN(n7221)
         );
  AOI21_X1 U9014 ( .B1(n10307), .B2(n7340), .A(n7221), .ZN(n7226) );
  NAND2_X1 U9015 ( .A1(n7222), .A2(n7223), .ZN(n7224) );
  XNOR2_X1 U9016 ( .A(n7224), .B(n8009), .ZN(n7331) );
  NAND2_X1 U9017 ( .A1(n7331), .A2(n8696), .ZN(n7225) );
  OAI211_X1 U9018 ( .C1(n7328), .C2(n10320), .A(n7226), .B(n7225), .ZN(
        P2_U3225) );
  OAI21_X1 U9019 ( .B1(n7228), .B2(n8764), .A(n7227), .ZN(n7229) );
  AOI21_X1 U9020 ( .B1(n7230), .B2(n8760), .A(n7229), .ZN(n10332) );
  NAND2_X1 U9021 ( .A1(n7564), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7231) );
  OAI21_X1 U9022 ( .B1(n10332), .B2(n7564), .A(n7231), .ZN(P2_U3465) );
  NOR2_X1 U9023 ( .A1(n7233), .A2(n7232), .ZN(n7235) );
  NOR2_X1 U9024 ( .A1(n7235), .A2(n7234), .ZN(n7239) );
  OR2_X1 U9025 ( .A1(n7254), .A2(n8966), .ZN(n7350) );
  NAND2_X1 U9026 ( .A1(n7254), .A2(n8966), .ZN(n7236) );
  NAND2_X1 U9027 ( .A1(n7350), .A2(n7236), .ZN(n7238) );
  INV_X1 U9028 ( .A(n7351), .ZN(n7237) );
  AOI21_X1 U9029 ( .B1(n7239), .B2(n7238), .A(n7237), .ZN(n7262) );
  INV_X1 U9030 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7240) );
  MUX2_X1 U9031 ( .A(n8966), .B(n7240), .S(n8489), .Z(n7241) );
  NAND2_X1 U9032 ( .A1(n7241), .A2(n7254), .ZN(n7353) );
  INV_X1 U9033 ( .A(n7241), .ZN(n7242) );
  NAND2_X1 U9034 ( .A1(n7242), .A2(n7363), .ZN(n7243) );
  NAND2_X1 U9035 ( .A1(n7353), .A2(n7243), .ZN(n7244) );
  AOI21_X1 U9036 ( .B1(n7246), .B2(n7245), .A(n7244), .ZN(n7360) );
  AND3_X1 U9037 ( .A1(n7246), .A2(n7245), .A3(n7244), .ZN(n7247) );
  OAI21_X1 U9038 ( .B1(n7360), .B2(n7247), .A(n8382), .ZN(n7261) );
  NAND2_X1 U9039 ( .A1(n7249), .A2(n7248), .ZN(n7251) );
  XNOR2_X1 U9040 ( .A(n7254), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7252) );
  OAI21_X1 U9041 ( .B1(n7253), .B2(n7252), .A(n7364), .ZN(n7259) );
  INV_X1 U9042 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U9043 ( .A1(n8450), .A2(n7254), .ZN(n7256) );
  AND2_X1 U9044 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7601) );
  INV_X1 U9045 ( .A(n7601), .ZN(n7255) );
  OAI211_X1 U9046 ( .C1(n7257), .C2(n8441), .A(n7256), .B(n7255), .ZN(n7258)
         );
  AOI21_X1 U9047 ( .B1(n7259), .B2(n8499), .A(n7258), .ZN(n7260) );
  OAI211_X1 U9048 ( .C1(n7262), .C2(n8501), .A(n7261), .B(n7260), .ZN(P2_U3194) );
  INV_X1 U9049 ( .A(n7263), .ZN(n7280) );
  OAI222_X1 U9050 ( .A1(n8874), .A2(n7280), .B1(n8878), .B2(n6162), .C1(n8037), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  OR2_X1 U9051 ( .A1(n7264), .A2(n7268), .ZN(n7265) );
  AND2_X1 U9052 ( .A1(n7266), .A2(n7265), .ZN(n10204) );
  XOR2_X1 U9053 ( .A(n7267), .B(n7268), .Z(n7269) );
  AOI222_X1 U9054 ( .A1(n9927), .A2(n7269), .B1(n9390), .B2(n10234), .C1(n9392), .C2(n9929), .ZN(n10219) );
  OAI211_X1 U9055 ( .C1(n5174), .C2(n7275), .A(n9932), .B(n7271), .ZN(n10214)
         );
  OAI211_X1 U9056 ( .C1(n10233), .C2(n10204), .A(n10219), .B(n10214), .ZN(
        n7277) );
  INV_X1 U9057 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7272) );
  OAI22_X1 U9058 ( .A1(n10000), .A2(n7275), .B1(n10289), .B2(n7272), .ZN(n7273) );
  AOI21_X1 U9059 ( .B1(n7277), .B2(n10289), .A(n7273), .ZN(n7274) );
  INV_X1 U9060 ( .A(n7274), .ZN(P1_U3465) );
  OAI22_X1 U9061 ( .A1(n9935), .A2(n7275), .B1(n10296), .B2(n5489), .ZN(n7276)
         );
  AOI21_X1 U9062 ( .B1(n7277), .B2(n10296), .A(n7276), .ZN(n7278) );
  INV_X1 U9063 ( .A(n7278), .ZN(P1_U3526) );
  OAI222_X1 U9064 ( .A1(P1_U3086), .A2(n7281), .B1(n8174), .B2(n7280), .C1(
        n7279), .C2(n10018), .ZN(P1_U3335) );
  XNOR2_X1 U9065 ( .A(n7282), .B(n7798), .ZN(n7286) );
  OR2_X1 U9066 ( .A1(n7323), .A2(n7826), .ZN(n7284) );
  NAND2_X1 U9067 ( .A1(n7483), .A2(n4419), .ZN(n7283) );
  NAND2_X1 U9068 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  NOR2_X1 U9069 ( .A1(n7286), .A2(n7285), .ZN(n7311) );
  NAND2_X1 U9070 ( .A1(n7288), .A2(n7287), .ZN(n7291) );
  INV_X1 U9071 ( .A(n7288), .ZN(n7290) );
  OAI21_X1 U9072 ( .B1(n7294), .B2(n7293), .A(n7313), .ZN(n7295) );
  NAND2_X1 U9073 ( .A1(n7295), .A2(n9352), .ZN(n7300) );
  NAND2_X1 U9074 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10107) );
  INV_X1 U9075 ( .A(n10107), .ZN(n7298) );
  OAI22_X1 U9076 ( .A1(n10199), .A2(n9364), .B1(n9370), .B2(n7296), .ZN(n7297)
         );
  AOI211_X1 U9077 ( .C1(n9372), .C2(n9930), .A(n7298), .B(n7297), .ZN(n7299)
         );
  OAI211_X1 U9078 ( .C1(n9374), .C2(n10193), .A(n7300), .B(n7299), .ZN(
        P1_U3239) );
  NAND2_X1 U9079 ( .A1(n7301), .A2(n7999), .ZN(n7302) );
  XNOR2_X1 U9080 ( .A(n7303), .B(n7999), .ZN(n7307) );
  OAI22_X1 U9081 ( .A1(n7403), .A2(n8671), .B1(n7623), .B2(n8673), .ZN(n7304)
         );
  AOI21_X1 U9082 ( .B1(n7305), .B2(n10299), .A(n7304), .ZN(n7306) );
  OAI21_X1 U9083 ( .B1(n8668), .B2(n7307), .A(n7306), .ZN(n7488) );
  NAND2_X1 U9084 ( .A1(n7488), .A2(n8678), .ZN(n7310) );
  OAI22_X1 U9085 ( .A1(n8678), .A2(n7033), .B1(n7430), .B2(n8683), .ZN(n7308)
         );
  AOI21_X1 U9086 ( .B1(n10307), .B2(n7490), .A(n7308), .ZN(n7309) );
  OAI211_X1 U9087 ( .C1(n7487), .C2(n10314), .A(n7310), .B(n7309), .ZN(
        P2_U3224) );
  INV_X1 U9088 ( .A(n7311), .ZN(n7312) );
  NAND2_X1 U9089 ( .A1(n9930), .A2(n4419), .ZN(n7314) );
  OAI21_X1 U9090 ( .B1(n7547), .B2(n7812), .A(n7314), .ZN(n7315) );
  XNOR2_X1 U9091 ( .A(n7315), .B(n7798), .ZN(n7318) );
  NAND2_X1 U9092 ( .A1(n9930), .A2(n7807), .ZN(n7316) );
  OAI21_X1 U9093 ( .B1(n7547), .B2(n6776), .A(n7316), .ZN(n7317) );
  NOR2_X1 U9094 ( .A1(n7318), .A2(n7317), .ZN(n7691) );
  NAND2_X1 U9095 ( .A1(n7318), .A2(n7317), .ZN(n7690) );
  INV_X1 U9096 ( .A(n7690), .ZN(n7319) );
  NOR2_X1 U9097 ( .A1(n7691), .A2(n7319), .ZN(n7320) );
  XNOR2_X1 U9098 ( .A(n7692), .B(n7320), .ZN(n7321) );
  NAND2_X1 U9099 ( .A1(n7321), .A2(n9352), .ZN(n7326) );
  INV_X1 U9100 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7322) );
  NOR2_X1 U9101 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7322), .ZN(n10047) );
  OAI22_X1 U9102 ( .A1(n7547), .A2(n9364), .B1(n9370), .B2(n7323), .ZN(n7324)
         );
  AOI211_X1 U9103 ( .C1(n9372), .C2(n9388), .A(n10047), .B(n7324), .ZN(n7325)
         );
  OAI211_X1 U9104 ( .C1(n9374), .C2(n7386), .A(n7326), .B(n7325), .ZN(P1_U3213) );
  INV_X1 U9105 ( .A(n6172), .ZN(n7334) );
  OAI222_X1 U9106 ( .A1(n8874), .A2(n7334), .B1(P2_U3151), .B2(n4855), .C1(
        n7327), .C2(n8878), .ZN(P2_U3274) );
  INV_X1 U9107 ( .A(n7340), .ZN(n7329) );
  OAI21_X1 U9108 ( .B1(n7329), .B2(n8764), .A(n7328), .ZN(n7330) );
  AOI21_X1 U9109 ( .B1(n8760), .B2(n7331), .A(n7330), .ZN(n10335) );
  NAND2_X1 U9110 ( .A1(n7564), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7332) );
  OAI21_X1 U9111 ( .B1(n10335), .B2(n7564), .A(n7332), .ZN(P2_U3467) );
  OAI222_X1 U9112 ( .A1(n7335), .A2(P1_U3086), .B1(n8174), .B2(n7334), .C1(
        n7333), .C2(n10018), .ZN(P1_U3334) );
  NAND2_X1 U9113 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  XNOR2_X1 U9114 ( .A(n6746), .B(n7340), .ZN(n7404) );
  INV_X1 U9115 ( .A(n7404), .ZN(n7423) );
  XNOR2_X1 U9116 ( .A(n7411), .B(n7423), .ZN(n7424) );
  XNOR2_X1 U9117 ( .A(n7424), .B(n8361), .ZN(n7348) );
  AOI21_X1 U9118 ( .B1(n8331), .B2(n8362), .A(n7339), .ZN(n7346) );
  NAND2_X1 U9119 ( .A1(n8353), .A2(n7340), .ZN(n7345) );
  INV_X1 U9120 ( .A(n7341), .ZN(n7342) );
  NAND2_X1 U9121 ( .A1(n8332), .A2(n7342), .ZN(n7344) );
  NAND2_X1 U9122 ( .A1(n8344), .A2(n7425), .ZN(n7343) );
  NAND4_X1 U9123 ( .A1(n7346), .A2(n7345), .A3(n7344), .A4(n7343), .ZN(n7347)
         );
  AOI21_X1 U9124 ( .B1(n7348), .B2(n8315), .A(n7347), .ZN(n7349) );
  INV_X1 U9125 ( .A(n7349), .ZN(P2_U3161) );
  NOR2_X1 U9126 ( .A1(n7354), .A2(n7352), .ZN(n7510) );
  AOI21_X1 U9127 ( .B1(n7354), .B2(n7352), .A(n7510), .ZN(n7374) );
  INV_X1 U9128 ( .A(n7353), .ZN(n7359) );
  MUX2_X1 U9129 ( .A(n7354), .B(n8754), .S(n8489), .Z(n7355) );
  NAND2_X1 U9130 ( .A1(n7355), .A2(n7509), .ZN(n7527) );
  INV_X1 U9131 ( .A(n7355), .ZN(n7356) );
  NAND2_X1 U9132 ( .A1(n7356), .A2(n7516), .ZN(n7357) );
  AND2_X1 U9133 ( .A1(n7527), .A2(n7357), .ZN(n7358) );
  OAI21_X1 U9134 ( .B1(n7360), .B2(n7359), .A(n7358), .ZN(n7528) );
  INV_X1 U9135 ( .A(n7528), .ZN(n7362) );
  NOR3_X1 U9136 ( .A1(n7360), .A2(n7359), .A3(n7358), .ZN(n7361) );
  OAI21_X1 U9137 ( .B1(n7362), .B2(n7361), .A(n8382), .ZN(n7373) );
  NAND2_X1 U9138 ( .A1(n7363), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7365) );
  NAND2_X1 U9139 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7366), .ZN(n7517) );
  OAI21_X1 U9140 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7366), .A(n7517), .ZN(
        n7371) );
  INV_X1 U9141 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U9142 ( .A1(n8450), .A2(n7509), .ZN(n7368) );
  AND2_X1 U9143 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7659) );
  INV_X1 U9144 ( .A(n7659), .ZN(n7367) );
  OAI211_X1 U9145 ( .C1(n7369), .C2(n8441), .A(n7368), .B(n7367), .ZN(n7370)
         );
  AOI21_X1 U9146 ( .B1(n7371), .B2(n8499), .A(n7370), .ZN(n7372) );
  OAI211_X1 U9147 ( .C1(n7374), .C2(n8501), .A(n7373), .B(n7372), .ZN(P2_U3195) );
  INV_X1 U9148 ( .A(n7375), .ZN(n7378) );
  OAI21_X1 U9149 ( .B1(n7378), .B2(n7377), .A(n7376), .ZN(n7379) );
  NOR2_X1 U9150 ( .A1(n7379), .A2(n7384), .ZN(n9921) );
  AOI21_X1 U9151 ( .B1(n7384), .B2(n7379), .A(n9921), .ZN(n7380) );
  NOR2_X1 U9152 ( .A1(n7380), .A2(n10283), .ZN(n7543) );
  INV_X1 U9153 ( .A(n7543), .ZN(n7394) );
  NAND2_X1 U9154 ( .A1(n7296), .A2(n10248), .ZN(n7382) );
  OAI21_X1 U9155 ( .B1(n7385), .B2(n7384), .A(n7457), .ZN(n7545) );
  OAI211_X1 U9156 ( .C1(n7477), .C2(n7547), .A(n9932), .B(n9931), .ZN(n7542)
         );
  NOR2_X1 U9157 ( .A1(n10205), .A2(n7386), .ZN(n7387) );
  AOI21_X1 U9158 ( .B1(n10220), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7387), .ZN(
        n7388) );
  OAI21_X1 U9159 ( .B1(n10198), .B2(n7547), .A(n7388), .ZN(n7389) );
  INV_X1 U9160 ( .A(n7389), .ZN(n7391) );
  INV_X1 U9161 ( .A(n9779), .ZN(n8065) );
  AOI22_X1 U9162 ( .A1(n9784), .A2(n9388), .B1(n8065), .B2(n9389), .ZN(n7390)
         );
  OAI211_X1 U9163 ( .C1(n7542), .C2(n10213), .A(n7391), .B(n7390), .ZN(n7392)
         );
  AOI21_X1 U9164 ( .B1(n7545), .B2(n10216), .A(n7392), .ZN(n7393) );
  OAI21_X1 U9165 ( .B1(n7394), .B2(n10220), .A(n7393), .ZN(P1_U3286) );
  OAI21_X1 U9166 ( .B1(n7395), .B2(n8007), .A(n7222), .ZN(n10303) );
  INV_X1 U9167 ( .A(n10303), .ZN(n10298) );
  NAND2_X1 U9168 ( .A1(n8361), .A2(n8685), .ZN(n10302) );
  OAI21_X1 U9169 ( .B1(n7396), .B2(n8764), .A(n10302), .ZN(n7401) );
  INV_X1 U9170 ( .A(n7214), .ZN(n7397) );
  AOI21_X1 U9171 ( .B1(n8007), .B2(n7398), .A(n7397), .ZN(n7400) );
  OAI22_X1 U9172 ( .A1(n7400), .A2(n8668), .B1(n7399), .B2(n8671), .ZN(n10297)
         );
  AOI211_X1 U9173 ( .C1(n10298), .C2(n8760), .A(n7401), .B(n10297), .ZN(n10334) );
  OR2_X1 U9174 ( .A1(n10334), .A2(n7564), .ZN(n7402) );
  OAI21_X1 U9175 ( .B1(n8772), .B2(n6808), .A(n7402), .ZN(P2_U3466) );
  XNOR2_X1 U9176 ( .A(n7490), .B(n6746), .ZN(n7426) );
  AOI22_X1 U9177 ( .A1(n7426), .A2(n7442), .B1(n7403), .B2(n7404), .ZN(n7410)
         );
  OAI21_X1 U9178 ( .B1(n7404), .B2(n7403), .A(n7442), .ZN(n7406) );
  INV_X1 U9179 ( .A(n7426), .ZN(n7405) );
  NAND2_X1 U9180 ( .A1(n7406), .A2(n7405), .ZN(n7408) );
  NAND3_X1 U9181 ( .A1(n7423), .A2(n7425), .A3(n8361), .ZN(n7407) );
  NAND2_X1 U9182 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  NAND2_X1 U9183 ( .A1(n7412), .A2(n7623), .ZN(n7595) );
  NAND2_X1 U9184 ( .A1(n4520), .A2(n7595), .ZN(n7413) );
  XNOR2_X1 U9185 ( .A(n7450), .B(n8106), .ZN(n7596) );
  XNOR2_X1 U9186 ( .A(n7413), .B(n7596), .ZN(n7421) );
  NAND2_X1 U9187 ( .A1(n7450), .A2(n8353), .ZN(n7419) );
  AOI21_X1 U9188 ( .B1(n8331), .B2(n7425), .A(n7414), .ZN(n7418) );
  INV_X1 U9189 ( .A(n7447), .ZN(n7415) );
  NAND2_X1 U9190 ( .A1(n8332), .A2(n7415), .ZN(n7417) );
  NAND2_X1 U9191 ( .A1(n8344), .A2(n8359), .ZN(n7416) );
  NAND4_X1 U9192 ( .A1(n7419), .A2(n7418), .A3(n7417), .A4(n7416), .ZN(n7420)
         );
  AOI21_X1 U9193 ( .B1(n7421), .B2(n8315), .A(n7420), .ZN(n7422) );
  INV_X1 U9194 ( .A(n7422), .ZN(P2_U3157) );
  OAI22_X1 U9195 ( .A1(n7424), .A2(n8361), .B1(n7411), .B2(n7423), .ZN(n7428)
         );
  XNOR2_X1 U9196 ( .A(n7426), .B(n7425), .ZN(n7427) );
  XNOR2_X1 U9197 ( .A(n7428), .B(n7427), .ZN(n7437) );
  AOI21_X1 U9198 ( .B1(n8331), .B2(n8361), .A(n7429), .ZN(n7435) );
  NAND2_X1 U9199 ( .A1(n8353), .A2(n7490), .ZN(n7434) );
  INV_X1 U9200 ( .A(n7430), .ZN(n7431) );
  NAND2_X1 U9201 ( .A1(n8332), .A2(n7431), .ZN(n7433) );
  NAND2_X1 U9202 ( .A1(n8344), .A2(n8360), .ZN(n7432) );
  NAND4_X1 U9203 ( .A1(n7435), .A2(n7434), .A3(n7433), .A4(n7432), .ZN(n7436)
         );
  AOI21_X1 U9204 ( .B1(n7437), .B2(n8315), .A(n7436), .ZN(n7438) );
  INV_X1 U9205 ( .A(n7438), .ZN(P2_U3171) );
  NAND2_X1 U9206 ( .A1(n7439), .A2(n7881), .ZN(n7440) );
  AND2_X1 U9207 ( .A1(n7897), .A2(n7895), .ZN(n8012) );
  XNOR2_X1 U9208 ( .A(n7440), .B(n8012), .ZN(n7471) );
  XOR2_X1 U9209 ( .A(n8012), .B(n7441), .Z(n7444) );
  OAI22_X1 U9210 ( .A1(n7442), .A2(n8671), .B1(n7599), .B2(n8673), .ZN(n7443)
         );
  AOI21_X1 U9211 ( .B1(n7444), .B2(n8690), .A(n7443), .ZN(n7445) );
  OAI21_X1 U9212 ( .B1(n7471), .B2(n7446), .A(n7445), .ZN(n7473) );
  NAND2_X1 U9213 ( .A1(n7473), .A2(n8678), .ZN(n7452) );
  OAI22_X1 U9214 ( .A1(n8678), .A2(n7448), .B1(n7447), .B2(n8683), .ZN(n7449)
         );
  AOI21_X1 U9215 ( .B1(n10307), .B2(n7450), .A(n7449), .ZN(n7451) );
  OAI211_X1 U9216 ( .C1(n7471), .C2(n10314), .A(n7452), .B(n7451), .ZN(
        P2_U3223) );
  NAND2_X1 U9217 ( .A1(n7454), .A2(n7453), .ZN(n7461) );
  OAI21_X1 U9218 ( .B1(n9921), .B2(n7455), .A(n7458), .ZN(n7456) );
  XOR2_X1 U9219 ( .A(n7461), .B(n7456), .Z(n7570) );
  INV_X1 U9220 ( .A(n9751), .ZN(n9789) );
  NAND2_X1 U9221 ( .A1(n7457), .A2(n4456), .ZN(n9920) );
  NAND2_X1 U9222 ( .A1(n7459), .A2(n7458), .ZN(n9925) );
  NAND2_X1 U9223 ( .A1(n9920), .A2(n9925), .ZN(n9919) );
  NAND2_X1 U9224 ( .A1(n9294), .A2(n4418), .ZN(n7460) );
  NAND2_X1 U9225 ( .A1(n9919), .A2(n7460), .ZN(n7462) );
  NAND2_X1 U9226 ( .A1(n7462), .A2(n7461), .ZN(n7582) );
  OAI21_X1 U9227 ( .B1(n7462), .B2(n7461), .A(n7582), .ZN(n7568) );
  AOI21_X1 U9228 ( .B1(n10234), .B2(n9387), .A(n7463), .ZN(n7566) );
  NOR2_X1 U9229 ( .A1(n9779), .A2(n9294), .ZN(n7466) );
  OAI22_X1 U9230 ( .A1(n10208), .A2(n7464), .B1(n9297), .B2(n10205), .ZN(n7465) );
  AOI211_X1 U9231 ( .C1(n10211), .C2(n4416), .A(n7466), .B(n7465), .ZN(n7467)
         );
  OAI21_X1 U9232 ( .B1(n7566), .B2(n10213), .A(n7467), .ZN(n7468) );
  AOI21_X1 U9233 ( .B1(n10216), .B2(n7568), .A(n7468), .ZN(n7469) );
  OAI21_X1 U9234 ( .B1(n7570), .B2(n9789), .A(n7469), .ZN(P1_U3284) );
  OAI22_X1 U9235 ( .A1(n7471), .A2(n7486), .B1(n7470), .B2(n8764), .ZN(n7472)
         );
  NOR2_X1 U9236 ( .A1(n7473), .A2(n7472), .ZN(n10339) );
  NAND2_X1 U9237 ( .A1(n7564), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7474) );
  OAI21_X1 U9238 ( .B1(n10339), .B2(n7564), .A(n7474), .ZN(P2_U3469) );
  OAI21_X1 U9239 ( .B1(n7476), .B2(n7479), .A(n7475), .ZN(n10201) );
  AOI211_X1 U9240 ( .C1(n7483), .C2(n7478), .A(n9778), .B(n7477), .ZN(n10192)
         );
  XNOR2_X1 U9241 ( .A(n7375), .B(n7479), .ZN(n7480) );
  AOI222_X1 U9242 ( .A1(n9927), .A2(n7480), .B1(n9930), .B2(n10234), .C1(n9390), .C2(n9929), .ZN(n10203) );
  INV_X1 U9243 ( .A(n10203), .ZN(n7481) );
  AOI211_X1 U9244 ( .C1(n10285), .C2(n10201), .A(n10192), .B(n7481), .ZN(n7485) );
  AOI22_X1 U9245 ( .A1(n9833), .A2(n7483), .B1(n5414), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7482) );
  OAI21_X1 U9246 ( .B1(n7485), .B2(n5414), .A(n7482), .ZN(P1_U3528) );
  AOI22_X1 U9247 ( .A1(n9955), .A2(n7483), .B1(n10287), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n7484) );
  OAI21_X1 U9248 ( .B1(n7485), .B2(n10287), .A(n7484), .ZN(P1_U3471) );
  NOR2_X1 U9249 ( .A1(n7487), .A2(n7486), .ZN(n7489) );
  AOI211_X1 U9250 ( .C1(n8766), .C2(n7490), .A(n7489), .B(n7488), .ZN(n10337)
         );
  OR2_X1 U9251 ( .A1(n10337), .A2(n7564), .ZN(n7491) );
  OAI21_X1 U9252 ( .B1(n8772), .B2(n7165), .A(n7491), .ZN(P2_U3468) );
  NAND2_X1 U9253 ( .A1(n7495), .A2(n10013), .ZN(n7493) );
  OAI211_X1 U9254 ( .C1(n7494), .C2(n10009), .A(n7493), .B(n7492), .ZN(
        P1_U3332) );
  NAND2_X1 U9255 ( .A1(n7495), .A2(n9175), .ZN(n7497) );
  NAND2_X1 U9256 ( .A1(n7496), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8045) );
  OAI211_X1 U9257 ( .C1(n7498), .C2(n8878), .A(n7497), .B(n8045), .ZN(P2_U3272) );
  XNOR2_X1 U9258 ( .A(n7499), .B(n7500), .ZN(n7562) );
  INV_X1 U9259 ( .A(n7562), .ZN(n7507) );
  XNOR2_X1 U9260 ( .A(n7501), .B(n8014), .ZN(n7502) );
  OAI222_X1 U9261 ( .A1(n8673), .A2(n7657), .B1(n8671), .B2(n7623), .C1(n7502), 
        .C2(n8668), .ZN(n7560) );
  NAND2_X1 U9262 ( .A1(n7560), .A2(n8678), .ZN(n7506) );
  OAI22_X1 U9263 ( .A1(n8678), .A2(n7503), .B1(n7627), .B2(n8683), .ZN(n7504)
         );
  AOI21_X1 U9264 ( .B1(n7633), .B2(n10307), .A(n7504), .ZN(n7505) );
  OAI211_X1 U9265 ( .C1(n7507), .C2(n8666), .A(n7506), .B(n7505), .ZN(P2_U3222) );
  NOR2_X1 U9266 ( .A1(n7509), .A2(n7508), .ZN(n7511) );
  NAND2_X1 U9267 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8371), .ZN(n7512) );
  OAI21_X1 U9268 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8371), .A(n7512), .ZN(
        n7513) );
  NOR2_X1 U9269 ( .A1(n7514), .A2(n7513), .ZN(n8369) );
  AOI21_X1 U9270 ( .B1(n7514), .B2(n7513), .A(n8369), .ZN(n7535) );
  AOI22_X1 U9271 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8371), .B1(n7522), .B2(
        n9020), .ZN(n7520) );
  NAND2_X1 U9272 ( .A1(n7516), .A2(n7515), .ZN(n7518) );
  OAI21_X1 U9273 ( .B1(n7520), .B2(n7519), .A(n8372), .ZN(n7533) );
  NAND2_X1 U9274 ( .A1(n8482), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U9275 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8217) );
  OAI211_X1 U9276 ( .C1(n8486), .C2(n8371), .A(n7521), .B(n8217), .ZN(n7532)
         );
  MUX2_X1 U9277 ( .A(n8677), .B(n9020), .S(n8489), .Z(n7523) );
  NAND2_X1 U9278 ( .A1(n7523), .A2(n7522), .ZN(n8375) );
  INV_X1 U9279 ( .A(n7523), .ZN(n7524) );
  NAND2_X1 U9280 ( .A1(n7524), .A2(n8371), .ZN(n7525) );
  NAND2_X1 U9281 ( .A1(n8375), .A2(n7525), .ZN(n7526) );
  AOI21_X1 U9282 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n8381) );
  INV_X1 U9283 ( .A(n8381), .ZN(n7530) );
  NAND3_X1 U9284 ( .A1(n7528), .A2(n7527), .A3(n7526), .ZN(n7529) );
  AOI21_X1 U9285 ( .B1(n7530), .B2(n7529), .A(n8494), .ZN(n7531) );
  AOI211_X1 U9286 ( .C1(n8499), .C2(n7533), .A(n7532), .B(n7531), .ZN(n7534)
         );
  OAI21_X1 U9287 ( .B1(n7535), .B2(n8501), .A(n7534), .ZN(P2_U3196) );
  INV_X1 U9288 ( .A(n7536), .ZN(n7539) );
  OAI222_X1 U9289 ( .A1(P1_U3086), .A2(n7538), .B1(n8174), .B2(n7539), .C1(
        n7537), .C2(n10018), .ZN(P1_U3333) );
  OAI222_X1 U9290 ( .A1(n8878), .A2(n7540), .B1(n8874), .B2(n7539), .C1(n4857), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  AOI22_X1 U9291 ( .A1(n9929), .A2(n9389), .B1(n9388), .B2(n10234), .ZN(n7541)
         );
  NAND2_X1 U9292 ( .A1(n7542), .A2(n7541), .ZN(n7544) );
  AOI211_X1 U9293 ( .C1(n10285), .C2(n7545), .A(n7544), .B(n7543), .ZN(n7552)
         );
  INV_X1 U9294 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7546) );
  OAI22_X1 U9295 ( .A1(n10000), .A2(n7547), .B1(n10289), .B2(n7546), .ZN(n7548) );
  INV_X1 U9296 ( .A(n7548), .ZN(n7549) );
  OAI21_X1 U9297 ( .B1(n7552), .B2(n10287), .A(n7549), .ZN(P1_U3474) );
  AOI22_X1 U9298 ( .A1(n9833), .A2(n7550), .B1(n5414), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7551) );
  OAI21_X1 U9299 ( .B1(n7552), .B2(n5414), .A(n7551), .ZN(P1_U3529) );
  XNOR2_X1 U9300 ( .A(n7553), .B(n6069), .ZN(n7554) );
  AOI222_X1 U9301 ( .A1(n8690), .A2(n7554), .B1(n8359), .B2(n8687), .C1(n8358), 
        .C2(n8685), .ZN(n8763) );
  OAI22_X1 U9302 ( .A1(n8678), .A2(n8966), .B1(n7603), .B2(n8683), .ZN(n7555)
         );
  AOI21_X1 U9303 ( .B1(n7906), .B2(n10307), .A(n7555), .ZN(n7559) );
  NAND2_X1 U9304 ( .A1(n7556), .A2(n7557), .ZN(n8759) );
  NAND3_X1 U9305 ( .A1(n8761), .A2(n8759), .A3(n8696), .ZN(n7558) );
  OAI211_X1 U9306 ( .C1(n8763), .C2(n10320), .A(n7559), .B(n7558), .ZN(
        P2_U3221) );
  AOI21_X1 U9307 ( .B1(n8766), .B2(n7633), .A(n7560), .ZN(n7565) );
  NAND2_X1 U9308 ( .A1(n10338), .A2(n8760), .ZN(n8851) );
  INV_X1 U9309 ( .A(n8851), .ZN(n8863) );
  AOI22_X1 U9310 ( .A1(n7562), .A2(n8863), .B1(P2_REG0_REG_11__SCAN_IN), .B2(
        n10341), .ZN(n7561) );
  OAI21_X1 U9311 ( .B1(n7565), .B2(n10341), .A(n7561), .ZN(P2_U3423) );
  NAND2_X1 U9312 ( .A1(n8772), .A2(n8760), .ZN(n8750) );
  INV_X1 U9313 ( .A(n8750), .ZN(n8756) );
  AOI22_X1 U9314 ( .A1(n7562), .A2(n8756), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n7564), .ZN(n7563) );
  OAI21_X1 U9315 ( .B1(n7565), .B2(n7564), .A(n7563), .ZN(P2_U3470) );
  OAI21_X1 U9316 ( .B1(n9294), .B2(n10273), .A(n7566), .ZN(n7567) );
  AOI21_X1 U9317 ( .B1(n7568), .B2(n10285), .A(n7567), .ZN(n7569) );
  OAI21_X1 U9318 ( .B1(n7570), .B2(n10283), .A(n7569), .ZN(n7576) );
  INV_X1 U9319 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7571) );
  OAI22_X1 U9320 ( .A1(n9935), .A2(n7699), .B1(n10296), .B2(n7571), .ZN(n7572)
         );
  AOI21_X1 U9321 ( .B1(n7576), .B2(n10296), .A(n7572), .ZN(n7573) );
  INV_X1 U9322 ( .A(n7573), .ZN(P1_U3531) );
  INV_X1 U9323 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7574) );
  OAI22_X1 U9324 ( .A1(n10000), .A2(n7699), .B1(n10289), .B2(n7574), .ZN(n7575) );
  AOI21_X1 U9325 ( .B1(n7576), .B2(n10289), .A(n7575), .ZN(n7577) );
  INV_X1 U9326 ( .A(n7577), .ZN(P1_U3480) );
  INV_X1 U9327 ( .A(n7578), .ZN(n7579) );
  AOI21_X1 U9328 ( .B1(n7583), .B2(n7580), .A(n7579), .ZN(n7640) );
  NAND2_X1 U9329 ( .A1(n9232), .A2(n7699), .ZN(n7581) );
  NAND2_X1 U9330 ( .A1(n7582), .A2(n7581), .ZN(n7584) );
  OAI21_X1 U9331 ( .B1(n7584), .B2(n7583), .A(n7609), .ZN(n7642) );
  NAND2_X1 U9332 ( .A1(n7642), .A2(n10216), .ZN(n7594) );
  NAND2_X1 U9333 ( .A1(n9784), .A2(n8119), .ZN(n7587) );
  INV_X1 U9334 ( .A(n7585), .ZN(n9210) );
  AOI22_X1 U9335 ( .A1(n9728), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9210), .B2(
        n10194), .ZN(n7586) );
  OAI211_X1 U9336 ( .C1(n9232), .C2(n9779), .A(n7587), .B(n7586), .ZN(n7592)
         );
  OAI21_X1 U9337 ( .B1(n7588), .B2(n7607), .A(n9932), .ZN(n7590) );
  OR2_X1 U9338 ( .A1(n7590), .A2(n7589), .ZN(n7638) );
  NOR2_X1 U9339 ( .A1(n7638), .A2(n10213), .ZN(n7591) );
  AOI211_X1 U9340 ( .C1(n10211), .C2(n9200), .A(n7592), .B(n7591), .ZN(n7593)
         );
  OAI211_X1 U9341 ( .C1(n7640), .C2(n9789), .A(n7594), .B(n7593), .ZN(P1_U3283) );
  XNOR2_X1 U9342 ( .A(n8014), .B(n6746), .ZN(n7629) );
  XOR2_X1 U9343 ( .A(n8106), .B(n7906), .Z(n7653) );
  XNOR2_X1 U9344 ( .A(n7653), .B(n7657), .ZN(n7598) );
  XNOR2_X1 U9345 ( .A(n4510), .B(n7598), .ZN(n7606) );
  NOR2_X1 U9346 ( .A1(n8342), .A2(n7599), .ZN(n7600) );
  AOI211_X1 U9347 ( .C1(n8344), .C2(n8358), .A(n7601), .B(n7600), .ZN(n7602)
         );
  OAI21_X1 U9348 ( .B1(n7603), .B2(n8346), .A(n7602), .ZN(n7604) );
  AOI21_X1 U9349 ( .B1(n7906), .B2(n8353), .A(n7604), .ZN(n7605) );
  OAI21_X1 U9350 ( .B1(n7606), .B2(n8348), .A(n7605), .ZN(P2_U3164) );
  NAND2_X1 U9351 ( .A1(n10254), .A2(n7607), .ZN(n7608) );
  XNOR2_X1 U9352 ( .A(n8121), .B(n7610), .ZN(n10261) );
  INV_X1 U9353 ( .A(n7589), .ZN(n7611) );
  AOI211_X1 U9354 ( .C1(n10257), .C2(n7611), .A(n9778), .B(n4516), .ZN(n10255)
         );
  INV_X1 U9355 ( .A(n10274), .ZN(n9386) );
  NOR2_X1 U9356 ( .A1(n9779), .A2(n10254), .ZN(n7614) );
  OAI22_X1 U9357 ( .A1(n10208), .A2(n7612), .B1(n9339), .B2(n10205), .ZN(n7613) );
  AOI211_X1 U9358 ( .C1(n9784), .C2(n9386), .A(n7614), .B(n7613), .ZN(n7615)
         );
  OAI21_X1 U9359 ( .B1(n8118), .B2(n10198), .A(n7615), .ZN(n7621) );
  AOI21_X1 U9360 ( .B1(n7617), .B2(n7616), .A(n10283), .ZN(n7619) );
  NAND2_X1 U9361 ( .A1(n7619), .A2(n7618), .ZN(n10258) );
  NOR2_X1 U9362 ( .A1(n10258), .A2(n10220), .ZN(n7620) );
  AOI211_X1 U9363 ( .C1(n10255), .C2(n10191), .A(n7621), .B(n7620), .ZN(n7622)
         );
  OAI21_X1 U9364 ( .B1(n10261), .B2(n9753), .A(n7622), .ZN(P1_U3282) );
  NOR2_X1 U9365 ( .A1(n8342), .A2(n7623), .ZN(n7624) );
  AOI211_X1 U9366 ( .C1(n8344), .C2(n8688), .A(n7625), .B(n7624), .ZN(n7626)
         );
  OAI21_X1 U9367 ( .B1(n7627), .B2(n8346), .A(n7626), .ZN(n7632) );
  AOI211_X1 U9368 ( .C1(n7630), .C2(n7629), .A(n8348), .B(n7628), .ZN(n7631)
         );
  AOI211_X1 U9369 ( .C1(n7633), .C2(n8353), .A(n7632), .B(n7631), .ZN(n7634)
         );
  INV_X1 U9370 ( .A(n7634), .ZN(P2_U3176) );
  INV_X1 U9371 ( .A(n7635), .ZN(n7652) );
  OAI222_X1 U9372 ( .A1(n7637), .A2(P1_U3086), .B1(n8174), .B2(n7652), .C1(
        n7636), .C2(n10018), .ZN(P1_U3331) );
  AOI22_X1 U9373 ( .A1(n9929), .A2(n9928), .B1(n8119), .B2(n10234), .ZN(n7639)
         );
  OAI211_X1 U9374 ( .C1(n7640), .C2(n10283), .A(n7639), .B(n7638), .ZN(n7641)
         );
  AOI21_X1 U9375 ( .B1(n7642), .B2(n10285), .A(n7641), .ZN(n7644) );
  MUX2_X1 U9376 ( .A(n5551), .B(n7644), .S(n10296), .Z(n7643) );
  OAI21_X1 U9377 ( .B1(n7607), .B2(n9935), .A(n7643), .ZN(P1_U3532) );
  INV_X1 U9378 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7645) );
  MUX2_X1 U9379 ( .A(n7645), .B(n7644), .S(n10289), .Z(n7646) );
  OAI21_X1 U9380 ( .B1(n7607), .B2(n10000), .A(n7646), .ZN(P1_U3483) );
  INV_X1 U9381 ( .A(n7647), .ZN(n8048) );
  OAI222_X1 U9382 ( .A1(n8874), .A2(n8048), .B1(P2_U3151), .B2(n7649), .C1(
        n7648), .C2(n8878), .ZN(P2_U3270) );
  OAI222_X1 U9383 ( .A1(n8874), .A2(n7652), .B1(P2_U3151), .B2(n7651), .C1(
        n7650), .C2(n8878), .ZN(P2_U3271) );
  XNOR2_X1 U9384 ( .A(n8861), .B(n8106), .ZN(n7654) );
  NOR2_X1 U9385 ( .A1(n7654), .A2(n8358), .ZN(n8071) );
  INV_X1 U9386 ( .A(n8071), .ZN(n7655) );
  NAND2_X1 U9387 ( .A1(n7654), .A2(n8358), .ZN(n8070) );
  NAND2_X1 U9388 ( .A1(n7655), .A2(n8070), .ZN(n7656) );
  XNOR2_X1 U9389 ( .A(n8072), .B(n7656), .ZN(n7663) );
  NOR2_X1 U9390 ( .A1(n8342), .A2(n7657), .ZN(n7658) );
  AOI211_X1 U9391 ( .C1(n8344), .C2(n8686), .A(n7659), .B(n7658), .ZN(n7660)
         );
  OAI21_X1 U9392 ( .B1(n8682), .B2(n8346), .A(n7660), .ZN(n7661) );
  AOI21_X1 U9393 ( .B1(n8861), .B2(n8353), .A(n7661), .ZN(n7662) );
  OAI21_X1 U9394 ( .B1(n7663), .B2(n8348), .A(n7662), .ZN(P2_U3174) );
  NAND3_X1 U9395 ( .A1(n7664), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9396 ( .A1(n10014), .A2(n9175), .ZN(n7666) );
  NAND2_X1 U9397 ( .A1(n9173), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7665) );
  OAI211_X1 U9398 ( .C1(n5902), .C2(n7667), .A(n7666), .B(n7665), .ZN(P2_U3264) );
  INV_X1 U9399 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7671) );
  INV_X1 U9400 ( .A(n7669), .ZN(n7670) );
  NAND2_X1 U9401 ( .A1(n7670), .A2(n10311), .ZN(n7688) );
  OAI21_X1 U9402 ( .B1(n8678), .B2(n7671), .A(n7688), .ZN(n7674) );
  NOR2_X1 U9403 ( .A1(n7672), .A2(n8666), .ZN(n7673) );
  AOI211_X1 U9404 ( .C1(n10307), .C2(n7675), .A(n7674), .B(n7673), .ZN(n7676)
         );
  OAI21_X1 U9405 ( .B1(n7668), .B2(n10310), .A(n7676), .ZN(P2_U3204) );
  NAND2_X1 U9406 ( .A1(n5943), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7681) );
  INV_X1 U9407 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7678) );
  OR2_X1 U9408 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  OAI211_X1 U9409 ( .C1(n9045), .C2(n6323), .A(n7681), .B(n7680), .ZN(n7682)
         );
  INV_X1 U9410 ( .A(n7682), .ZN(n7683) );
  NAND2_X1 U9411 ( .A1(n7684), .A2(n7683), .ZN(n8355) );
  INV_X1 U9412 ( .A(n7685), .ZN(n7686) );
  NAND2_X1 U9413 ( .A1(n8355), .A2(n7686), .ZN(n8700) );
  NOR2_X1 U9414 ( .A1(n8700), .A2(n10341), .ZN(n8774) );
  AOI21_X1 U9415 ( .B1(n10341), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8774), .ZN(
        n7687) );
  OAI21_X1 U9416 ( .B1(n8699), .B2(n8835), .A(n7687), .ZN(P2_U3458) );
  AOI21_X1 U9417 ( .B1(n7688), .B2(n8700), .A(n10320), .ZN(n8503) );
  AOI21_X1 U9418 ( .B1(n10320), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8503), .ZN(
        n7689) );
  OAI21_X1 U9419 ( .B1(n8699), .B2(n8633), .A(n7689), .ZN(P2_U3202) );
  OR2_X1 U9420 ( .A1(n9294), .A2(n7826), .ZN(n7694) );
  NAND2_X1 U9421 ( .A1(n10184), .A2(n7808), .ZN(n7693) );
  NAND2_X1 U9422 ( .A1(n7694), .A2(n7693), .ZN(n7701) );
  INV_X1 U9423 ( .A(n7701), .ZN(n9229) );
  OAI22_X1 U9424 ( .A1(n9294), .A2(n6776), .B1(n4418), .B2(n7812), .ZN(n7695)
         );
  XNOR2_X1 U9425 ( .A(n7695), .B(n7798), .ZN(n9289) );
  INV_X1 U9426 ( .A(n9289), .ZN(n9227) );
  NAND2_X1 U9427 ( .A1(n4416), .A2(n7821), .ZN(n7697) );
  OAI21_X1 U9428 ( .B1(n9232), .B2(n6776), .A(n7697), .ZN(n7698) );
  XNOR2_X1 U9429 ( .A(n7698), .B(n6924), .ZN(n9291) );
  OAI22_X1 U9430 ( .A1(n9232), .A2(n7826), .B1(n7699), .B2(n6776), .ZN(n7700)
         );
  INV_X1 U9431 ( .A(n7700), .ZN(n9290) );
  OAI22_X1 U9432 ( .A1(n9229), .A2(n9227), .B1(n9291), .B2(n9290), .ZN(n7705)
         );
  OAI21_X1 U9433 ( .B1(n9289), .B2(n7701), .A(n7700), .ZN(n7703) );
  NOR3_X1 U9434 ( .A1(n9289), .A2(n7701), .A3(n7700), .ZN(n7702) );
  AOI21_X1 U9435 ( .B1(n9291), .B2(n7703), .A(n7702), .ZN(n7704) );
  AOI22_X1 U9436 ( .A1(n10257), .A2(n7821), .B1(n4419), .B2(n8119), .ZN(n7706)
         );
  XOR2_X1 U9437 ( .A(n7798), .B(n7706), .Z(n9335) );
  OR2_X1 U9438 ( .A1(n8118), .A2(n6776), .ZN(n7708) );
  OR2_X1 U9439 ( .A1(n9794), .A2(n7826), .ZN(n7707) );
  NAND2_X1 U9440 ( .A1(n7708), .A2(n7707), .ZN(n7717) );
  NAND2_X1 U9441 ( .A1(n9200), .A2(n7808), .ZN(n7710) );
  OR2_X1 U9442 ( .A1(n10254), .A2(n7826), .ZN(n7709) );
  NAND2_X1 U9443 ( .A1(n7710), .A2(n7709), .ZN(n9205) );
  NAND2_X1 U9444 ( .A1(n9200), .A2(n7821), .ZN(n7712) );
  OR2_X1 U9445 ( .A1(n10254), .A2(n6776), .ZN(n7711) );
  NAND2_X1 U9446 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  XNOR2_X1 U9447 ( .A(n7713), .B(n7798), .ZN(n9331) );
  OAI22_X1 U9448 ( .A1(n9335), .A2(n7717), .B1(n9205), .B2(n9331), .ZN(n7714)
         );
  NOR2_X1 U9449 ( .A1(n9204), .A2(n7714), .ZN(n7722) );
  INV_X1 U9450 ( .A(n7717), .ZN(n9334) );
  NAND2_X1 U9451 ( .A1(n9331), .A2(n9205), .ZN(n7716) );
  INV_X1 U9452 ( .A(n9335), .ZN(n7715) );
  AOI21_X1 U9453 ( .B1(n9334), .B2(n7716), .A(n7715), .ZN(n7720) );
  INV_X1 U9454 ( .A(n7716), .ZN(n7718) );
  NOR2_X1 U9455 ( .A1(n7722), .A2(n7721), .ZN(n9247) );
  OAI22_X1 U9456 ( .A1(n10269), .A2(n7812), .B1(n10274), .B2(n6776), .ZN(n7723) );
  XNOR2_X1 U9457 ( .A(n7723), .B(n7798), .ZN(n7725) );
  OAI22_X1 U9458 ( .A1(n10269), .A2(n6776), .B1(n10274), .B2(n7826), .ZN(n7724) );
  NOR2_X1 U9459 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  AOI21_X1 U9460 ( .B1(n7725), .B2(n7724), .A(n7726), .ZN(n9246) );
  NAND2_X1 U9461 ( .A1(n9247), .A2(n9246), .ZN(n9245) );
  INV_X1 U9462 ( .A(n7726), .ZN(n7727) );
  NAND2_X1 U9463 ( .A1(n9245), .A2(n7727), .ZN(n9314) );
  NAND2_X1 U9464 ( .A1(n10279), .A2(n7821), .ZN(n7729) );
  OR2_X1 U9465 ( .A1(n9911), .A2(n6776), .ZN(n7728) );
  NAND2_X1 U9466 ( .A1(n7729), .A2(n7728), .ZN(n7730) );
  XNOR2_X1 U9467 ( .A(n7730), .B(n7798), .ZN(n7731) );
  INV_X1 U9468 ( .A(n9911), .ZN(n9385) );
  AOI22_X1 U9469 ( .A1(n10279), .A2(n7808), .B1(n7807), .B2(n9385), .ZN(n7732)
         );
  XNOR2_X1 U9470 ( .A(n7731), .B(n7732), .ZN(n9315) );
  INV_X1 U9471 ( .A(n7731), .ZN(n7733) );
  NAND2_X1 U9472 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  NAND2_X1 U9473 ( .A1(n9313), .A2(n7734), .ZN(n7737) );
  OAI22_X1 U9474 ( .A1(n8122), .A2(n7812), .B1(n10276), .B2(n6776), .ZN(n7735)
         );
  XOR2_X1 U9475 ( .A(n7798), .B(n7735), .Z(n7736) );
  OAI22_X1 U9476 ( .A1(n8122), .A2(n6776), .B1(n10276), .B2(n7826), .ZN(n9182)
         );
  INV_X1 U9477 ( .A(n9182), .ZN(n7738) );
  AOI22_X1 U9478 ( .A1(n9747), .A2(n7821), .B1(n4419), .B2(n9893), .ZN(n7740)
         );
  XNOR2_X1 U9479 ( .A(n7740), .B(n7798), .ZN(n7742) );
  INV_X1 U9480 ( .A(n7741), .ZN(n7744) );
  INV_X1 U9481 ( .A(n7742), .ZN(n7743) );
  OAI22_X1 U9482 ( .A1(n9905), .A2(n6776), .B1(n9912), .B2(n7826), .ZN(n9367)
         );
  NAND2_X1 U9483 ( .A1(n9725), .A2(n7821), .ZN(n7748) );
  OR2_X1 U9484 ( .A1(n9712), .A2(n6776), .ZN(n7747) );
  NAND2_X1 U9485 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  XNOR2_X1 U9486 ( .A(n7749), .B(n6924), .ZN(n7754) );
  INV_X1 U9487 ( .A(n7754), .ZN(n7752) );
  NOR2_X1 U9488 ( .A1(n9712), .A2(n7826), .ZN(n7750) );
  AOI21_X1 U9489 ( .B1(n9725), .B2(n7808), .A(n7750), .ZN(n7753) );
  INV_X1 U9490 ( .A(n7753), .ZN(n7751) );
  NAND2_X1 U9491 ( .A1(n7752), .A2(n7751), .ZN(n9264) );
  NAND2_X1 U9492 ( .A1(n9888), .A2(n7821), .ZN(n7756) );
  NAND2_X1 U9493 ( .A1(n9892), .A2(n7808), .ZN(n7755) );
  NAND2_X1 U9494 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  XNOR2_X1 U9495 ( .A(n7757), .B(n6924), .ZN(n9273) );
  AND2_X1 U9496 ( .A1(n9892), .A2(n7807), .ZN(n7758) );
  AOI21_X1 U9497 ( .B1(n9888), .B2(n4419), .A(n7758), .ZN(n7759) );
  INV_X1 U9498 ( .A(n9273), .ZN(n7760) );
  INV_X1 U9499 ( .A(n7759), .ZN(n9272) );
  OAI22_X1 U9500 ( .A1(n9874), .A2(n7812), .B1(n9662), .B2(n6776), .ZN(n7761)
         );
  XNOR2_X1 U9501 ( .A(n7761), .B(n7798), .ZN(n9217) );
  OR2_X1 U9502 ( .A1(n9874), .A2(n6776), .ZN(n7763) );
  OR2_X1 U9503 ( .A1(n9662), .A2(n7826), .ZN(n7762) );
  NAND2_X1 U9504 ( .A1(n7763), .A2(n7762), .ZN(n9215) );
  NAND2_X1 U9505 ( .A1(n9217), .A2(n9215), .ZN(n9302) );
  INV_X1 U9506 ( .A(n9302), .ZN(n7769) );
  NAND2_X1 U9507 ( .A1(n9701), .A2(n7821), .ZN(n7765) );
  OR2_X1 U9508 ( .A1(n9713), .A2(n6776), .ZN(n7764) );
  NAND2_X1 U9509 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  XNOR2_X1 U9510 ( .A(n7766), .B(n6924), .ZN(n9213) );
  NOR2_X1 U9511 ( .A1(n9713), .A2(n7826), .ZN(n7767) );
  AOI21_X1 U9512 ( .B1(n9701), .B2(n7808), .A(n7767), .ZN(n9346) );
  INV_X1 U9513 ( .A(n9217), .ZN(n7774) );
  INV_X1 U9514 ( .A(n9213), .ZN(n9212) );
  INV_X1 U9515 ( .A(n9346), .ZN(n7770) );
  OAI21_X1 U9516 ( .B1(n9212), .B2(n7770), .A(n9215), .ZN(n7773) );
  NOR3_X1 U9517 ( .A1(n9215), .A2(n9212), .A3(n7770), .ZN(n7772) );
  AOI22_X1 U9518 ( .A1(n9867), .A2(n7821), .B1(n4419), .B2(n9870), .ZN(n7771)
         );
  XOR2_X1 U9519 ( .A(n7798), .B(n7771), .Z(n7775) );
  INV_X1 U9520 ( .A(n9867), .ZN(n9666) );
  OAI22_X1 U9521 ( .A1(n9666), .A2(n6776), .B1(n9654), .B2(n7826), .ZN(n7776)
         );
  NOR2_X1 U9522 ( .A1(n7775), .A2(n7776), .ZN(n9305) );
  AOI211_X1 U9523 ( .C1(n7774), .C2(n7773), .A(n7772), .B(n9305), .ZN(n7779)
         );
  INV_X1 U9524 ( .A(n7775), .ZN(n7778) );
  INV_X1 U9525 ( .A(n7776), .ZN(n7777) );
  NOR2_X1 U9526 ( .A1(n7778), .A2(n7777), .ZN(n9304) );
  AOI22_X1 U9527 ( .A1(n9650), .A2(n7821), .B1(n4419), .B2(n9384), .ZN(n7780)
         );
  XNOR2_X1 U9528 ( .A(n7780), .B(n7798), .ZN(n7782) );
  OAI22_X1 U9529 ( .A1(n7781), .A2(n6776), .B1(n9664), .B2(n7826), .ZN(n7783)
         );
  XNOR2_X1 U9530 ( .A(n7782), .B(n7783), .ZN(n9238) );
  OAI22_X1 U9531 ( .A1(n9967), .A2(n4426), .B1(n9631), .B2(n6776), .ZN(n7786)
         );
  XNOR2_X1 U9532 ( .A(n7786), .B(n7798), .ZN(n9191) );
  OAI22_X1 U9533 ( .A1(n9967), .A2(n6776), .B1(n9631), .B2(n7826), .ZN(n7792)
         );
  OAI22_X1 U9534 ( .A1(n9636), .A2(n7812), .B1(n9841), .B2(n6776), .ZN(n7787)
         );
  XNOR2_X1 U9535 ( .A(n7787), .B(n7798), .ZN(n7791) );
  OR2_X1 U9536 ( .A1(n9841), .A2(n7826), .ZN(n7788) );
  AOI22_X1 U9537 ( .A1(n9191), .A2(n7792), .B1(n7791), .B2(n9324), .ZN(n7790)
         );
  INV_X1 U9538 ( .A(n9324), .ZN(n7794) );
  INV_X1 U9539 ( .A(n7792), .ZN(n9190) );
  AOI21_X1 U9540 ( .B1(n9189), .B2(n7794), .A(n9190), .ZN(n7793) );
  NAND3_X1 U9541 ( .A1(n9190), .A2(n9189), .A3(n7794), .ZN(n7795) );
  OAI22_X1 U9542 ( .A1(n9604), .A2(n6776), .B1(n9842), .B2(n7826), .ZN(n7800)
         );
  OAI22_X1 U9543 ( .A1(n9604), .A2(n7812), .B1(n9842), .B2(n6776), .ZN(n7799)
         );
  XNOR2_X1 U9544 ( .A(n7799), .B(n7798), .ZN(n7801) );
  XOR2_X1 U9545 ( .A(n7800), .B(n7801), .Z(n9281) );
  NAND2_X1 U9546 ( .A1(n9280), .A2(n9281), .ZN(n7803) );
  NAND2_X1 U9547 ( .A1(n9956), .A2(n7821), .ZN(n7805) );
  NAND2_X1 U9548 ( .A1(n9821), .A2(n7808), .ZN(n7804) );
  NAND2_X1 U9549 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  XNOR2_X1 U9550 ( .A(n7806), .B(n7798), .ZN(n7809) );
  AOI22_X1 U9551 ( .A1(n9956), .A2(n7808), .B1(n7807), .B2(n9821), .ZN(n7810)
         );
  XNOR2_X1 U9552 ( .A(n7809), .B(n7810), .ZN(n9256) );
  INV_X1 U9553 ( .A(n7809), .ZN(n7811) );
  AOI22_X1 U9554 ( .A1(n9255), .A2(n9256), .B1(n7811), .B2(n7810), .ZN(n9355)
         );
  OAI22_X1 U9555 ( .A1(n9824), .A2(n6776), .B1(n9576), .B2(n7826), .ZN(n7814)
         );
  OAI22_X1 U9556 ( .A1(n9824), .A2(n4426), .B1(n9576), .B2(n6776), .ZN(n7813)
         );
  XNOR2_X1 U9557 ( .A(n7813), .B(n7798), .ZN(n7815) );
  XOR2_X1 U9558 ( .A(n7814), .B(n7815), .Z(n9354) );
  NAND2_X1 U9559 ( .A1(n9355), .A2(n9354), .ZN(n9353) );
  NAND2_X1 U9560 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  NOR2_X1 U9561 ( .A1(n9527), .A2(n7826), .ZN(n7817) );
  AOI21_X1 U9562 ( .B1(n9946), .B2(n4419), .A(n7817), .ZN(n7831) );
  NAND2_X1 U9563 ( .A1(n9946), .A2(n7821), .ZN(n7819) );
  OR2_X1 U9564 ( .A1(n9527), .A2(n6776), .ZN(n7818) );
  NAND2_X1 U9565 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  XNOR2_X1 U9566 ( .A(n7820), .B(n7798), .ZN(n7830) );
  XOR2_X1 U9567 ( .A(n7831), .B(n7830), .Z(n8194) );
  NAND2_X1 U9568 ( .A1(n9814), .A2(n7821), .ZN(n7823) );
  OR2_X1 U9569 ( .A1(n9548), .A2(n6776), .ZN(n7822) );
  NAND2_X1 U9570 ( .A1(n7823), .A2(n7822), .ZN(n7824) );
  XNOR2_X1 U9571 ( .A(n7824), .B(n7798), .ZN(n7828) );
  NAND2_X1 U9572 ( .A1(n9814), .A2(n4419), .ZN(n7825) );
  OAI21_X1 U9573 ( .B1(n9548), .B2(n7826), .A(n7825), .ZN(n7827) );
  XNOR2_X1 U9574 ( .A(n7828), .B(n7827), .ZN(n7837) );
  INV_X1 U9575 ( .A(n7837), .ZN(n7829) );
  NAND2_X1 U9576 ( .A1(n7829), .A2(n9352), .ZN(n7842) );
  INV_X1 U9577 ( .A(n7830), .ZN(n7832) );
  NAND2_X1 U9578 ( .A1(n7832), .A2(n7831), .ZN(n7836) );
  NAND4_X1 U9579 ( .A1(n8196), .A2(n9352), .A3(n7837), .A4(n7836), .ZN(n7841)
         );
  INV_X1 U9580 ( .A(n7833), .ZN(n9534) );
  NAND2_X1 U9581 ( .A1(n9361), .A2(n9534), .ZN(n7835) );
  INV_X1 U9582 ( .A(n9527), .ZN(n9822) );
  AOI22_X1 U9583 ( .A1(n9357), .A2(n9822), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7834) );
  OAI211_X1 U9584 ( .C1(n9528), .C2(n9359), .A(n7835), .B(n7834), .ZN(n7839)
         );
  NOR3_X1 U9585 ( .A1(n7837), .A2(n9378), .A3(n7836), .ZN(n7838) );
  AOI211_X1 U9586 ( .C1(n9814), .C2(n9376), .A(n7839), .B(n7838), .ZN(n7840)
         );
  OAI211_X1 U9587 ( .C1(n8196), .C2(n7842), .A(n7841), .B(n7840), .ZN(P1_U3220) );
  MUX2_X1 U9588 ( .A(n8517), .B(n8779), .S(n7973), .Z(n7966) );
  INV_X1 U9589 ( .A(n8855), .ZN(n7914) );
  INV_X1 U9590 ( .A(n7843), .ZN(n7844) );
  OR2_X1 U9591 ( .A1(n7915), .A2(n7844), .ZN(n8675) );
  NOR2_X1 U9592 ( .A1(n6280), .A2(n7845), .ZN(n7854) );
  INV_X1 U9593 ( .A(n7849), .ZN(n7853) );
  INV_X1 U9594 ( .A(n5930), .ZN(n7851) );
  AOI21_X1 U9595 ( .B1(n7849), .B2(n7848), .A(n7851), .ZN(n7850) );
  NAND2_X1 U9596 ( .A1(n7866), .A2(n7855), .ZN(n7858) );
  OAI21_X1 U9597 ( .B1(n7856), .B2(n4421), .A(n7863), .ZN(n7857) );
  MUX2_X1 U9598 ( .A(n7858), .B(n7857), .S(n7977), .Z(n7860) );
  AOI21_X1 U9599 ( .B1(n7865), .B2(n7864), .A(n7872), .ZN(n7876) );
  INV_X1 U9600 ( .A(n7866), .ZN(n7869) );
  OAI211_X1 U9601 ( .C1(n7870), .C2(n7869), .A(n7868), .B(n7867), .ZN(n7875)
         );
  NOR2_X1 U9602 ( .A1(n4832), .A2(n7872), .ZN(n7874) );
  INV_X1 U9603 ( .A(n7877), .ZN(n7878) );
  AOI22_X1 U9604 ( .A1(n7879), .A2(n8007), .B1(n7973), .B2(n7878), .ZN(n7894)
         );
  NAND2_X1 U9605 ( .A1(n7881), .A2(n7880), .ZN(n7883) );
  NAND2_X1 U9606 ( .A1(n7886), .A2(n7885), .ZN(n7882) );
  MUX2_X1 U9607 ( .A(n7883), .B(n7882), .S(n7973), .Z(n7893) );
  AOI21_X1 U9608 ( .B1(n7885), .B2(n7884), .A(n7893), .ZN(n7889) );
  INV_X1 U9609 ( .A(n7886), .ZN(n7888) );
  INV_X1 U9610 ( .A(n7895), .ZN(n7887) );
  NOR3_X1 U9611 ( .A1(n7889), .A2(n7888), .A3(n7887), .ZN(n7890) );
  MUX2_X1 U9612 ( .A(n7891), .B(n7890), .S(n7977), .Z(n7892) );
  OAI21_X1 U9613 ( .B1(n7894), .B2(n7893), .A(n7892), .ZN(n7899) );
  NAND3_X1 U9614 ( .A1(n7899), .A2(n7895), .A3(n7900), .ZN(n7896) );
  NAND3_X1 U9615 ( .A1(n7899), .A2(n7898), .A3(n7897), .ZN(n7901) );
  INV_X1 U9616 ( .A(n7902), .ZN(n7903) );
  OR2_X1 U9617 ( .A1(n7904), .A2(n7903), .ZN(n8016) );
  INV_X1 U9618 ( .A(n7905), .ZN(n7908) );
  INV_X1 U9619 ( .A(n7906), .ZN(n8765) );
  NOR2_X1 U9620 ( .A1(n8765), .A2(n8688), .ZN(n7907) );
  MUX2_X1 U9621 ( .A(n7908), .B(n7907), .S(n7977), .Z(n7909) );
  MUX2_X1 U9622 ( .A(n7911), .B(n7910), .S(n7973), .Z(n7912) );
  INV_X1 U9623 ( .A(n7912), .ZN(n7913) );
  INV_X1 U9624 ( .A(n8658), .ZN(n8019) );
  INV_X1 U9625 ( .A(n7915), .ZN(n7917) );
  OAI211_X1 U9626 ( .C1(n8658), .C2(n7917), .A(n7923), .B(n7916), .ZN(n7918)
         );
  MUX2_X1 U9627 ( .A(n7919), .B(n7918), .S(n7973), .Z(n7920) );
  AOI211_X1 U9628 ( .C1(n7921), .C2(n8019), .A(n4754), .B(n7920), .ZN(n7922)
         );
  NOR2_X1 U9629 ( .A1(n7922), .A2(n8635), .ZN(n7926) );
  NAND2_X1 U9630 ( .A1(n7926), .A2(n7923), .ZN(n7928) );
  INV_X1 U9631 ( .A(n7930), .ZN(n7931) );
  OAI21_X1 U9632 ( .B1(n7932), .B2(n7931), .A(n7997), .ZN(n7942) );
  INV_X1 U9633 ( .A(n7933), .ZN(n7936) );
  NOR2_X1 U9634 ( .A1(n7934), .A2(n7936), .ZN(n7935) );
  MUX2_X1 U9635 ( .A(n7936), .B(n7935), .S(n7973), .Z(n7941) );
  NAND2_X1 U9636 ( .A1(n7997), .A2(n7937), .ZN(n7938) );
  OAI211_X1 U9637 ( .C1(n7939), .C2(n7938), .A(n8595), .B(n7998), .ZN(n7940)
         );
  AOI22_X1 U9638 ( .A1(n7942), .A2(n7977), .B1(n7941), .B2(n7940), .ZN(n7948)
         );
  AOI21_X1 U9639 ( .B1(n7945), .B2(n7943), .A(n7973), .ZN(n7947) );
  MUX2_X1 U9640 ( .A(n7945), .B(n7944), .S(n7977), .Z(n7946) );
  NAND2_X1 U9641 ( .A1(n7996), .A2(n8552), .ZN(n7952) );
  MUX2_X1 U9642 ( .A(n7952), .B(n7951), .S(n7977), .Z(n7953) );
  INV_X1 U9643 ( .A(n7995), .ZN(n7954) );
  MUX2_X1 U9644 ( .A(n7955), .B(n7954), .S(n7973), .Z(n7956) );
  MUX2_X1 U9645 ( .A(n7958), .B(n7957), .S(n7973), .Z(n7959) );
  MUX2_X1 U9646 ( .A(n4436), .B(n7960), .S(n7973), .Z(n7962) );
  INV_X1 U9647 ( .A(n7961), .ZN(n7964) );
  MUX2_X1 U9648 ( .A(n7964), .B(n7963), .S(n7973), .Z(n7965) );
  AOI21_X1 U9649 ( .B1(n4632), .B2(n7966), .A(n7967), .ZN(n7975) );
  NAND2_X1 U9650 ( .A1(n8114), .A2(n7968), .ZN(n7970) );
  OR2_X1 U9651 ( .A1(n5952), .A2(n8115), .ZN(n7969) );
  NAND2_X1 U9652 ( .A1(n8703), .A2(n7976), .ZN(n8031) );
  NAND2_X1 U9653 ( .A1(n8031), .A2(n7971), .ZN(n7986) );
  NOR2_X1 U9654 ( .A1(n7978), .A2(n7986), .ZN(n7972) );
  NAND2_X1 U9655 ( .A1(n8699), .A2(n8355), .ZN(n8033) );
  OAI211_X1 U9656 ( .C1(n7975), .C2(n8517), .A(n7972), .B(n8033), .ZN(n7984)
         );
  INV_X1 U9657 ( .A(n7976), .ZN(n8356) );
  OAI21_X1 U9658 ( .B1(n7976), .B2(n7973), .A(n8703), .ZN(n7974) );
  OAI211_X1 U9659 ( .C1(n7977), .C2(n8356), .A(n8033), .B(n7974), .ZN(n7983)
         );
  INV_X1 U9660 ( .A(n7975), .ZN(n7980) );
  OR2_X1 U9661 ( .A1(n8703), .A2(n7976), .ZN(n8030) );
  NAND3_X1 U9662 ( .A1(n8030), .A2(n7977), .A3(n7985), .ZN(n7979) );
  AOI211_X1 U9663 ( .C1(n7981), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7982)
         );
  INV_X1 U9664 ( .A(n7985), .ZN(n7989) );
  INV_X1 U9665 ( .A(n7986), .ZN(n7988) );
  OAI21_X1 U9666 ( .B1(n8355), .B2(n8703), .A(n8699), .ZN(n7987) );
  OAI211_X1 U9667 ( .C1(n7990), .C2(n7989), .A(n7988), .B(n7987), .ZN(n7993)
         );
  INV_X1 U9668 ( .A(n8030), .ZN(n7992) );
  NAND2_X1 U9669 ( .A1(n8552), .A2(n8550), .ZN(n8558) );
  AND4_X1 U9670 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(n8008)
         );
  NOR2_X1 U9671 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  NAND4_X1 U9672 ( .A1(n8008), .A2(n8007), .A3(n4427), .A4(n8006), .ZN(n8010)
         );
  NOR2_X1 U9673 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  NAND3_X1 U9674 ( .A1(n8012), .A2(n6030), .A3(n8011), .ZN(n8013) );
  NOR2_X1 U9675 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  NAND3_X1 U9676 ( .A1(n8016), .A2(n8015), .A3(n6069), .ZN(n8017) );
  NOR2_X1 U9677 ( .A1(n8675), .A2(n8017), .ZN(n8018) );
  NAND3_X1 U9678 ( .A1(n8645), .A2(n8019), .A3(n8018), .ZN(n8020) );
  NOR2_X1 U9679 ( .A1(n8635), .A2(n8020), .ZN(n8021) );
  NAND4_X1 U9680 ( .A1(n8595), .A2(n8604), .A3(n6149), .A4(n8021), .ZN(n8022)
         );
  NOR2_X1 U9681 ( .A1(n8582), .A2(n8022), .ZN(n8023) );
  NAND2_X1 U9682 ( .A1(n8568), .A2(n8023), .ZN(n8024) );
  NOR2_X1 U9683 ( .A1(n8558), .A2(n8024), .ZN(n8025) );
  NAND3_X1 U9684 ( .A1(n8533), .A2(n8553), .A3(n8025), .ZN(n8026) );
  NOR2_X1 U9685 ( .A1(n8524), .A2(n8026), .ZN(n8027) );
  NAND3_X1 U9686 ( .A1(n8515), .A2(n8506), .A3(n8027), .ZN(n8028) );
  NOR2_X1 U9687 ( .A1(n8029), .A2(n8028), .ZN(n8032) );
  NAND4_X1 U9688 ( .A1(n8033), .A2(n8032), .A3(n8031), .A4(n8030), .ZN(n8035)
         );
  NAND3_X1 U9689 ( .A1(n8041), .A2(n8040), .A3(n8489), .ZN(n8042) );
  OAI211_X1 U9690 ( .C1(n8043), .C2(n8045), .A(n8042), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8044) );
  OAI21_X1 U9691 ( .B1(n8046), .B2(n8045), .A(n8044), .ZN(P2_U3296) );
  OAI222_X1 U9692 ( .A1(n8049), .A2(P1_U3086), .B1(n8174), .B2(n8048), .C1(
        n8047), .C2(n10009), .ZN(P1_U3330) );
  AOI21_X1 U9693 ( .B1(n10191), .B2(n9932), .A(n10211), .ZN(n8057) );
  NAND4_X1 U9694 ( .A1(n10237), .A2(n8051), .A3(n8050), .A4(n10208), .ZN(n8053) );
  NAND2_X1 U9695 ( .A1(n10220), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8052) );
  OAI211_X1 U9696 ( .C1(n5462), .C2(n10205), .A(n8053), .B(n8052), .ZN(n8054)
         );
  AOI21_X1 U9697 ( .B1(n9784), .B2(n6777), .A(n8054), .ZN(n8055) );
  OAI21_X1 U9698 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(P1_U3293) );
  AOI22_X1 U9699 ( .A1(n9728), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10194), .ZN(n8058) );
  OAI21_X1 U9700 ( .B1(n10198), .B2(n8059), .A(n8058), .ZN(n8064) );
  INV_X1 U9701 ( .A(n9784), .ZN(n8061) );
  OAI22_X1 U9702 ( .A1(n8062), .A2(n10213), .B1(n8061), .B2(n8060), .ZN(n8063)
         );
  AOI211_X1 U9703 ( .C1(n8065), .C2(n6777), .A(n8064), .B(n8063), .ZN(n8068)
         );
  NAND2_X1 U9704 ( .A1(n8066), .A2(n9751), .ZN(n8067) );
  OAI211_X1 U9705 ( .C1(n8069), .C2(n9753), .A(n8068), .B(n8067), .ZN(P1_U3291) );
  XNOR2_X1 U9706 ( .A(n8855), .B(n8106), .ZN(n8073) );
  XNOR2_X1 U9707 ( .A(n8073), .B(n8686), .ZN(n8216) );
  XNOR2_X1 U9708 ( .A(n8848), .B(n8106), .ZN(n8075) );
  XNOR2_X1 U9709 ( .A(n8075), .B(n8357), .ZN(n8350) );
  INV_X1 U9710 ( .A(n8075), .ZN(n8076) );
  XNOR2_X1 U9711 ( .A(n8842), .B(n8106), .ZN(n8263) );
  XNOR2_X1 U9712 ( .A(n8631), .B(n6746), .ZN(n8077) );
  NAND2_X1 U9713 ( .A1(n8077), .A2(n8647), .ZN(n8271) );
  NOR2_X1 U9714 ( .A1(n8077), .A2(n8647), .ZN(n8273) );
  XNOR2_X1 U9715 ( .A(n8737), .B(n8106), .ZN(n8078) );
  XOR2_X1 U9716 ( .A(n8637), .B(n8078), .Z(n8323) );
  INV_X1 U9717 ( .A(n8078), .ZN(n8079) );
  XNOR2_X1 U9718 ( .A(n8829), .B(n8106), .ZN(n8080) );
  XOR2_X1 U9719 ( .A(n8615), .B(n8080), .Z(n8231) );
  INV_X1 U9720 ( .A(n8080), .ZN(n8081) );
  XNOR2_X1 U9721 ( .A(n8596), .B(n8106), .ZN(n8082) );
  XOR2_X1 U9722 ( .A(n8579), .B(n8082), .Z(n8297) );
  XNOR2_X1 U9723 ( .A(n8251), .B(n8106), .ZN(n8084) );
  XOR2_X1 U9724 ( .A(n8589), .B(n8084), .Z(n8247) );
  INV_X1 U9725 ( .A(n8084), .ZN(n8086) );
  NAND2_X1 U9726 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  XNOR2_X1 U9727 ( .A(n8815), .B(n8106), .ZN(n8090) );
  XNOR2_X1 U9728 ( .A(n8090), .B(n8560), .ZN(n8303) );
  INV_X1 U9729 ( .A(n8303), .ZN(n8088) );
  XOR2_X1 U9730 ( .A(n8106), .B(n8803), .Z(n8286) );
  XNOR2_X1 U9731 ( .A(n8809), .B(n6746), .ZN(n8093) );
  OAI22_X1 U9732 ( .A1(n8286), .A2(n8285), .B1(n8307), .B2(n8093), .ZN(n8089)
         );
  INV_X1 U9733 ( .A(n8089), .ZN(n8091) );
  NAND2_X1 U9734 ( .A1(n8090), .A2(n8560), .ZN(n8224) );
  AND2_X1 U9735 ( .A1(n8091), .A2(n8224), .ZN(n8092) );
  NAND2_X1 U9736 ( .A1(n8223), .A2(n8092), .ZN(n8097) );
  OAI21_X1 U9737 ( .B1(n8283), .B2(n8570), .A(n8561), .ZN(n8095) );
  NOR3_X1 U9738 ( .A1(n8283), .A2(n8570), .A3(n8561), .ZN(n8094) );
  AOI21_X1 U9739 ( .B1(n8286), .B2(n8095), .A(n8094), .ZN(n8096) );
  NAND2_X1 U9740 ( .A1(n8097), .A2(n8096), .ZN(n8254) );
  XNOR2_X1 U9741 ( .A(n8797), .B(n8106), .ZN(n8098) );
  XOR2_X1 U9742 ( .A(n8545), .B(n8098), .Z(n8255) );
  NAND2_X1 U9743 ( .A1(n8254), .A2(n8255), .ZN(n8100) );
  XNOR2_X1 U9744 ( .A(n8791), .B(n8106), .ZN(n8102) );
  XNOR2_X1 U9745 ( .A(n8101), .B(n8102), .ZN(n8330) );
  INV_X1 U9746 ( .A(n8101), .ZN(n8103) );
  XNOR2_X1 U9747 ( .A(n8785), .B(n8106), .ZN(n8104) );
  NAND2_X1 U9748 ( .A1(n8104), .A2(n8526), .ZN(n8105) );
  OAI21_X1 U9749 ( .B1(n8104), .B2(n8526), .A(n8105), .ZN(n8206) );
  XOR2_X1 U9750 ( .A(n8106), .B(n8506), .Z(n8107) );
  XNOR2_X1 U9751 ( .A(n8108), .B(n8107), .ZN(n8113) );
  NAND2_X1 U9752 ( .A1(n8508), .A2(n8344), .ZN(n8110) );
  AOI22_X1 U9753 ( .A1(n8511), .A2(n8332), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8109) );
  OAI211_X1 U9754 ( .C1(n8336), .C2(n8342), .A(n8110), .B(n8109), .ZN(n8111)
         );
  AOI21_X1 U9755 ( .B1(n8779), .B2(n8353), .A(n8111), .ZN(n8112) );
  OAI21_X1 U9756 ( .B1(n8113), .B2(n8348), .A(n8112), .ZN(P2_U3160) );
  INV_X1 U9757 ( .A(n8114), .ZN(n8173) );
  OAI222_X1 U9758 ( .A1(n8878), .A2(n8115), .B1(n8874), .B2(n8173), .C1(
        P2_U3151), .C2(n5904), .ZN(P2_U3265) );
  INV_X1 U9759 ( .A(n8116), .ZN(n8880) );
  OAI222_X1 U9760 ( .A1(n8117), .A2(P1_U3086), .B1(n8174), .B2(n8880), .C1(
        n9074), .C2(n10018), .ZN(P1_U3329) );
  INV_X1 U9761 ( .A(n9712), .ZN(n9901) );
  NAND2_X1 U9762 ( .A1(n10257), .A2(n8119), .ZN(n8120) );
  OAI22_X1 U9763 ( .A1(n9775), .A2(n9774), .B1(n10279), .B2(n9385), .ZN(n9757)
         );
  NOR2_X1 U9764 ( .A1(n9905), .A2(n9912), .ZN(n8123) );
  OAI22_X1 U9765 ( .A1(n9735), .A2(n8123), .B1(n9893), .B2(n9747), .ZN(n9720)
         );
  NAND2_X1 U9766 ( .A1(n9888), .A2(n9892), .ZN(n8124) );
  NAND2_X1 U9767 ( .A1(n9874), .A2(n9662), .ZN(n8127) );
  NOR2_X1 U9768 ( .A1(n9874), .A2(n9662), .ZN(n8126) );
  NAND2_X1 U9769 ( .A1(n9867), .A2(n9870), .ZN(n8129) );
  NOR2_X1 U9770 ( .A1(n9867), .A2(n9870), .ZN(n8128) );
  NAND2_X1 U9771 ( .A1(n7781), .A2(n9664), .ZN(n9588) );
  NAND2_X1 U9772 ( .A1(n9636), .A2(n9841), .ZN(n9610) );
  NAND2_X1 U9773 ( .A1(n9967), .A2(n9631), .ZN(n8130) );
  AND2_X1 U9774 ( .A1(n9588), .A2(n8132), .ZN(n8131) );
  INV_X1 U9775 ( .A(n8132), .ZN(n8136) );
  NAND2_X1 U9776 ( .A1(n9650), .A2(n9384), .ZN(n9625) );
  NAND2_X1 U9777 ( .A1(n9854), .A2(n9857), .ZN(n8133) );
  INV_X1 U9778 ( .A(n9591), .ZN(n8134) );
  AND2_X1 U9779 ( .A1(n9589), .A2(n8134), .ZN(n8135) );
  INV_X1 U9780 ( .A(n8138), .ZN(n8139) );
  NOR2_X1 U9781 ( .A1(n9956), .A2(n9821), .ZN(n8141) );
  NAND2_X1 U9782 ( .A1(n9575), .A2(n9821), .ZN(n8140) );
  NOR2_X1 U9783 ( .A1(n9824), .A2(n9576), .ZN(n8143) );
  NAND2_X1 U9784 ( .A1(n9824), .A2(n9576), .ZN(n8142) );
  NAND2_X1 U9785 ( .A1(n8144), .A2(n9527), .ZN(n8145) );
  INV_X1 U9786 ( .A(n9814), .ZN(n9536) );
  AND2_X1 U9787 ( .A1(n10296), .A2(n10285), .ZN(n9816) );
  NAND2_X1 U9788 ( .A1(n8186), .A2(n9816), .ZN(n8171) );
  INV_X1 U9789 ( .A(n9661), .ZN(n8149) );
  INV_X1 U9790 ( .A(n9648), .ZN(n8150) );
  NOR2_X1 U9791 ( .A1(n9867), .A2(n9654), .ZN(n9645) );
  NOR2_X1 U9792 ( .A1(n9613), .A2(n8152), .ZN(n8153) );
  NAND2_X2 U9793 ( .A1(n9574), .A2(n9575), .ZN(n9573) );
  INV_X1 U9794 ( .A(n8156), .ZN(n9558) );
  NOR2_X1 U9795 ( .A1(n9557), .A2(n9558), .ZN(n8157) );
  NAND2_X1 U9796 ( .A1(n9550), .A2(n8160), .ZN(n9522) );
  NAND2_X1 U9797 ( .A1(n9522), .A2(n9532), .ZN(n9526) );
  NAND2_X1 U9798 ( .A1(n9526), .A2(n8161), .ZN(n8163) );
  XNOR2_X1 U9799 ( .A(n8163), .B(n4714), .ZN(n8167) );
  AOI22_X1 U9800 ( .A1(n9929), .A2(n8146), .B1(n9381), .B2(n8164), .ZN(n8165)
         );
  AOI21_X2 U9801 ( .B1(n8167), .B2(n9927), .A(n8166), .ZN(n8180) );
  INV_X1 U9802 ( .A(n8188), .ZN(n8179) );
  OAI211_X1 U9803 ( .C1(n8179), .C2(n4606), .A(n9932), .B(n9515), .ZN(n8175)
         );
  NAND2_X1 U9804 ( .A1(n8180), .A2(n8175), .ZN(n8187) );
  NAND2_X1 U9805 ( .A1(n8171), .A2(n8170), .ZN(P1_U3551) );
  OAI222_X1 U9806 ( .A1(n5376), .A2(P1_U3086), .B1(n8174), .B2(n8173), .C1(
        n8172), .C2(n10009), .ZN(P1_U3325) );
  NAND2_X1 U9807 ( .A1(n8186), .A2(n10216), .ZN(n8185) );
  INV_X1 U9808 ( .A(n8175), .ZN(n8183) );
  INV_X1 U9809 ( .A(n8176), .ZN(n8177) );
  AOI22_X1 U9810 ( .A1(n10220), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8177), .B2(
        n10194), .ZN(n8178) );
  OAI21_X1 U9811 ( .B1(n8179), .B2(n10198), .A(n8178), .ZN(n8182) );
  NOR2_X1 U9812 ( .A1(n8180), .A2(n10220), .ZN(n8181) );
  NAND2_X1 U9813 ( .A1(n8185), .A2(n8184), .ZN(P1_U3356) );
  AND2_X1 U9814 ( .A1(n10289), .A2(n10285), .ZN(n9943) );
  NAND2_X1 U9815 ( .A1(n8186), .A2(n9943), .ZN(n8191) );
  NAND2_X1 U9816 ( .A1(n8191), .A2(n8190), .ZN(P1_U3519) );
  INV_X1 U9817 ( .A(n8192), .ZN(n8870) );
  OAI222_X1 U9818 ( .A1(n10018), .A2(n8193), .B1(P1_U3086), .B2(n5377), .C1(
        n8870), .C2(n8174), .ZN(P1_U3326) );
  NAND2_X1 U9819 ( .A1(n8195), .A2(n8194), .ZN(n8197) );
  INV_X1 U9820 ( .A(n8198), .ZN(n9544) );
  NOR2_X1 U9821 ( .A1(n9359), .A2(n9548), .ZN(n8201) );
  OAI22_X1 U9822 ( .A1(n9370), .A2(n9576), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8199), .ZN(n8200) );
  AOI211_X1 U9823 ( .C1(n9544), .C2(n9361), .A(n8201), .B(n8200), .ZN(n8203)
         );
  NAND2_X1 U9824 ( .A1(n9946), .A2(n9376), .ZN(n8202) );
  OAI211_X1 U9825 ( .C1(n8204), .C2(n9378), .A(n8203), .B(n8202), .ZN(P1_U3214) );
  AOI21_X1 U9826 ( .B1(n8205), .B2(n8206), .A(n8348), .ZN(n8208) );
  NAND2_X1 U9827 ( .A1(n8208), .A2(n8207), .ZN(n8213) );
  INV_X1 U9828 ( .A(n8520), .ZN(n8210) );
  AOI22_X1 U9829 ( .A1(n8535), .A2(n8331), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8209) );
  OAI21_X1 U9830 ( .B1(n8210), .B2(n8346), .A(n8209), .ZN(n8211) );
  AOI21_X1 U9831 ( .B1(n8344), .B2(n8517), .A(n8211), .ZN(n8212) );
  OAI211_X1 U9832 ( .C1(n8214), .C2(n8311), .A(n8213), .B(n8212), .ZN(P2_U3154) );
  XOR2_X1 U9833 ( .A(n8216), .B(n8215), .Z(n8222) );
  OAI21_X1 U9834 ( .B1(n8335), .B2(n8672), .A(n8217), .ZN(n8218) );
  AOI21_X1 U9835 ( .B1(n8331), .B2(n8358), .A(n8218), .ZN(n8219) );
  OAI21_X1 U9836 ( .B1(n8676), .B2(n8346), .A(n8219), .ZN(n8220) );
  AOI21_X1 U9837 ( .B1(n8855), .B2(n8353), .A(n8220), .ZN(n8221) );
  OAI21_X1 U9838 ( .B1(n8222), .B2(n8348), .A(n8221), .ZN(P2_U3155) );
  NAND2_X1 U9839 ( .A1(n8223), .A2(n8224), .ZN(n8282) );
  XNOR2_X1 U9840 ( .A(n8282), .B(n8283), .ZN(n8284) );
  XNOR2_X1 U9841 ( .A(n8284), .B(n8307), .ZN(n8229) );
  AOI22_X1 U9842 ( .A1(n8331), .A2(n8560), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8226) );
  NAND2_X1 U9843 ( .A1(n8332), .A2(n8564), .ZN(n8225) );
  OAI211_X1 U9844 ( .C1(n8285), .C2(n8335), .A(n8226), .B(n8225), .ZN(n8227)
         );
  AOI21_X1 U9845 ( .B1(n8809), .B2(n8353), .A(n8227), .ZN(n8228) );
  OAI21_X1 U9846 ( .B1(n8229), .B2(n8348), .A(n8228), .ZN(P2_U3156) );
  INV_X1 U9847 ( .A(n8829), .ZN(n8238) );
  OAI211_X1 U9848 ( .C1(n8232), .C2(n8231), .A(n8230), .B(n8315), .ZN(n8237)
         );
  NAND2_X1 U9849 ( .A1(n8344), .A2(n8605), .ZN(n8233) );
  NAND2_X1 U9850 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8483) );
  OAI211_X1 U9851 ( .C1(n8234), .C2(n8342), .A(n8233), .B(n8483), .ZN(n8235)
         );
  AOI21_X1 U9852 ( .B1(n8608), .B2(n8332), .A(n8235), .ZN(n8236) );
  OAI211_X1 U9853 ( .C1(n8238), .C2(n8311), .A(n8237), .B(n8236), .ZN(P2_U3159) );
  XNOR2_X1 U9854 ( .A(n8240), .B(n8239), .ZN(n8241) );
  NAND2_X1 U9855 ( .A1(n8241), .A2(n8315), .ZN(n8245) );
  AOI22_X1 U9856 ( .A1(n8331), .A2(n6690), .B1(n8353), .B2(n8767), .ZN(n8244)
         );
  NAND2_X1 U9857 ( .A1(n8317), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U9858 ( .A1(n8344), .A2(n8366), .ZN(n8242) );
  NAND4_X1 U9859 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(
        P2_U3162) );
  XOR2_X1 U9860 ( .A(n8246), .B(n8247), .Z(n8253) );
  AOI22_X1 U9861 ( .A1(n8344), .A2(n8560), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8249) );
  NAND2_X1 U9862 ( .A1(n8332), .A2(n8580), .ZN(n8248) );
  OAI211_X1 U9863 ( .C1(n8579), .C2(n8342), .A(n8249), .B(n8248), .ZN(n8250)
         );
  AOI21_X1 U9864 ( .B1(n8251), .B2(n8353), .A(n8250), .ZN(n8252) );
  OAI21_X1 U9865 ( .B1(n8253), .B2(n8348), .A(n8252), .ZN(P2_U3163) );
  XOR2_X1 U9866 ( .A(n8255), .B(n8254), .Z(n8261) );
  AOI22_X1 U9867 ( .A1(n8561), .A2(n8331), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8257) );
  NAND2_X1 U9868 ( .A1(n8537), .A2(n8332), .ZN(n8256) );
  OAI211_X1 U9869 ( .C1(n8258), .C2(n8335), .A(n8257), .B(n8256), .ZN(n8259)
         );
  AOI21_X1 U9870 ( .B1(n8797), .B2(n8353), .A(n8259), .ZN(n8260) );
  OAI21_X1 U9871 ( .B1(n8261), .B2(n8348), .A(n8260), .ZN(P2_U3165) );
  XNOR2_X1 U9872 ( .A(n8263), .B(n8659), .ZN(n8264) );
  XNOR2_X1 U9873 ( .A(n8265), .B(n8264), .ZN(n8270) );
  OR2_X1 U9874 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6112), .ZN(n8405) );
  OAI21_X1 U9875 ( .B1(n8342), .B2(n8672), .A(n8405), .ZN(n8266) );
  AOI21_X1 U9876 ( .B1(n8344), .B2(n8616), .A(n8266), .ZN(n8267) );
  OAI21_X1 U9877 ( .B1(n8652), .B2(n8346), .A(n8267), .ZN(n8268) );
  AOI21_X1 U9878 ( .B1(n8842), .B2(n8353), .A(n8268), .ZN(n8269) );
  OAI21_X1 U9879 ( .B1(n8270), .B2(n8348), .A(n8269), .ZN(P2_U3166) );
  INV_X1 U9880 ( .A(n8271), .ZN(n8272) );
  NOR2_X1 U9881 ( .A1(n8273), .A2(n8272), .ZN(n8274) );
  XNOR2_X1 U9882 ( .A(n8275), .B(n8274), .ZN(n8281) );
  NAND2_X1 U9883 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8427) );
  OAI21_X1 U9884 ( .B1(n8342), .B2(n8276), .A(n8427), .ZN(n8277) );
  AOI21_X1 U9885 ( .B1(n8344), .B2(n8637), .A(n8277), .ZN(n8278) );
  OAI21_X1 U9886 ( .B1(n8632), .B2(n8346), .A(n8278), .ZN(n8279) );
  AOI21_X1 U9887 ( .B1(n8631), .B2(n8353), .A(n8279), .ZN(n8280) );
  OAI21_X1 U9888 ( .B1(n8281), .B2(n8348), .A(n8280), .ZN(P2_U3168) );
  OAI22_X1 U9889 ( .A1(n8284), .A2(n8570), .B1(n8283), .B2(n8282), .ZN(n8288)
         );
  XNOR2_X1 U9890 ( .A(n8286), .B(n8285), .ZN(n8287) );
  XNOR2_X1 U9891 ( .A(n8288), .B(n8287), .ZN(n8293) );
  AOI22_X1 U9892 ( .A1(n8545), .A2(n8344), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8290) );
  NAND2_X1 U9893 ( .A1(n8548), .A2(n8332), .ZN(n8289) );
  OAI211_X1 U9894 ( .C1(n8307), .C2(n8342), .A(n8290), .B(n8289), .ZN(n8291)
         );
  AOI21_X1 U9895 ( .B1(n8803), .B2(n8353), .A(n8291), .ZN(n8292) );
  OAI21_X1 U9896 ( .B1(n8293), .B2(n8348), .A(n8292), .ZN(P2_U3169) );
  INV_X1 U9897 ( .A(n8295), .ZN(n8296) );
  AOI21_X1 U9898 ( .B1(n8297), .B2(n8294), .A(n8296), .ZN(n8302) );
  AOI22_X1 U9899 ( .A1(n8344), .A2(n8589), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8299) );
  NAND2_X1 U9900 ( .A1(n8332), .A2(n8597), .ZN(n8298) );
  OAI211_X1 U9901 ( .C1(n8591), .C2(n8342), .A(n8299), .B(n8298), .ZN(n8300)
         );
  AOI21_X1 U9902 ( .B1(n8596), .B2(n8353), .A(n8300), .ZN(n8301) );
  OAI21_X1 U9903 ( .B1(n8302), .B2(n8348), .A(n8301), .ZN(P2_U3173) );
  INV_X1 U9904 ( .A(n8815), .ZN(n8312) );
  AOI21_X1 U9905 ( .B1(n8304), .B2(n8303), .A(n8348), .ZN(n8305) );
  NAND2_X1 U9906 ( .A1(n8305), .A2(n8223), .ZN(n8310) );
  AOI22_X1 U9907 ( .A1(n8331), .A2(n8589), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8306) );
  OAI21_X1 U9908 ( .B1(n8307), .B2(n8335), .A(n8306), .ZN(n8308) );
  AOI21_X1 U9909 ( .B1(n8573), .B2(n8332), .A(n8308), .ZN(n8309) );
  OAI211_X1 U9910 ( .C1(n8312), .C2(n8311), .A(n8310), .B(n8309), .ZN(P2_U3175) );
  XNOR2_X1 U9911 ( .A(n8313), .B(n8314), .ZN(n8316) );
  NAND2_X1 U9912 ( .A1(n8316), .A2(n8315), .ZN(n8321) );
  AOI22_X1 U9913 ( .A1(n8331), .A2(n8367), .B1(n8353), .B2(n4421), .ZN(n8320)
         );
  NAND2_X1 U9914 ( .A1(n8317), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U9915 ( .A1(n8344), .A2(n8365), .ZN(n8318) );
  NAND4_X1 U9916 ( .A1(n8321), .A2(n8320), .A3(n8319), .A4(n8318), .ZN(
        P2_U3177) );
  XOR2_X1 U9917 ( .A(n8322), .B(n8323), .Z(n8329) );
  NAND2_X1 U9918 ( .A1(n8344), .A2(n8615), .ZN(n8325) );
  NAND2_X1 U9919 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8439) );
  OAI211_X1 U9920 ( .C1(n8647), .C2(n8342), .A(n8325), .B(n8439), .ZN(n8326)
         );
  AOI21_X1 U9921 ( .B1(n8619), .B2(n8332), .A(n8326), .ZN(n8328) );
  NAND2_X1 U9922 ( .A1(n8737), .A2(n8353), .ZN(n8327) );
  OAI211_X1 U9923 ( .C1(n8329), .C2(n8348), .A(n8328), .B(n8327), .ZN(P2_U3178) );
  XNOR2_X1 U9924 ( .A(n8330), .B(n8535), .ZN(n8339) );
  AOI22_X1 U9925 ( .A1(n8545), .A2(n8331), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8334) );
  NAND2_X1 U9926 ( .A1(n8529), .A2(n8332), .ZN(n8333) );
  OAI211_X1 U9927 ( .C1(n8336), .C2(n8335), .A(n8334), .B(n8333), .ZN(n8337)
         );
  AOI21_X1 U9928 ( .B1(n8791), .B2(n8353), .A(n8337), .ZN(n8338) );
  OAI21_X1 U9929 ( .B1(n8339), .B2(n8348), .A(n8338), .ZN(P2_U3180) );
  NOR2_X1 U9930 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8340), .ZN(n8385) );
  NOR2_X1 U9931 ( .A1(n8342), .A2(n8341), .ZN(n8343) );
  AOI211_X1 U9932 ( .C1(n8344), .C2(n8659), .A(n8385), .B(n8343), .ZN(n8345)
         );
  OAI21_X1 U9933 ( .B1(n8662), .B2(n8346), .A(n8345), .ZN(n8352) );
  AOI211_X1 U9934 ( .C1(n8350), .C2(n8349), .A(n8348), .B(n8347), .ZN(n8351)
         );
  AOI211_X1 U9935 ( .C1(n8848), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8354)
         );
  INV_X1 U9936 ( .A(n8354), .ZN(P2_U3181) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8355), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9938 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8356), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8508), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8517), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8526), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8535), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8545), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8561), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8570), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8560), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9947 ( .A(n8589), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8368), .Z(
        P2_U3512) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9949 ( .A(n8615), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8368), .Z(
        P2_U3510) );
  MUX2_X1 U9950 ( .A(n8637), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8368), .Z(
        P2_U3509) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8616), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9952 ( .A(n8659), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8368), .Z(
        P2_U3507) );
  MUX2_X1 U9953 ( .A(n8357), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8368), .Z(
        P2_U3506) );
  MUX2_X1 U9954 ( .A(n8686), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8368), .Z(
        P2_U3505) );
  MUX2_X1 U9955 ( .A(n8358), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8368), .Z(
        P2_U3504) );
  MUX2_X1 U9956 ( .A(n8688), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8368), .Z(
        P2_U3503) );
  MUX2_X1 U9957 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8359), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9958 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8360), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8361), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8362), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9961 ( .A(n8363), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8368), .Z(
        P2_U3497) );
  MUX2_X1 U9962 ( .A(n8364), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8368), .Z(
        P2_U3496) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8365), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9964 ( .A(n8366), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8368), .Z(
        P2_U3493) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8367), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9966 ( .A(n6690), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8368), .Z(
        P2_U3491) );
  AOI21_X1 U9967 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8371), .A(n8369), .ZN(
        n8392) );
  XNOR2_X1 U9968 ( .A(n8393), .B(n8392), .ZN(n8370) );
  AOI21_X1 U9969 ( .B1(n8661), .B2(n8370), .A(n8394), .ZN(n8391) );
  NAND2_X1 U9970 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9971 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8374), .ZN(n8401) );
  OAI21_X1 U9972 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8374), .A(n8401), .ZN(
        n8389) );
  INV_X1 U9973 ( .A(n8375), .ZN(n8380) );
  MUX2_X1 U9974 ( .A(n8661), .B(n9107), .S(n8489), .Z(n8376) );
  NAND2_X1 U9975 ( .A1(n8376), .A2(n8393), .ZN(n8412) );
  INV_X1 U9976 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U9977 ( .A1(n8377), .A2(n8400), .ZN(n8378) );
  AND2_X1 U9978 ( .A1(n8412), .A2(n8378), .ZN(n8379) );
  OAI21_X1 U9979 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8413) );
  INV_X1 U9980 ( .A(n8413), .ZN(n8384) );
  NOR3_X1 U9981 ( .A1(n8381), .A2(n8380), .A3(n8379), .ZN(n8383) );
  OAI21_X1 U9982 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8387) );
  AOI21_X1 U9983 ( .B1(n8482), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8385), .ZN(
        n8386) );
  OAI211_X1 U9984 ( .C1(n8486), .C2(n8400), .A(n8387), .B(n8386), .ZN(n8388)
         );
  AOI21_X1 U9985 ( .B1(n8499), .B2(n8389), .A(n8388), .ZN(n8390) );
  OAI21_X1 U9986 ( .B1(n8391), .B2(n8501), .A(n8390), .ZN(P2_U3197) );
  NOR2_X1 U9987 ( .A1(n8393), .A2(n8392), .ZN(n8395) );
  NOR2_X1 U9988 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  NAND2_X1 U9989 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8422), .ZN(n8396) );
  OAI21_X1 U9990 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8422), .A(n8396), .ZN(
        n8397) );
  NOR2_X1 U9991 ( .A1(n8398), .A2(n8397), .ZN(n8421) );
  AOI21_X1 U9992 ( .B1(n8398), .B2(n8397), .A(n8421), .ZN(n8420) );
  AOI22_X1 U9993 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8422), .B1(n8425), .B2(
        n8745), .ZN(n8404) );
  NAND2_X1 U9994 ( .A1(n8400), .A2(n8399), .ZN(n8402) );
  NAND2_X1 U9995 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  NAND2_X1 U9996 ( .A1(n8404), .A2(n8403), .ZN(n8424) );
  OAI21_X1 U9997 ( .B1(n8404), .B2(n8403), .A(n8424), .ZN(n8418) );
  INV_X1 U9998 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U9999 ( .A1(n8450), .A2(n8425), .ZN(n8406) );
  OAI211_X1 U10000 ( .C1(n8407), .C2(n8441), .A(n8406), .B(n8405), .ZN(n8417)
         );
  MUX2_X1 U10001 ( .A(n8651), .B(n8745), .S(n8489), .Z(n8408) );
  NAND2_X1 U10002 ( .A1(n8408), .A2(n8425), .ZN(n8429) );
  INV_X1 U10003 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U10004 ( .A1(n8409), .A2(n8422), .ZN(n8410) );
  NAND2_X1 U10005 ( .A1(n8429), .A2(n8410), .ZN(n8411) );
  AOI21_X1 U10006 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8432) );
  INV_X1 U10007 ( .A(n8432), .ZN(n8415) );
  NAND3_X1 U10008 ( .A1(n8413), .A2(n8412), .A3(n8411), .ZN(n8414) );
  AOI21_X1 U10009 ( .B1(n8415), .B2(n8414), .A(n8494), .ZN(n8416) );
  AOI211_X1 U10010 ( .C1(n8418), .C2(n8499), .A(n8417), .B(n8416), .ZN(n8419)
         );
  OAI21_X1 U10011 ( .B1(n8420), .B2(n8501), .A(n8419), .ZN(P2_U3198) );
  AOI21_X1 U10012 ( .B1(n9059), .B2(n8423), .A(n8451), .ZN(n8438) );
  OAI21_X1 U10013 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8426), .A(n8465), .ZN(
        n8436) );
  NAND2_X1 U10014 ( .A1(n8450), .A2(n8452), .ZN(n8428) );
  OAI211_X1 U10015 ( .C1(n9148), .C2(n8441), .A(n8428), .B(n8427), .ZN(n8435)
         );
  INV_X1 U10016 ( .A(n8429), .ZN(n8431) );
  MUX2_X1 U10017 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8489), .Z(n8443) );
  XNOR2_X1 U10018 ( .A(n8443), .B(n8452), .ZN(n8430) );
  OAI21_X1 U10019 ( .B1(n8432), .B2(n8431), .A(n8430), .ZN(n8442) );
  OR3_X1 U10020 ( .A1(n8432), .A2(n8431), .A3(n8430), .ZN(n8433) );
  AOI21_X1 U10021 ( .B1(n8442), .B2(n8433), .A(n8494), .ZN(n8434) );
  AOI211_X1 U10022 ( .C1(n8436), .C2(n8499), .A(n8435), .B(n8434), .ZN(n8437)
         );
  OAI21_X1 U10023 ( .B1(n8438), .B2(n8501), .A(n8437), .ZN(P2_U3199) );
  INV_X1 U10024 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8440) );
  OAI21_X1 U10025 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8449) );
  OAI21_X1 U10026 ( .B1(n8443), .B2(n8460), .A(n8442), .ZN(n8444) );
  MUX2_X1 U10027 ( .A(n8621), .B(n8462), .S(n8489), .Z(n8445) );
  NAND2_X1 U10028 ( .A1(n8444), .A2(n8445), .ZN(n8488) );
  INV_X1 U10029 ( .A(n8444), .ZN(n8447) );
  INV_X1 U10030 ( .A(n8445), .ZN(n8446) );
  NAND2_X1 U10031 ( .A1(n8447), .A2(n8446), .ZN(n8468) );
  AOI211_X1 U10032 ( .C1(n8488), .C2(n8468), .A(n8467), .B(n8494), .ZN(n8448)
         );
  AOI211_X1 U10033 ( .C1(n8450), .C2(n8467), .A(n8449), .B(n8448), .ZN(n8473)
         );
  OR2_X1 U10034 ( .A1(n8453), .A2(n8452), .ZN(n8456) );
  OR2_X1 U10035 ( .A1(n8467), .A2(n8621), .ZN(n8474) );
  NAND2_X1 U10036 ( .A1(n8467), .A2(n8621), .ZN(n8454) );
  NAND2_X1 U10037 ( .A1(n8474), .A2(n8454), .ZN(n8455) );
  AND3_X1 U10038 ( .A1(n8457), .A2(n8456), .A3(n8455), .ZN(n8459) );
  OAI21_X1 U10039 ( .B1(n8476), .B2(n8459), .A(n8458), .ZN(n8472) );
  NAND2_X1 U10040 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  XNOR2_X1 U10041 ( .A(n8467), .B(n8462), .ZN(n8464) );
  AND3_X1 U10042 ( .A1(n8465), .A2(n8464), .A3(n8463), .ZN(n8466) );
  OAI21_X1 U10043 ( .B1(n8479), .B2(n8466), .A(n8499), .ZN(n8471) );
  NAND2_X1 U10044 ( .A1(n8468), .A2(n8467), .ZN(n8487) );
  INV_X1 U10045 ( .A(n8487), .ZN(n8469) );
  NAND3_X1 U10046 ( .A1(n8488), .A2(P2_U3893), .A3(n8469), .ZN(n8470) );
  NAND4_X1 U10047 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(
        P2_U3200) );
  INV_X1 U10048 ( .A(n8474), .ZN(n8475) );
  NOR2_X1 U10049 ( .A1(n8476), .A2(n8475), .ZN(n8478) );
  XNOR2_X1 U10050 ( .A(n8485), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8491) );
  INV_X1 U10051 ( .A(n8491), .ZN(n8477) );
  XNOR2_X1 U10052 ( .A(n8478), .B(n8477), .ZN(n8502) );
  AOI21_X1 U10053 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8480), .A(n8479), .ZN(
        n8481) );
  XNOR2_X1 U10054 ( .A(n8485), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8490) );
  XNOR2_X1 U10055 ( .A(n8481), .B(n8490), .ZN(n8498) );
  NAND2_X1 U10056 ( .A1(n8482), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8484) );
  OAI211_X1 U10057 ( .C1(n8486), .C2(n8485), .A(n8484), .B(n8483), .ZN(n8497)
         );
  NAND2_X1 U10058 ( .A1(n8488), .A2(n8487), .ZN(n8493) );
  MUX2_X1 U10059 ( .A(n8491), .B(n8490), .S(n8489), .Z(n8492) );
  XNOR2_X1 U10060 ( .A(n8493), .B(n8492), .ZN(n8495) );
  NOR2_X1 U10061 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  AOI211_X1 U10062 ( .C1(n8499), .C2(n8498), .A(n8497), .B(n8496), .ZN(n8500)
         );
  OAI21_X1 U10063 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(P2_U3201) );
  INV_X1 U10064 ( .A(n8703), .ZN(n8776) );
  AOI21_X1 U10065 ( .B1(n10320), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8503), .ZN(
        n8504) );
  OAI21_X1 U10066 ( .B1(n8776), .B2(n8633), .A(n8504), .ZN(P2_U3203) );
  INV_X1 U10067 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8510) );
  XNOR2_X1 U10068 ( .A(n8507), .B(n8506), .ZN(n8509) );
  AOI222_X1 U10069 ( .A1(n8690), .A2(n8509), .B1(n8508), .B2(n8685), .C1(n8526), .C2(n8687), .ZN(n8777) );
  MUX2_X1 U10070 ( .A(n8510), .B(n8777), .S(n8678), .Z(n8513) );
  AOI22_X1 U10071 ( .A1(n8779), .A2(n10307), .B1(n10311), .B2(n8511), .ZN(
        n8512) );
  OAI211_X1 U10072 ( .C1(n8782), .C2(n8666), .A(n8513), .B(n8512), .ZN(
        P2_U3205) );
  XNOR2_X1 U10073 ( .A(n8514), .B(n8515), .ZN(n8788) );
  INV_X1 U10074 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8519) );
  XNOR2_X1 U10075 ( .A(n8516), .B(n8515), .ZN(n8518) );
  AOI222_X1 U10076 ( .A1(n8690), .A2(n8518), .B1(n8517), .B2(n8685), .C1(n8535), .C2(n8687), .ZN(n8783) );
  MUX2_X1 U10077 ( .A(n8519), .B(n8783), .S(n8678), .Z(n8522) );
  AOI22_X1 U10078 ( .A1(n8785), .A2(n10307), .B1(n10311), .B2(n8520), .ZN(
        n8521) );
  OAI211_X1 U10079 ( .C1(n8788), .C2(n8666), .A(n8522), .B(n8521), .ZN(
        P2_U3206) );
  XNOR2_X1 U10080 ( .A(n8523), .B(n8524), .ZN(n8794) );
  XNOR2_X1 U10081 ( .A(n8525), .B(n8524), .ZN(n8527) );
  AOI222_X1 U10082 ( .A1(n8690), .A2(n8527), .B1(n8545), .B2(n8687), .C1(n8526), .C2(n8685), .ZN(n8789) );
  MUX2_X1 U10083 ( .A(n8528), .B(n8789), .S(n8678), .Z(n8531) );
  AOI22_X1 U10084 ( .A1(n8791), .A2(n10307), .B1(n10311), .B2(n8529), .ZN(
        n8530) );
  OAI211_X1 U10085 ( .C1(n8794), .C2(n8666), .A(n8531), .B(n8530), .ZN(
        P2_U3207) );
  XNOR2_X1 U10086 ( .A(n8532), .B(n8533), .ZN(n8800) );
  XNOR2_X1 U10087 ( .A(n8534), .B(n8533), .ZN(n8536) );
  AOI222_X1 U10088 ( .A1(n8690), .A2(n8536), .B1(n8561), .B2(n8687), .C1(n8535), .C2(n8685), .ZN(n8795) );
  INV_X1 U10089 ( .A(n8795), .ZN(n8541) );
  INV_X1 U10090 ( .A(n8797), .ZN(n8539) );
  INV_X1 U10091 ( .A(n8537), .ZN(n8538) );
  OAI22_X1 U10092 ( .A1(n8539), .A2(n8547), .B1(n8538), .B2(n8683), .ZN(n8540)
         );
  OAI21_X1 U10093 ( .B1(n8541), .B2(n8540), .A(n8678), .ZN(n8543) );
  NAND2_X1 U10094 ( .A1(n10320), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8542) );
  OAI211_X1 U10095 ( .C1(n8800), .C2(n8666), .A(n8543), .B(n8542), .ZN(
        P2_U3208) );
  XNOR2_X1 U10096 ( .A(n8544), .B(n8553), .ZN(n8546) );
  AOI222_X1 U10097 ( .A1(n8690), .A2(n8546), .B1(n8545), .B2(n8685), .C1(n8570), .C2(n8687), .ZN(n8801) );
  INV_X1 U10098 ( .A(n8547), .ZN(n8693) );
  AOI22_X1 U10099 ( .A1(n8803), .A2(n8693), .B1(n10311), .B2(n8548), .ZN(n8549) );
  AOI21_X1 U10100 ( .B1(n8801), .B2(n8549), .A(n10320), .ZN(n8556) );
  INV_X1 U10101 ( .A(n8550), .ZN(n8551) );
  AOI21_X1 U10102 ( .B1(n8557), .B2(n8552), .A(n8551), .ZN(n8554) );
  XNOR2_X1 U10103 ( .A(n8554), .B(n8553), .ZN(n8806) );
  OAI22_X1 U10104 ( .A1(n8806), .A2(n8666), .B1(n9001), .B2(n8678), .ZN(n8555)
         );
  OR2_X1 U10105 ( .A1(n8556), .A2(n8555), .ZN(P2_U3209) );
  XNOR2_X1 U10106 ( .A(n8557), .B(n8558), .ZN(n8812) );
  XNOR2_X1 U10107 ( .A(n8559), .B(n8558), .ZN(n8562) );
  AOI222_X1 U10108 ( .A1(n8690), .A2(n8562), .B1(n8561), .B2(n8685), .C1(n8560), .C2(n8687), .ZN(n8807) );
  MUX2_X1 U10109 ( .A(n8563), .B(n8807), .S(n8678), .Z(n8566) );
  AOI22_X1 U10110 ( .A1(n8809), .A2(n10307), .B1(n10311), .B2(n8564), .ZN(
        n8565) );
  OAI211_X1 U10111 ( .C1(n8812), .C2(n8666), .A(n8566), .B(n8565), .ZN(
        P2_U3210) );
  XNOR2_X1 U10112 ( .A(n8567), .B(n8568), .ZN(n8818) );
  XNOR2_X1 U10113 ( .A(n8569), .B(n8568), .ZN(n8571) );
  AOI222_X1 U10114 ( .A1(n8690), .A2(n8571), .B1(n8570), .B2(n8685), .C1(n8589), .C2(n8687), .ZN(n8813) );
  MUX2_X1 U10115 ( .A(n8572), .B(n8813), .S(n8678), .Z(n8575) );
  AOI22_X1 U10116 ( .A1(n8815), .A2(n10307), .B1(n10311), .B2(n8573), .ZN(
        n8574) );
  OAI211_X1 U10117 ( .C1(n8818), .C2(n8666), .A(n8575), .B(n8574), .ZN(
        P2_U3211) );
  XOR2_X1 U10118 ( .A(n8582), .B(n8576), .Z(n8577) );
  OAI222_X1 U10119 ( .A1(n8671), .A2(n8579), .B1(n8673), .B2(n8578), .C1(n8668), .C2(n8577), .ZN(n8819) );
  AOI21_X1 U10120 ( .B1(n10311), .B2(n8580), .A(n8819), .ZN(n8587) );
  INV_X1 U10121 ( .A(n8582), .ZN(n8583) );
  XNOR2_X1 U10122 ( .A(n8581), .B(n8583), .ZN(n8725) );
  OAI22_X1 U10123 ( .A1(n8820), .A2(n8633), .B1(n8584), .B2(n8678), .ZN(n8585)
         );
  AOI21_X1 U10124 ( .B1(n8725), .B2(n8696), .A(n8585), .ZN(n8586) );
  OAI21_X1 U10125 ( .B1(n8587), .B2(n10320), .A(n8586), .ZN(P2_U3212) );
  XNOR2_X1 U10126 ( .A(n8588), .B(n8595), .ZN(n8593) );
  NAND2_X1 U10127 ( .A1(n8589), .A2(n8685), .ZN(n8590) );
  OAI21_X1 U10128 ( .B1(n8591), .B2(n8671), .A(n8590), .ZN(n8592) );
  AOI21_X1 U10129 ( .B1(n8593), .B2(n8690), .A(n8592), .ZN(n8730) );
  XNOR2_X1 U10130 ( .A(n8594), .B(n8595), .ZN(n8728) );
  INV_X1 U10131 ( .A(n8596), .ZN(n8827) );
  AOI22_X1 U10132 ( .A1(n10320), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n10311), 
        .B2(n8597), .ZN(n8598) );
  OAI21_X1 U10133 ( .B1(n8827), .B2(n8633), .A(n8598), .ZN(n8599) );
  AOI21_X1 U10134 ( .B1(n8728), .B2(n8696), .A(n8599), .ZN(n8600) );
  OAI21_X1 U10135 ( .B1(n8730), .B2(n10320), .A(n8600), .ZN(P2_U3213) );
  NAND2_X1 U10136 ( .A1(n8736), .A2(n8601), .ZN(n8602) );
  XNOR2_X1 U10137 ( .A(n8602), .B(n8604), .ZN(n8832) );
  INV_X1 U10138 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8607) );
  XOR2_X1 U10139 ( .A(n8604), .B(n8603), .Z(n8606) );
  AOI222_X1 U10140 ( .A1(n8690), .A2(n8606), .B1(n8637), .B2(n8687), .C1(n8605), .C2(n8685), .ZN(n8828) );
  MUX2_X1 U10141 ( .A(n8607), .B(n8828), .S(n8678), .Z(n8610) );
  AOI22_X1 U10142 ( .A1(n8829), .A2(n10307), .B1(n10311), .B2(n8608), .ZN(
        n8609) );
  OAI211_X1 U10143 ( .C1(n8832), .C2(n8666), .A(n8610), .B(n8609), .ZN(
        P2_U3214) );
  NAND2_X1 U10144 ( .A1(n8649), .A2(n8611), .ZN(n8636) );
  NAND2_X1 U10145 ( .A1(n8636), .A2(n8635), .ZN(n8634) );
  NAND2_X1 U10146 ( .A1(n8634), .A2(n8612), .ZN(n8613) );
  XNOR2_X1 U10147 ( .A(n8613), .B(n6149), .ZN(n8614) );
  NAND2_X1 U10148 ( .A1(n8614), .A2(n8690), .ZN(n8618) );
  AOI22_X1 U10149 ( .A1(n8616), .A2(n8687), .B1(n8685), .B2(n8615), .ZN(n8617)
         );
  NAND2_X1 U10150 ( .A1(n8618), .A2(n8617), .ZN(n8741) );
  INV_X1 U10151 ( .A(n8741), .ZN(n8627) );
  INV_X1 U10152 ( .A(n8619), .ZN(n8620) );
  OAI22_X1 U10153 ( .A1(n8678), .A2(n8621), .B1(n8620), .B2(n8683), .ZN(n8622)
         );
  AOI21_X1 U10154 ( .B1(n8737), .B2(n10307), .A(n8622), .ZN(n8626) );
  NAND2_X1 U10155 ( .A1(n8624), .A2(n8623), .ZN(n8735) );
  NAND3_X1 U10156 ( .A1(n8736), .A2(n8696), .A3(n8735), .ZN(n8625) );
  OAI211_X1 U10157 ( .C1(n8627), .C2(n10320), .A(n8626), .B(n8625), .ZN(
        P2_U3215) );
  INV_X1 U10158 ( .A(n8629), .ZN(n8630) );
  AOI21_X1 U10159 ( .B1(n8635), .B2(n8628), .A(n8630), .ZN(n8837) );
  INV_X1 U10160 ( .A(n8837), .ZN(n8642) );
  INV_X1 U10161 ( .A(n8631), .ZN(n8836) );
  OAI22_X1 U10162 ( .A1(n8836), .A2(n8633), .B1(n8632), .B2(n8683), .ZN(n8641)
         );
  OAI211_X1 U10163 ( .C1(n8636), .C2(n8635), .A(n8634), .B(n8690), .ZN(n8639)
         );
  AOI22_X1 U10164 ( .A1(n8685), .A2(n8637), .B1(n8659), .B2(n8687), .ZN(n8638)
         );
  NAND2_X1 U10165 ( .A1(n8639), .A2(n8638), .ZN(n8834) );
  MUX2_X1 U10166 ( .A(n8834), .B(P2_REG2_REG_17__SCAN_IN), .S(n10320), .Z(
        n8640) );
  AOI211_X1 U10167 ( .C1(n8696), .C2(n8642), .A(n8641), .B(n8640), .ZN(n8643)
         );
  INV_X1 U10168 ( .A(n8643), .ZN(P2_U3216) );
  XNOR2_X1 U10169 ( .A(n8644), .B(n8645), .ZN(n8845) );
  AOI21_X1 U10170 ( .B1(n8646), .B2(n8645), .A(n8668), .ZN(n8650) );
  OAI22_X1 U10171 ( .A1(n8672), .A2(n8671), .B1(n8647), .B2(n8673), .ZN(n8648)
         );
  AOI21_X1 U10172 ( .B1(n8650), .B2(n8649), .A(n8648), .ZN(n8841) );
  MUX2_X1 U10173 ( .A(n8841), .B(n8651), .S(n10320), .Z(n8655) );
  INV_X1 U10174 ( .A(n8652), .ZN(n8653) );
  AOI22_X1 U10175 ( .A1(n8842), .A2(n10307), .B1(n10311), .B2(n8653), .ZN(
        n8654) );
  OAI211_X1 U10176 ( .C1(n8845), .C2(n8666), .A(n8655), .B(n8654), .ZN(
        P2_U3217) );
  XNOR2_X1 U10177 ( .A(n8656), .B(n8658), .ZN(n8852) );
  XNOR2_X1 U10178 ( .A(n8657), .B(n8658), .ZN(n8660) );
  AOI222_X1 U10179 ( .A1(n8690), .A2(n8660), .B1(n8659), .B2(n8685), .C1(n8686), .C2(n8687), .ZN(n8846) );
  MUX2_X1 U10180 ( .A(n8661), .B(n8846), .S(n8678), .Z(n8665) );
  INV_X1 U10181 ( .A(n8662), .ZN(n8663) );
  AOI22_X1 U10182 ( .A1(n8848), .A2(n10307), .B1(n10311), .B2(n8663), .ZN(
        n8664) );
  OAI211_X1 U10183 ( .C1(n8852), .C2(n8666), .A(n8665), .B(n8664), .ZN(
        P2_U3218) );
  XNOR2_X1 U10184 ( .A(n8667), .B(n8675), .ZN(n8669) );
  OAI222_X1 U10185 ( .A1(n8673), .A2(n8672), .B1(n8671), .B2(n8670), .C1(n8669), .C2(n8668), .ZN(n8751) );
  AOI21_X1 U10186 ( .B1(n8693), .B2(n8855), .A(n8751), .ZN(n8681) );
  XNOR2_X1 U10187 ( .A(n8674), .B(n8675), .ZN(n8856) );
  OAI22_X1 U10188 ( .A1(n8678), .A2(n8677), .B1(n8676), .B2(n8683), .ZN(n8679)
         );
  AOI21_X1 U10189 ( .B1(n8856), .B2(n8696), .A(n8679), .ZN(n8680) );
  OAI21_X1 U10190 ( .B1(n8681), .B2(n10320), .A(n8680), .ZN(P2_U3219) );
  NOR2_X1 U10191 ( .A1(n8683), .A2(n8682), .ZN(n8692) );
  XNOR2_X1 U10192 ( .A(n8684), .B(n8695), .ZN(n8689) );
  AOI222_X1 U10193 ( .A1(n8690), .A2(n8689), .B1(n8688), .B2(n8687), .C1(n8686), .C2(n8685), .ZN(n8859) );
  INV_X1 U10194 ( .A(n8859), .ZN(n8691) );
  AOI211_X1 U10195 ( .C1(n8693), .C2(n8861), .A(n8692), .B(n8691), .ZN(n8698)
         );
  XNOR2_X1 U10196 ( .A(n8694), .B(n8695), .ZN(n8864) );
  AOI22_X1 U10197 ( .A1(n8864), .A2(n8696), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10320), .ZN(n8697) );
  OAI21_X1 U10198 ( .B1(n8698), .B2(n10310), .A(n8697), .ZN(P2_U3220) );
  NAND2_X1 U10199 ( .A1(n7991), .A2(n8755), .ZN(n8702) );
  INV_X1 U10200 ( .A(n8700), .ZN(n8701) );
  NAND2_X1 U10201 ( .A1(n8701), .A2(n8772), .ZN(n8704) );
  OAI211_X1 U10202 ( .C1(n8772), .C2(n7678), .A(n8702), .B(n8704), .ZN(
        P2_U3490) );
  NAND2_X1 U10203 ( .A1(n8703), .A2(n8755), .ZN(n8705) );
  OAI211_X1 U10204 ( .C1(n8772), .C2(n6320), .A(n8705), .B(n8704), .ZN(
        P2_U3489) );
  MUX2_X1 U10205 ( .A(n9003), .B(n8777), .S(n8772), .Z(n8707) );
  NAND2_X1 U10206 ( .A1(n8779), .A2(n8755), .ZN(n8706) );
  OAI211_X1 U10207 ( .C1(n8782), .C2(n8750), .A(n8707), .B(n8706), .ZN(
        P2_U3487) );
  MUX2_X1 U10208 ( .A(n8708), .B(n8783), .S(n8772), .Z(n8710) );
  NAND2_X1 U10209 ( .A1(n8785), .A2(n8755), .ZN(n8709) );
  OAI211_X1 U10210 ( .C1(n8788), .C2(n8750), .A(n8710), .B(n8709), .ZN(
        P2_U3486) );
  INV_X1 U10211 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8711) );
  MUX2_X1 U10212 ( .A(n8711), .B(n8789), .S(n8772), .Z(n8713) );
  NAND2_X1 U10213 ( .A1(n8791), .A2(n8755), .ZN(n8712) );
  OAI211_X1 U10214 ( .C1(n8750), .C2(n8794), .A(n8713), .B(n8712), .ZN(
        P2_U3485) );
  MUX2_X1 U10215 ( .A(n9016), .B(n8795), .S(n8772), .Z(n8715) );
  NAND2_X1 U10216 ( .A1(n8797), .A2(n8755), .ZN(n8714) );
  OAI211_X1 U10217 ( .C1(n8800), .C2(n8750), .A(n8715), .B(n8714), .ZN(
        P2_U3484) );
  INV_X1 U10218 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U10219 ( .A(n8716), .B(n8801), .S(n8772), .Z(n8718) );
  NAND2_X1 U10220 ( .A1(n8803), .A2(n8755), .ZN(n8717) );
  OAI211_X1 U10221 ( .C1(n8750), .C2(n8806), .A(n8718), .B(n8717), .ZN(
        P2_U3483) );
  INV_X1 U10222 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8719) );
  MUX2_X1 U10223 ( .A(n8719), .B(n8807), .S(n8772), .Z(n8721) );
  NAND2_X1 U10224 ( .A1(n8809), .A2(n8755), .ZN(n8720) );
  OAI211_X1 U10225 ( .C1(n8812), .C2(n8750), .A(n8721), .B(n8720), .ZN(
        P2_U3482) );
  INV_X1 U10226 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8722) );
  MUX2_X1 U10227 ( .A(n8722), .B(n8813), .S(n8772), .Z(n8724) );
  NAND2_X1 U10228 ( .A1(n8815), .A2(n8755), .ZN(n8723) );
  OAI211_X1 U10229 ( .C1(n8818), .C2(n8750), .A(n8724), .B(n8723), .ZN(
        P2_U3481) );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8819), .S(n8772), .Z(n8727) );
  INV_X1 U10231 ( .A(n8725), .ZN(n8821) );
  OAI22_X1 U10232 ( .A1(n8821), .A2(n8750), .B1(n8820), .B2(n8742), .ZN(n8726)
         );
  OR2_X1 U10233 ( .A1(n8727), .A2(n8726), .ZN(P2_U3480) );
  INV_X1 U10234 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U10235 ( .A1(n8728), .A2(n8760), .ZN(n8729) );
  AND2_X1 U10236 ( .A1(n8730), .A2(n8729), .ZN(n8824) );
  MUX2_X1 U10237 ( .A(n8949), .B(n8824), .S(n8772), .Z(n8731) );
  OAI21_X1 U10238 ( .B1(n8827), .B2(n8742), .A(n8731), .ZN(P2_U3479) );
  MUX2_X1 U10239 ( .A(n8732), .B(n8828), .S(n8772), .Z(n8734) );
  NAND2_X1 U10240 ( .A1(n8829), .A2(n8755), .ZN(n8733) );
  OAI211_X1 U10241 ( .C1(n8832), .C2(n8750), .A(n8734), .B(n8733), .ZN(
        P2_U3478) );
  NAND3_X1 U10242 ( .A1(n8736), .A2(n8760), .A3(n8735), .ZN(n8739) );
  NAND2_X1 U10243 ( .A1(n8737), .A2(n8766), .ZN(n8738) );
  NAND2_X1 U10244 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8833), .S(n8772), .Z(
        P2_U3477) );
  MUX2_X1 U10246 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8834), .S(n8772), .Z(n8744) );
  OAI22_X1 U10247 ( .A1(n8837), .A2(n8750), .B1(n8836), .B2(n8742), .ZN(n8743)
         );
  OR2_X1 U10248 ( .A1(n8744), .A2(n8743), .ZN(P2_U3476) );
  MUX2_X1 U10249 ( .A(n8745), .B(n8841), .S(n8772), .Z(n8747) );
  NAND2_X1 U10250 ( .A1(n8842), .A2(n8755), .ZN(n8746) );
  OAI211_X1 U10251 ( .C1(n8845), .C2(n8750), .A(n8747), .B(n8746), .ZN(
        P2_U3475) );
  MUX2_X1 U10252 ( .A(n9107), .B(n8846), .S(n8772), .Z(n8749) );
  NAND2_X1 U10253 ( .A1(n8848), .A2(n8755), .ZN(n8748) );
  OAI211_X1 U10254 ( .C1(n8750), .C2(n8852), .A(n8749), .B(n8748), .ZN(
        P2_U3474) );
  INV_X1 U10255 ( .A(n8751), .ZN(n8853) );
  MUX2_X1 U10256 ( .A(n9020), .B(n8853), .S(n8772), .Z(n8753) );
  AOI22_X1 U10257 ( .A1(n8856), .A2(n8756), .B1(n8755), .B2(n8855), .ZN(n8752)
         );
  NAND2_X1 U10258 ( .A1(n8753), .A2(n8752), .ZN(P2_U3473) );
  MUX2_X1 U10259 ( .A(n8754), .B(n8859), .S(n8772), .Z(n8758) );
  AOI22_X1 U10260 ( .A1(n8864), .A2(n8756), .B1(n8755), .B2(n8861), .ZN(n8757)
         );
  NAND2_X1 U10261 ( .A1(n8758), .A2(n8757), .ZN(P2_U3472) );
  NAND3_X1 U10262 ( .A1(n8761), .A2(n8760), .A3(n8759), .ZN(n8762) );
  OAI211_X1 U10263 ( .C1(n8765), .C2(n8764), .A(n8763), .B(n8762), .ZN(n8867)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8867), .S(n8772), .Z(
        P2_U3471) );
  AOI22_X1 U10265 ( .A1(n8769), .A2(n8768), .B1(n8767), .B2(n8766), .ZN(n8770)
         );
  AND2_X1 U10266 ( .A1(n8771), .A2(n8770), .ZN(n10323) );
  INV_X1 U10267 ( .A(n10323), .ZN(n8773) );
  MUX2_X1 U10268 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8773), .S(n8772), .Z(
        P2_U3460) );
  AOI21_X1 U10269 ( .B1(n10341), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8774), .ZN(
        n8775) );
  OAI21_X1 U10270 ( .B1(n8776), .B2(n8835), .A(n8775), .ZN(P2_U3457) );
  INV_X1 U10271 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8778) );
  MUX2_X1 U10272 ( .A(n8778), .B(n8777), .S(n10338), .Z(n8781) );
  NAND2_X1 U10273 ( .A1(n8779), .A2(n8862), .ZN(n8780) );
  OAI211_X1 U10274 ( .C1(n8782), .C2(n8851), .A(n8781), .B(n8780), .ZN(
        P2_U3455) );
  INV_X1 U10275 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8784) );
  MUX2_X1 U10276 ( .A(n8784), .B(n8783), .S(n10338), .Z(n8787) );
  NAND2_X1 U10277 ( .A1(n8785), .A2(n8862), .ZN(n8786) );
  OAI211_X1 U10278 ( .C1(n8788), .C2(n8851), .A(n8787), .B(n8786), .ZN(
        P2_U3454) );
  INV_X1 U10279 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8790) );
  MUX2_X1 U10280 ( .A(n8790), .B(n8789), .S(n10338), .Z(n8793) );
  NAND2_X1 U10281 ( .A1(n8791), .A2(n8862), .ZN(n8792) );
  OAI211_X1 U10282 ( .C1(n8794), .C2(n8851), .A(n8793), .B(n8792), .ZN(
        P2_U3453) );
  INV_X1 U10283 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8796) );
  MUX2_X1 U10284 ( .A(n8796), .B(n8795), .S(n10338), .Z(n8799) );
  NAND2_X1 U10285 ( .A1(n8797), .A2(n8862), .ZN(n8798) );
  OAI211_X1 U10286 ( .C1(n8800), .C2(n8851), .A(n8799), .B(n8798), .ZN(
        P2_U3452) );
  INV_X1 U10287 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10288 ( .A(n8802), .B(n8801), .S(n10338), .Z(n8805) );
  NAND2_X1 U10289 ( .A1(n8803), .A2(n8862), .ZN(n8804) );
  OAI211_X1 U10290 ( .C1(n8806), .C2(n8851), .A(n8805), .B(n8804), .ZN(
        P2_U3451) );
  INV_X1 U10291 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8808) );
  MUX2_X1 U10292 ( .A(n8808), .B(n8807), .S(n10338), .Z(n8811) );
  NAND2_X1 U10293 ( .A1(n8809), .A2(n8862), .ZN(n8810) );
  OAI211_X1 U10294 ( .C1(n8812), .C2(n8851), .A(n8811), .B(n8810), .ZN(
        P2_U3450) );
  INV_X1 U10295 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U10296 ( .A(n8814), .B(n8813), .S(n10338), .Z(n8817) );
  NAND2_X1 U10297 ( .A1(n8815), .A2(n8862), .ZN(n8816) );
  OAI211_X1 U10298 ( .C1(n8818), .C2(n8851), .A(n8817), .B(n8816), .ZN(
        P2_U3449) );
  MUX2_X1 U10299 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8819), .S(n10338), .Z(
        n8823) );
  OAI22_X1 U10300 ( .A1(n8821), .A2(n8851), .B1(n8820), .B2(n8835), .ZN(n8822)
         );
  OR2_X1 U10301 ( .A1(n8823), .A2(n8822), .ZN(P2_U3448) );
  INV_X1 U10302 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8825) );
  MUX2_X1 U10303 ( .A(n8825), .B(n8824), .S(n10338), .Z(n8826) );
  OAI21_X1 U10304 ( .B1(n8827), .B2(n8835), .A(n8826), .ZN(P2_U3447) );
  MUX2_X1 U10305 ( .A(n9134), .B(n8828), .S(n10338), .Z(n8831) );
  NAND2_X1 U10306 ( .A1(n8829), .A2(n8862), .ZN(n8830) );
  OAI211_X1 U10307 ( .C1(n8832), .C2(n8851), .A(n8831), .B(n8830), .ZN(
        P2_U3446) );
  MUX2_X1 U10308 ( .A(n8833), .B(P2_REG0_REG_18__SCAN_IN), .S(n10341), .Z(
        P2_U3444) );
  MUX2_X1 U10309 ( .A(n8834), .B(P2_REG0_REG_17__SCAN_IN), .S(n10341), .Z(
        n8839) );
  OAI22_X1 U10310 ( .A1(n8837), .A2(n8851), .B1(n8836), .B2(n8835), .ZN(n8838)
         );
  OR2_X1 U10311 ( .A1(n8839), .A2(n8838), .ZN(P2_U3441) );
  INV_X1 U10312 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U10313 ( .A(n8841), .B(n8840), .S(n10341), .Z(n8844) );
  NAND2_X1 U10314 ( .A1(n8842), .A2(n8862), .ZN(n8843) );
  OAI211_X1 U10315 ( .C1(n8845), .C2(n8851), .A(n8844), .B(n8843), .ZN(
        P2_U3438) );
  INV_X1 U10316 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10317 ( .A(n8847), .B(n8846), .S(n10338), .Z(n8850) );
  NAND2_X1 U10318 ( .A1(n8848), .A2(n8862), .ZN(n8849) );
  OAI211_X1 U10319 ( .C1(n8852), .C2(n8851), .A(n8850), .B(n8849), .ZN(
        P2_U3435) );
  INV_X1 U10320 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U10321 ( .A(n8854), .B(n8853), .S(n10338), .Z(n8858) );
  AOI22_X1 U10322 ( .A1(n8856), .A2(n8863), .B1(n8862), .B2(n8855), .ZN(n8857)
         );
  NAND2_X1 U10323 ( .A1(n8858), .A2(n8857), .ZN(P2_U3432) );
  INV_X1 U10324 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8860) );
  MUX2_X1 U10325 ( .A(n8860), .B(n8859), .S(n10338), .Z(n8866) );
  AOI22_X1 U10326 ( .A1(n8864), .A2(n8863), .B1(n8862), .B2(n8861), .ZN(n8865)
         );
  NAND2_X1 U10327 ( .A1(n8866), .A2(n8865), .ZN(P2_U3429) );
  MUX2_X1 U10328 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8867), .S(n10338), .Z(
        P2_U3426) );
  OAI222_X1 U10329 ( .A1(n8874), .A2(n8870), .B1(n8869), .B2(P2_U3151), .C1(
        n8868), .C2(n8878), .ZN(P2_U3266) );
  INV_X1 U10330 ( .A(n8871), .ZN(n10017) );
  AOI21_X1 U10331 ( .B1(n9173), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8872), .ZN(
        n8873) );
  OAI21_X1 U10332 ( .B1(n10017), .B2(n8874), .A(n8873), .ZN(P2_U3267) );
  INV_X1 U10333 ( .A(n8875), .ZN(n10020) );
  AOI21_X1 U10334 ( .B1(n9173), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8876), .ZN(
        n8877) );
  OAI21_X1 U10335 ( .B1(n10020), .B2(n8874), .A(n8877), .ZN(P2_U3268) );
  OAI222_X1 U10336 ( .A1(n8874), .A2(n8880), .B1(P2_U3151), .B2(n8879), .C1(
        n9007), .C2(n8878), .ZN(P2_U3269) );
  NAND2_X1 U10337 ( .A1(keyinput1), .A2(keyinput12), .ZN(n8882) );
  NOR3_X1 U10338 ( .A1(keyinput105), .A2(keyinput71), .A3(n8882), .ZN(n8883)
         );
  NAND3_X1 U10339 ( .A1(keyinput3), .A2(keyinput114), .A3(n8883), .ZN(n8897)
         );
  NOR2_X1 U10340 ( .A1(keyinput123), .A2(keyinput96), .ZN(n8884) );
  NAND3_X1 U10341 ( .A1(keyinput41), .A2(keyinput115), .A3(n8884), .ZN(n8885)
         );
  NOR3_X1 U10342 ( .A1(keyinput67), .A2(keyinput122), .A3(n8885), .ZN(n8895)
         );
  INV_X1 U10343 ( .A(keyinput78), .ZN(n8886) );
  NAND4_X1 U10344 ( .A1(keyinput99), .A2(keyinput46), .A3(keyinput25), .A4(
        n8886), .ZN(n8893) );
  NOR2_X1 U10345 ( .A1(keyinput34), .A2(keyinput112), .ZN(n8887) );
  NAND3_X1 U10346 ( .A1(keyinput45), .A2(keyinput62), .A3(n8887), .ZN(n8892)
         );
  INV_X1 U10347 ( .A(keyinput103), .ZN(n8888) );
  NAND4_X1 U10348 ( .A1(keyinput57), .A2(keyinput33), .A3(keyinput22), .A4(
        n8888), .ZN(n8891) );
  NOR2_X1 U10349 ( .A1(keyinput91), .A2(keyinput110), .ZN(n8889) );
  NAND3_X1 U10350 ( .A1(keyinput74), .A2(keyinput65), .A3(n8889), .ZN(n8890)
         );
  NOR4_X1 U10351 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n8894)
         );
  NAND4_X1 U10352 ( .A1(keyinput89), .A2(keyinput93), .A3(n8895), .A4(n8894), 
        .ZN(n8896) );
  NOR4_X1 U10353 ( .A1(keyinput23), .A2(keyinput39), .A3(n8897), .A4(n8896), 
        .ZN(n8947) );
  NOR4_X1 U10354 ( .A1(keyinput44), .A2(keyinput6), .A3(keyinput24), .A4(
        keyinput68), .ZN(n8903) );
  NAND2_X1 U10355 ( .A1(keyinput47), .A2(keyinput29), .ZN(n8898) );
  NOR3_X1 U10356 ( .A1(keyinput50), .A2(keyinput107), .A3(n8898), .ZN(n8902)
         );
  INV_X1 U10357 ( .A(keyinput58), .ZN(n8899) );
  NOR4_X1 U10358 ( .A1(keyinput48), .A2(keyinput63), .A3(keyinput8), .A4(n8899), .ZN(n8901) );
  NOR4_X1 U10359 ( .A1(keyinput52), .A2(keyinput69), .A3(keyinput95), .A4(
        keyinput76), .ZN(n8900) );
  NAND4_X1 U10360 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8945)
         );
  INV_X1 U10361 ( .A(keyinput4), .ZN(n8906) );
  INV_X1 U10362 ( .A(keyinput88), .ZN(n8904) );
  NAND4_X1 U10363 ( .A1(keyinput26), .A2(keyinput54), .A3(keyinput59), .A4(
        n8904), .ZN(n8905) );
  NOR4_X1 U10364 ( .A1(keyinput113), .A2(keyinput121), .A3(n8906), .A4(n8905), 
        .ZN(n8911) );
  INV_X1 U10365 ( .A(keyinput66), .ZN(n8907) );
  NOR4_X1 U10366 ( .A1(keyinput81), .A2(keyinput2), .A3(keyinput87), .A4(n8907), .ZN(n8910) );
  NAND2_X1 U10367 ( .A1(keyinput111), .A2(keyinput31), .ZN(n8908) );
  NOR3_X1 U10368 ( .A1(keyinput75), .A2(keyinput17), .A3(n8908), .ZN(n8909) );
  NAND3_X1 U10369 ( .A1(n8911), .A2(n8910), .A3(n8909), .ZN(n8944) );
  INV_X1 U10370 ( .A(keyinput14), .ZN(n8912) );
  NAND4_X1 U10371 ( .A1(keyinput97), .A2(keyinput109), .A3(keyinput11), .A4(
        n8912), .ZN(n8913) );
  NOR3_X1 U10372 ( .A1(keyinput124), .A2(keyinput18), .A3(n8913), .ZN(n8927)
         );
  NAND2_X1 U10373 ( .A1(keyinput20), .A2(keyinput125), .ZN(n8914) );
  NOR3_X1 U10374 ( .A1(keyinput36), .A2(keyinput80), .A3(n8914), .ZN(n8915) );
  NAND3_X1 U10375 ( .A1(keyinput32), .A2(keyinput51), .A3(n8915), .ZN(n8925)
         );
  NAND2_X1 U10376 ( .A1(keyinput72), .A2(keyinput92), .ZN(n8916) );
  NOR3_X1 U10377 ( .A1(keyinput77), .A2(keyinput117), .A3(n8916), .ZN(n8923)
         );
  INV_X1 U10378 ( .A(keyinput35), .ZN(n8917) );
  NOR4_X1 U10379 ( .A1(keyinput16), .A2(keyinput30), .A3(keyinput53), .A4(
        n8917), .ZN(n8922) );
  NAND2_X1 U10380 ( .A1(keyinput120), .A2(keyinput56), .ZN(n8918) );
  NOR3_X1 U10381 ( .A1(keyinput27), .A2(keyinput61), .A3(n8918), .ZN(n8921) );
  NAND2_X1 U10382 ( .A1(keyinput85), .A2(keyinput118), .ZN(n8919) );
  NOR3_X1 U10383 ( .A1(keyinput49), .A2(keyinput126), .A3(n8919), .ZN(n8920)
         );
  NAND4_X1 U10384 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n8924)
         );
  NOR4_X1 U10385 ( .A1(keyinput79), .A2(keyinput104), .A3(n8925), .A4(n8924), 
        .ZN(n8926) );
  NAND4_X1 U10386 ( .A1(keyinput40), .A2(keyinput106), .A3(n8927), .A4(n8926), 
        .ZN(n8943) );
  NOR2_X1 U10387 ( .A1(keyinput90), .A2(keyinput19), .ZN(n8928) );
  NAND3_X1 U10388 ( .A1(keyinput42), .A2(keyinput102), .A3(n8928), .ZN(n8929)
         );
  NOR3_X1 U10389 ( .A1(keyinput7), .A2(keyinput94), .A3(n8929), .ZN(n8941) );
  NAND2_X1 U10390 ( .A1(keyinput43), .A2(keyinput119), .ZN(n8930) );
  NOR3_X1 U10391 ( .A1(keyinput70), .A2(keyinput127), .A3(n8930), .ZN(n8931)
         );
  NAND3_X1 U10392 ( .A1(keyinput55), .A2(keyinput21), .A3(n8931), .ZN(n8939)
         );
  AND4_X1 U10393 ( .A1(keyinput13), .A2(keyinput98), .A3(keyinput73), .A4(
        keyinput108), .ZN(n8937) );
  NAND2_X1 U10394 ( .A1(keyinput10), .A2(keyinput101), .ZN(n8932) );
  NOR3_X1 U10395 ( .A1(keyinput38), .A2(keyinput60), .A3(n8932), .ZN(n8936) );
  NAND3_X1 U10396 ( .A1(keyinput84), .A2(keyinput15), .A3(keyinput0), .ZN(
        n8933) );
  NOR2_X1 U10397 ( .A1(keyinput64), .A2(n8933), .ZN(n8935) );
  NOR4_X1 U10398 ( .A1(keyinput9), .A2(keyinput86), .A3(keyinput83), .A4(
        keyinput28), .ZN(n8934) );
  NAND4_X1 U10399 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), .ZN(n8938)
         );
  NOR4_X1 U10400 ( .A1(keyinput5), .A2(keyinput116), .A3(n8939), .A4(n8938), 
        .ZN(n8940) );
  NAND4_X1 U10401 ( .A1(keyinput37), .A2(keyinput82), .A3(n8941), .A4(n8940), 
        .ZN(n8942) );
  NOR4_X1 U10402 ( .A1(n8945), .A2(n8944), .A3(n8943), .A4(n8942), .ZN(n8946)
         );
  AOI21_X1 U10403 ( .B1(n8947), .B2(n8946), .A(keyinput100), .ZN(n9171) );
  AOI22_X1 U10404 ( .A1(n9800), .A2(keyinput101), .B1(n8949), .B2(keyinput13), 
        .ZN(n8948) );
  OAI221_X1 U10405 ( .B1(n9800), .B2(keyinput101), .C1(n8949), .C2(keyinput13), 
        .A(n8948), .ZN(n8959) );
  INV_X1 U10406 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8951) );
  AOI22_X1 U10407 ( .A1(n8952), .A2(keyinput98), .B1(keyinput73), .B2(n8951), 
        .ZN(n8950) );
  OAI221_X1 U10408 ( .B1(n8952), .B2(keyinput98), .C1(n8951), .C2(keyinput73), 
        .A(n8950), .ZN(n8958) );
  AOI22_X1 U10409 ( .A1(n8954), .A2(keyinput108), .B1(keyinput60), .B2(n7178), 
        .ZN(n8953) );
  OAI221_X1 U10410 ( .B1(n8954), .B2(keyinput108), .C1(n7178), .C2(keyinput60), 
        .A(n8953), .ZN(n8957) );
  AOI22_X1 U10411 ( .A1(n10165), .A2(keyinput10), .B1(n5931), .B2(keyinput37), 
        .ZN(n8955) );
  OAI221_X1 U10412 ( .B1(n10165), .B2(keyinput10), .C1(n5931), .C2(keyinput37), 
        .A(n8955), .ZN(n8956) );
  NOR4_X1 U10413 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8998)
         );
  INV_X1 U10414 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10328) );
  INV_X1 U10415 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8961) );
  AOI22_X1 U10416 ( .A1(n10328), .A2(keyinput82), .B1(keyinput7), .B2(n8961), 
        .ZN(n8960) );
  OAI221_X1 U10417 ( .B1(n10328), .B2(keyinput82), .C1(n8961), .C2(keyinput7), 
        .A(n8960), .ZN(n8970) );
  AOI22_X1 U10418 ( .A1(n10037), .A2(keyinput94), .B1(keyinput90), .B2(n10078), 
        .ZN(n8962) );
  OAI221_X1 U10419 ( .B1(n10037), .B2(keyinput94), .C1(n10078), .C2(keyinput90), .A(n8962), .ZN(n8969) );
  AOI22_X1 U10420 ( .A1(n5471), .A2(keyinput42), .B1(n8964), .B2(keyinput19), 
        .ZN(n8963) );
  OAI221_X1 U10421 ( .B1(n5471), .B2(keyinput42), .C1(n8964), .C2(keyinput19), 
        .A(n8963), .ZN(n8968) );
  INV_X1 U10422 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U10423 ( .A1(n8966), .A2(keyinput102), .B1(keyinput5), .B2(n10221), 
        .ZN(n8965) );
  OAI221_X1 U10424 ( .B1(n8966), .B2(keyinput102), .C1(n10221), .C2(keyinput5), 
        .A(n8965), .ZN(n8967) );
  NOR4_X1 U10425 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n8997)
         );
  INV_X1 U10426 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U10427 ( .A1(n10109), .A2(keyinput116), .B1(n8972), .B2(keyinput55), 
        .ZN(n8971) );
  OAI221_X1 U10428 ( .B1(n10109), .B2(keyinput116), .C1(n8972), .C2(keyinput55), .A(n8971), .ZN(n8981) );
  INV_X1 U10429 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U10430 ( .A1(n8974), .A2(keyinput21), .B1(keyinput119), .B2(n10265), 
        .ZN(n8973) );
  OAI221_X1 U10431 ( .B1(n8974), .B2(keyinput21), .C1(n10265), .C2(keyinput119), .A(n8973), .ZN(n8980) );
  AOI22_X1 U10432 ( .A1(n8976), .A2(keyinput127), .B1(keyinput70), .B2(n6710), 
        .ZN(n8975) );
  OAI221_X1 U10433 ( .B1(n8976), .B2(keyinput127), .C1(n6710), .C2(keyinput70), 
        .A(n8975), .ZN(n8979) );
  INV_X1 U10434 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10322) );
  INV_X1 U10435 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U10436 ( .A1(n10322), .A2(keyinput43), .B1(keyinput9), .B2(n10229), 
        .ZN(n8977) );
  OAI221_X1 U10437 ( .B1(n10322), .B2(keyinput43), .C1(n10229), .C2(keyinput9), 
        .A(n8977), .ZN(n8978) );
  NOR4_X1 U10438 ( .A1(n8981), .A2(n8980), .A3(n8979), .A4(n8978), .ZN(n8996)
         );
  INV_X1 U10439 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8983) );
  AOI22_X1 U10440 ( .A1(n8984), .A2(keyinput0), .B1(keyinput84), .B2(n8983), 
        .ZN(n8982) );
  OAI221_X1 U10441 ( .B1(n8984), .B2(keyinput0), .C1(n8983), .C2(keyinput84), 
        .A(n8982), .ZN(n8994) );
  INV_X1 U10442 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8986) );
  INV_X1 U10443 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U10444 ( .A1(n8986), .A2(keyinput28), .B1(keyinput15), .B2(n10336), 
        .ZN(n8985) );
  OAI221_X1 U10445 ( .B1(n8986), .B2(keyinput28), .C1(n10336), .C2(keyinput15), 
        .A(n8985), .ZN(n8993) );
  AOI22_X1 U10446 ( .A1(n8988), .A2(keyinput64), .B1(keyinput23), .B2(P1_U3086), .ZN(n8987) );
  OAI221_X1 U10447 ( .B1(n8988), .B2(keyinput64), .C1(P1_U3086), .C2(
        keyinput23), .A(n8987), .ZN(n8992) );
  XOR2_X1 U10448 ( .A(n7612), .B(keyinput83), .Z(n8990) );
  XNOR2_X1 U10449 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput86), .ZN(n8989) );
  NAND2_X1 U10450 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NOR4_X1 U10451 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n8991), .ZN(n8995)
         );
  NAND4_X1 U10452 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n9169)
         );
  INV_X1 U10453 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9001) );
  AOI22_X1 U10454 ( .A1(n9001), .A2(keyinput39), .B1(keyinput12), .B2(n9000), 
        .ZN(n8999) );
  OAI221_X1 U10455 ( .B1(n9001), .B2(keyinput39), .C1(n9000), .C2(keyinput12), 
        .A(n8999), .ZN(n9014) );
  AOI22_X1 U10456 ( .A1(n9004), .A2(keyinput71), .B1(keyinput3), .B2(n9003), 
        .ZN(n9002) );
  OAI221_X1 U10457 ( .B1(n9004), .B2(keyinput71), .C1(n9003), .C2(keyinput3), 
        .A(n9002), .ZN(n9013) );
  AOI22_X1 U10458 ( .A1(n9007), .A2(keyinput114), .B1(n9006), .B2(keyinput105), 
        .ZN(n9005) );
  OAI221_X1 U10459 ( .B1(n9007), .B2(keyinput114), .C1(n9006), .C2(keyinput105), .A(n9005), .ZN(n9012) );
  AOI22_X1 U10460 ( .A1(n9010), .A2(keyinput1), .B1(keyinput45), .B2(n9009), 
        .ZN(n9008) );
  OAI221_X1 U10461 ( .B1(n9010), .B2(keyinput1), .C1(n9009), .C2(keyinput45), 
        .A(n9008), .ZN(n9011) );
  NOR4_X1 U10462 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n9057)
         );
  AOI22_X1 U10463 ( .A1(n9017), .A2(keyinput25), .B1(keyinput91), .B2(n9016), 
        .ZN(n9015) );
  OAI221_X1 U10464 ( .B1(n9017), .B2(keyinput25), .C1(n9016), .C2(keyinput91), 
        .A(n9015), .ZN(n9018) );
  INV_X1 U10465 ( .A(n9018), .ZN(n9029) );
  AOI22_X1 U10466 ( .A1(n9020), .A2(keyinput99), .B1(keyinput78), .B2(n9194), 
        .ZN(n9019) );
  OAI221_X1 U10467 ( .B1(n9020), .B2(keyinput99), .C1(n9194), .C2(keyinput78), 
        .A(n9019), .ZN(n9021) );
  INV_X1 U10468 ( .A(n9021), .ZN(n9028) );
  XNOR2_X1 U10469 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput46), .ZN(n9024) );
  XNOR2_X1 U10470 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput112), .ZN(n9023) );
  XNOR2_X1 U10471 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput34), .ZN(n9022) );
  AND3_X1 U10472 ( .A1(n9024), .A2(n9023), .A3(n9022), .ZN(n9027) );
  INV_X1 U10473 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10224) );
  INV_X1 U10474 ( .A(keyinput62), .ZN(n9025) );
  XNOR2_X1 U10475 ( .A(n10224), .B(n9025), .ZN(n9026) );
  AND4_X1 U10476 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(n9056)
         );
  INV_X1 U10477 ( .A(SI_15_), .ZN(n9032) );
  AOI22_X1 U10478 ( .A1(n9032), .A2(keyinput74), .B1(n9031), .B2(keyinput110), 
        .ZN(n9030) );
  OAI221_X1 U10479 ( .B1(n9032), .B2(keyinput74), .C1(n9031), .C2(keyinput110), 
        .A(n9030), .ZN(n9042) );
  INV_X1 U10480 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9034) );
  AOI22_X1 U10481 ( .A1(n9034), .A2(keyinput65), .B1(keyinput33), .B2(n7464), 
        .ZN(n9033) );
  OAI221_X1 U10482 ( .B1(n9034), .B2(keyinput65), .C1(n7464), .C2(keyinput33), 
        .A(n9033), .ZN(n9041) );
  INV_X1 U10483 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U10484 ( .A1(n9036), .A2(keyinput57), .B1(keyinput22), .B2(n9469), 
        .ZN(n9035) );
  OAI221_X1 U10485 ( .B1(n9036), .B2(keyinput57), .C1(n9469), .C2(keyinput22), 
        .A(n9035), .ZN(n9040) );
  AOI22_X1 U10486 ( .A1(n9038), .A2(keyinput103), .B1(keyinput89), .B2(n5513), 
        .ZN(n9037) );
  OAI221_X1 U10487 ( .B1(n9038), .B2(keyinput103), .C1(n5513), .C2(keyinput89), 
        .A(n9037), .ZN(n9039) );
  NOR4_X1 U10488 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n9055)
         );
  AOI22_X1 U10489 ( .A1(n9744), .A2(keyinput113), .B1(keyinput122), .B2(n10349), .ZN(n9043) );
  OAI221_X1 U10490 ( .B1(n9744), .B2(keyinput113), .C1(n10349), .C2(
        keyinput122), .A(n9043), .ZN(n9053) );
  INV_X1 U10491 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9045) );
  AOI22_X1 U10492 ( .A1(n9046), .A2(keyinput96), .B1(keyinput123), .B2(n9045), 
        .ZN(n9044) );
  OAI221_X1 U10493 ( .B1(n9046), .B2(keyinput96), .C1(n9045), .C2(keyinput123), 
        .A(n9044), .ZN(n9052) );
  XOR2_X1 U10494 ( .A(n5555), .B(keyinput93), .Z(n9050) );
  XNOR2_X1 U10495 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput41), .ZN(n9049) );
  XNOR2_X1 U10496 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput67), .ZN(n9048) );
  XNOR2_X1 U10497 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput115), .ZN(n9047) );
  NAND4_X1 U10498 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n9051)
         );
  NOR3_X1 U10499 ( .A1(n9053), .A2(n9052), .A3(n9051), .ZN(n9054) );
  NAND4_X1 U10500 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9168)
         );
  INV_X1 U10501 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U10502 ( .A1(n9059), .A2(keyinput125), .B1(keyinput80), .B2(n10330), 
        .ZN(n9058) );
  OAI221_X1 U10503 ( .B1(n9059), .B2(keyinput125), .C1(n10330), .C2(keyinput80), .A(n9058), .ZN(n9067) );
  AOI22_X1 U10504 ( .A1(n7080), .A2(keyinput51), .B1(n8651), .B2(keyinput36), 
        .ZN(n9060) );
  OAI221_X1 U10505 ( .B1(n7080), .B2(keyinput51), .C1(n8651), .C2(keyinput36), 
        .A(n9060), .ZN(n9066) );
  INV_X1 U10506 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U10507 ( .A1(n6708), .A2(keyinput104), .B1(keyinput40), .B2(n10228), 
        .ZN(n9061) );
  OAI221_X1 U10508 ( .B1(n6708), .B2(keyinput104), .C1(n10228), .C2(keyinput40), .A(n9061), .ZN(n9065) );
  INV_X1 U10509 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U10510 ( .A1(n10227), .A2(keyinput20), .B1(n9063), .B2(keyinput79), 
        .ZN(n9062) );
  OAI221_X1 U10511 ( .B1(n10227), .B2(keyinput20), .C1(n9063), .C2(keyinput79), 
        .A(n9062), .ZN(n9064) );
  NOR4_X1 U10512 ( .A1(n9067), .A2(n9066), .A3(n9065), .A4(n9064), .ZN(n9105)
         );
  AOI22_X1 U10513 ( .A1(n9069), .A2(keyinput117), .B1(keyinput32), .B2(n10207), 
        .ZN(n9068) );
  OAI221_X1 U10514 ( .B1(n9069), .B2(keyinput117), .C1(n10207), .C2(keyinput32), .A(n9068), .ZN(n9080) );
  AOI22_X1 U10515 ( .A1(n7220), .A2(keyinput35), .B1(n9071), .B2(keyinput30), 
        .ZN(n9070) );
  OAI221_X1 U10516 ( .B1(n7220), .B2(keyinput35), .C1(n9071), .C2(keyinput30), 
        .A(n9070), .ZN(n9079) );
  AOI22_X1 U10517 ( .A1(n9074), .A2(keyinput77), .B1(keyinput72), .B2(n9073), 
        .ZN(n9072) );
  OAI221_X1 U10518 ( .B1(n9074), .B2(keyinput77), .C1(n9073), .C2(keyinput72), 
        .A(n9072), .ZN(n9078) );
  XNOR2_X1 U10519 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput92), .ZN(n9076) );
  XNOR2_X1 U10520 ( .A(P2_REG0_REG_11__SCAN_IN), .B(keyinput53), .ZN(n9075) );
  NAND2_X1 U10521 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  NOR4_X1 U10522 ( .A1(n9080), .A2(n9079), .A3(n9078), .A4(n9077), .ZN(n9104)
         );
  INV_X1 U10523 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U10524 ( .A1(n6104), .A2(keyinput61), .B1(keyinput38), .B2(n10151), 
        .ZN(n9081) );
  OAI221_X1 U10525 ( .B1(n6104), .B2(keyinput61), .C1(n10151), .C2(keyinput38), 
        .A(n9081), .ZN(n9090) );
  INV_X1 U10526 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U10527 ( .A1(n9083), .A2(keyinput49), .B1(keyinput85), .B2(n10333), 
        .ZN(n9082) );
  OAI221_X1 U10528 ( .B1(n9083), .B2(keyinput49), .C1(n10333), .C2(keyinput85), 
        .A(n9082), .ZN(n9089) );
  INV_X1 U10529 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U10530 ( .A1(n10225), .A2(keyinput56), .B1(n7664), .B2(keyinput120), 
        .ZN(n9084) );
  OAI221_X1 U10531 ( .B1(n10225), .B2(keyinput56), .C1(n7664), .C2(keyinput120), .A(n9084), .ZN(n9088) );
  XOR2_X1 U10532 ( .A(n6112), .B(keyinput27), .Z(n9086) );
  XNOR2_X1 U10533 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput126), .ZN(n9085) );
  NAND2_X1 U10534 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  NOR4_X1 U10535 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9103)
         );
  AOI22_X1 U10536 ( .A1(n9092), .A2(keyinput106), .B1(keyinput109), .B2(n5462), 
        .ZN(n9091) );
  OAI221_X1 U10537 ( .B1(n9092), .B2(keyinput106), .C1(n5462), .C2(keyinput109), .A(n9091), .ZN(n9101) );
  AOI22_X1 U10538 ( .A1(n10154), .A2(keyinput97), .B1(keyinput124), .B2(n9094), 
        .ZN(n9093) );
  OAI221_X1 U10539 ( .B1(n10154), .B2(keyinput97), .C1(n9094), .C2(keyinput124), .A(n9093), .ZN(n9100) );
  XOR2_X1 U10540 ( .A(n6181), .B(keyinput118), .Z(n9098) );
  XNOR2_X1 U10541 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput11), .ZN(n9097) );
  XNOR2_X1 U10542 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput18), .ZN(n9096) );
  XNOR2_X1 U10543 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput14), .ZN(n9095) );
  NAND4_X1 U10544 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9099)
         );
  NOR3_X1 U10545 ( .A1(n9101), .A2(n9100), .A3(n9099), .ZN(n9102) );
  NAND4_X1 U10546 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n9167)
         );
  AOI22_X1 U10547 ( .A1(n9107), .A2(keyinput31), .B1(keyinput17), .B2(n9696), 
        .ZN(n9106) );
  OAI221_X1 U10548 ( .B1(n9107), .B2(keyinput31), .C1(n9696), .C2(keyinput17), 
        .A(n9106), .ZN(n9117) );
  AOI22_X1 U10549 ( .A1(n10179), .A2(keyinput87), .B1(n10222), .B2(keyinput50), 
        .ZN(n9108) );
  OAI221_X1 U10550 ( .B1(n10179), .B2(keyinput87), .C1(n10222), .C2(keyinput50), .A(n9108), .ZN(n9116) );
  INV_X1 U10551 ( .A(P1_B_REG_SCAN_IN), .ZN(n9110) );
  AOI22_X1 U10552 ( .A1(n9111), .A2(keyinput2), .B1(keyinput66), .B2(n9110), 
        .ZN(n9109) );
  OAI221_X1 U10553 ( .B1(n9111), .B2(keyinput2), .C1(n9110), .C2(keyinput66), 
        .A(n9109), .ZN(n9115) );
  XNOR2_X1 U10554 ( .A(P2_REG1_REG_19__SCAN_IN), .B(keyinput81), .ZN(n9113) );
  XNOR2_X1 U10555 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput111), .ZN(n9112) );
  NAND2_X1 U10556 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  NOR4_X1 U10557 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n9165)
         );
  INV_X1 U10558 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9119) );
  AOI22_X1 U10559 ( .A1(n9120), .A2(keyinput121), .B1(keyinput88), .B2(n9119), 
        .ZN(n9118) );
  OAI221_X1 U10560 ( .B1(n9120), .B2(keyinput121), .C1(n9119), .C2(keyinput88), 
        .A(n9118), .ZN(n9124) );
  NAND2_X1 U10561 ( .A1(n5967), .A2(keyinput4), .ZN(n9121) );
  OAI221_X1 U10562 ( .B1(n8881), .B2(keyinput100), .C1(n5967), .C2(keyinput4), 
        .A(n9121), .ZN(n9123) );
  XOR2_X1 U10563 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput26), .Z(n9122) );
  OR3_X1 U10564 ( .A1(n9124), .A2(n9123), .A3(n9122), .ZN(n9129) );
  AOI22_X1 U10565 ( .A1(n9126), .A2(keyinput59), .B1(keyinput75), .B2(n10226), 
        .ZN(n9125) );
  OAI221_X1 U10566 ( .B1(n9126), .B2(keyinput59), .C1(n10226), .C2(keyinput75), 
        .A(n9125), .ZN(n9128) );
  XNOR2_X1 U10567 ( .A(n10223), .B(keyinput54), .ZN(n9127) );
  NOR3_X1 U10568 ( .A1(n9129), .A2(n9128), .A3(n9127), .ZN(n9164) );
  AOI22_X1 U10569 ( .A1(n9132), .A2(keyinput76), .B1(n9131), .B2(keyinput48), 
        .ZN(n9130) );
  OAI221_X1 U10570 ( .B1(n9132), .B2(keyinput76), .C1(n9131), .C2(keyinput48), 
        .A(n9130), .ZN(n9144) );
  AOI22_X1 U10571 ( .A1(n9135), .A2(keyinput69), .B1(keyinput95), .B2(n9134), 
        .ZN(n9133) );
  OAI221_X1 U10572 ( .B1(n9135), .B2(keyinput69), .C1(n9134), .C2(keyinput95), 
        .A(n9133), .ZN(n9143) );
  AOI22_X1 U10573 ( .A1(n9138), .A2(keyinput8), .B1(keyinput16), .B2(n9137), 
        .ZN(n9136) );
  OAI221_X1 U10574 ( .B1(n9138), .B2(keyinput8), .C1(n9137), .C2(keyinput16), 
        .A(n9136), .ZN(n9142) );
  INV_X1 U10575 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9140) );
  AOI22_X1 U10576 ( .A1(n9140), .A2(keyinput58), .B1(keyinput63), .B2(n10230), 
        .ZN(n9139) );
  OAI221_X1 U10577 ( .B1(n9140), .B2(keyinput58), .C1(n10230), .C2(keyinput63), 
        .A(n9139), .ZN(n9141) );
  NOR4_X1 U10578 ( .A1(n9144), .A2(n9143), .A3(n9142), .A4(n9141), .ZN(n9163)
         );
  AOI22_X1 U10579 ( .A1(n9147), .A2(keyinput107), .B1(keyinput52), .B2(n9146), 
        .ZN(n9145) );
  OAI221_X1 U10580 ( .B1(n9147), .B2(keyinput107), .C1(n9146), .C2(keyinput52), 
        .A(n9145), .ZN(n9152) );
  XNOR2_X1 U10581 ( .A(n9148), .B(keyinput68), .ZN(n9151) );
  XNOR2_X1 U10582 ( .A(n9149), .B(keyinput47), .ZN(n9150) );
  OR3_X1 U10583 ( .A1(n9152), .A2(n9151), .A3(n9150), .ZN(n9161) );
  INV_X1 U10584 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9154) );
  AOI22_X1 U10585 ( .A1(n9155), .A2(keyinput6), .B1(n9154), .B2(keyinput24), 
        .ZN(n9153) );
  OAI221_X1 U10586 ( .B1(n9155), .B2(keyinput6), .C1(n9154), .C2(keyinput24), 
        .A(n9153), .ZN(n9160) );
  INV_X1 U10587 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9158) );
  INV_X1 U10588 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9157) );
  AOI22_X1 U10589 ( .A1(n9158), .A2(keyinput29), .B1(keyinput44), .B2(n9157), 
        .ZN(n9156) );
  OAI221_X1 U10590 ( .B1(n9158), .B2(keyinput29), .C1(n9157), .C2(keyinput44), 
        .A(n9156), .ZN(n9159) );
  NOR3_X1 U10591 ( .A1(n9161), .A2(n9160), .A3(n9159), .ZN(n9162) );
  NAND4_X1 U10592 ( .A1(n9165), .A2(n9164), .A3(n9163), .A4(n9162), .ZN(n9166)
         );
  NOR4_X1 U10593 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9170)
         );
  OAI21_X1 U10594 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(n9171), .A(n9170), .ZN(
        n9178) );
  INV_X1 U10595 ( .A(n9172), .ZN(n9176) );
  AOI222_X1 U10596 ( .A1(n9176), .A2(n9175), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9174), .C1(P1_DATAO_REG_10__SCAN_IN), .C2(n9173), .ZN(n9177) );
  XOR2_X1 U10597 ( .A(n9178), .B(n9177), .Z(P2_U3285) );
  INV_X1 U10598 ( .A(n9179), .ZN(n9180) );
  MUX2_X1 U10599 ( .A(n9180), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10600 ( .B1(n9182), .B2(n9181), .A(n4497), .ZN(n9187) );
  NAND2_X1 U10601 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10149)
         );
  OAI21_X1 U10602 ( .B1(n9370), .B2(n9911), .A(n10149), .ZN(n9183) );
  AOI21_X1 U10603 ( .B1(n9372), .B2(n9893), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10604 ( .B1(n9374), .B2(n9758), .A(n9184), .ZN(n9185) );
  AOI21_X1 U10605 ( .B1(n9914), .B2(n9376), .A(n9185), .ZN(n9186) );
  OAI21_X1 U10606 ( .B1(n9187), .B2(n9378), .A(n9186), .ZN(P1_U3215) );
  XNOR2_X1 U10607 ( .A(n9191), .B(n9190), .ZN(n9192) );
  XNOR2_X1 U10608 ( .A(n9193), .B(n9192), .ZN(n9199) );
  OAI22_X1 U10609 ( .A1(n9359), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9194), .ZN(n9195) );
  AOI21_X1 U10610 ( .B1(n9357), .B2(n9857), .A(n9195), .ZN(n9196) );
  OAI21_X1 U10611 ( .B1(n9374), .B2(n9615), .A(n9196), .ZN(n9197) );
  AOI21_X1 U10612 ( .B1(n9622), .B2(n9376), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10613 ( .B1(n9199), .B2(n9378), .A(n9198), .ZN(P1_U3216) );
  NAND2_X1 U10614 ( .A1(n9372), .A2(n8119), .ZN(n9203) );
  NAND2_X1 U10615 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10035)
         );
  NAND2_X1 U10616 ( .A1(n9376), .A2(n9200), .ZN(n9202) );
  NAND2_X1 U10617 ( .A1(n9357), .A2(n9928), .ZN(n9201) );
  NAND4_X1 U10618 ( .A1(n9203), .A2(n10035), .A3(n9202), .A4(n9201), .ZN(n9209) );
  XOR2_X1 U10619 ( .A(n9204), .B(n9331), .Z(n9206) );
  NOR2_X1 U10620 ( .A1(n9206), .A2(n9205), .ZN(n9332) );
  AOI21_X1 U10621 ( .B1(n9206), .B2(n9205), .A(n9332), .ZN(n9207) );
  NOR2_X1 U10622 ( .A1(n9207), .A2(n9378), .ZN(n9208) );
  AOI211_X1 U10623 ( .C1(n9210), .C2(n9361), .A(n9209), .B(n9208), .ZN(n9211)
         );
  INV_X1 U10624 ( .A(n9211), .ZN(P1_U3217) );
  XNOR2_X1 U10625 ( .A(n9214), .B(n9212), .ZN(n9345) );
  NAND2_X1 U10626 ( .A1(n9345), .A2(n9346), .ZN(n9344) );
  NAND2_X1 U10627 ( .A1(n9214), .A2(n9213), .ZN(n9218) );
  AND2_X1 U10628 ( .A1(n9344), .A2(n9218), .ZN(n9220) );
  INV_X1 U10629 ( .A(n9215), .ZN(n9216) );
  XNOR2_X1 U10630 ( .A(n9217), .B(n9216), .ZN(n9219) );
  NAND3_X1 U10631 ( .A1(n9344), .A2(n9219), .A3(n9218), .ZN(n9303) );
  OAI211_X1 U10632 ( .C1(n9220), .C2(n9219), .A(n9352), .B(n9303), .ZN(n9225)
         );
  NOR2_X1 U10633 ( .A1(n9221), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9509) );
  AOI21_X1 U10634 ( .B1(n9372), .B2(n9870), .A(n9509), .ZN(n9222) );
  OAI21_X1 U10635 ( .B1(n9713), .B2(n9370), .A(n9222), .ZN(n9223) );
  AOI21_X1 U10636 ( .B1(n9678), .B2(n9361), .A(n9223), .ZN(n9224) );
  OAI211_X1 U10637 ( .C1(n9874), .C2(n9364), .A(n9225), .B(n9224), .ZN(
        P1_U3219) );
  XNOR2_X1 U10638 ( .A(n9226), .B(n9227), .ZN(n9228) );
  NAND2_X1 U10639 ( .A1(n9228), .A2(n9229), .ZN(n9288) );
  OAI21_X1 U10640 ( .B1(n9229), .B2(n9228), .A(n9288), .ZN(n9230) );
  NAND2_X1 U10641 ( .A1(n9230), .A2(n9352), .ZN(n9235) );
  NAND2_X1 U10642 ( .A1(n9357), .A2(n9930), .ZN(n9231) );
  NAND2_X1 U10643 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10061) );
  OAI211_X1 U10644 ( .C1(n9232), .C2(n9359), .A(n9231), .B(n10061), .ZN(n9233)
         );
  AOI21_X1 U10645 ( .B1(n10184), .B2(n9376), .A(n9233), .ZN(n9234) );
  OAI211_X1 U10646 ( .C1(n9374), .C2(n10181), .A(n9235), .B(n9234), .ZN(
        P1_U3221) );
  OAI21_X1 U10647 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9239) );
  NAND2_X1 U10648 ( .A1(n9239), .A2(n9352), .ZN(n9244) );
  OAI22_X1 U10649 ( .A1(n9359), .A2(n9841), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9240), .ZN(n9242) );
  NOR2_X1 U10650 ( .A1(n9374), .A2(n9651), .ZN(n9241) );
  AOI211_X1 U10651 ( .C1(n9357), .C2(n9870), .A(n9242), .B(n9241), .ZN(n9243)
         );
  OAI211_X1 U10652 ( .C1(n7781), .C2(n9364), .A(n9244), .B(n9243), .ZN(
        P1_U3223) );
  OAI21_X1 U10653 ( .B1(n9247), .B2(n9246), .A(n9245), .ZN(n9248) );
  NAND2_X1 U10654 ( .A1(n9248), .A2(n9352), .ZN(n9254) );
  INV_X1 U10655 ( .A(n9799), .ZN(n9252) );
  AOI21_X1 U10656 ( .B1(n9357), .B2(n8119), .A(n9249), .ZN(n9250) );
  OAI21_X1 U10657 ( .B1(n9911), .B2(n9359), .A(n9250), .ZN(n9251) );
  AOI21_X1 U10658 ( .B1(n9252), .B2(n9361), .A(n9251), .ZN(n9253) );
  OAI211_X1 U10659 ( .C1(n10269), .C2(n9364), .A(n9254), .B(n9253), .ZN(
        P1_U3224) );
  XOR2_X1 U10660 ( .A(n9256), .B(n9255), .Z(n9262) );
  INV_X1 U10661 ( .A(n9257), .ZN(n9582) );
  NAND2_X1 U10662 ( .A1(n9361), .A2(n9582), .ZN(n9259) );
  INV_X1 U10663 ( .A(n9576), .ZN(n9382) );
  AOI22_X1 U10664 ( .A1(n9372), .A2(n9382), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9258) );
  OAI211_X1 U10665 ( .C1(n9842), .C2(n9370), .A(n9259), .B(n9258), .ZN(n9260)
         );
  AOI21_X1 U10666 ( .B1(n9956), .B2(n9376), .A(n9260), .ZN(n9261) );
  OAI21_X1 U10667 ( .B1(n9262), .B2(n9378), .A(n9261), .ZN(P1_U3225) );
  NAND2_X1 U10668 ( .A1(n4444), .A2(n9264), .ZN(n9265) );
  XNOR2_X1 U10669 ( .A(n9263), .B(n9265), .ZN(n9270) );
  NAND2_X1 U10670 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9461) );
  OAI21_X1 U10671 ( .B1(n9359), .B2(n9699), .A(n9461), .ZN(n9266) );
  AOI21_X1 U10672 ( .B1(n9357), .B2(n9893), .A(n9266), .ZN(n9267) );
  OAI21_X1 U10673 ( .B1(n9374), .B2(n9726), .A(n9267), .ZN(n9268) );
  AOI21_X1 U10674 ( .B1(n9725), .B2(n9376), .A(n9268), .ZN(n9269) );
  OAI21_X1 U10675 ( .B1(n9270), .B2(n9378), .A(n9269), .ZN(P1_U3226) );
  XNOR2_X1 U10676 ( .A(n9273), .B(n9272), .ZN(n9274) );
  XNOR2_X1 U10677 ( .A(n9271), .B(n9274), .ZN(n9279) );
  INV_X1 U10678 ( .A(n9713), .ZN(n9871) );
  NAND2_X1 U10679 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10177)
         );
  OAI21_X1 U10680 ( .B1(n9370), .B2(n9712), .A(n10177), .ZN(n9275) );
  AOI21_X1 U10681 ( .B1(n9372), .B2(n9871), .A(n9275), .ZN(n9276) );
  OAI21_X1 U10682 ( .B1(n9374), .B2(n9707), .A(n9276), .ZN(n9277) );
  AOI21_X1 U10683 ( .B1(n9888), .B2(n9376), .A(n9277), .ZN(n9278) );
  OAI21_X1 U10684 ( .B1(n9279), .B2(n9378), .A(n9278), .ZN(P1_U3228) );
  XOR2_X1 U10685 ( .A(n9281), .B(n9280), .Z(n9287) );
  INV_X1 U10686 ( .A(n9631), .ZN(n9383) );
  OAI22_X1 U10687 ( .A1(n9359), .A2(n9566), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9282), .ZN(n9283) );
  AOI21_X1 U10688 ( .B1(n9357), .B2(n9383), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10689 ( .B1(n9374), .B2(n9600), .A(n9284), .ZN(n9285) );
  AOI21_X1 U10690 ( .B1(n9838), .B2(n9376), .A(n9285), .ZN(n9286) );
  OAI21_X1 U10691 ( .B1(n9287), .B2(n9378), .A(n9286), .ZN(P1_U3229) );
  OAI21_X1 U10692 ( .B1(n9289), .B2(n9226), .A(n9288), .ZN(n9293) );
  XNOR2_X1 U10693 ( .A(n9291), .B(n9290), .ZN(n9292) );
  XNOR2_X1 U10694 ( .A(n9293), .B(n9292), .ZN(n9301) );
  NAND2_X1 U10695 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10076) );
  OAI21_X1 U10696 ( .B1(n9370), .B2(n9294), .A(n10076), .ZN(n9295) );
  AOI21_X1 U10697 ( .B1(n9372), .B2(n9387), .A(n9295), .ZN(n9296) );
  OAI21_X1 U10698 ( .B1(n9374), .B2(n9297), .A(n9296), .ZN(n9298) );
  AOI21_X1 U10699 ( .B1(n4416), .B2(n9376), .A(n9298), .ZN(n9300) );
  OAI21_X1 U10700 ( .B1(n9301), .B2(n9378), .A(n9300), .ZN(P1_U3231) );
  NAND2_X1 U10701 ( .A1(n9303), .A2(n9302), .ZN(n9307) );
  NOR2_X1 U10702 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  XNOR2_X1 U10703 ( .A(n9307), .B(n9306), .ZN(n9312) );
  NOR2_X1 U10704 ( .A1(n9374), .A2(n9668), .ZN(n9310) );
  AOI22_X1 U10705 ( .A1(n9372), .A2(n9384), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9308) );
  OAI21_X1 U10706 ( .B1(n9662), .B2(n9370), .A(n9308), .ZN(n9309) );
  AOI211_X1 U10707 ( .C1(n9867), .C2(n9376), .A(n9310), .B(n9309), .ZN(n9311)
         );
  OAI21_X1 U10708 ( .B1(n9312), .B2(n9378), .A(n9311), .ZN(P1_U3233) );
  OAI21_X1 U10709 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9316) );
  NAND2_X1 U10710 ( .A1(n9316), .A2(n9352), .ZN(n9322) );
  INV_X1 U10711 ( .A(n9780), .ZN(n9320) );
  INV_X1 U10712 ( .A(n10276), .ZN(n9902) );
  NOR2_X1 U10713 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9317), .ZN(n10136) );
  AOI21_X1 U10714 ( .B1(n9372), .B2(n9902), .A(n10136), .ZN(n9318) );
  OAI21_X1 U10715 ( .B1(n10274), .B2(n9370), .A(n9318), .ZN(n9319) );
  AOI21_X1 U10716 ( .B1(n9320), .B2(n9361), .A(n9319), .ZN(n9321) );
  OAI211_X1 U10717 ( .C1(n4604), .C2(n9364), .A(n9322), .B(n9321), .ZN(
        P1_U3234) );
  AOI21_X1 U10718 ( .B1(n9325), .B2(n9324), .A(n9323), .ZN(n9330) );
  AOI22_X1 U10719 ( .A1(n9372), .A2(n9383), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9327) );
  NAND2_X1 U10720 ( .A1(n9357), .A2(n9384), .ZN(n9326) );
  OAI211_X1 U10721 ( .C1(n9374), .C2(n9637), .A(n9327), .B(n9326), .ZN(n9328)
         );
  AOI21_X1 U10722 ( .B1(n9854), .B2(n9376), .A(n9328), .ZN(n9329) );
  OAI21_X1 U10723 ( .B1(n9330), .B2(n9378), .A(n9329), .ZN(P1_U3235) );
  INV_X1 U10724 ( .A(n9331), .ZN(n9333) );
  AOI21_X1 U10725 ( .B1(n9333), .B2(n9204), .A(n9332), .ZN(n9337) );
  XNOR2_X1 U10726 ( .A(n9335), .B(n9334), .ZN(n9336) );
  XNOR2_X1 U10727 ( .A(n9337), .B(n9336), .ZN(n9343) );
  NAND2_X1 U10728 ( .A1(n9357), .A2(n9387), .ZN(n9338) );
  NAND2_X1 U10729 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10123)
         );
  OAI211_X1 U10730 ( .C1(n10274), .C2(n9359), .A(n9338), .B(n10123), .ZN(n9341) );
  NOR2_X1 U10731 ( .A1(n9374), .A2(n9339), .ZN(n9340) );
  AOI211_X1 U10732 ( .C1(n10257), .C2(n9376), .A(n9341), .B(n9340), .ZN(n9342)
         );
  OAI21_X1 U10733 ( .B1(n9343), .B2(n9378), .A(n9342), .ZN(P1_U3236) );
  OAI21_X1 U10734 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9347) );
  NAND2_X1 U10735 ( .A1(n9347), .A2(n9352), .ZN(n9351) );
  INV_X1 U10736 ( .A(n9662), .ZN(n9879) );
  NAND2_X1 U10737 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9490) );
  OAI21_X1 U10738 ( .B1(n9370), .B2(n9699), .A(n9490), .ZN(n9349) );
  NOR2_X1 U10739 ( .A1(n9374), .A2(n9695), .ZN(n9348) );
  AOI211_X1 U10740 ( .C1(n9372), .C2(n9879), .A(n9349), .B(n9348), .ZN(n9350)
         );
  OAI211_X1 U10741 ( .C1(n9882), .C2(n9364), .A(n9351), .B(n9350), .ZN(
        P1_U3238) );
  OAI211_X1 U10742 ( .C1(n9355), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9363)
         );
  INV_X1 U10743 ( .A(n9356), .ZN(n9564) );
  AOI22_X1 U10744 ( .A1(n9357), .A2(n9821), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9358) );
  OAI21_X1 U10745 ( .B1(n9527), .B2(n9359), .A(n9358), .ZN(n9360) );
  AOI21_X1 U10746 ( .B1(n9564), .B2(n9361), .A(n9360), .ZN(n9362) );
  OAI211_X1 U10747 ( .C1(n9824), .C2(n9364), .A(n9363), .B(n9362), .ZN(
        P1_U3240) );
  INV_X1 U10748 ( .A(n9365), .ZN(n9366) );
  AOI21_X1 U10749 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9379) );
  AND2_X1 U10750 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U10751 ( .A1(n9370), .A2(n10276), .ZN(n9371) );
  AOI211_X1 U10752 ( .C1(n9372), .C2(n9901), .A(n10162), .B(n9371), .ZN(n9373)
         );
  OAI21_X1 U10753 ( .B1(n9374), .B2(n9743), .A(n9373), .ZN(n9375) );
  AOI21_X1 U10754 ( .B1(n9747), .B2(n9376), .A(n9375), .ZN(n9377) );
  OAI21_X1 U10755 ( .B1(n9379), .B2(n9378), .A(n9377), .ZN(P1_U3241) );
  MUX2_X1 U10756 ( .A(n9380), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9394), .Z(
        P1_U3585) );
  MUX2_X1 U10757 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9381), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8146), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10759 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9822), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10760 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9382), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10761 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9821), .S(P1_U3973), .Z(
        P1_U3579) );
  INV_X1 U10762 ( .A(n9842), .ZN(n9614) );
  MUX2_X1 U10763 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9614), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10764 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9383), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10765 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9857), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10766 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9384), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10767 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9879), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10768 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9871), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10769 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9892), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10770 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9901), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10771 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9893), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10772 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9902), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10773 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9385), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10774 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9386), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10775 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8119), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10776 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9387), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10777 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9928), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10778 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9388), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10779 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9389), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10780 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9390), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10781 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9391), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10782 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9392), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10783 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9393), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10784 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6777), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10785 ( .A(n9395), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9394), .Z(
        P1_U3554) );
  OAI211_X1 U10786 ( .C1(n9397), .C2(n9407), .A(n10175), .B(n9396), .ZN(n9405)
         );
  OAI211_X1 U10787 ( .C1(n9400), .C2(n9399), .A(n10174), .B(n9398), .ZN(n9404)
         );
  AOI22_X1 U10788 ( .A1(n10138), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9403) );
  NAND2_X1 U10789 ( .A1(n10171), .A2(n9401), .ZN(n9402) );
  NAND4_X1 U10790 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(
        P1_U3244) );
  MUX2_X1 U10791 ( .A(n9407), .B(n9406), .S(n10021), .Z(n9409) );
  NAND2_X1 U10792 ( .A1(n9409), .A2(n9408), .ZN(n9410) );
  OAI211_X1 U10793 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9411), .A(n9410), .B(
        P1_U3973), .ZN(n9453) );
  NAND2_X1 U10794 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U10795 ( .A1(n10138), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9412) );
  OAI211_X1 U10796 ( .C1(n10121), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9415)
         );
  INV_X1 U10797 ( .A(n9415), .ZN(n9424) );
  OAI211_X1 U10798 ( .C1(n9418), .C2(n9417), .A(n10174), .B(n9416), .ZN(n9423)
         );
  OAI211_X1 U10799 ( .C1(n9421), .C2(n9420), .A(n10175), .B(n9419), .ZN(n9422)
         );
  NAND4_X1 U10800 ( .A1(n9453), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(
        P1_U3245) );
  INV_X1 U10801 ( .A(n9425), .ZN(n9429) );
  INV_X1 U10802 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9427) );
  OAI21_X1 U10803 ( .B1(n10180), .B2(n9427), .A(n9426), .ZN(n9428) );
  AOI21_X1 U10804 ( .B1(n9429), .B2(n10171), .A(n9428), .ZN(n9438) );
  OAI211_X1 U10805 ( .C1(n9432), .C2(n9431), .A(n10174), .B(n9430), .ZN(n9437)
         );
  OAI211_X1 U10806 ( .C1(n9435), .C2(n9434), .A(n10175), .B(n9433), .ZN(n9436)
         );
  NAND3_X1 U10807 ( .A1(n9438), .A2(n9437), .A3(n9436), .ZN(P1_U3246) );
  NAND2_X1 U10808 ( .A1(n10138), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9441) );
  INV_X1 U10809 ( .A(n9439), .ZN(n9440) );
  OAI211_X1 U10810 ( .C1(n10121), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  INV_X1 U10811 ( .A(n9443), .ZN(n9452) );
  OAI211_X1 U10812 ( .C1(n9446), .C2(n9445), .A(n10175), .B(n9444), .ZN(n9451)
         );
  OAI211_X1 U10813 ( .C1(n9449), .C2(n9448), .A(n10174), .B(n9447), .ZN(n9450)
         );
  NAND4_X1 U10814 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(
        P1_U3247) );
  OAI21_X1 U10815 ( .B1(n9463), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9454), .ZN(
        n10128) );
  MUX2_X1 U10816 ( .A(n9455), .B(P1_REG1_REG_13__SCAN_IN), .S(n10134), .Z(
        n10127) );
  NOR2_X1 U10817 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  AOI21_X1 U10818 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10134), .A(n10126), 
        .ZN(n10145) );
  XNOR2_X1 U10819 ( .A(n10148), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U10820 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  AOI21_X1 U10821 ( .B1(n10148), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10143), 
        .ZN(n9456) );
  NOR2_X1 U10822 ( .A1(n9456), .A2(n9465), .ZN(n9457) );
  XNOR2_X1 U10823 ( .A(n9465), .B(n9456), .ZN(n10155) );
  NOR2_X1 U10824 ( .A1(n10154), .A2(n10155), .ZN(n10153) );
  NOR2_X1 U10825 ( .A1(n9457), .A2(n10153), .ZN(n9459) );
  AOI22_X1 U10826 ( .A1(n9485), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9899), .B2(
        n9468), .ZN(n9458) );
  NAND2_X1 U10827 ( .A1(n9458), .A2(n9459), .ZN(n9484) );
  OAI21_X1 U10828 ( .B1(n9459), .B2(n9458), .A(n9484), .ZN(n9474) );
  NAND2_X1 U10829 ( .A1(n10138), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9460) );
  OAI211_X1 U10830 ( .C1(n10121), .C2(n9468), .A(n9461), .B(n9460), .ZN(n9473)
         );
  OAI21_X1 U10831 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9463), .A(n9462), .ZN(
        n10131) );
  XNOR2_X1 U10832 ( .A(n10134), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U10833 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  AOI22_X1 U10834 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9464), .B1(n10148), 
        .B2(n9759), .ZN(n10141) );
  NOR2_X1 U10835 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  NOR2_X1 U10836 ( .A1(n9744), .A2(n10158), .ZN(n10157) );
  NOR2_X1 U10837 ( .A1(n9467), .A2(n10157), .ZN(n9471) );
  AOI22_X1 U10838 ( .A1(n9485), .A2(n9469), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9468), .ZN(n9470) );
  NOR2_X1 U10839 ( .A1(n9471), .A2(n9470), .ZN(n9478) );
  AOI211_X1 U10840 ( .C1(n9471), .C2(n9470), .A(n9478), .B(n10156), .ZN(n9472)
         );
  AOI211_X1 U10841 ( .C1(n10174), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9475)
         );
  INV_X1 U10842 ( .A(n9475), .ZN(P1_U3259) );
  NAND2_X1 U10843 ( .A1(n9476), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9501) );
  OR2_X1 U10844 ( .A1(n9476), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U10845 ( .A1(n9501), .A2(n9477), .ZN(n9483) );
  AOI21_X1 U10846 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9485), .A(n9478), .ZN(
        n10168) );
  OR2_X1 U10847 ( .A1(n10172), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U10848 ( .A1(n10172), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9479) );
  AND2_X1 U10849 ( .A1(n9480), .A2(n9479), .ZN(n10167) );
  NAND2_X1 U10850 ( .A1(n10168), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U10851 ( .A1(n10166), .A2(n9480), .ZN(n9482) );
  INV_X1 U10852 ( .A(n9502), .ZN(n9481) );
  AOI211_X1 U10853 ( .C1(n9483), .C2(n9482), .A(n10156), .B(n9481), .ZN(n9496)
         );
  OAI21_X1 U10854 ( .B1(n9485), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9484), .ZN(
        n10170) );
  XNOR2_X1 U10855 ( .A(n10172), .B(n9486), .ZN(n10169) );
  AOI22_X1 U10856 ( .A1(n10170), .A2(n10169), .B1(n9487), .B2(n9486), .ZN(
        n9489) );
  NOR2_X1 U10857 ( .A1(n9494), .A2(n9885), .ZN(n9497) );
  AOI21_X1 U10858 ( .B1(n9885), .B2(n9494), .A(n9497), .ZN(n9488) );
  NAND2_X1 U10859 ( .A1(n9489), .A2(n9488), .ZN(n9499) );
  OAI211_X1 U10860 ( .C1(n9489), .C2(n9488), .A(n9499), .B(n10174), .ZN(n9493)
         );
  INV_X1 U10861 ( .A(n9490), .ZN(n9491) );
  AOI21_X1 U10862 ( .B1(n10138), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9491), .ZN(
        n9492) );
  OAI211_X1 U10863 ( .C1(n10121), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OR2_X1 U10864 ( .A1(n9496), .A2(n9495), .ZN(P1_U3261) );
  INV_X1 U10865 ( .A(n9497), .ZN(n9498) );
  NAND2_X1 U10866 ( .A1(n9499), .A2(n9498), .ZN(n9500) );
  XNOR2_X1 U10867 ( .A(n9500), .B(n9877), .ZN(n9505) );
  NAND2_X1 U10868 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  XNOR2_X1 U10869 ( .A(n9503), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U10870 ( .A1(n9507), .A2(n10175), .ZN(n9504) );
  INV_X1 U10871 ( .A(n9505), .ZN(n9506) );
  OAI22_X1 U10872 ( .A1(n9507), .A2(n10156), .B1(n9506), .B2(n10152), .ZN(
        n9508) );
  NAND2_X1 U10873 ( .A1(n9510), .A2(n10191), .ZN(n9513) );
  INV_X1 U10874 ( .A(n9511), .ZN(n9807) );
  NOR2_X1 U10875 ( .A1(n9807), .A2(n10220), .ZN(n9518) );
  AOI21_X1 U10876 ( .B1(n10220), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9518), .ZN(
        n9512) );
  OAI211_X1 U10877 ( .C1(n9514), .C2(n10198), .A(n9513), .B(n9512), .ZN(
        P1_U3263) );
  NOR2_X1 U10878 ( .A1(n10208), .A2(n9517), .ZN(n9519) );
  AOI211_X1 U10879 ( .C1(n9520), .C2(n10211), .A(n9519), .B(n9518), .ZN(n9521)
         );
  OAI21_X1 U10880 ( .B1(n9808), .B2(n10213), .A(n9521), .ZN(P1_U3264) );
  INV_X1 U10881 ( .A(n9522), .ZN(n9524) );
  INV_X1 U10882 ( .A(n9532), .ZN(n9523) );
  NAND3_X1 U10883 ( .A1(n9526), .A2(n9927), .A3(n9525), .ZN(n9531) );
  NOR2_X1 U10884 ( .A1(n9527), .A2(n10273), .ZN(n9529) );
  NOR2_X1 U10885 ( .A1(n9529), .A2(n4999), .ZN(n9530) );
  NAND2_X1 U10886 ( .A1(n9533), .A2(n9532), .ZN(n9811) );
  NAND3_X1 U10887 ( .A1(n9812), .A2(n9811), .A3(n10216), .ZN(n9539) );
  AOI211_X1 U10888 ( .C1(n9814), .C2(n9543), .A(n9778), .B(n4606), .ZN(n9813)
         );
  AOI22_X1 U10889 ( .A1(n10220), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9534), 
        .B2(n10194), .ZN(n9535) );
  OAI21_X1 U10890 ( .B1(n9536), .B2(n10198), .A(n9535), .ZN(n9537) );
  AOI21_X1 U10891 ( .B1(n9813), .B2(n10191), .A(n9537), .ZN(n9538) );
  OAI211_X1 U10892 ( .C1(n10220), .C2(n9540), .A(n9539), .B(n9538), .ZN(
        P1_U3265) );
  OAI211_X1 U10893 ( .C1(n9542), .C2(n8144), .A(n9932), .B(n9543), .ZN(n9817)
         );
  INV_X1 U10894 ( .A(n9817), .ZN(n9554) );
  AOI22_X1 U10895 ( .A1(n9728), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9544), .B2(
        n10194), .ZN(n9545) );
  OAI21_X1 U10896 ( .B1(n8144), .B2(n10198), .A(n9545), .ZN(n9553) );
  AOI21_X1 U10897 ( .B1(n9547), .B2(n9546), .A(n10283), .ZN(n9551) );
  OAI22_X1 U10898 ( .A1(n9548), .A2(n10275), .B1(n9576), .B2(n10273), .ZN(
        n9549) );
  AOI21_X1 U10899 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(n9818) );
  NOR2_X1 U10900 ( .A1(n9818), .A2(n10220), .ZN(n9552) );
  AOI211_X1 U10901 ( .C1(n9554), .C2(n10191), .A(n9553), .B(n9552), .ZN(n9555)
         );
  OAI21_X1 U10902 ( .B1(n9948), .B2(n9753), .A(n9555), .ZN(P1_U3266) );
  INV_X1 U10903 ( .A(n9573), .ZN(n9559) );
  OAI21_X1 U10904 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9561) );
  NAND2_X1 U10905 ( .A1(n9561), .A2(n9560), .ZN(n9827) );
  INV_X1 U10906 ( .A(n9581), .ZN(n9562) );
  AOI211_X1 U10907 ( .C1(n9563), .C2(n9562), .A(n9778), .B(n9542), .ZN(n9826)
         );
  NAND2_X1 U10908 ( .A1(n9826), .A2(n10191), .ZN(n9569) );
  AOI22_X1 U10909 ( .A1(n10220), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9564), 
        .B2(n10194), .ZN(n9565) );
  OAI21_X1 U10910 ( .B1(n9779), .B2(n9566), .A(n9565), .ZN(n9567) );
  AOI21_X1 U10911 ( .B1(n9784), .B2(n9822), .A(n9567), .ZN(n9568) );
  OAI211_X1 U10912 ( .C1(n9824), .C2(n10198), .A(n9569), .B(n9568), .ZN(n9570)
         );
  AOI21_X1 U10913 ( .B1(n9827), .B2(n9751), .A(n9570), .ZN(n9571) );
  OAI21_X1 U10914 ( .B1(n9952), .B2(n9753), .A(n9571), .ZN(P1_U3267) );
  XNOR2_X1 U10915 ( .A(n9572), .B(n9575), .ZN(n9959) );
  OAI211_X1 U10916 ( .C1(n9575), .C2(n9574), .A(n9573), .B(n9927), .ZN(n9578)
         );
  OR2_X1 U10917 ( .A1(n9576), .A2(n10275), .ZN(n9577) );
  OAI211_X1 U10918 ( .C1(n9842), .C2(n10273), .A(n9578), .B(n9577), .ZN(n9831)
         );
  INV_X1 U10919 ( .A(n9956), .ZN(n9585) );
  NAND2_X1 U10920 ( .A1(n9598), .A2(n9956), .ZN(n9579) );
  NAND2_X1 U10921 ( .A1(n9579), .A2(n9932), .ZN(n9580) );
  NOR2_X1 U10922 ( .A1(n9581), .A2(n9580), .ZN(n9830) );
  NAND2_X1 U10923 ( .A1(n9830), .A2(n10191), .ZN(n9584) );
  AOI22_X1 U10924 ( .A1(n9728), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9582), .B2(
        n10194), .ZN(n9583) );
  OAI211_X1 U10925 ( .C1(n9585), .C2(n10198), .A(n9584), .B(n9583), .ZN(n9586)
         );
  AOI21_X1 U10926 ( .B1(n9831), .B2(n10208), .A(n9586), .ZN(n9587) );
  OAI21_X1 U10927 ( .B1(n9959), .B2(n9753), .A(n9587), .ZN(P1_U3268) );
  NAND2_X1 U10928 ( .A1(n9643), .A2(n9588), .ZN(n9626) );
  NAND2_X1 U10929 ( .A1(n9626), .A2(n9589), .ZN(n9611) );
  AND2_X1 U10930 ( .A1(n9611), .A2(n9590), .ZN(n9592) );
  NOR2_X1 U10931 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  XNOR2_X1 U10932 ( .A(n9593), .B(n4448), .ZN(n9963) );
  OAI211_X1 U10933 ( .C1(n9595), .C2(n4448), .A(n9594), .B(n9927), .ZN(n9597)
         );
  NAND2_X1 U10934 ( .A1(n9821), .A2(n10234), .ZN(n9596) );
  OAI211_X1 U10935 ( .C1(n9631), .C2(n10273), .A(n9597), .B(n9596), .ZN(n9836)
         );
  INV_X1 U10936 ( .A(n9598), .ZN(n9599) );
  AOI211_X1 U10937 ( .C1(n9838), .C2(n9619), .A(n9778), .B(n9599), .ZN(n9837)
         );
  NAND2_X1 U10938 ( .A1(n9837), .A2(n10191), .ZN(n9603) );
  INV_X1 U10939 ( .A(n9600), .ZN(n9601) );
  AOI22_X1 U10940 ( .A1(n10220), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9601), 
        .B2(n10194), .ZN(n9602) );
  OAI211_X1 U10941 ( .C1(n9604), .C2(n10198), .A(n9603), .B(n9602), .ZN(n9605)
         );
  AOI21_X1 U10942 ( .B1(n9836), .B2(n10208), .A(n9605), .ZN(n9606) );
  OAI21_X1 U10943 ( .B1(n9963), .B2(n9753), .A(n9606), .ZN(P1_U3269) );
  NAND2_X1 U10944 ( .A1(n9607), .A2(n9608), .ZN(n9609) );
  AOI21_X1 U10945 ( .B1(n9613), .B2(n9609), .A(n4461), .ZN(n9846) );
  AND2_X1 U10946 ( .A1(n9611), .A2(n9610), .ZN(n9612) );
  XOR2_X1 U10947 ( .A(n9613), .B(n9612), .Z(n9848) );
  NAND2_X1 U10948 ( .A1(n9848), .A2(n10216), .ZN(n9624) );
  NAND2_X1 U10949 ( .A1(n9784), .A2(n9614), .ZN(n9618) );
  INV_X1 U10950 ( .A(n9615), .ZN(n9616) );
  AOI22_X1 U10951 ( .A1(n9728), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9616), .B2(
        n10194), .ZN(n9617) );
  OAI211_X1 U10952 ( .C1(n9841), .C2(n9779), .A(n9618), .B(n9617), .ZN(n9621)
         );
  OAI211_X1 U10953 ( .C1(n9634), .C2(n9967), .A(n9932), .B(n9619), .ZN(n9844)
         );
  NOR2_X1 U10954 ( .A1(n9844), .A2(n10213), .ZN(n9620) );
  AOI211_X1 U10955 ( .C1(n10211), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9623)
         );
  OAI211_X1 U10956 ( .C1(n9846), .C2(n9789), .A(n9624), .B(n9623), .ZN(
        P1_U3270) );
  NAND2_X1 U10957 ( .A1(n9626), .A2(n9625), .ZN(n9628) );
  XNOR2_X1 U10958 ( .A(n9628), .B(n9627), .ZN(n9971) );
  OAI211_X1 U10959 ( .C1(n9630), .C2(n9629), .A(n9607), .B(n9927), .ZN(n9633)
         );
  OR2_X1 U10960 ( .A1(n9631), .A2(n10275), .ZN(n9632) );
  OAI211_X1 U10961 ( .C1(n9664), .C2(n10273), .A(n9633), .B(n9632), .ZN(n9852)
         );
  INV_X1 U10962 ( .A(n9634), .ZN(n9635) );
  OAI211_X1 U10963 ( .C1(n9636), .C2(n5001), .A(n9635), .B(n9932), .ZN(n9851)
         );
  OAI22_X1 U10964 ( .A1(n10208), .A2(n9638), .B1(n9637), .B2(n10205), .ZN(
        n9639) );
  AOI21_X1 U10965 ( .B1(n9854), .B2(n10211), .A(n9639), .ZN(n9640) );
  OAI21_X1 U10966 ( .B1(n9851), .B2(n10213), .A(n9640), .ZN(n9641) );
  AOI21_X1 U10967 ( .B1(n9852), .B2(n10208), .A(n9641), .ZN(n9642) );
  OAI21_X1 U10968 ( .B1(n9971), .B2(n9753), .A(n9642), .ZN(P1_U3271) );
  XOR2_X1 U10969 ( .A(n9643), .B(n9648), .Z(n9975) );
  NOR2_X1 U10970 ( .A1(n9646), .A2(n9645), .ZN(n9649) );
  OAI21_X1 U10971 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9861) );
  AOI211_X1 U10972 ( .C1(n9650), .C2(n4493), .A(n9778), .B(n5001), .ZN(n9860)
         );
  NAND2_X1 U10973 ( .A1(n9860), .A2(n10191), .ZN(n9657) );
  INV_X1 U10974 ( .A(n9651), .ZN(n9652) );
  AOI22_X1 U10975 ( .A1(n9728), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9652), .B2(
        n10194), .ZN(n9653) );
  OAI21_X1 U10976 ( .B1(n9779), .B2(n9654), .A(n9653), .ZN(n9655) );
  AOI21_X1 U10977 ( .B1(n9784), .B2(n9857), .A(n9655), .ZN(n9656) );
  OAI211_X1 U10978 ( .C1(n7781), .C2(n10198), .A(n9657), .B(n9656), .ZN(n9658)
         );
  AOI21_X1 U10979 ( .B1(n9751), .B2(n9861), .A(n9658), .ZN(n9659) );
  OAI21_X1 U10980 ( .B1(n9975), .B2(n9753), .A(n9659), .ZN(P1_U3272) );
  XOR2_X1 U10981 ( .A(n9660), .B(n9661), .Z(n9979) );
  XNOR2_X1 U10982 ( .A(n8148), .B(n9661), .ZN(n9663) );
  OAI222_X1 U10983 ( .A1(n10275), .A2(n9664), .B1(n9663), .B2(n10283), .C1(
        n10273), .C2(n9662), .ZN(n9865) );
  INV_X1 U10984 ( .A(n9665), .ZN(n9667) );
  OAI211_X1 U10985 ( .C1(n9667), .C2(n9666), .A(n9932), .B(n4493), .ZN(n9864)
         );
  INV_X1 U10986 ( .A(n9668), .ZN(n9669) );
  AOI22_X1 U10987 ( .A1(n9728), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9669), .B2(
        n10194), .ZN(n9671) );
  NAND2_X1 U10988 ( .A1(n9867), .A2(n10211), .ZN(n9670) );
  OAI211_X1 U10989 ( .C1(n9864), .C2(n10213), .A(n9671), .B(n9670), .ZN(n9672)
         );
  AOI21_X1 U10990 ( .B1(n9865), .B2(n10208), .A(n9672), .ZN(n9673) );
  OAI21_X1 U10991 ( .B1(n9979), .B2(n9753), .A(n9673), .ZN(P1_U3273) );
  XOR2_X1 U10992 ( .A(n9674), .B(n9675), .Z(n9983) );
  XNOR2_X1 U10993 ( .A(n9676), .B(n9675), .ZN(n9876) );
  OAI211_X1 U10994 ( .C1(n9677), .C2(n9874), .A(n9932), .B(n9665), .ZN(n9873)
         );
  NAND2_X1 U10995 ( .A1(n9784), .A2(n9870), .ZN(n9680) );
  AOI22_X1 U10996 ( .A1(n9728), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9678), .B2(
        n10194), .ZN(n9679) );
  OAI211_X1 U10997 ( .C1(n9713), .C2(n9779), .A(n9680), .B(n9679), .ZN(n9681)
         );
  AOI21_X1 U10998 ( .B1(n9682), .B2(n10211), .A(n9681), .ZN(n9683) );
  OAI21_X1 U10999 ( .B1(n9873), .B2(n10213), .A(n9683), .ZN(n9684) );
  AOI21_X1 U11000 ( .B1(n9876), .B2(n9751), .A(n9684), .ZN(n9685) );
  OAI21_X1 U11001 ( .B1(n9983), .B2(n9753), .A(n9685), .ZN(P1_U3274) );
  OAI21_X1 U11002 ( .B1(n9688), .B2(n9687), .A(n9686), .ZN(n9987) );
  AND2_X1 U11003 ( .A1(n9689), .A2(n9690), .ZN(n9693) );
  OAI21_X1 U11004 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(n9884) );
  INV_X1 U11005 ( .A(n9677), .ZN(n9694) );
  OAI211_X1 U11006 ( .C1(n9882), .C2(n4494), .A(n9694), .B(n9932), .ZN(n9881)
         );
  OAI22_X1 U11007 ( .A1(n10208), .A2(n9696), .B1(n9695), .B2(n10205), .ZN(
        n9697) );
  AOI21_X1 U11008 ( .B1(n9784), .B2(n9879), .A(n9697), .ZN(n9698) );
  OAI21_X1 U11009 ( .B1(n9699), .B2(n9779), .A(n9698), .ZN(n9700) );
  AOI21_X1 U11010 ( .B1(n9701), .B2(n10211), .A(n9700), .ZN(n9702) );
  OAI21_X1 U11011 ( .B1(n9881), .B2(n10213), .A(n9702), .ZN(n9703) );
  AOI21_X1 U11012 ( .B1(n9884), .B2(n9751), .A(n9703), .ZN(n9704) );
  OAI21_X1 U11013 ( .B1(n9987), .B2(n9753), .A(n9704), .ZN(P1_U3275) );
  XNOR2_X1 U11014 ( .A(n9706), .B(n9705), .ZN(n9891) );
  AOI211_X1 U11015 ( .C1(n9888), .C2(n5008), .A(n9778), .B(n4494), .ZN(n9887)
         );
  INV_X1 U11016 ( .A(n9707), .ZN(n9708) );
  AOI22_X1 U11017 ( .A1(n9728), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9708), .B2(
        n10194), .ZN(n9709) );
  OAI21_X1 U11018 ( .B1(n4602), .B2(n10198), .A(n9709), .ZN(n9717) );
  AOI21_X1 U11019 ( .B1(n9711), .B2(n9710), .A(n10283), .ZN(n9715) );
  OAI22_X1 U11020 ( .A1(n9713), .A2(n10275), .B1(n9712), .B2(n10273), .ZN(
        n9714) );
  AOI21_X1 U11021 ( .B1(n9715), .B2(n9689), .A(n9714), .ZN(n9890) );
  NOR2_X1 U11022 ( .A1(n9890), .A2(n10220), .ZN(n9716) );
  AOI211_X1 U11023 ( .C1(n9887), .C2(n10191), .A(n9717), .B(n9716), .ZN(n9718)
         );
  OAI21_X1 U11024 ( .B1(n9891), .B2(n9753), .A(n9718), .ZN(P1_U3276) );
  AOI21_X1 U11025 ( .B1(n9722), .B2(n9720), .A(n9719), .ZN(n9721) );
  INV_X1 U11026 ( .A(n9721), .ZN(n9992) );
  XNOR2_X1 U11027 ( .A(n9723), .B(n9722), .ZN(n9898) );
  INV_X1 U11028 ( .A(n9725), .ZN(n9895) );
  INV_X1 U11029 ( .A(n5008), .ZN(n9724) );
  AOI211_X1 U11030 ( .C1(n9725), .C2(n9742), .A(n9778), .B(n9724), .ZN(n9896)
         );
  NAND2_X1 U11031 ( .A1(n9896), .A2(n10191), .ZN(n9732) );
  INV_X1 U11032 ( .A(n9726), .ZN(n9727) );
  AOI22_X1 U11033 ( .A1(n9728), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9727), .B2(
        n10194), .ZN(n9729) );
  OAI21_X1 U11034 ( .B1(n9779), .B2(n9912), .A(n9729), .ZN(n9730) );
  AOI21_X1 U11035 ( .B1(n9784), .B2(n9892), .A(n9730), .ZN(n9731) );
  OAI211_X1 U11036 ( .C1(n9895), .C2(n10198), .A(n9732), .B(n9731), .ZN(n9733)
         );
  AOI21_X1 U11037 ( .B1(n9751), .B2(n9898), .A(n9733), .ZN(n9734) );
  OAI21_X1 U11038 ( .B1(n9992), .B2(n9753), .A(n9734), .ZN(P1_U3277) );
  XNOR2_X1 U11039 ( .A(n9735), .B(n9737), .ZN(n9997) );
  INV_X1 U11040 ( .A(n9736), .ZN(n9739) );
  OAI21_X1 U11041 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9741) );
  NAND2_X1 U11042 ( .A1(n9741), .A2(n9740), .ZN(n9907) );
  OAI211_X1 U11043 ( .C1(n9762), .C2(n9905), .A(n9742), .B(n9932), .ZN(n9904)
         );
  NOR2_X1 U11044 ( .A1(n9779), .A2(n10276), .ZN(n9746) );
  OAI22_X1 U11045 ( .A1(n10208), .A2(n9744), .B1(n9743), .B2(n10205), .ZN(
        n9745) );
  AOI211_X1 U11046 ( .C1(n9784), .C2(n9901), .A(n9746), .B(n9745), .ZN(n9749)
         );
  NAND2_X1 U11047 ( .A1(n9747), .A2(n10211), .ZN(n9748) );
  OAI211_X1 U11048 ( .C1(n9904), .C2(n10213), .A(n9749), .B(n9748), .ZN(n9750)
         );
  AOI21_X1 U11049 ( .B1(n9907), .B2(n9751), .A(n9750), .ZN(n9752) );
  OAI21_X1 U11050 ( .B1(n9997), .B2(n9753), .A(n9752), .ZN(P1_U3278) );
  AOI21_X1 U11051 ( .B1(n9754), .B2(n9756), .A(n10283), .ZN(n9755) );
  NAND2_X1 U11052 ( .A1(n9755), .A2(n9736), .ZN(n9916) );
  XNOR2_X1 U11053 ( .A(n9757), .B(n9756), .ZN(n9910) );
  NAND2_X1 U11054 ( .A1(n9910), .A2(n10216), .ZN(n9768) );
  OAI22_X1 U11055 ( .A1(n10208), .A2(n9759), .B1(n9758), .B2(n10205), .ZN(
        n9760) );
  AOI21_X1 U11056 ( .B1(n9784), .B2(n9893), .A(n9760), .ZN(n9761) );
  OAI21_X1 U11057 ( .B1(n9911), .B2(n9779), .A(n9761), .ZN(n9766) );
  INV_X1 U11058 ( .A(n9762), .ZN(n9764) );
  AOI21_X1 U11059 ( .B1(n9776), .B2(n9914), .A(n9778), .ZN(n9763) );
  NAND2_X1 U11060 ( .A1(n9764), .A2(n9763), .ZN(n9915) );
  NOR2_X1 U11061 ( .A1(n9915), .A2(n10213), .ZN(n9765) );
  AOI211_X1 U11062 ( .C1(n10211), .C2(n9914), .A(n9766), .B(n9765), .ZN(n9767)
         );
  OAI211_X1 U11063 ( .C1(n10220), .C2(n9916), .A(n9768), .B(n9767), .ZN(
        P1_U3279) );
  INV_X1 U11064 ( .A(n9769), .ZN(n9773) );
  AOI21_X1 U11065 ( .B1(n9770), .B2(n9771), .A(n9774), .ZN(n9772) );
  NOR2_X1 U11066 ( .A1(n9773), .A2(n9772), .ZN(n10282) );
  XNOR2_X1 U11067 ( .A(n9775), .B(n9774), .ZN(n10286) );
  NAND2_X1 U11068 ( .A1(n10286), .A2(n10216), .ZN(n9788) );
  INV_X1 U11069 ( .A(n9776), .ZN(n9777) );
  AOI211_X1 U11070 ( .C1(n10279), .C2(n9801), .A(n9778), .B(n9777), .ZN(n10277) );
  NOR2_X1 U11071 ( .A1(n9779), .A2(n10274), .ZN(n9783) );
  OAI22_X1 U11072 ( .A1(n10208), .A2(n9781), .B1(n9780), .B2(n10205), .ZN(
        n9782) );
  AOI211_X1 U11073 ( .C1(n9784), .C2(n9902), .A(n9783), .B(n9782), .ZN(n9785)
         );
  OAI21_X1 U11074 ( .B1(n4604), .B2(n10198), .A(n9785), .ZN(n9786) );
  AOI21_X1 U11075 ( .B1(n10277), .B2(n10191), .A(n9786), .ZN(n9787) );
  OAI211_X1 U11076 ( .C1(n10282), .C2(n9789), .A(n9788), .B(n9787), .ZN(
        P1_U3280) );
  INV_X1 U11077 ( .A(n9790), .ZN(n9791) );
  NOR2_X1 U11078 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  AOI21_X1 U11079 ( .B1(n7618), .B2(n9793), .A(n10283), .ZN(n9796) );
  OAI22_X1 U11080 ( .A1(n9911), .A2(n10275), .B1(n9794), .B2(n10273), .ZN(
        n9795) );
  AOI21_X1 U11081 ( .B1(n9770), .B2(n9796), .A(n9795), .ZN(n10267) );
  XNOR2_X1 U11082 ( .A(n9798), .B(n9797), .ZN(n10271) );
  NAND2_X1 U11083 ( .A1(n10271), .A2(n10216), .ZN(n9806) );
  OAI22_X1 U11084 ( .A1(n10208), .A2(n9800), .B1(n9799), .B2(n10205), .ZN(
        n9803) );
  OAI211_X1 U11085 ( .C1(n4516), .C2(n10269), .A(n9932), .B(n9801), .ZN(n10266) );
  NOR2_X1 U11086 ( .A1(n10266), .A2(n10213), .ZN(n9802) );
  AOI211_X1 U11087 ( .C1(n10211), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9805)
         );
  OAI211_X1 U11088 ( .C1(n10220), .C2(n10267), .A(n9806), .B(n9805), .ZN(
        P1_U3281) );
  INV_X1 U11089 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9809) );
  MUX2_X1 U11090 ( .A(n9939), .B(n9809), .S(n5414), .Z(n9810) );
  OAI21_X1 U11091 ( .B1(n9941), .B2(n9935), .A(n9810), .ZN(P1_U3552) );
  NAND3_X1 U11092 ( .A1(n9812), .A2(n9811), .A3(n10285), .ZN(n9815) );
  NAND2_X1 U11093 ( .A1(n9815), .A2(n4489), .ZN(n9942) );
  MUX2_X1 U11094 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9942), .S(n10296), .Z(
        P1_U3550) );
  NAND2_X1 U11095 ( .A1(n9818), .A2(n9817), .ZN(n9944) );
  MUX2_X1 U11096 ( .A(n9944), .B(P1_REG1_REG_27__SCAN_IN), .S(n5414), .Z(n9819) );
  AOI21_X1 U11097 ( .B1(n9833), .B2(n9946), .A(n9819), .ZN(n9820) );
  OAI21_X1 U11098 ( .B1(n9948), .B2(n9909), .A(n9820), .ZN(P1_U3549) );
  AOI22_X1 U11099 ( .A1(n9822), .A2(n10234), .B1(n9929), .B2(n9821), .ZN(n9823) );
  OAI21_X1 U11100 ( .B1(n9824), .B2(n10268), .A(n9823), .ZN(n9825) );
  AOI211_X1 U11101 ( .C1(n9827), .C2(n9927), .A(n9826), .B(n9825), .ZN(n9949)
         );
  MUX2_X1 U11102 ( .A(n9828), .B(n9949), .S(n10296), .Z(n9829) );
  OAI21_X1 U11103 ( .B1(n9952), .B2(n9909), .A(n9829), .ZN(P1_U3548) );
  NOR2_X1 U11104 ( .A1(n9831), .A2(n9830), .ZN(n9954) );
  MUX2_X1 U11105 ( .A(n9954), .B(n9832), .S(n5414), .Z(n9835) );
  NAND2_X1 U11106 ( .A1(n9956), .A2(n9833), .ZN(n9834) );
  OAI211_X1 U11107 ( .C1(n9959), .C2(n9909), .A(n9835), .B(n9834), .ZN(
        P1_U3547) );
  AOI211_X1 U11108 ( .C1(n10280), .C2(n9838), .A(n9837), .B(n9836), .ZN(n9960)
         );
  MUX2_X1 U11109 ( .A(n9839), .B(n9960), .S(n10296), .Z(n9840) );
  OAI21_X1 U11110 ( .B1(n9963), .B2(n9909), .A(n9840), .ZN(P1_U3546) );
  OAI22_X1 U11111 ( .A1(n9842), .A2(n10275), .B1(n9841), .B2(n10273), .ZN(
        n9843) );
  INV_X1 U11112 ( .A(n9843), .ZN(n9845) );
  OAI211_X1 U11113 ( .C1(n9846), .C2(n10283), .A(n9845), .B(n9844), .ZN(n9847)
         );
  AOI21_X1 U11114 ( .B1(n9848), .B2(n10285), .A(n9847), .ZN(n9964) );
  MUX2_X1 U11115 ( .A(n9849), .B(n9964), .S(n10296), .Z(n9850) );
  OAI21_X1 U11116 ( .B1(n9967), .B2(n9935), .A(n9850), .ZN(P1_U3545) );
  INV_X1 U11117 ( .A(n9851), .ZN(n9853) );
  AOI211_X1 U11118 ( .C1(n10280), .C2(n9854), .A(n9853), .B(n9852), .ZN(n9968)
         );
  MUX2_X1 U11119 ( .A(n9855), .B(n9968), .S(n10296), .Z(n9856) );
  OAI21_X1 U11120 ( .B1(n9971), .B2(n9909), .A(n9856), .ZN(P1_U3544) );
  AOI22_X1 U11121 ( .A1(n9857), .A2(n10234), .B1(n9929), .B2(n9870), .ZN(n9858) );
  OAI21_X1 U11122 ( .B1(n7781), .B2(n10268), .A(n9858), .ZN(n9859) );
  AOI211_X1 U11123 ( .C1(n9861), .C2(n9927), .A(n9860), .B(n9859), .ZN(n9972)
         );
  MUX2_X1 U11124 ( .A(n9862), .B(n9972), .S(n10296), .Z(n9863) );
  OAI21_X1 U11125 ( .B1(n9975), .B2(n9909), .A(n9863), .ZN(P1_U3543) );
  INV_X1 U11126 ( .A(n9864), .ZN(n9866) );
  AOI211_X1 U11127 ( .C1(n10280), .C2(n9867), .A(n9866), .B(n9865), .ZN(n9976)
         );
  MUX2_X1 U11128 ( .A(n9868), .B(n9976), .S(n10296), .Z(n9869) );
  OAI21_X1 U11129 ( .B1(n9979), .B2(n9909), .A(n9869), .ZN(P1_U3542) );
  AOI22_X1 U11130 ( .A1(n9871), .A2(n9929), .B1(n10234), .B2(n9870), .ZN(n9872) );
  OAI211_X1 U11131 ( .C1(n9874), .C2(n10268), .A(n9873), .B(n9872), .ZN(n9875)
         );
  AOI21_X1 U11132 ( .B1(n9876), .B2(n9927), .A(n9875), .ZN(n9980) );
  MUX2_X1 U11133 ( .A(n9877), .B(n9980), .S(n10296), .Z(n9878) );
  OAI21_X1 U11134 ( .B1(n9983), .B2(n9909), .A(n9878), .ZN(P1_U3541) );
  AOI22_X1 U11135 ( .A1(n9879), .A2(n10234), .B1(n9929), .B2(n9892), .ZN(n9880) );
  OAI211_X1 U11136 ( .C1(n9882), .C2(n10268), .A(n9881), .B(n9880), .ZN(n9883)
         );
  AOI21_X1 U11137 ( .B1(n9884), .B2(n9927), .A(n9883), .ZN(n9984) );
  MUX2_X1 U11138 ( .A(n9885), .B(n9984), .S(n10296), .Z(n9886) );
  OAI21_X1 U11139 ( .B1(n9987), .B2(n9909), .A(n9886), .ZN(P1_U3540) );
  AOI21_X1 U11140 ( .B1(n10280), .B2(n9888), .A(n9887), .ZN(n9889) );
  OAI211_X1 U11141 ( .C1(n9891), .C2(n10233), .A(n9890), .B(n9889), .ZN(n9988)
         );
  MUX2_X1 U11142 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9988), .S(n10296), .Z(
        P1_U3539) );
  AOI22_X1 U11143 ( .A1(n9893), .A2(n9929), .B1(n10234), .B2(n9892), .ZN(n9894) );
  OAI21_X1 U11144 ( .B1(n9895), .B2(n10268), .A(n9894), .ZN(n9897) );
  AOI211_X1 U11145 ( .C1(n9898), .C2(n9927), .A(n9897), .B(n9896), .ZN(n9989)
         );
  MUX2_X1 U11146 ( .A(n9899), .B(n9989), .S(n10296), .Z(n9900) );
  OAI21_X1 U11147 ( .B1(n9992), .B2(n9909), .A(n9900), .ZN(P1_U3538) );
  AOI22_X1 U11148 ( .A1(n9929), .A2(n9902), .B1(n9901), .B2(n10234), .ZN(n9903) );
  OAI211_X1 U11149 ( .C1(n9905), .C2(n10268), .A(n9904), .B(n9903), .ZN(n9906)
         );
  AOI21_X1 U11150 ( .B1(n9907), .B2(n9927), .A(n9906), .ZN(n9993) );
  MUX2_X1 U11151 ( .A(n10154), .B(n9993), .S(n10296), .Z(n9908) );
  OAI21_X1 U11152 ( .B1(n9997), .B2(n9909), .A(n9908), .ZN(P1_U3537) );
  NAND2_X1 U11153 ( .A1(n9910), .A2(n10285), .ZN(n9918) );
  OAI22_X1 U11154 ( .A1(n9912), .A2(n10275), .B1(n9911), .B2(n10273), .ZN(
        n9913) );
  AOI21_X1 U11155 ( .B1(n9914), .B2(n10280), .A(n9913), .ZN(n9917) );
  NAND4_X1 U11156 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9998)
         );
  MUX2_X1 U11157 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9998), .S(n10296), .Z(
        P1_U3536) );
  OAI21_X1 U11158 ( .B1(n9920), .B2(n9925), .A(n9919), .ZN(n10188) );
  INV_X1 U11159 ( .A(n10188), .ZN(n9934) );
  INV_X1 U11160 ( .A(n9921), .ZN(n9923) );
  NAND2_X1 U11161 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  XOR2_X1 U11162 ( .A(n9925), .B(n9924), .Z(n9926) );
  AOI222_X1 U11163 ( .A1(n9930), .A2(n9929), .B1(n9928), .B2(n10234), .C1(
        n9927), .C2(n9926), .ZN(n10190) );
  INV_X1 U11164 ( .A(n9931), .ZN(n9933) );
  OAI211_X1 U11165 ( .C1(n9933), .C2(n4418), .A(n9932), .B(n5009), .ZN(n10186)
         );
  OAI211_X1 U11166 ( .C1(n10233), .C2(n9934), .A(n10190), .B(n10186), .ZN(
        n10002) );
  OAI22_X1 U11167 ( .A1(n9935), .A2(n4418), .B1(n10296), .B2(n6637), .ZN(n9936) );
  AOI21_X1 U11168 ( .B1(n10002), .B2(n10296), .A(n9936), .ZN(n9937) );
  INV_X1 U11169 ( .A(n9937), .ZN(P1_U3530) );
  INV_X1 U11170 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9938) );
  MUX2_X1 U11171 ( .A(n9939), .B(n9938), .S(n10287), .Z(n9940) );
  OAI21_X1 U11172 ( .B1(n9941), .B2(n10000), .A(n9940), .ZN(P1_U3520) );
  MUX2_X1 U11173 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9942), .S(n10289), .Z(
        P1_U3518) );
  MUX2_X1 U11174 ( .A(n9944), .B(P1_REG0_REG_27__SCAN_IN), .S(n10287), .Z(
        n9945) );
  AOI21_X1 U11175 ( .B1(n9955), .B2(n9946), .A(n9945), .ZN(n9947) );
  OAI21_X1 U11176 ( .B1(n9948), .B2(n9996), .A(n9947), .ZN(P1_U3517) );
  MUX2_X1 U11177 ( .A(n9950), .B(n9949), .S(n10289), .Z(n9951) );
  OAI21_X1 U11178 ( .B1(n9952), .B2(n9996), .A(n9951), .ZN(P1_U3516) );
  MUX2_X1 U11179 ( .A(n9954), .B(n9953), .S(n10287), .Z(n9958) );
  NAND2_X1 U11180 ( .A1(n9956), .A2(n9955), .ZN(n9957) );
  OAI211_X1 U11181 ( .C1(n9959), .C2(n9996), .A(n9958), .B(n9957), .ZN(
        P1_U3515) );
  MUX2_X1 U11182 ( .A(n9961), .B(n9960), .S(n10289), .Z(n9962) );
  OAI21_X1 U11183 ( .B1(n9963), .B2(n9996), .A(n9962), .ZN(P1_U3514) );
  MUX2_X1 U11184 ( .A(n9965), .B(n9964), .S(n10289), .Z(n9966) );
  OAI21_X1 U11185 ( .B1(n9967), .B2(n10000), .A(n9966), .ZN(P1_U3513) );
  INV_X1 U11186 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9969) );
  MUX2_X1 U11187 ( .A(n9969), .B(n9968), .S(n10289), .Z(n9970) );
  OAI21_X1 U11188 ( .B1(n9971), .B2(n9996), .A(n9970), .ZN(P1_U3512) );
  MUX2_X1 U11189 ( .A(n9973), .B(n9972), .S(n10289), .Z(n9974) );
  OAI21_X1 U11190 ( .B1(n9975), .B2(n9996), .A(n9974), .ZN(P1_U3511) );
  MUX2_X1 U11191 ( .A(n9977), .B(n9976), .S(n10289), .Z(n9978) );
  OAI21_X1 U11192 ( .B1(n9979), .B2(n9996), .A(n9978), .ZN(P1_U3510) );
  MUX2_X1 U11193 ( .A(n9981), .B(n9980), .S(n10289), .Z(n9982) );
  OAI21_X1 U11194 ( .B1(n9983), .B2(n9996), .A(n9982), .ZN(P1_U3509) );
  INV_X1 U11195 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9985) );
  MUX2_X1 U11196 ( .A(n9985), .B(n9984), .S(n10289), .Z(n9986) );
  OAI21_X1 U11197 ( .B1(n9987), .B2(n9996), .A(n9986), .ZN(P1_U3507) );
  MUX2_X1 U11198 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9988), .S(n10289), .Z(
        P1_U3504) );
  MUX2_X1 U11199 ( .A(n9990), .B(n9989), .S(n10289), .Z(n9991) );
  OAI21_X1 U11200 ( .B1(n9992), .B2(n9996), .A(n9991), .ZN(P1_U3501) );
  INV_X1 U11201 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9994) );
  MUX2_X1 U11202 ( .A(n9994), .B(n9993), .S(n10289), .Z(n9995) );
  OAI21_X1 U11203 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(P1_U3498) );
  MUX2_X1 U11204 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9998), .S(n10289), .Z(
        P1_U3495) );
  INV_X1 U11205 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9999) );
  OAI22_X1 U11206 ( .A1(n10000), .A2(n4418), .B1(n10289), .B2(n9999), .ZN(
        n10001) );
  AOI21_X1 U11207 ( .B1(n10002), .B2(n10289), .A(n10001), .ZN(n10003) );
  INV_X1 U11208 ( .A(n10003), .ZN(P1_U3477) );
  MUX2_X1 U11209 ( .A(P1_D_REG_1__SCAN_IN), .B(n10006), .S(n10231), .Z(
        P1_U3440) );
  MUX2_X1 U11210 ( .A(P1_D_REG_0__SCAN_IN), .B(n10007), .S(n10231), .Z(
        P1_U3439) );
  NAND3_X1 U11211 ( .A1(n5374), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10011) );
  OAI22_X1 U11212 ( .A1(n10008), .A2(n10011), .B1(n10010), .B2(n10009), .ZN(
        n10012) );
  AOI21_X1 U11213 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10015) );
  INV_X1 U11214 ( .A(n10015), .ZN(P1_U3324) );
  OAI222_X1 U11215 ( .A1(n5381), .A2(P1_U3086), .B1(n8174), .B2(n10017), .C1(
        n10016), .C2(n10018), .ZN(P1_U3327) );
  OAI222_X1 U11216 ( .A1(P1_U3086), .A2(n10021), .B1(n8174), .B2(n10020), .C1(
        n10019), .C2(n10018), .ZN(P1_U3328) );
  MUX2_X1 U11217 ( .A(n10022), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U11218 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10026) );
  NAND2_X1 U11219 ( .A1(n10175), .A2(n10026), .ZN(n10032) );
  AOI21_X1 U11220 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10030) );
  NAND2_X1 U11221 ( .A1(n10174), .A2(n10030), .ZN(n10031) );
  OAI211_X1 U11222 ( .C1(n10121), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        n10034) );
  INV_X1 U11223 ( .A(n10034), .ZN(n10036) );
  OAI211_X1 U11224 ( .C1(n10180), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        P1_U3253) );
  AOI211_X1 U11225 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10152), .ZN(
        n10044) );
  AOI211_X1 U11226 ( .C1(n10042), .C2(n4454), .A(n10041), .B(n10156), .ZN(
        n10043) );
  AOI211_X1 U11227 ( .C1(n10171), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10046) );
  INV_X1 U11228 ( .A(n10046), .ZN(n10048) );
  AOI211_X1 U11229 ( .C1(n10138), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n10048), .B(
        n10047), .ZN(n10049) );
  INV_X1 U11230 ( .A(n10049), .ZN(P1_U3250) );
  INV_X1 U11231 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10063) );
  INV_X1 U11232 ( .A(n10050), .ZN(n10060) );
  INV_X1 U11233 ( .A(n10051), .ZN(n10055) );
  INV_X1 U11234 ( .A(n10052), .ZN(n10054) );
  AOI211_X1 U11235 ( .C1(n10055), .C2(n10054), .A(n10053), .B(n10152), .ZN(
        n10059) );
  AOI211_X1 U11236 ( .C1(n10057), .C2(n4524), .A(n10056), .B(n10156), .ZN(
        n10058) );
  AOI211_X1 U11237 ( .C1(n10171), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10062) );
  OAI211_X1 U11238 ( .C1(n10180), .C2(n10063), .A(n10062), .B(n10061), .ZN(
        P1_U3251) );
  OAI21_X1 U11239 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10067) );
  NAND2_X1 U11240 ( .A1(n10175), .A2(n10067), .ZN(n10073) );
  OAI21_X1 U11241 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10071) );
  NAND2_X1 U11242 ( .A1(n10174), .A2(n10071), .ZN(n10072) );
  OAI211_X1 U11243 ( .C1(n10121), .C2(n10074), .A(n10073), .B(n10072), .ZN(
        n10075) );
  INV_X1 U11244 ( .A(n10075), .ZN(n10077) );
  OAI211_X1 U11245 ( .C1(n10180), .C2(n10078), .A(n10077), .B(n10076), .ZN(
        P1_U3252) );
  XNOR2_X1 U11246 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U11247 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10094) );
  INV_X1 U11248 ( .A(n10079), .ZN(n10083) );
  INV_X1 U11249 ( .A(n10080), .ZN(n10082) );
  AOI211_X1 U11250 ( .C1(n10083), .C2(n10082), .A(n10081), .B(n10152), .ZN(
        n10090) );
  INV_X1 U11251 ( .A(n10084), .ZN(n10088) );
  INV_X1 U11252 ( .A(n10085), .ZN(n10087) );
  AOI211_X1 U11253 ( .C1(n10088), .C2(n10087), .A(n10086), .B(n10156), .ZN(
        n10089) );
  AOI211_X1 U11254 ( .C1(n10171), .C2(n10091), .A(n10090), .B(n10089), .ZN(
        n10093) );
  OAI211_X1 U11255 ( .C1(n10180), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        P1_U3248) );
  AOI21_X1 U11256 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10098) );
  NAND2_X1 U11257 ( .A1(n10175), .A2(n10098), .ZN(n10104) );
  AOI21_X1 U11258 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10102) );
  NAND2_X1 U11259 ( .A1(n10174), .A2(n10102), .ZN(n10103) );
  OAI211_X1 U11260 ( .C1(n10121), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10106) );
  INV_X1 U11261 ( .A(n10106), .ZN(n10108) );
  OAI211_X1 U11262 ( .C1(n10180), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        P1_U3249) );
  INV_X1 U11263 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10125) );
  AOI21_X1 U11264 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n10113) );
  NAND2_X1 U11265 ( .A1(n10175), .A2(n10113), .ZN(n10119) );
  AOI21_X1 U11266 ( .B1(n10116), .B2(n10115), .A(n10114), .ZN(n10117) );
  NAND2_X1 U11267 ( .A1(n10174), .A2(n10117), .ZN(n10118) );
  OAI211_X1 U11268 ( .C1(n10121), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10122) );
  INV_X1 U11269 ( .A(n10122), .ZN(n10124) );
  OAI211_X1 U11270 ( .C1(n10180), .C2(n10125), .A(n10124), .B(n10123), .ZN(
        P1_U3254) );
  AOI211_X1 U11271 ( .C1(n10128), .C2(n10127), .A(n10152), .B(n10126), .ZN(
        n10133) );
  AOI211_X1 U11272 ( .C1(n10131), .C2(n10130), .A(n10156), .B(n10129), .ZN(
        n10132) );
  AOI211_X1 U11273 ( .C1(n10171), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10135) );
  INV_X1 U11274 ( .A(n10135), .ZN(n10137) );
  AOI211_X1 U11275 ( .C1(n10138), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10137), 
        .B(n10136), .ZN(n10139) );
  INV_X1 U11276 ( .A(n10139), .ZN(P1_U3256) );
  AOI211_X1 U11277 ( .C1(n10142), .C2(n10141), .A(n10140), .B(n10156), .ZN(
        n10147) );
  AOI211_X1 U11278 ( .C1(n10145), .C2(n10144), .A(n10152), .B(n10143), .ZN(
        n10146) );
  AOI211_X1 U11279 ( .C1(n10171), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  OAI211_X1 U11280 ( .C1(n10180), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        P1_U3257) );
  AOI211_X1 U11281 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10160) );
  AOI211_X1 U11282 ( .C1(n10158), .C2(n9744), .A(n10157), .B(n10156), .ZN(
        n10159) );
  AOI211_X1 U11283 ( .C1(n10171), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10164) );
  INV_X1 U11284 ( .A(n10162), .ZN(n10163) );
  OAI211_X1 U11285 ( .C1(n10180), .C2(n10165), .A(n10164), .B(n10163), .ZN(
        P1_U3258) );
  OAI21_X1 U11286 ( .B1(n10168), .B2(n10167), .A(n10166), .ZN(n10176) );
  XNOR2_X1 U11287 ( .A(n10170), .B(n10169), .ZN(n10173) );
  AOI222_X1 U11288 ( .A1(n10176), .A2(n10175), .B1(n10174), .B2(n10173), .C1(
        n10172), .C2(n10171), .ZN(n10178) );
  OAI211_X1 U11289 ( .C1(n10180), .C2(n10179), .A(n10178), .B(n10177), .ZN(
        P1_U3260) );
  OAI22_X1 U11290 ( .A1(n10208), .A2(n10182), .B1(n10181), .B2(n10205), .ZN(
        n10183) );
  AOI21_X1 U11291 ( .B1(n10211), .B2(n10184), .A(n10183), .ZN(n10185) );
  OAI21_X1 U11292 ( .B1(n10186), .B2(n10213), .A(n10185), .ZN(n10187) );
  AOI21_X1 U11293 ( .B1(n10188), .B2(n10216), .A(n10187), .ZN(n10189) );
  OAI21_X1 U11294 ( .B1(n10220), .B2(n10190), .A(n10189), .ZN(P1_U3285) );
  NAND2_X1 U11295 ( .A1(n10192), .A2(n10191), .ZN(n10197) );
  INV_X1 U11296 ( .A(n10193), .ZN(n10195) );
  AOI22_X1 U11297 ( .A1(n9728), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10195), .B2(
        n10194), .ZN(n10196) );
  OAI211_X1 U11298 ( .C1(n10199), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10200) );
  AOI21_X1 U11299 ( .B1(n10216), .B2(n10201), .A(n10200), .ZN(n10202) );
  OAI21_X1 U11300 ( .B1(n10220), .B2(n10203), .A(n10202), .ZN(P1_U3287) );
  INV_X1 U11301 ( .A(n10204), .ZN(n10217) );
  OAI22_X1 U11302 ( .A1(n10208), .A2(n10207), .B1(n10206), .B2(n10205), .ZN(
        n10209) );
  AOI21_X1 U11303 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10212) );
  OAI21_X1 U11304 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10215) );
  AOI21_X1 U11305 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10218) );
  OAI21_X1 U11306 ( .B1(n10220), .B2(n10219), .A(n10218), .ZN(P1_U3289) );
  NOR2_X1 U11307 ( .A1(n10231), .A2(n10221), .ZN(P1_U3294) );
  AND2_X1 U11308 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10232), .ZN(P1_U3295) );
  NOR2_X1 U11309 ( .A1(n10231), .A2(n10222), .ZN(P1_U3296) );
  AND2_X1 U11310 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10232), .ZN(P1_U3297) );
  NOR2_X1 U11311 ( .A1(n10231), .A2(n10223), .ZN(P1_U3298) );
  AND2_X1 U11312 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10232), .ZN(P1_U3299) );
  AND2_X1 U11313 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10232), .ZN(P1_U3300) );
  AND2_X1 U11314 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10232), .ZN(P1_U3301) );
  NOR2_X1 U11315 ( .A1(n10231), .A2(n10224), .ZN(P1_U3302) );
  AND2_X1 U11316 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10232), .ZN(P1_U3303) );
  AND2_X1 U11317 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10232), .ZN(P1_U3304) );
  AND2_X1 U11318 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10232), .ZN(P1_U3305) );
  NOR2_X1 U11319 ( .A1(n10231), .A2(n10225), .ZN(P1_U3306) );
  AND2_X1 U11320 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10232), .ZN(P1_U3307) );
  AND2_X1 U11321 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10232), .ZN(P1_U3308) );
  AND2_X1 U11322 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10232), .ZN(P1_U3309) );
  NOR2_X1 U11323 ( .A1(n10231), .A2(n10226), .ZN(P1_U3310) );
  AND2_X1 U11324 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10232), .ZN(P1_U3311) );
  NOR2_X1 U11325 ( .A1(n10231), .A2(n10227), .ZN(P1_U3312) );
  NOR2_X1 U11326 ( .A1(n10231), .A2(n10228), .ZN(P1_U3313) );
  AND2_X1 U11327 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10232), .ZN(P1_U3314) );
  NOR2_X1 U11328 ( .A1(n10231), .A2(n10229), .ZN(P1_U3315) );
  NOR2_X1 U11329 ( .A1(n10231), .A2(n10230), .ZN(P1_U3316) );
  AND2_X1 U11330 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10232), .ZN(P1_U3317) );
  AND2_X1 U11331 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10232), .ZN(P1_U3318) );
  AND2_X1 U11332 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10232), .ZN(P1_U3319) );
  AND2_X1 U11333 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10232), .ZN(P1_U3320) );
  AND2_X1 U11334 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10232), .ZN(P1_U3321) );
  AND2_X1 U11335 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10232), .ZN(P1_U3322) );
  AND2_X1 U11336 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10232), .ZN(P1_U3323) );
  NAND2_X1 U11337 ( .A1(n10233), .A2(n10283), .ZN(n10238) );
  AOI222_X1 U11338 ( .A1(n10238), .A2(n10237), .B1(n10236), .B2(n10235), .C1(
        n6777), .C2(n10234), .ZN(n10290) );
  INV_X1 U11339 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11340 ( .A1(n10289), .A2(n10290), .B1(n10239), .B2(n10287), .ZN(
        P1_U3453) );
  INV_X1 U11341 ( .A(n10260), .ZN(n10240) );
  NAND2_X1 U11342 ( .A1(n10241), .A2(n10240), .ZN(n10243) );
  OAI211_X1 U11343 ( .C1(n5468), .C2(n10268), .A(n10243), .B(n10242), .ZN(
        n10244) );
  NOR2_X1 U11344 ( .A1(n10245), .A2(n10244), .ZN(n10291) );
  INV_X1 U11345 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U11346 ( .A1(n10289), .A2(n10291), .B1(n10246), .B2(n10287), .ZN(
        P1_U3456) );
  OAI21_X1 U11347 ( .B1(n10248), .B2(n10268), .A(n10247), .ZN(n10249) );
  AOI21_X1 U11348 ( .B1(n10250), .B2(n10285), .A(n10249), .ZN(n10251) );
  AND2_X1 U11349 ( .A1(n10252), .A2(n10251), .ZN(n10292) );
  INV_X1 U11350 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U11351 ( .A1(n10289), .A2(n10292), .B1(n10253), .B2(n10287), .ZN(
        P1_U3468) );
  INV_X1 U11352 ( .A(n10261), .ZN(n10263) );
  OAI22_X1 U11353 ( .A1(n10274), .A2(n10275), .B1(n10254), .B2(n10273), .ZN(
        n10256) );
  AOI211_X1 U11354 ( .C1(n10280), .C2(n10257), .A(n10256), .B(n10255), .ZN(
        n10259) );
  OAI211_X1 U11355 ( .C1(n10261), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        n10262) );
  AOI21_X1 U11356 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10293) );
  AOI22_X1 U11357 ( .A1(n10289), .A2(n10293), .B1(n10265), .B2(n10287), .ZN(
        P1_U3486) );
  OAI211_X1 U11358 ( .C1(n10269), .C2(n10268), .A(n10267), .B(n10266), .ZN(
        n10270) );
  AOI21_X1 U11359 ( .B1(n10271), .B2(n10285), .A(n10270), .ZN(n10294) );
  INV_X1 U11360 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U11361 ( .A1(n10289), .A2(n10294), .B1(n10272), .B2(n10287), .ZN(
        P1_U3489) );
  OAI22_X1 U11362 ( .A1(n10276), .A2(n10275), .B1(n10274), .B2(n10273), .ZN(
        n10278) );
  AOI211_X1 U11363 ( .C1(n10280), .C2(n10279), .A(n10278), .B(n10277), .ZN(
        n10281) );
  OAI21_X1 U11364 ( .B1(n10283), .B2(n10282), .A(n10281), .ZN(n10284) );
  AOI21_X1 U11365 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(n10295) );
  INV_X1 U11366 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U11367 ( .A1(n10289), .A2(n10295), .B1(n10288), .B2(n10287), .ZN(
        P1_U3492) );
  AOI22_X1 U11368 ( .A1(n10296), .A2(n10290), .B1(n5463), .B2(n5414), .ZN(
        P1_U3522) );
  AOI22_X1 U11369 ( .A1(n10296), .A2(n10291), .B1(n5457), .B2(n5414), .ZN(
        P1_U3523) );
  AOI22_X1 U11370 ( .A1(n10296), .A2(n10292), .B1(n5503), .B2(n5414), .ZN(
        P1_U3527) );
  AOI22_X1 U11371 ( .A1(n10296), .A2(n10293), .B1(n6643), .B2(n5414), .ZN(
        P1_U3533) );
  AOI22_X1 U11372 ( .A1(n10296), .A2(n10294), .B1(n5563), .B2(n5414), .ZN(
        P1_U3534) );
  AOI22_X1 U11373 ( .A1(n10296), .A2(n10295), .B1(n9455), .B2(n5414), .ZN(
        P1_U3535) );
  AOI21_X1 U11374 ( .B1(n10299), .B2(n10298), .A(n10297), .ZN(n10309) );
  AOI22_X1 U11375 ( .A1(n10320), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n10311), 
        .B2(n10300), .ZN(n10301) );
  OAI21_X1 U11376 ( .B1(n10320), .B2(n10302), .A(n10301), .ZN(n10305) );
  NOR2_X1 U11377 ( .A1(n10303), .A2(n10314), .ZN(n10304) );
  AOI211_X1 U11378 ( .C1(n10307), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10308) );
  OAI21_X1 U11379 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(P2_U3226) );
  AOI22_X1 U11380 ( .A1(n10313), .A2(n10312), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10311), .ZN(n10318) );
  INV_X1 U11381 ( .A(n10314), .ZN(n10315) );
  AOI22_X1 U11382 ( .A1(n10316), .A2(n10315), .B1(P2_REG2_REG_2__SCAN_IN), 
        .B2(n10320), .ZN(n10317) );
  OAI221_X1 U11383 ( .B1(n10320), .B2(n10319), .C1(n10320), .C2(n10318), .A(
        n10317), .ZN(P2_U3231) );
  AOI22_X1 U11384 ( .A1(n10341), .A2(n10322), .B1(n10321), .B2(n10338), .ZN(
        P2_U3390) );
  INV_X1 U11385 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U11386 ( .A1(n10341), .A2(n10324), .B1(n10323), .B2(n10338), .ZN(
        P2_U3393) );
  INV_X1 U11387 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11388 ( .A1(n10341), .A2(n10326), .B1(n10325), .B2(n10338), .ZN(
        P2_U3396) );
  AOI22_X1 U11389 ( .A1(n10341), .A2(n10328), .B1(n10327), .B2(n10338), .ZN(
        P2_U3399) );
  AOI22_X1 U11390 ( .A1(n10341), .A2(n10330), .B1(n10329), .B2(n10338), .ZN(
        P2_U3402) );
  AOI22_X1 U11391 ( .A1(n10341), .A2(n5967), .B1(n10331), .B2(n10338), .ZN(
        P2_U3405) );
  AOI22_X1 U11392 ( .A1(n10341), .A2(n10333), .B1(n10332), .B2(n10338), .ZN(
        P2_U3408) );
  AOI22_X1 U11393 ( .A1(n10341), .A2(n5988), .B1(n10334), .B2(n10338), .ZN(
        P2_U3411) );
  AOI22_X1 U11394 ( .A1(n10341), .A2(n10336), .B1(n10335), .B2(n10338), .ZN(
        P2_U3414) );
  AOI22_X1 U11395 ( .A1(n10341), .A2(n6023), .B1(n10337), .B2(n10338), .ZN(
        P2_U3417) );
  INV_X1 U11396 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U11397 ( .A1(n10341), .A2(n10340), .B1(n10339), .B2(n10338), .ZN(
        P2_U3420) );
  OAI222_X1 U11398 ( .A1(n10346), .A2(n10345), .B1(n10346), .B2(n10344), .C1(
        n10343), .C2(n10342), .ZN(ADD_1068_U5) );
  AOI21_X1 U11399 ( .B1(n10349), .B2(n10348), .A(n10347), .ZN(ADD_1068_U46) );
  OAI21_X1 U11400 ( .B1(n10352), .B2(n10351), .A(n10350), .ZN(n10353) );
  XNOR2_X1 U11401 ( .A(n10353), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11402 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(ADD_1068_U56) );
  OAI21_X1 U11403 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1068_U57) );
  OAI21_X1 U11404 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1068_U58) );
  OAI21_X1 U11405 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(ADD_1068_U59) );
  OAI21_X1 U11406 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(ADD_1068_U60) );
  OAI21_X1 U11407 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(ADD_1068_U61) );
  OAI21_X1 U11408 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(ADD_1068_U62) );
  OAI21_X1 U11409 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(ADD_1068_U63) );
  OAI21_X1 U11410 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(ADD_1068_U50) );
  OAI21_X1 U11411 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(ADD_1068_U51) );
  OAI21_X1 U11412 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(ADD_1068_U47) );
  OAI21_X1 U11413 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(ADD_1068_U49) );
  OAI21_X1 U11414 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(ADD_1068_U48) );
  AOI21_X1 U11415 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(ADD_1068_U54) );
  AOI21_X1 U11416 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(ADD_1068_U53) );
  OAI21_X1 U11417 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4938 ( .A(n7696), .Z(n7821) );
  AND2_X1 U4944 ( .A1(n6665), .A2(n6664), .ZN(n6924) );
  CLKBUF_X1 U4996 ( .A(n5479), .Z(n5708) );
  CLKBUF_X1 U5746 ( .A(n9299), .Z(n4416) );
  CLKBUF_X1 U5996 ( .A(n10310), .Z(n10320) );
endmodule

