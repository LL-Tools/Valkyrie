

module b21_C_gen_AntiSAT_k_256_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4474, n4475, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550;

  INV_X2 U4979 ( .A(n6149), .ZN(n6185) );
  CLKBUF_X2 U4980 ( .A(n4482), .Z(n8841) );
  INV_X2 U4981 ( .A(n5634), .ZN(n5951) );
  CLKBUF_X2 U4982 ( .A(n5282), .Z(n8851) );
  BUF_X2 U4983 ( .A(n6326), .Z(n7867) );
  NAND2_X1 U4984 ( .A1(n5905), .A2(n5154), .ZN(n5978) );
  XNOR2_X1 U4985 ( .A(n5124), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5130) );
  INV_X1 U4986 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5453) );
  AND2_X2 U4987 ( .A1(n6811), .A2(n5978), .ZN(n5953) );
  OR2_X1 U4988 ( .A1(n9471), .A2(n9448), .ZN(n9443) );
  OR2_X1 U4989 ( .A1(n8590), .A2(n8073), .ZN(n7949) );
  INV_X2 U4990 ( .A(n6815), .ZN(n5327) );
  AND2_X1 U4991 ( .A1(n9174), .A2(n8905), .ZN(n9630) );
  INV_X1 U4992 ( .A(n7660), .ZN(n7723) );
  INV_X1 U4993 ( .A(n6869), .ZN(n10011) );
  INV_X1 U4994 ( .A(n6040), .ZN(n5320) );
  MUX2_X1 U4995 ( .A(n6445), .B(P2_REG2_REG_1__SCAN_IN), .S(n7120), .Z(n6452)
         );
  NAND2_X1 U4996 ( .A1(n4808), .A2(n4574), .ZN(n9333) );
  AOI211_X1 U4997 ( .C1(n8499), .C2(n8524), .A(n8261), .B(n8260), .ZN(n8262)
         );
  AND3_X1 U4998 ( .A1(n6022), .A2(n6021), .A3(n4610), .ZN(n4474) );
  AND4_X1 U4999 ( .A1(n5987), .A2(n6232), .A3(n6163), .A4(n6286), .ZN(n4475)
         );
  OAI21_X2 U5000 ( .B1(n9159), .B2(n5069), .A(n5066), .ZN(n5065) );
  AOI21_X2 U5002 ( .B1(n7280), .B2(P2_REG2_REG_10__SCAN_IN), .A(n4516), .ZN(
        n8102) );
  NOR2_X2 U5003 ( .A1(n7485), .A2(n10072), .ZN(n7537) );
  AND2_X2 U5004 ( .A1(n5456), .A2(n5455), .ZN(n9668) );
  OAI21_X2 U5005 ( .B1(n8390), .B2(n7839), .A(n7978), .ZN(n8357) );
  AND3_X2 U5006 ( .A1(n5193), .A2(n5192), .A3(n5191), .ZN(n6801) );
  XNOR2_X2 U5007 ( .A(n7619), .B(n7617), .ZN(n7788) );
  NAND2_X2 U5008 ( .A1(n7752), .A2(n7613), .ZN(n7619) );
  OAI222_X1 U5009 ( .A1(n9595), .A2(n10273), .B1(n7594), .B2(n6489), .C1(
        P1_U3084), .C2(n6610), .ZN(P1_U3346) );
  NAND2_X2 U5010 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6015) );
  OAI21_X2 U5011 ( .B1(n7293), .B2(n8041), .A(n7292), .ZN(n7377) );
  NAND2_X1 U5012 ( .A1(n7243), .A2(n7918), .ZN(n7293) );
  INV_X1 U5013 ( .A(n6850), .ZN(n6939) );
  NAND4_X2 U5014 ( .A1(n5221), .A2(n5220), .A3(n5219), .A4(n5218), .ZN(n6850)
         );
  NAND2_X4 U5015 ( .A1(n6020), .A2(n6018), .ZN(n6085) );
  XNOR2_X2 U5016 ( .A(n5503), .B(n5502), .ZN(n6637) );
  NAND2_X2 U5017 ( .A1(n4986), .A2(n4985), .ZN(n5503) );
  AOI21_X2 U5018 ( .B1(n7171), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7199), .ZN(
        n7212) );
  AND2_X1 U5019 ( .A1(n5953), .A2(n5160), .ZN(n4477) );
  XNOR2_X2 U5020 ( .A(n5556), .B(n5552), .ZN(n6700) );
  AND2_X1 U5021 ( .A1(n4727), .A2(n4726), .ZN(n5974) );
  XNOR2_X1 U5022 ( .A(n7626), .B(n7624), .ZN(n7704) );
  OR2_X1 U5023 ( .A1(n9348), .A2(n9158), .ZN(n4808) );
  NAND2_X1 U5024 ( .A1(n6230), .A2(n7460), .ZN(n7544) );
  NOR3_X2 U5025 ( .A1(n9409), .A2(n4706), .A3(n9542), .ZN(n9349) );
  AOI21_X1 U5026 ( .B1(n7255), .B2(n8999), .A(n7254), .ZN(n7256) );
  NOR2_X1 U5027 ( .A1(n7312), .A2(n8872), .ZN(n7265) );
  INV_X1 U5028 ( .A(n8031), .ZN(n4478) );
  INV_X2 U5029 ( .A(n6952), .ZN(n9900) );
  NAND4_X1 U5030 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n8088)
         );
  NAND2_X1 U5031 ( .A1(n5291), .A2(n5290), .ZN(n5316) );
  CLKBUF_X2 U5032 ( .A(n6855), .Z(n4483) );
  BUF_X1 U5033 ( .A(n5235), .Z(n4482) );
  CLKBUF_X2 U5034 ( .A(n5217), .Z(n5958) );
  CLKBUF_X2 U5035 ( .A(n6115), .Z(n7737) );
  INV_X4 U5036 ( .A(n5377), .ZN(n8838) );
  NOR2_X1 U5037 ( .A1(n5129), .A2(n5130), .ZN(n5235) );
  INV_X2 U5038 ( .A(n6274), .ZN(n7637) );
  INV_X1 U5039 ( .A(n8848), .ZN(n5347) );
  INV_X2 U5040 ( .A(n5292), .ZN(n5377) );
  NAND2_X1 U5041 ( .A1(n5159), .A2(n5158), .ZN(n9327) );
  INV_X2 U5042 ( .A(n9980), .ZN(n8275) );
  OAI21_X1 U5043 ( .B1(n9499), .B2(n9660), .A(n4782), .ZN(n9573) );
  NAND2_X1 U5044 ( .A1(n4783), .A2(n9214), .ZN(n9499) );
  AOI21_X1 U5045 ( .B1(n5020), .B2(n5970), .A(n5019), .ZN(n5018) );
  NAND2_X1 U5046 ( .A1(n5974), .A2(n5973), .ZN(n5022) );
  AOI21_X1 U5047 ( .B1(n8245), .B2(n10004), .A(n8244), .ZN(n8520) );
  NAND2_X1 U5048 ( .A1(n9236), .A2(n9238), .ZN(n5081) );
  NAND2_X1 U5049 ( .A1(n4810), .A2(n4814), .ZN(n9247) );
  OR2_X1 U5050 ( .A1(n9290), .A2(n4523), .ZN(n4810) );
  OR2_X1 U5051 ( .A1(n9290), .A2(n9165), .ZN(n4824) );
  NAND2_X1 U5052 ( .A1(n7630), .A2(n4529), .ZN(n7760) );
  OR2_X1 U5053 ( .A1(n9159), .A2(n5071), .ZN(n9533) );
  AND2_X1 U5054 ( .A1(n5667), .A2(n5666), .ZN(n8740) );
  OAI21_X1 U5055 ( .B1(n4941), .B2(n4935), .A(n4932), .ZN(n9239) );
  NOR2_X1 U5056 ( .A1(n9363), .A2(n9366), .ZN(n9365) );
  AND2_X1 U5057 ( .A1(n8692), .A2(n4583), .ZN(n8738) );
  NAND2_X1 U5058 ( .A1(n4601), .A2(n4600), .ZN(n8341) );
  OAI21_X1 U5059 ( .B1(n7709), .B2(n4968), .A(n4966), .ZN(n7752) );
  NOR2_X1 U5060 ( .A1(n9193), .A2(n9192), .ZN(n9292) );
  NOR2_X1 U5061 ( .A1(n9367), .A2(n9186), .ZN(n9356) );
  AOI21_X1 U5062 ( .B1(n9400), .B2(n9185), .A(n9184), .ZN(n9367) );
  NOR3_X2 U5063 ( .A1(n8393), .A2(n4775), .A3(n8543), .ZN(n4777) );
  OR2_X2 U5064 ( .A1(n8403), .A2(n8567), .ZN(n8393) );
  AND2_X1 U5065 ( .A1(n9349), .A2(n9339), .ZN(n9334) );
  NAND2_X1 U5066 ( .A1(n5086), .A2(n5084), .ZN(n9142) );
  AND2_X1 U5067 ( .A1(n6280), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U5068 ( .A1(n7335), .A2(n5386), .ZN(n5035) );
  NAND2_X1 U5069 ( .A1(n9829), .A2(n7444), .ZN(n5086) );
  OR2_X1 U5070 ( .A1(n7407), .A2(n7408), .ZN(n7462) );
  NOR2_X1 U5071 ( .A1(n7837), .A2(n8429), .ZN(n4874) );
  AND2_X1 U5072 ( .A1(n7521), .A2(n6250), .ZN(n4965) );
  INV_X1 U5073 ( .A(n4741), .ZN(n4740) );
  OAI21_X1 U5074 ( .B1(n7438), .B2(n4912), .A(n4910), .ZN(n9631) );
  NAND2_X1 U5075 ( .A1(n5305), .A2(n7006), .ZN(n5037) );
  AND2_X1 U5076 ( .A1(n8665), .A2(n5471), .ZN(n5033) );
  NAND2_X1 U5077 ( .A1(n5701), .A2(n5700), .ZN(n9537) );
  NAND2_X1 U5078 ( .A1(n5596), .A2(n5595), .ZN(n9561) );
  NAND2_X1 U5079 ( .A1(n5563), .A2(n5562), .ZN(n9565) );
  OAI21_X1 U5080 ( .B1(n9854), .B2(n9865), .A(n7097), .ZN(n7309) );
  NAND2_X1 U5081 ( .A1(n5511), .A2(n5510), .ZN(n9452) );
  OR2_X1 U5082 ( .A1(n9643), .A2(n9143), .ZN(n9174) );
  AOI21_X1 U5083 ( .B1(n4915), .B2(n4918), .A(n8889), .ZN(n4913) );
  NAND2_X1 U5084 ( .A1(n6254), .A2(n6253), .ZN(n7540) );
  NAND2_X1 U5085 ( .A1(n5485), .A2(n5484), .ZN(n9471) );
  AND2_X1 U5086 ( .A1(n9172), .A2(n9171), .ZN(n4494) );
  NAND2_X1 U5087 ( .A1(n6238), .A2(n6237), .ZN(n10072) );
  NAND2_X1 U5088 ( .A1(n6217), .A2(n6216), .ZN(n7483) );
  NAND2_X1 U5089 ( .A1(n4662), .A2(n5501), .ZN(n5526) );
  NAND2_X1 U5090 ( .A1(n4789), .A2(n9633), .ZN(n9172) );
  NOR2_X1 U5091 ( .A1(n7030), .A2(n4979), .ZN(n4978) );
  OR2_X1 U5092 ( .A1(n5503), .A2(n5502), .ZN(n4662) );
  OR2_X1 U5093 ( .A1(n8089), .A2(n4762), .ZN(n4761) );
  AND2_X1 U5094 ( .A1(n7913), .A2(n7908), .ZN(n8035) );
  INV_X1 U5095 ( .A(n10041), .ZN(n7924) );
  AND2_X1 U5096 ( .A1(n4764), .A2(n4763), .ZN(n8089) );
  AND3_X1 U5097 ( .A1(n6170), .A2(n6169), .A3(n6168), .ZN(n10041) );
  OR2_X1 U5098 ( .A1(n5422), .A2(n4799), .ZN(n4987) );
  NAND2_X1 U5099 ( .A1(n5380), .A2(n5379), .ZN(n7440) );
  NAND3_X1 U5100 ( .A1(n4794), .A2(n4793), .A3(n4795), .ZN(n6496) );
  OR2_X1 U5101 ( .A1(n9855), .A2(n8882), .ZN(n7312) );
  OR2_X1 U5103 ( .A1(n5392), .A2(n4562), .ZN(n4794) );
  OAI211_X1 U5104 ( .C1(n5377), .C2(n10323), .A(n5324), .B(n5323), .ZN(n8882)
         );
  OR2_X1 U5105 ( .A1(n5352), .A2(n5351), .ZN(n8872) );
  NAND2_X2 U5106 ( .A1(n6888), .A2(n8451), .ZN(n9993) );
  XNOR2_X1 U5107 ( .A(n6802), .B(n6801), .ZN(n6818) );
  BUF_X1 U5108 ( .A(n6802), .Z(n4480) );
  INV_X1 U5109 ( .A(n9975), .ZN(n7041) );
  INV_X1 U5110 ( .A(n6759), .ZN(n6884) );
  NOR2_X1 U5111 ( .A1(n6961), .A2(n4698), .ZN(n9857) );
  OAI211_X1 U5112 ( .C1(n6149), .C2(n6476), .A(n6110), .B(n6109), .ZN(n9975)
         );
  NAND2_X1 U5113 ( .A1(n4474), .A2(n4490), .ZN(n6759) );
  NAND2_X1 U5114 ( .A1(n5316), .A2(n5315), .ZN(n5319) );
  XNOR2_X1 U5115 ( .A(n5316), .B(n5315), .ZN(n6476) );
  AND4_X1 U5116 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n6901)
         );
  AND4_X1 U5117 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6870)
         );
  OAI22_X1 U5118 ( .A1(n4796), .A2(n4798), .B1(n5105), .B2(n4801), .ZN(n4795)
         );
  NAND2_X2 U5119 ( .A1(n5178), .A2(n6811), .ZN(n6815) );
  OR2_X1 U5120 ( .A1(n9063), .A2(n5886), .ZN(n5160) );
  AND2_X1 U5121 ( .A1(n7593), .A2(n5130), .ZN(n5282) );
  OAI211_X1 U5122 ( .C1(n5347), .C2(n6478), .A(n5246), .B(n5245), .ZN(n6964)
         );
  AND2_X2 U5123 ( .A1(n6059), .A2(n4479), .ZN(n6326) );
  NAND2_X1 U5124 ( .A1(n6059), .A2(n6468), .ZN(n6149) );
  NOR2_X2 U5125 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  NAND2_X2 U5126 ( .A1(n8619), .A2(n6017), .ZN(n7648) );
  XNOR2_X1 U5127 ( .A(n5145), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U5128 ( .A1(n7069), .A2(n8979), .ZN(n6811) );
  BUF_X1 U5129 ( .A(n6017), .Z(n8616) );
  MUX2_X1 U5130 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5125), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5126) );
  AOI21_X1 U5131 ( .B1(n4653), .B2(n5342), .A(n4652), .ZN(n4651) );
  OAI21_X1 U5132 ( .B1(n5158), .B2(P1_IR_REG_20__SCAN_IN), .A(n4543), .ZN(
        n5143) );
  NAND2_X1 U5133 ( .A1(n5171), .A2(n5164), .ZN(n9688) );
  NAND2_X1 U5134 ( .A1(n5158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5140) );
  OR2_X1 U5135 ( .A1(n5127), .A2(n5453), .ZN(n5124) );
  NAND2_X2 U5136 ( .A1(n5167), .A2(n5166), .ZN(n5923) );
  AND2_X2 U5137 ( .A1(n6013), .A2(n6014), .ZN(n8619) );
  AOI21_X1 U5138 ( .B1(n5343), .B2(n4654), .A(n4542), .ZN(n4653) );
  MUX2_X1 U5139 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5165), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5167) );
  MUX2_X1 U5140 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6010), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6013) );
  XNOR2_X1 U5141 ( .A(n5206), .B(n5188), .ZN(n5205) );
  NOR2_X1 U5142 ( .A1(n5374), .A2(n5135), .ZN(n4749) );
  NAND3_X1 U5143 ( .A1(n5094), .A2(n4907), .A3(n5123), .ZN(n5164) );
  NAND2_X1 U5144 ( .A1(n4751), .A2(n4750), .ZN(n5374) );
  AND2_X1 U5145 ( .A1(n5121), .A2(n5095), .ZN(n5094) );
  NAND2_X2 U5146 ( .A1(n6468), .A2(P2_U3152), .ZN(n6488) );
  NOR2_X1 U5147 ( .A1(n5136), .A2(n5120), .ZN(n5121) );
  INV_X2 U5148 ( .A(n5320), .ZN(n4479) );
  INV_X1 U5149 ( .A(n6040), .ZN(n6468) );
  AND2_X1 U5150 ( .A1(n6108), .A2(n4973), .ZN(n4875) );
  AND4_X1 U5151 ( .A1(n10247), .A2(n10479), .A3(n5114), .A4(n5619), .ZN(n5115)
         );
  AND2_X2 U5152 ( .A1(n6067), .A2(n5988), .ZN(n6108) );
  AND2_X1 U5153 ( .A1(n5989), .A2(n4971), .ZN(n4973) );
  AND4_X1 U5154 ( .A1(n5113), .A2(n5530), .A3(n5622), .A4(n5112), .ZN(n5116)
         );
  AND4_X1 U5155 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n4487)
         );
  AND2_X1 U5156 ( .A1(n5990), .A2(n5991), .ZN(n5063) );
  INV_X1 U5157 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6163) );
  INV_X1 U5158 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10454) );
  INV_X1 U5159 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5619) );
  INV_X1 U5160 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6286) );
  NOR2_X1 U5161 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5113) );
  NOR2_X2 U5162 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6067) );
  INV_X1 U5163 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9129) );
  INV_X4 U5164 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5165 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10479) );
  INV_X1 U5166 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4725) );
  NOR2_X2 U5167 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5210) );
  NOR2_X1 U5168 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5983) );
  NOR2_X1 U5169 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5984) );
  NOR2_X1 U5170 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5985) );
  NOR2_X1 U5171 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5986) );
  BUF_X2 U5172 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9960) );
  INV_X1 U5173 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5989) );
  NOR2_X1 U5174 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5988) );
  NOR2_X1 U5175 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5987) );
  INV_X1 U5176 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10247) );
  NOR2_X1 U5177 ( .A1(n6803), .A2(n6852), .ZN(n6819) );
  NAND4_X2 U5178 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n6803)
         );
  NAND3_X1 U5179 ( .A1(n5185), .A2(n5184), .A3(n5183), .ZN(n6802) );
  INV_X1 U5180 ( .A(n6818), .ZN(n8995) );
  NAND2_X1 U5181 ( .A1(n6020), .A2(n8619), .ZN(n4481) );
  NAND2_X4 U5182 ( .A1(n6020), .A2(n8619), .ZN(n6274) );
  AND3_X2 U5183 ( .A1(n5210), .A2(n4695), .A3(n4725), .ZN(n5263) );
  AND2_X1 U5184 ( .A1(n5106), .A2(n4664), .ZN(n4663) );
  NAND2_X1 U5185 ( .A1(n5502), .A2(n5501), .ZN(n4664) );
  OR2_X1 U5186 ( .A1(n8540), .A2(n8285), .ZN(n7990) );
  OAI22_X1 U5187 ( .A1(n9261), .A2(n5951), .B1(n9279), .B2(n5882), .ZN(n5837)
         );
  OR2_X1 U5188 ( .A1(n9501), .A2(n9168), .ZN(n9221) );
  NAND2_X1 U5189 ( .A1(n4688), .A2(n4693), .ZN(n5789) );
  NAND2_X1 U5190 ( .A1(n4676), .A2(n4672), .ZN(n5723) );
  INV_X1 U5191 ( .A(n4673), .ZN(n4672) );
  OAI21_X1 U5192 ( .B1(n4675), .B2(n4674), .A(n5692), .ZN(n4673) );
  NAND2_X1 U5193 ( .A1(n4596), .A2(n4508), .ZN(n4764) );
  NOR2_X1 U5194 ( .A1(n9163), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U5195 ( .A1(n5070), .A2(n9164), .ZN(n5069) );
  NAND2_X1 U5196 ( .A1(n9261), .A2(n9279), .ZN(n4825) );
  AOI21_X1 U5197 ( .B1(n4682), .B2(n5646), .A(n5668), .ZN(n4681) );
  OAI21_X1 U5198 ( .B1(n8190), .B2(n4893), .A(n7856), .ZN(n4892) );
  NAND2_X1 U5199 ( .A1(n4520), .A2(n4893), .ZN(n4891) );
  INV_X1 U5200 ( .A(n8619), .ZN(n6018) );
  OR2_X1 U5201 ( .A1(n7680), .A2(n7677), .ZN(n7736) );
  OR2_X1 U5202 ( .A1(n8517), .A2(n8218), .ZN(n7845) );
  NOR2_X1 U5203 ( .A1(n8523), .A2(n8529), .ZN(n4772) );
  NAND2_X1 U5204 ( .A1(n8339), .A2(n8359), .ZN(n4627) );
  OR2_X1 U5205 ( .A1(n8549), .A2(n8359), .ZN(n7841) );
  OR2_X1 U5206 ( .A1(n10072), .A2(n8075), .ZN(n7941) );
  NOR2_X1 U5207 ( .A1(n10055), .A2(n7463), .ZN(n4638) );
  NAND2_X1 U5208 ( .A1(n8083), .A2(n7041), .ZN(n7902) );
  AND2_X1 U5209 ( .A1(n5041), .A2(n8032), .ZN(n4613) );
  NAND2_X1 U5210 ( .A1(n4478), .A2(n6902), .ZN(n5041) );
  INV_X1 U5211 ( .A(n6086), .ZN(n6115) );
  NAND2_X1 U5212 ( .A1(n8459), .A2(n8197), .ZN(n4635) );
  NAND2_X1 U5213 ( .A1(n5051), .A2(n5053), .ZN(n5047) );
  AND2_X1 U5214 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  OR2_X1 U5215 ( .A1(n9287), .A2(n5951), .ZN(n5805) );
  AND2_X1 U5216 ( .A1(n8674), .A2(n8700), .ZN(n5030) );
  INV_X1 U5217 ( .A(n5080), .ZN(n5078) );
  INV_X1 U5218 ( .A(n9253), .ZN(n4936) );
  NAND2_X1 U5219 ( .A1(n9517), .A2(n9294), .ZN(n8941) );
  OR2_X1 U5220 ( .A1(n9532), .A2(n9160), .ZN(n8987) );
  OR2_X1 U5221 ( .A1(n8969), .A2(n5909), .ZN(n7504) );
  NAND2_X1 U5222 ( .A1(n5867), .A2(n5866), .ZN(n5944) );
  NAND2_X1 U5223 ( .A1(n5011), .A2(n5009), .ZN(n5867) );
  AOI21_X1 U5224 ( .B1(n5012), .B2(n4566), .A(n5010), .ZN(n5009) );
  AND2_X1 U5225 ( .A1(n5724), .A2(n5699), .ZN(n5722) );
  AOI21_X1 U5226 ( .B1(n4658), .B2(n4661), .A(n5003), .ZN(n4655) );
  NOR2_X1 U5227 ( .A1(n5587), .A2(n5006), .ZN(n5005) );
  INV_X1 U5228 ( .A(n5554), .ZN(n5006) );
  NOR2_X1 U5229 ( .A1(n6422), .A2(n4970), .ZN(n4969) );
  INV_X1 U5230 ( .A(n6419), .ZN(n4970) );
  OAI21_X1 U5231 ( .B1(n8019), .B2(n8018), .A(n8023), .ZN(n8025) );
  INV_X1 U5232 ( .A(n6085), .ZN(n4828) );
  NAND2_X1 U5233 ( .A1(n4828), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6091) );
  INV_X1 U5234 ( .A(n8090), .ZN(n4763) );
  INV_X1 U5235 ( .A(n4609), .ZN(n4608) );
  OAI21_X1 U5236 ( .B1(n5055), .B2(n8234), .A(n8219), .ZN(n4609) );
  INV_X1 U5237 ( .A(n7998), .ZN(n4859) );
  NAND2_X1 U5238 ( .A1(n8529), .A2(n8286), .ZN(n7998) );
  XNOR2_X1 U5239 ( .A(n8523), .B(n8241), .ZN(n8256) );
  INV_X1 U5240 ( .A(n4623), .ZN(n4622) );
  AND2_X1 U5241 ( .A1(n4620), .A2(n8326), .ZN(n4619) );
  NAND2_X1 U5242 ( .A1(n4623), .A2(n4621), .ZN(n4620) );
  INV_X1 U5243 ( .A(n4624), .ZN(n4621) );
  AND2_X1 U5244 ( .A1(n7960), .A2(n7962), .ZN(n8430) );
  INV_X2 U5245 ( .A(n6059), .ZN(n6404) );
  NAND2_X1 U5246 ( .A1(n7600), .A2(n7599), .ZN(n8540) );
  NAND2_X1 U5247 ( .A1(n5811), .A2(n5787), .ZN(n8637) );
  INV_X1 U5248 ( .A(n5099), .ZN(n4745) );
  INV_X1 U5249 ( .A(n8655), .ZN(n4746) );
  NOR2_X1 U5250 ( .A1(n5026), .A2(n4531), .ZN(n5025) );
  INV_X1 U5251 ( .A(n5028), .ZN(n5026) );
  AND2_X1 U5252 ( .A1(n6808), .A2(n6721), .ZN(n6676) );
  INV_X1 U5253 ( .A(n9055), .ZN(n4649) );
  AND2_X1 U5254 ( .A1(n5858), .A2(n5857), .ZN(n9167) );
  OR2_X1 U5255 ( .A1(n8753), .A2(n5852), .ZN(n5858) );
  NAND2_X1 U5256 ( .A1(n8776), .A2(n8775), .ZN(n9492) );
  NOR2_X1 U5257 ( .A1(n9166), .A2(n4823), .ZN(n4822) );
  INV_X1 U5258 ( .A(n5102), .ZN(n4823) );
  AND2_X1 U5259 ( .A1(n5759), .A2(n5758), .ZN(n9325) );
  NAND2_X1 U5260 ( .A1(n4790), .A2(n4486), .ZN(n5088) );
  NAND2_X1 U5261 ( .A1(n7104), .A2(n7103), .ZN(n4898) );
  INV_X1 U5262 ( .A(n9632), .ZN(n9871) );
  NOR2_X1 U5263 ( .A1(n9491), .A2(n4899), .ZN(n4699) );
  AND2_X1 U5264 ( .A1(n9492), .A2(n9647), .ZN(n4899) );
  NAND2_X1 U5265 ( .A1(n5947), .A2(n5946), .ZN(n9495) );
  NAND2_X1 U5266 ( .A1(n4692), .A2(n5763), .ZN(n5772) );
  XNOR2_X1 U5267 ( .A(n5156), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9063) );
  INV_X1 U5268 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5111) );
  INV_X1 U5269 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4788) );
  AOI21_X1 U5270 ( .B1(n9231), .B2(n9840), .A(n9230), .ZN(n9498) );
  NAND2_X1 U5271 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U5272 ( .A1(n5081), .A2(n5080), .ZN(n9214) );
  NAND2_X1 U5273 ( .A1(n5079), .A2(n9197), .ZN(n4783) );
  NAND2_X1 U5274 ( .A1(n5081), .A2(n5083), .ZN(n5079) );
  MUX2_X1 U5275 ( .A(n7883), .B(n7882), .S(n8017), .Z(n7897) );
  MUX2_X1 U5276 ( .A(n7934), .B(n7933), .S(n8017), .Z(n7939) );
  INV_X1 U5277 ( .A(n4846), .ZN(n4842) );
  NAND2_X1 U5278 ( .A1(n7955), .A2(n7954), .ZN(n4845) );
  NAND2_X1 U5279 ( .A1(n9042), .A2(n8971), .ZN(n4669) );
  AND2_X1 U5280 ( .A1(n5063), .A2(n4980), .ZN(n5062) );
  NAND2_X1 U5281 ( .A1(n5764), .A2(n5763), .ZN(n4694) );
  NOR2_X1 U5282 ( .A1(n5135), .A2(n5141), .ZN(n5039) );
  INV_X1 U5283 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U5284 ( .A1(n5555), .A2(n5008), .ZN(n5007) );
  INV_X1 U5285 ( .A(n5527), .ZN(n5008) );
  INV_X1 U5286 ( .A(n5552), .ZN(n5555) );
  NAND2_X1 U5287 ( .A1(n4965), .A2(n4963), .ZN(n4962) );
  INV_X1 U5288 ( .A(n6246), .ZN(n4963) );
  NAND2_X1 U5289 ( .A1(n5000), .A2(n4998), .ZN(n8021) );
  NOR2_X1 U5290 ( .A1(n7874), .A2(n4999), .ZN(n4998) );
  INV_X1 U5291 ( .A(n7868), .ZN(n4999) );
  NAND2_X1 U5292 ( .A1(n8021), .A2(n8013), .ZN(n8059) );
  OR2_X1 U5293 ( .A1(n8183), .A2(n8071), .ZN(n8011) );
  OR2_X1 U5294 ( .A1(n8535), .A2(n8212), .ZN(n7995) );
  NOR2_X1 U5295 ( .A1(n8265), .A2(n8264), .ZN(n7844) );
  NAND2_X1 U5296 ( .A1(n7995), .A2(n7993), .ZN(n8211) );
  NAND2_X1 U5297 ( .A1(n4619), .A2(n4622), .ZN(n4616) );
  NOR2_X1 U5298 ( .A1(n8555), .A2(n8560), .ZN(n4776) );
  INV_X1 U5299 ( .A(n8356), .ZN(n4600) );
  OR2_X1 U5300 ( .A1(n8560), .A2(n8392), .ZN(n7978) );
  NAND2_X1 U5301 ( .A1(n4872), .A2(n4873), .ZN(n4870) );
  NAND2_X1 U5302 ( .A1(n4874), .A2(n4872), .ZN(n4871) );
  NOR2_X1 U5303 ( .A1(n8590), .A2(n8585), .ZN(n4779) );
  NOR2_X1 U5304 ( .A1(n7940), .A2(n4884), .ZN(n4883) );
  INV_X1 U5305 ( .A(n7938), .ZN(n4884) );
  INV_X1 U5306 ( .A(n7913), .ZN(n4863) );
  AND2_X1 U5307 ( .A1(n8307), .A2(n8293), .ZN(n8271) );
  NOR2_X1 U5308 ( .A1(n8320), .A2(n8540), .ZN(n8307) );
  NAND2_X1 U5309 ( .A1(n7958), .A2(n7956), .ZN(n8443) );
  MUX2_X1 U5310 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6037), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6039) );
  AND2_X1 U5311 ( .A1(n5063), .A2(n4973), .ZN(n4972) );
  AOI21_X1 U5312 ( .B1(n4506), .B2(n5099), .A(n4568), .ZN(n4747) );
  OR2_X1 U5313 ( .A1(n9505), .A2(n9167), .ZN(n9196) );
  OR2_X1 U5314 ( .A1(n9517), .A2(n9294), .ZN(n8942) );
  OR2_X1 U5315 ( .A1(n9525), .A2(n9325), .ZN(n9191) );
  NOR3_X1 U5316 ( .A1(n9328), .A2(n4925), .A3(n4517), .ZN(n4924) );
  OR2_X1 U5317 ( .A1(n9537), .A2(n9324), .ZN(n9189) );
  NAND2_X1 U5318 ( .A1(n4931), .A2(n9187), .ZN(n4930) );
  INV_X1 U5319 ( .A(n9354), .ZN(n4931) );
  NAND2_X1 U5320 ( .A1(n4905), .A2(n4903), .ZN(n4902) );
  INV_X1 U5321 ( .A(n9178), .ZN(n4903) );
  NOR2_X1 U5322 ( .A1(n9436), .A2(n4906), .ZN(n4905) );
  INV_X1 U5323 ( .A(n9179), .ZN(n4906) );
  NAND2_X1 U5324 ( .A1(n5334), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5359) );
  INV_X1 U5325 ( .A(n5336), .ZN(n5334) );
  AND2_X1 U5326 ( .A1(n9063), .A2(n9327), .ZN(n5917) );
  XNOR2_X1 U5327 ( .A(n7860), .B(n7859), .ZN(n7857) );
  NAND2_X1 U5328 ( .A1(n4992), .A2(n4991), .ZN(n7853) );
  AOI21_X1 U5329 ( .B1(n4994), .B2(n4996), .A(n4591), .ZN(n4991) );
  NAND2_X1 U5330 ( .A1(n5944), .A2(n4994), .ZN(n4992) );
  NOR2_X1 U5331 ( .A1(n4687), .A2(n5815), .ZN(n4684) );
  AOI21_X1 U5332 ( .B1(n4693), .B2(n4690), .A(n5017), .ZN(n4689) );
  INV_X1 U5333 ( .A(n5763), .ZN(n4690) );
  INV_X1 U5334 ( .A(n4689), .ZN(n4687) );
  NOR2_X1 U5335 ( .A1(n4693), .A2(n5815), .ZN(n4686) );
  NAND2_X1 U5336 ( .A1(n5743), .A2(n5742), .ZN(n5765) );
  INV_X1 U5337 ( .A(n4681), .ZN(n4680) );
  AOI21_X1 U5338 ( .B1(n4681), .B2(n4679), .A(n4580), .ZN(n4678) );
  INV_X1 U5339 ( .A(n5646), .ZN(n4679) );
  AND2_X1 U5340 ( .A1(n5616), .A2(n5592), .ZN(n5614) );
  NAND2_X1 U5341 ( .A1(n5586), .A2(n5560), .ZN(n5587) );
  NAND2_X1 U5342 ( .A1(n4657), .A2(n4663), .ZN(n5528) );
  AOI21_X1 U5343 ( .B1(n5105), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5344 ( .A(n5451), .ZN(n4989) );
  NAND2_X1 U5345 ( .A1(n4800), .A2(n4804), .ZN(n5422) );
  NAND2_X1 U5346 ( .A1(n5390), .A2(n5373), .ZN(n5391) );
  AOI21_X1 U5347 ( .B1(n4949), .B2(n7811), .A(n4571), .ZN(n4948) );
  NAND2_X1 U5348 ( .A1(n4960), .A2(n4959), .ZN(n4958) );
  INV_X1 U5349 ( .A(n6071), .ZN(n4959) );
  AOI21_X1 U5350 ( .B1(n4948), .B2(n4950), .A(n4946), .ZN(n4945) );
  INV_X1 U5351 ( .A(n7726), .ZN(n4946) );
  INV_X1 U5352 ( .A(n4948), .ZN(n4947) );
  AND2_X1 U5353 ( .A1(n8024), .A2(n8275), .ZN(n8066) );
  INV_X1 U5354 ( .A(n6780), .ZN(n4952) );
  INV_X1 U5355 ( .A(n6134), .ZN(n4979) );
  INV_X1 U5356 ( .A(n6131), .ZN(n4976) );
  INV_X1 U5357 ( .A(n6154), .ZN(n4975) );
  NAND2_X1 U5358 ( .A1(n7709), .A2(n4969), .ZN(n7750) );
  AOI21_X1 U5359 ( .B1(n4524), .B2(n4894), .A(n4890), .ZN(n4889) );
  AOI21_X1 U5360 ( .B1(n8235), .B2(n7742), .A(n7685), .ZN(n8218) );
  NAND2_X1 U5361 ( .A1(n7737), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n4827) );
  AND4_X1 U5362 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n7077)
         );
  OR2_X1 U5363 ( .A1(n7223), .A2(n4525), .ZN(n4757) );
  NAND2_X1 U5364 ( .A1(n4757), .A2(n4756), .ZN(n4599) );
  INV_X1 U5365 ( .A(n7125), .ZN(n4756) );
  OR2_X1 U5366 ( .A1(n7188), .A2(n7187), .ZN(n4596) );
  AND2_X1 U5367 ( .A1(n8093), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4762) );
  NOR2_X1 U5368 ( .A1(n8190), .A2(n8226), .ZN(n8189) );
  NAND2_X1 U5369 ( .A1(n8238), .A2(n8221), .ZN(n4607) );
  NAND2_X1 U5370 ( .A1(n4608), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U5371 ( .A1(n8234), .A2(n7848), .ZN(n4604) );
  INV_X1 U5372 ( .A(n5056), .ZN(n5055) );
  OAI21_X1 U5373 ( .B1(n8256), .B2(n5057), .A(n8217), .ZN(n5056) );
  INV_X1 U5374 ( .A(n8215), .ZN(n5057) );
  NOR2_X1 U5375 ( .A1(n8256), .A2(n8267), .ZN(n5059) );
  NAND2_X1 U5376 ( .A1(n8296), .A2(n8210), .ZN(n8281) );
  NAND2_X1 U5377 ( .A1(n6662), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7601) );
  INV_X1 U5378 ( .A(n6663), .ZN(n6662) );
  NAND2_X1 U5379 ( .A1(n8543), .A2(n8346), .ZN(n8302) );
  AND2_X1 U5380 ( .A1(n4627), .A2(n4628), .ZN(n4624) );
  NAND2_X1 U5381 ( .A1(n4552), .A2(n4627), .ZN(n4623) );
  NAND2_X1 U5382 ( .A1(n4628), .A2(n8208), .ZN(n4626) );
  NAND2_X1 U5383 ( .A1(n7985), .A2(n8302), .ZN(n8326) );
  NAND2_X1 U5384 ( .A1(n7841), .A2(n7974), .ZN(n8343) );
  NOR2_X1 U5385 ( .A1(n8366), .A2(n8345), .ZN(n8208) );
  NAND2_X1 U5386 ( .A1(n8366), .A2(n8345), .ZN(n4628) );
  NOR2_X1 U5387 ( .A1(n8393), .A2(n8560), .ZN(n8370) );
  AOI21_X1 U5388 ( .B1(n8402), .B2(n8202), .A(n8201), .ZN(n8385) );
  NOR2_X1 U5389 ( .A1(n8200), .A2(n8570), .ZN(n8201) );
  OAI21_X1 U5390 ( .B1(n8441), .B2(n4869), .A(n7960), .ZN(n4868) );
  INV_X1 U5391 ( .A(n4874), .ZN(n4869) );
  NAND2_X1 U5392 ( .A1(n4867), .A2(n4870), .ZN(n8409) );
  CLKBUF_X1 U5393 ( .A(n8428), .Z(n8441) );
  AOI21_X1 U5394 ( .B1(n4633), .B2(n8467), .A(n4551), .ZN(n4632) );
  NAND2_X1 U5395 ( .A1(n4635), .A2(n4633), .ZN(n8440) );
  NAND2_X1 U5396 ( .A1(n8481), .A2(n4779), .ZN(n8460) );
  OR2_X1 U5397 ( .A1(n8590), .A2(n8470), .ZN(n8195) );
  OAI21_X1 U5398 ( .B1(n7395), .B2(n4639), .A(n4547), .ZN(n7532) );
  NAND2_X1 U5399 ( .A1(n4642), .A2(n4640), .ZN(n4639) );
  INV_X1 U5400 ( .A(n8043), .ZN(n4640) );
  AND4_X1 U5401 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n8073)
         );
  NAND2_X1 U5402 ( .A1(n4550), .A2(n7936), .ZN(n4882) );
  INV_X1 U5403 ( .A(n7941), .ZN(n4885) );
  NAND2_X1 U5404 ( .A1(n7478), .A2(n4883), .ZN(n4881) );
  INV_X1 U5405 ( .A(n8045), .ZN(n7475) );
  AND2_X1 U5406 ( .A1(n7941), .A2(n7936), .ZN(n8045) );
  OAI21_X1 U5407 ( .B1(n7395), .B2(n8043), .A(n4636), .ZN(n7396) );
  INV_X1 U5408 ( .A(n4638), .ZN(n4636) );
  NAND2_X1 U5409 ( .A1(n7396), .A2(n7399), .ZN(n7474) );
  NAND2_X1 U5410 ( .A1(n8082), .A2(n6989), .ZN(n5052) );
  NAND2_X1 U5411 ( .A1(n7917), .A2(n7918), .ZN(n8040) );
  AOI21_X1 U5412 ( .B1(n8030), .B2(n4614), .A(n4539), .ZN(n4612) );
  NAND2_X1 U5413 ( .A1(n4613), .A2(n5042), .ZN(n6987) );
  NAND2_X1 U5414 ( .A1(n6886), .A2(n6885), .ZN(n6887) );
  NAND2_X1 U5415 ( .A1(n6887), .A2(n8029), .ZN(n6900) );
  AND2_X1 U5416 ( .A1(n8027), .A2(n7876), .ZN(n8486) );
  NAND2_X1 U5417 ( .A1(n7597), .A2(n7596), .ZN(n8523) );
  INV_X1 U5418 ( .A(n6904), .ZN(n10023) );
  AND3_X1 U5419 ( .A1(n4875), .A2(n4475), .A3(n4487), .ZN(n6029) );
  NAND2_X1 U5420 ( .A1(n8674), .A2(n5029), .ZN(n5028) );
  INV_X1 U5421 ( .A(n5814), .ZN(n5029) );
  AND2_X1 U5422 ( .A1(n5814), .A2(n5810), .ZN(n8700) );
  AOI21_X1 U5423 ( .B1(n5033), .B2(n7514), .A(n4538), .ZN(n5031) );
  AOI21_X1 U5424 ( .B1(n4740), .B2(n4742), .A(n4739), .ZN(n4738) );
  INV_X1 U5425 ( .A(n7427), .ZN(n4739) );
  AND2_X1 U5426 ( .A1(n5880), .A2(n5879), .ZN(n9168) );
  AND2_X1 U5427 ( .A1(n5929), .A2(n5957), .ZN(n9217) );
  INV_X1 U5428 ( .A(n4812), .ZN(n4811) );
  OAI21_X1 U5429 ( .B1(n4814), .B2(n4507), .A(n5082), .ZN(n4812) );
  NAND2_X1 U5430 ( .A1(n4541), .A2(n8984), .ZN(n4938) );
  XNOR2_X1 U5431 ( .A(n9505), .B(n9167), .ZN(n9253) );
  AOI21_X1 U5432 ( .B1(n4822), .B2(n9165), .A(n4496), .ZN(n4821) );
  INV_X1 U5433 ( .A(n9313), .ZN(n9280) );
  NAND2_X1 U5434 ( .A1(n9328), .A2(n5072), .ZN(n5071) );
  AND2_X1 U5435 ( .A1(n9537), .A2(n9358), .ZN(n4807) );
  INV_X1 U5436 ( .A(n9189), .ZN(n4925) );
  NAND2_X1 U5437 ( .A1(n9356), .A2(n4928), .ZN(n4926) );
  NOR2_X1 U5438 ( .A1(n4579), .A2(n5092), .ZN(n5091) );
  NAND2_X1 U5439 ( .A1(n9650), .A2(n9449), .ZN(n5089) );
  NAND3_X1 U5440 ( .A1(n9145), .A2(n9144), .A3(n4495), .ZN(n4790) );
  NAND2_X1 U5441 ( .A1(n9444), .A2(n9178), .ZN(n9441) );
  NOR2_X1 U5442 ( .A1(n8999), .A2(n4897), .ZN(n4896) );
  INV_X1 U5443 ( .A(n8806), .ZN(n4897) );
  INV_X1 U5444 ( .A(n9074), .ZN(n9868) );
  AND2_X1 U5445 ( .A1(n6817), .A2(n9060), .ZN(n9632) );
  AND2_X1 U5446 ( .A1(n6817), .A2(n5923), .ZN(n9635) );
  NAND2_X1 U5447 ( .A1(n5874), .A2(n5873), .ZN(n9501) );
  INV_X1 U5448 ( .A(n9251), .ZN(n9505) );
  NAND2_X1 U5449 ( .A1(n5676), .A2(n5675), .ZN(n9542) );
  INV_X1 U5450 ( .A(n5169), .ZN(n5168) );
  NOR2_X1 U5451 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5098) );
  XNOR2_X1 U5452 ( .A(n5865), .B(n5864), .ZN(n7643) );
  OAI21_X1 U5453 ( .B1(n5789), .B2(n4566), .A(n5012), .ZN(n5865) );
  XNOR2_X1 U5454 ( .A(n5841), .B(n5840), .ZN(n7631) );
  NAND2_X1 U5455 ( .A1(n5015), .A2(n5818), .ZN(n5841) );
  NAND2_X1 U5456 ( .A1(n5789), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U5457 ( .A1(n4997), .A2(n5724), .ZN(n5739) );
  NAND2_X1 U5458 ( .A1(n4749), .A2(n5040), .ZN(n5158) );
  INV_X1 U5459 ( .A(SI_7_), .ZN(n5346) );
  INV_X1 U5460 ( .A(n5318), .ZN(n4654) );
  NOR2_X1 U5461 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4695) );
  XNOR2_X1 U5462 ( .A(n5238), .B(n5209), .ZN(n5236) );
  INV_X1 U5463 ( .A(SI_2_), .ZN(n5209) );
  AND2_X1 U5464 ( .A1(n7654), .A2(n7653), .ZN(n8286) );
  AND4_X1 U5465 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n8492)
         );
  INV_X1 U5466 ( .A(n8324), .ZN(n8543) );
  NAND2_X1 U5467 ( .A1(n6406), .A2(n6405), .ZN(n8567) );
  NAND3_X2 U5468 ( .A1(n6041), .A2(n6042), .A3(n4861), .ZN(n6769) );
  OR2_X1 U5469 ( .A1(n6149), .A2(n6482), .ZN(n4861) );
  INV_X1 U5470 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5471 ( .B1(n4969), .B2(n4968), .A(n7748), .ZN(n4967) );
  INV_X1 U5472 ( .A(n7606), .ZN(n4968) );
  AND4_X1 U5473 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n7548)
         );
  OR2_X1 U5474 ( .A1(n7781), .A2(n7778), .ZN(n4595) );
  AND4_X1 U5475 ( .A1(n6298), .A2(n6297), .A3(n6296), .A4(n6295), .ZN(n8435)
         );
  INV_X1 U5476 ( .A(n8378), .ZN(n8412) );
  NAND2_X1 U5477 ( .A1(n8028), .A2(n8027), .ZN(n4984) );
  OR2_X1 U5478 ( .A1(n8025), .A2(n4983), .ZN(n4982) );
  OR2_X1 U5479 ( .A1(n8027), .A2(n8033), .ZN(n4983) );
  NAND2_X1 U5480 ( .A1(n7666), .A2(n7665), .ZN(n8241) );
  AND4_X1 U5481 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .ZN(n8075)
         );
  AND4_X1 U5482 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n7050)
         );
  NAND2_X1 U5483 ( .A1(n8328), .A2(n4565), .ZN(n8298) );
  NAND2_X1 U5484 ( .A1(n5775), .A2(n5774), .ZN(n9522) );
  NOR2_X1 U5485 ( .A1(n4498), .A2(n8749), .ZN(n4726) );
  INV_X1 U5486 ( .A(n9462), .ZN(n9143) );
  AND3_X1 U5487 ( .A1(n5731), .A2(n5730), .A3(n5729), .ZN(n9160) );
  NAND2_X1 U5488 ( .A1(n4748), .A2(n5024), .ZN(n5108) );
  NAND2_X1 U5489 ( .A1(n5762), .A2(n5761), .ZN(n8726) );
  INV_X1 U5490 ( .A(n9309), .ZN(n9525) );
  INV_X1 U5491 ( .A(n9073), .ZN(n8868) );
  AND2_X1 U5492 ( .A1(n5833), .A2(n5832), .ZN(n9279) );
  AND2_X1 U5493 ( .A1(n5911), .A2(n9847), .ZN(n8760) );
  AND2_X1 U5494 ( .A1(n5907), .A2(n6676), .ZN(n8751) );
  NOR2_X1 U5495 ( .A1(n7069), .A2(n4649), .ZN(n4648) );
  OR2_X1 U5496 ( .A1(n9058), .A2(n9057), .ZN(n4647) );
  INV_X1 U5497 ( .A(n4645), .ZN(n4644) );
  OAI21_X1 U5498 ( .B1(n9059), .B2(n5909), .A(n9061), .ZN(n4645) );
  INV_X1 U5499 ( .A(n9279), .ZN(n9254) );
  INV_X1 U5500 ( .A(n9492), .ZN(n9209) );
  INV_X1 U5501 ( .A(n5075), .ZN(n5074) );
  NAND2_X1 U5502 ( .A1(n4900), .A2(n9205), .ZN(n9491) );
  NAND2_X1 U5503 ( .A1(n4901), .A2(n9840), .ZN(n4900) );
  INV_X1 U5504 ( .A(n9501), .ZN(n9237) );
  INV_X1 U5505 ( .A(n9327), .ZN(n9863) );
  OR2_X1 U5506 ( .A1(n9376), .A2(n9934), .ZN(n9455) );
  NAND2_X1 U5507 ( .A1(n6810), .A2(n9847), .ZN(n9874) );
  INV_X1 U5508 ( .A(n9455), .ZN(n9833) );
  AND2_X1 U5509 ( .A1(n9497), .A2(n9498), .ZN(n4782) );
  OAI211_X1 U5510 ( .C1(n7897), .C2(n7885), .A(n7884), .B(n7913), .ZN(n7886)
         );
  OAI21_X1 U5511 ( .B1(n7907), .B2(n7906), .A(n7905), .ZN(n7909) );
  INV_X1 U5512 ( .A(n7919), .ZN(n4833) );
  AND2_X1 U5513 ( .A1(n7925), .A2(n7922), .ZN(n4838) );
  NAND2_X1 U5514 ( .A1(n4837), .A2(n7923), .ZN(n4836) );
  INV_X1 U5515 ( .A(n7925), .ZN(n4837) );
  NAND2_X1 U5516 ( .A1(n4834), .A2(n4835), .ZN(n7930) );
  NAND2_X1 U5517 ( .A1(n7920), .A2(n4832), .ZN(n4834) );
  AND2_X1 U5518 ( .A1(n7921), .A2(n4836), .ZN(n4835) );
  NOR2_X1 U5519 ( .A1(n4838), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5520 ( .A1(n8480), .A2(n7947), .ZN(n4846) );
  NOR2_X1 U5521 ( .A1(n4528), .A2(n4845), .ZN(n4843) );
  NAND2_X1 U5522 ( .A1(n4666), .A2(n8969), .ZN(n4665) );
  NAND2_X1 U5523 ( .A1(n4668), .A2(n8941), .ZN(n4667) );
  INV_X1 U5524 ( .A(n9194), .ZN(n4668) );
  OAI21_X1 U5525 ( .B1(n4830), .B2(n4829), .A(n4576), .ZN(n7981) );
  NAND2_X1 U5526 ( .A1(n7978), .A2(n7977), .ZN(n4829) );
  AOI21_X1 U5527 ( .B1(n7976), .B2(n8387), .A(n4831), .ZN(n4830) );
  AOI21_X1 U5528 ( .B1(n4851), .B2(n8000), .A(n7999), .ZN(n4849) );
  OAI21_X1 U5529 ( .B1(n7994), .B2(n4540), .A(n7996), .ZN(n4851) );
  NAND2_X1 U5530 ( .A1(n4852), .A2(n8000), .ZN(n4850) );
  AND2_X1 U5531 ( .A1(n4853), .A2(n7992), .ZN(n4852) );
  INV_X1 U5532 ( .A(n7994), .ZN(n4853) );
  INV_X1 U5533 ( .A(n5693), .ZN(n4677) );
  INV_X1 U5534 ( .A(n8012), .ZN(n4893) );
  OR2_X1 U5535 ( .A1(n8585), .A2(n8490), .ZN(n7953) );
  NAND2_X1 U5536 ( .A1(n7045), .A2(n7902), .ZN(n7883) );
  OR2_X1 U5537 ( .A1(n8580), .A2(n8435), .ZN(n7958) );
  NAND2_X1 U5538 ( .A1(n5050), .A2(n5051), .ZN(n5049) );
  INV_X1 U5539 ( .A(n5052), .ZN(n5050) );
  INV_X1 U5540 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5991) );
  INV_X1 U5541 ( .A(n8656), .ZN(n4744) );
  NOR2_X1 U5542 ( .A1(n4720), .A2(n5525), .ZN(n4713) );
  NAND2_X1 U5543 ( .A1(n4671), .A2(n4670), .ZN(n9042) );
  NAND2_X1 U5544 ( .A1(n8942), .A2(n8778), .ZN(n4671) );
  AND2_X1 U5545 ( .A1(n8941), .A2(n8983), .ZN(n4670) );
  OR2_X1 U5546 ( .A1(n9495), .A2(n9203), .ZN(n8961) );
  NOR2_X1 U5547 ( .A1(n9517), .A2(n9522), .ZN(n4704) );
  OAI21_X1 U5548 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(n7860) );
  INV_X1 U5549 ( .A(n4995), .ZN(n4994) );
  OAI21_X1 U5550 ( .B1(n5943), .B2(n4996), .A(n7585), .ZN(n4995) );
  INV_X1 U5551 ( .A(n5945), .ZN(n4996) );
  NOR2_X1 U5552 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n4491), .ZN(n4908) );
  INV_X1 U5553 ( .A(n5864), .ZN(n5010) );
  INV_X1 U5554 ( .A(n4678), .ZN(n4675) );
  NAND2_X1 U5555 ( .A1(n4680), .A2(n4677), .ZN(n4674) );
  AND2_X1 U5556 ( .A1(n4659), .A2(n4556), .ZN(n4658) );
  NAND2_X1 U5557 ( .A1(n4663), .A2(n4660), .ZN(n4659) );
  INV_X1 U5558 ( .A(n5501), .ZN(n4660) );
  INV_X1 U5559 ( .A(n4663), .ZN(n4661) );
  NAND2_X1 U5560 ( .A1(n5391), .A2(n5390), .ZN(n4806) );
  NAND2_X1 U5561 ( .A1(n5425), .A2(n5424), .ZN(n5451) );
  INV_X1 U5562 ( .A(n5365), .ZN(n4652) );
  INV_X1 U5563 ( .A(n8022), .ZN(n4890) );
  NOR2_X1 U5564 ( .A1(n4520), .A2(n7856), .ZN(n4894) );
  NOR2_X1 U5565 ( .A1(n8155), .A2(n4752), .ZN(n8165) );
  AND2_X1 U5566 ( .A1(n8156), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4752) );
  OR2_X1 U5567 ( .A1(n8529), .A2(n8286), .ZN(n7996) );
  NAND2_X1 U5568 ( .A1(n4776), .A2(n8339), .ZN(n4775) );
  OR2_X1 U5569 ( .A1(n8555), .A2(n8345), .ZN(n7980) );
  NAND2_X1 U5570 ( .A1(n4642), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U5571 ( .A1(n5061), .A2(n7531), .ZN(n4641) );
  AND2_X1 U5572 ( .A1(n7399), .A2(n7531), .ZN(n4642) );
  NAND2_X1 U5573 ( .A1(n6218), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6239) );
  INV_X1 U5574 ( .A(n6220), .ZN(n6218) );
  INV_X1 U5575 ( .A(n7883), .ZN(n7904) );
  INV_X1 U5576 ( .A(n6986), .ZN(n4614) );
  OR2_X1 U5577 ( .A1(n7484), .A2(n7483), .ZN(n7485) );
  AND2_X1 U5578 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  OAI21_X1 U5579 ( .B1(n5034), .B2(n4742), .A(n7428), .ZN(n4741) );
  INV_X1 U5580 ( .A(n5419), .ZN(n4742) );
  NAND2_X1 U5581 ( .A1(n4712), .A2(n4711), .ZN(n4719) );
  NAND2_X1 U5582 ( .A1(n4484), .A2(n5582), .ZN(n4711) );
  AOI21_X1 U5583 ( .B1(n4484), .B2(n4714), .A(n4713), .ZN(n4712) );
  NOR2_X1 U5584 ( .A1(n4720), .A2(n5033), .ZN(n4714) );
  INV_X1 U5585 ( .A(n4721), .ZN(n4717) );
  OR2_X1 U5586 ( .A1(n5928), .A2(n5927), .ZN(n5957) );
  NAND2_X1 U5587 ( .A1(n9501), .A2(n9168), .ZN(n8958) );
  NAND2_X1 U5588 ( .A1(n4704), .A2(n9261), .ZN(n4703) );
  INV_X1 U5589 ( .A(n4825), .ZN(n4816) );
  INV_X1 U5590 ( .A(n4821), .ZN(n4820) );
  NAND2_X1 U5591 ( .A1(n4815), .A2(n4825), .ZN(n4814) );
  INV_X1 U5592 ( .A(n4818), .ZN(n4815) );
  AOI21_X1 U5593 ( .B1(n4821), .B2(n4819), .A(n9013), .ZN(n4818) );
  INV_X1 U5594 ( .A(n4822), .ZN(n4819) );
  AND2_X1 U5595 ( .A1(n4920), .A2(n4558), .ZN(n4919) );
  NAND2_X1 U5596 ( .A1(n4924), .A2(n9190), .ZN(n4920) );
  INV_X1 U5597 ( .A(n9311), .ZN(n4927) );
  INV_X1 U5598 ( .A(n4924), .ZN(n4921) );
  INV_X1 U5599 ( .A(n5071), .ZN(n5070) );
  NOR2_X1 U5600 ( .A1(n5068), .A2(n5100), .ZN(n5067) );
  INV_X1 U5601 ( .A(n9164), .ZN(n5068) );
  NAND2_X1 U5602 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  INV_X1 U5603 ( .A(n4710), .ZN(n4708) );
  INV_X1 U5604 ( .A(n9154), .ZN(n5092) );
  OR2_X1 U5605 ( .A1(n9555), .A2(n9561), .ZN(n4710) );
  INV_X1 U5606 ( .A(n9148), .ZN(n5090) );
  NAND2_X1 U5607 ( .A1(n5541), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5565) );
  OR2_X1 U5608 ( .A1(n5513), .A2(n5512), .ZN(n5542) );
  AND2_X1 U5609 ( .A1(n9831), .A2(n4522), .ZN(n4696) );
  INV_X1 U5610 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U5611 ( .A1(n5358), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5403) );
  INV_X1 U5612 ( .A(n5359), .ZN(n5358) );
  NAND2_X1 U5613 ( .A1(n5308), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U5614 ( .A1(n6861), .A2(n6860), .ZN(n8802) );
  NOR2_X1 U5615 ( .A1(n9305), .A2(n4702), .ZN(n9281) );
  INV_X1 U5616 ( .A(n4704), .ZN(n4702) );
  NOR2_X1 U5617 ( .A1(n9305), .A2(n9522), .ZN(n9295) );
  NAND2_X1 U5618 ( .A1(n9171), .A2(n4913), .ZN(n4912) );
  AND2_X1 U5619 ( .A1(n4911), .A2(n9172), .ZN(n4910) );
  INV_X1 U5620 ( .A(n5818), .ZN(n5014) );
  INV_X1 U5621 ( .A(n5013), .ZN(n5012) );
  OAI21_X1 U5622 ( .B1(n5016), .B2(n4566), .A(n5839), .ZN(n5013) );
  NOR2_X1 U5623 ( .A1(n5819), .A2(n5017), .ZN(n5016) );
  NOR2_X1 U5624 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5095) );
  NOR2_X1 U5625 ( .A1(n5374), .A2(n5038), .ZN(n5142) );
  NAND2_X1 U5626 ( .A1(n5040), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5627 ( .A1(n5723), .A2(n5722), .ZN(n4997) );
  INV_X1 U5628 ( .A(n5643), .ZN(n4682) );
  XNOR2_X1 U5629 ( .A(n5553), .B(n10248), .ZN(n5552) );
  NAND2_X1 U5630 ( .A1(n5501), .A2(n5480), .ZN(n5502) );
  AOI21_X1 U5631 ( .B1(n4493), .B2(n4799), .A(n4549), .ZN(n4985) );
  INV_X1 U5632 ( .A(n5428), .ZN(n5431) );
  NOR2_X1 U5633 ( .A1(n4798), .A2(n5105), .ZN(n4797) );
  AOI21_X1 U5634 ( .B1(n4804), .B2(n4802), .A(n4990), .ZN(n4801) );
  INV_X1 U5635 ( .A(n5390), .ZN(n4802) );
  INV_X1 U5636 ( .A(n4801), .ZN(n4798) );
  NOR2_X1 U5637 ( .A1(n4804), .A2(n5105), .ZN(n4796) );
  INV_X1 U5638 ( .A(SI_5_), .ZN(n10357) );
  INV_X1 U5639 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5110) );
  MUX2_X1 U5640 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5320), .Z(n5238) );
  INV_X1 U5641 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4785) );
  INV_X1 U5642 ( .A(n4965), .ZN(n4964) );
  NAND3_X1 U5643 ( .A1(n4954), .A2(n4956), .A3(n6746), .ZN(n4953) );
  INV_X1 U5644 ( .A(n6712), .ZN(n4956) );
  INV_X1 U5645 ( .A(n4958), .ZN(n4951) );
  OR2_X1 U5646 ( .A1(n10008), .A2(n6032), .ZN(n7877) );
  OR2_X1 U5647 ( .A1(n6239), .A2(n10485), .ZN(n6255) );
  OR2_X1 U5648 ( .A1(n6255), .A2(n7286), .ZN(n6272) );
  NAND2_X1 U5649 ( .A1(n7544), .A2(n6246), .ZN(n7553) );
  AND3_X1 U5650 ( .A1(n8063), .A2(n8062), .A3(n8061), .ZN(n5104) );
  AND3_X1 U5651 ( .A1(n7640), .A2(n7639), .A3(n7638), .ZN(n8212) );
  AND4_X1 U5652 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n7379)
         );
  OR2_X1 U5653 ( .A1(n4481), .A2(n7133), .ZN(n4610) );
  NOR2_X1 U5654 ( .A1(n6452), .A2(n4769), .ZN(n7119) );
  NAND2_X1 U5655 ( .A1(n9960), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U5656 ( .A1(n4597), .A2(n7122), .ZN(n4759) );
  INV_X1 U5657 ( .A(n7146), .ZN(n4597) );
  NOR2_X1 U5658 ( .A1(n7328), .A2(n4768), .ZN(n7284) );
  NOR2_X1 U5659 ( .A1(n7276), .A2(n7481), .ZN(n4768) );
  NAND2_X1 U5660 ( .A1(n7352), .A2(n4767), .ZN(n7354) );
  OR2_X1 U5661 ( .A1(n7353), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4767) );
  OR2_X1 U5662 ( .A1(n8134), .A2(n4755), .ZN(n4754) );
  AND2_X1 U5663 ( .A1(n8135), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U5664 ( .A1(n8613), .A2(n6185), .ZN(n5000) );
  NAND2_X1 U5665 ( .A1(n8271), .A2(n4577), .ZN(n8226) );
  NAND2_X1 U5666 ( .A1(n7855), .A2(n7854), .ZN(n8190) );
  AOI21_X1 U5667 ( .B1(n8239), .B2(n8234), .A(n8005), .ZN(n8220) );
  AND2_X1 U5668 ( .A1(n7736), .A2(n7681), .ZN(n8235) );
  NAND2_X1 U5669 ( .A1(n8271), .A2(n8182), .ZN(n8272) );
  NAND2_X1 U5670 ( .A1(n8271), .A2(n4772), .ZN(n8250) );
  INV_X1 U5671 ( .A(n8256), .ZN(n8249) );
  AND3_X1 U5672 ( .A1(n7605), .A2(n7604), .A3(n7603), .ZN(n8285) );
  INV_X1 U5673 ( .A(n8211), .ZN(n8283) );
  AND2_X1 U5674 ( .A1(n8301), .A2(n8302), .ZN(n7842) );
  NAND2_X1 U5675 ( .A1(n4617), .A2(n4536), .ZN(n8296) );
  AND2_X1 U5676 ( .A1(n7990), .A2(n7989), .ZN(n8301) );
  NOR2_X1 U5677 ( .A1(n8393), .A2(n4774), .ZN(n8360) );
  INV_X1 U5678 ( .A(n4776), .ZN(n4774) );
  INV_X1 U5679 ( .A(n8317), .ZN(n8359) );
  NAND2_X1 U5680 ( .A1(n7978), .A2(n7979), .ZN(n8376) );
  OR2_X1 U5681 ( .A1(n8567), .A2(n8378), .ZN(n8203) );
  OR2_X1 U5682 ( .A1(n6407), .A2(n10426), .ZN(n6425) );
  AND4_X1 U5683 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n8392)
         );
  NOR2_X1 U5684 ( .A1(n4866), .A2(n8384), .ZN(n4865) );
  NAND2_X1 U5685 ( .A1(n4870), .A2(n8387), .ZN(n4866) );
  AOI21_X1 U5686 ( .B1(n4632), .B2(n4634), .A(n4573), .ZN(n4631) );
  AND2_X1 U5687 ( .A1(n8481), .A2(n4778), .ZN(n8421) );
  AND2_X1 U5688 ( .A1(n4492), .A2(n8422), .ZN(n4778) );
  NAND2_X1 U5689 ( .A1(n8481), .A2(n4492), .ZN(n8438) );
  NAND2_X1 U5690 ( .A1(n4488), .A2(n4879), .ZN(n4876) );
  NAND2_X1 U5691 ( .A1(n7478), .A2(n7938), .ZN(n4886) );
  INV_X1 U5692 ( .A(n8078), .ZN(n7463) );
  OR2_X1 U5693 ( .A1(n6202), .A2(n10470), .ZN(n6220) );
  NAND2_X1 U5694 ( .A1(n6177), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6202) );
  INV_X1 U5695 ( .A(n6179), .ZN(n6177) );
  AND2_X1 U5696 ( .A1(n7300), .A2(n7370), .ZN(n7384) );
  AOI21_X1 U5697 ( .B1(n7298), .B2(n8041), .A(n7297), .ZN(n7299) );
  NOR2_X1 U5698 ( .A1(n7236), .A2(n7924), .ZN(n7300) );
  INV_X1 U5699 ( .A(n7917), .ZN(n4864) );
  OR2_X1 U5700 ( .A1(n7018), .A2(n10033), .ZN(n7236) );
  NOR2_X1 U5701 ( .A1(n6931), .A2(n6904), .ZN(n7042) );
  AND4_X1 U5702 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n6988)
         );
  INV_X1 U5703 ( .A(n6899), .ZN(n5046) );
  NOR2_X1 U5704 ( .A1(n6769), .A2(n6768), .ZN(n6889) );
  NAND2_X1 U5705 ( .A1(n6871), .A2(n7888), .ZN(n6764) );
  NAND2_X1 U5706 ( .A1(n6764), .A2(n6760), .ZN(n6886) );
  NAND2_X1 U5707 ( .A1(n6384), .A2(n6383), .ZN(n8560) );
  INV_X1 U5708 ( .A(n10065), .ZN(n10074) );
  OR2_X1 U5709 ( .A1(n10008), .A2(n8033), .ZN(n10065) );
  INV_X1 U5710 ( .A(n10063), .ZN(n10073) );
  AND2_X1 U5711 ( .A1(n7559), .A2(n6341), .ZN(n9995) );
  AND2_X1 U5712 ( .A1(n4560), .A2(n5996), .ZN(n4629) );
  CLKBUF_X1 U5713 ( .A(n6368), .Z(n6454) );
  XNOR2_X1 U5714 ( .A(n6035), .B(n6034), .ZN(n7567) );
  NAND2_X1 U5715 ( .A1(n6033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6035) );
  XNOR2_X1 U5716 ( .A(n4981), .B(n4980), .ZN(n8062) );
  OR2_X1 U5717 ( .A1(n6025), .A2(n6195), .ZN(n4981) );
  INV_X1 U5718 ( .A(n6025), .ZN(n6027) );
  OR2_X1 U5719 ( .A1(n6166), .A2(n6165), .ZN(n6186) );
  AND2_X1 U5720 ( .A1(n8710), .A2(n5691), .ZN(n8647) );
  AND2_X1 U5721 ( .A1(n5030), .A2(n8748), .ZN(n4729) );
  NOR2_X1 U5722 ( .A1(n7083), .A2(n7084), .ZN(n4734) );
  NAND2_X1 U5723 ( .A1(n7083), .A2(n7084), .ZN(n4735) );
  NOR2_X1 U5724 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  INV_X1 U5725 ( .A(n7056), .ZN(n4733) );
  NAND2_X1 U5726 ( .A1(n5486), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5513) );
  INV_X1 U5727 ( .A(n5488), .ZN(n5486) );
  OR2_X1 U5728 ( .A1(n5565), .A2(n5564), .ZN(n5598) );
  NAND2_X1 U5729 ( .A1(n5597), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5628) );
  INV_X1 U5730 ( .A(n5598), .ZN(n5597) );
  NAND2_X1 U5731 ( .A1(n5793), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5826) );
  INV_X1 U5732 ( .A(n5795), .ZN(n5793) );
  OR2_X1 U5733 ( .A1(n5752), .A2(n8729), .ZN(n5778) );
  OR2_X1 U5734 ( .A1(n5436), .A2(n5435), .ZN(n5459) );
  NAND2_X1 U5735 ( .A1(n5457), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5488) );
  INV_X1 U5736 ( .A(n5459), .ZN(n5457) );
  INV_X1 U5737 ( .A(n5642), .ZN(n4730) );
  NAND2_X1 U5738 ( .A1(n8692), .A2(n5642), .ZN(n5667) );
  CLKBUF_X1 U5739 ( .A(n5348), .Z(n5982) );
  NOR2_X1 U5740 ( .A1(n5078), .A2(n4507), .ZN(n5076) );
  OAI21_X1 U5741 ( .B1(n5078), .B2(n5082), .A(n5077), .ZN(n5075) );
  AOI21_X1 U5742 ( .B1(n5080), .B2(n9235), .A(n4537), .ZN(n5077) );
  XNOR2_X1 U5743 ( .A(n9200), .B(n9199), .ZN(n4901) );
  NOR2_X2 U5744 ( .A1(n9248), .A2(n9501), .ZN(n9241) );
  AND2_X1 U5745 ( .A1(n9222), .A2(n5083), .ZN(n5080) );
  NAND2_X1 U5746 ( .A1(n9237), .A2(n9168), .ZN(n5083) );
  AOI21_X1 U5747 ( .B1(n4934), .B2(n4940), .A(n4933), .ZN(n4932) );
  INV_X1 U5748 ( .A(n9196), .ZN(n4933) );
  INV_X1 U5749 ( .A(n8941), .ZN(n9262) );
  AND2_X1 U5750 ( .A1(n9189), .A2(n8988), .ZN(n9342) );
  AND2_X1 U5751 ( .A1(n9548), .A2(n9389), .ZN(n4809) );
  OR2_X1 U5752 ( .A1(n5628), .A2(n5627), .ZN(n5655) );
  AND2_X1 U5753 ( .A1(n9187), .A2(n8990), .ZN(n9366) );
  AND2_X1 U5754 ( .A1(n5107), .A2(n5089), .ZN(n5087) );
  INV_X1 U5755 ( .A(n4905), .ZN(n4904) );
  OR2_X1 U5756 ( .A1(n9450), .A2(n9150), .ZN(n9428) );
  AND3_X1 U5757 ( .A1(n4696), .A2(n9668), .A3(n9663), .ZN(n9465) );
  NAND2_X1 U5758 ( .A1(n9831), .A2(n4522), .ZN(n9625) );
  NOR2_X1 U5759 ( .A1(n4494), .A2(n5085), .ZN(n5084) );
  INV_X1 U5760 ( .A(n7446), .ZN(n5085) );
  NAND2_X1 U5761 ( .A1(n9831), .A2(n9933), .ZN(n9830) );
  NAND2_X1 U5762 ( .A1(n4916), .A2(n8809), .ZN(n9835) );
  NAND2_X1 U5763 ( .A1(n4917), .A2(n8895), .ZN(n4916) );
  INV_X1 U5764 ( .A(n7438), .ZN(n4917) );
  INV_X1 U5765 ( .A(n7315), .ZN(n7098) );
  AND2_X1 U5766 ( .A1(n8878), .A2(n8863), .ZN(n7315) );
  AND4_X1 U5767 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6945)
         );
  NAND2_X1 U5768 ( .A1(n4697), .A2(n9894), .ZN(n6963) );
  INV_X1 U5769 ( .A(n6961), .ZN(n4697) );
  NAND2_X1 U5770 ( .A1(n8799), .A2(n8800), .ZN(n6857) );
  NAND2_X1 U5771 ( .A1(n5825), .A2(n5824), .ZN(n9511) );
  AND2_X1 U5772 ( .A1(n6813), .A2(n7069), .ZN(n9856) );
  AND2_X1 U5773 ( .A1(n6813), .A2(n5886), .ZN(n9647) );
  INV_X1 U5774 ( .A(n7440), .ZN(n9927) );
  XNOR2_X1 U5775 ( .A(n7853), .B(n7591), .ZN(n8774) );
  XNOR2_X1 U5776 ( .A(n7586), .B(n7585), .ZN(n7719) );
  NAND2_X1 U5777 ( .A1(n4993), .A2(n5945), .ZN(n7586) );
  XNOR2_X1 U5778 ( .A(n5944), .B(n5943), .ZN(n7595) );
  OAI211_X1 U5779 ( .C1(n5765), .C2(n4509), .A(n4685), .B(n4683), .ZN(n7598)
         );
  OAI22_X1 U5780 ( .A1(n4687), .A2(n4686), .B1(n5815), .B2(n4689), .ZN(n4685)
         );
  OAI21_X1 U5781 ( .B1(n5647), .B2(n4680), .A(n4678), .ZN(n5694) );
  NAND2_X1 U5782 ( .A1(n5002), .A2(n5586), .ZN(n5615) );
  NAND2_X1 U5783 ( .A1(n5001), .A2(n5005), .ZN(n5002) );
  NAND2_X1 U5784 ( .A1(n5001), .A2(n5554), .ZN(n5588) );
  AND2_X1 U5785 ( .A1(n5508), .A2(n5483), .ZN(n9094) );
  NAND2_X1 U5786 ( .A1(n4987), .A2(n4988), .ZN(n5475) );
  NAND2_X1 U5787 ( .A1(n4803), .A2(n5390), .ZN(n5420) );
  NAND2_X1 U5788 ( .A1(n5319), .A2(n5318), .ZN(n5344) );
  XNOR2_X1 U5789 ( .A(n5289), .B(n5261), .ZN(n5287) );
  XNOR2_X1 U5790 ( .A(n5258), .B(n5241), .ZN(n5256) );
  INV_X1 U5791 ( .A(SI_3_), .ZN(n5241) );
  AND4_X1 U5792 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n7295)
         );
  NAND2_X1 U5793 ( .A1(n6974), .A2(n4978), .ZN(n7073) );
  NAND2_X1 U5794 ( .A1(n6974), .A2(n6134), .ZN(n7031) );
  NAND2_X1 U5795 ( .A1(n4944), .A2(n4948), .ZN(n7727) );
  AND2_X1 U5796 ( .A1(n6201), .A2(n6200), .ZN(n10055) );
  NAND2_X1 U5797 ( .A1(n4957), .A2(n4958), .ZN(n6747) );
  OR2_X1 U5798 ( .A1(n6713), .A2(n6712), .ZN(n4957) );
  AOI21_X1 U5799 ( .B1(n4945), .B2(n4947), .A(n4578), .ZN(n4943) );
  OAI21_X1 U5800 ( .B1(n7812), .B2(n4947), .A(n4945), .ZN(n7734) );
  INV_X1 U5801 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U5802 ( .A1(n7633), .A2(n7632), .ZN(n8535) );
  NAND2_X1 U5803 ( .A1(n4955), .A2(n4953), .ZN(n6782) );
  AOI21_X1 U5804 ( .B1(n4978), .B2(n4976), .A(n4975), .ZN(n4974) );
  INV_X1 U5805 ( .A(n4978), .ZN(n4977) );
  NAND2_X1 U5806 ( .A1(n7709), .A2(n6419), .ZN(n6421) );
  NAND2_X1 U5807 ( .A1(n7553), .A2(n4965), .ZN(n7690) );
  NAND2_X1 U5808 ( .A1(n7616), .A2(n7615), .ZN(n8549) );
  OAI211_X1 U5809 ( .C1(n6149), .C2(n6472), .A(n6070), .B(n6069), .ZN(n6869)
         );
  AND2_X1 U5810 ( .A1(n6685), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7805) );
  INV_X1 U5811 ( .A(n7745), .ZN(n7830) );
  OR2_X1 U5812 ( .A1(n6697), .A2(n8434), .ZN(n7829) );
  NAND2_X1 U5813 ( .A1(n6403), .A2(n7796), .ZN(n7800) );
  NAND2_X1 U5814 ( .A1(n6438), .A2(n6131), .ZN(n6974) );
  INV_X1 U5815 ( .A(n7805), .ZN(n7828) );
  AND2_X1 U5816 ( .A1(n4827), .A2(n4826), .ZN(n6665) );
  INV_X1 U5817 ( .A(n7295), .ZN(n8080) );
  INV_X1 U5818 ( .A(n7077), .ZN(n8081) );
  INV_X1 U5819 ( .A(n6988), .ZN(n8083) );
  OR2_X1 U5820 ( .A1(n6086), .A2(n6049), .ZN(n6053) );
  AOI21_X1 U5821 ( .B1(n9607), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9603), .ZN(
        n7148) );
  AND2_X1 U5822 ( .A1(n4759), .A2(n4758), .ZN(n7223) );
  INV_X1 U5823 ( .A(n7224), .ZN(n4758) );
  INV_X1 U5824 ( .A(n4759), .ZN(n7225) );
  INV_X1 U5825 ( .A(n4599), .ZN(n7159) );
  INV_X1 U5826 ( .A(n4757), .ZN(n7126) );
  NAND2_X1 U5827 ( .A1(n7173), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4598) );
  AOI21_X1 U5828 ( .B1(n7213), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7210), .ZN(
        n7188) );
  INV_X1 U5829 ( .A(n4596), .ZN(n7186) );
  INV_X1 U5830 ( .A(n4764), .ZN(n8091) );
  INV_X1 U5831 ( .A(n7165), .ZN(n4760) );
  INV_X1 U5832 ( .A(n4761), .ZN(n7166) );
  AND2_X1 U5833 ( .A1(n4754), .A2(n4753), .ZN(n8155) );
  INV_X1 U5834 ( .A(n8137), .ZN(n4753) );
  INV_X1 U5835 ( .A(n4754), .ZN(n8138) );
  OAI21_X1 U5836 ( .B1(n8221), .B2(n4608), .A(n4603), .ZN(n4602) );
  NAND2_X1 U5837 ( .A1(n5058), .A2(n4497), .ZN(n4605) );
  NAND2_X1 U5838 ( .A1(n8243), .A2(n8242), .ZN(n8244) );
  XNOR2_X1 U5839 ( .A(n8233), .B(n8234), .ZN(n8522) );
  NAND2_X1 U5840 ( .A1(n8266), .A2(n7998), .ZN(n8255) );
  INV_X1 U5841 ( .A(n8535), .ZN(n8293) );
  AND2_X1 U5842 ( .A1(n7623), .A2(n7622), .ZN(n8324) );
  OR2_X1 U5843 ( .A1(n8353), .A2(n4622), .ZN(n4615) );
  NAND2_X1 U5844 ( .A1(n4618), .A2(n4623), .ZN(n8327) );
  NAND2_X1 U5845 ( .A1(n8353), .A2(n4624), .ZN(n4618) );
  NAND2_X1 U5846 ( .A1(n4625), .A2(n4628), .ZN(n8333) );
  OR2_X1 U5847 ( .A1(n8353), .A2(n8208), .ZN(n4625) );
  INV_X1 U5848 ( .A(n4868), .ZN(n8411) );
  NAND2_X1 U5849 ( .A1(n8440), .A2(n4513), .ZN(n8420) );
  NAND2_X1 U5850 ( .A1(n8481), .A2(n8485), .ZN(n8462) );
  NAND2_X1 U5851 ( .A1(n9993), .A2(n9974), .ZN(n9988) );
  NAND2_X1 U5852 ( .A1(n8194), .A2(n4515), .ZN(n8479) );
  NAND2_X1 U5853 ( .A1(n4881), .A2(n4882), .ZN(n7528) );
  NAND2_X1 U5854 ( .A1(n7474), .A2(n4514), .ZN(n7476) );
  NAND2_X1 U5855 ( .A1(n5048), .A2(n5051), .ZN(n7239) );
  NAND2_X1 U5856 ( .A1(n7017), .A2(n5052), .ZN(n5048) );
  NAND2_X1 U5857 ( .A1(n7040), .A2(n8030), .ZN(n7039) );
  NAND2_X1 U5858 ( .A1(n6987), .A2(n6986), .ZN(n7040) );
  NAND2_X1 U5859 ( .A1(n6924), .A2(n8031), .ZN(n6923) );
  NAND2_X1 U5860 ( .A1(n6900), .A2(n6899), .ZN(n6924) );
  NAND2_X1 U5861 ( .A1(n9996), .A2(n6361), .ZN(n8451) );
  INV_X1 U5862 ( .A(n7385), .ZN(n8427) );
  INV_X1 U5863 ( .A(n8062), .ZN(n7890) );
  XNOR2_X1 U5864 ( .A(n6031), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9980) );
  OR3_X1 U5865 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9960), .ZN(n6078) );
  NAND2_X1 U5866 ( .A1(n9960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U5867 ( .A1(n7416), .A2(n5419), .ZN(n7430) );
  AND2_X1 U5868 ( .A1(n5976), .A2(n8751), .ZN(n5977) );
  INV_X1 U5869 ( .A(n5022), .ZN(n5020) );
  NOR2_X1 U5870 ( .A1(n8708), .A2(n5721), .ZN(n8657) );
  NOR2_X1 U5871 ( .A1(n8657), .A2(n8656), .ZN(n8655) );
  NAND2_X1 U5872 ( .A1(n7515), .A2(n5033), .ZN(n8664) );
  NAND2_X1 U5873 ( .A1(n8699), .A2(n5814), .ZN(n8672) );
  AND2_X1 U5874 ( .A1(n5027), .A2(n5028), .ZN(n8673) );
  NAND2_X1 U5875 ( .A1(n5036), .A2(n5307), .ZN(n7004) );
  AND2_X1 U5876 ( .A1(n5307), .A2(n5305), .ZN(n7005) );
  INV_X1 U5877 ( .A(n5037), .ZN(n5036) );
  NAND2_X1 U5878 ( .A1(n5035), .A2(n5389), .ZN(n7418) );
  NAND2_X1 U5879 ( .A1(n4724), .A2(n5033), .ZN(n4723) );
  INV_X1 U5880 ( .A(n9634), .ZN(n9448) );
  AND2_X1 U5881 ( .A1(n6676), .A2(n5936), .ZN(n8757) );
  NAND2_X1 U5882 ( .A1(n5027), .A2(n5025), .ZN(n8747) );
  INV_X1 U5883 ( .A(n8760), .ZN(n8770) );
  NAND4_X1 U5884 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n9073)
         );
  OR2_X1 U5885 ( .A1(n6580), .A2(n6579), .ZN(n6582) );
  NAND2_X1 U5886 ( .A1(n8850), .A2(n8849), .ZN(n9482) );
  NAND2_X1 U5887 ( .A1(n8840), .A2(n8839), .ZN(n9486) );
  NAND2_X1 U5888 ( .A1(n4937), .A2(n4938), .ZN(n9252) );
  NAND2_X1 U5889 ( .A1(n4941), .A2(n4939), .ZN(n4937) );
  AND2_X1 U5890 ( .A1(n5847), .A2(n5846), .ZN(n9251) );
  NAND2_X1 U5891 ( .A1(n4817), .A2(n4821), .ZN(n9260) );
  NAND2_X1 U5892 ( .A1(n9290), .A2(n4822), .ZN(n4817) );
  NAND2_X1 U5893 ( .A1(n4824), .A2(n5102), .ZN(n9275) );
  INV_X1 U5894 ( .A(n9522), .ZN(n9301) );
  AND2_X1 U5895 ( .A1(n5751), .A2(n5750), .ZN(n9309) );
  NAND2_X1 U5896 ( .A1(n9533), .A2(n5100), .ZN(n9304) );
  NAND2_X1 U5897 ( .A1(n4926), .A2(n4922), .ZN(n9322) );
  NAND2_X1 U5898 ( .A1(n5726), .A2(n5725), .ZN(n9532) );
  NAND2_X1 U5899 ( .A1(n5088), .A2(n5089), .ZN(n9408) );
  NAND2_X1 U5900 ( .A1(n9441), .A2(n9179), .ZN(n9424) );
  AND2_X1 U5901 ( .A1(n4790), .A2(n4791), .ZN(n9149) );
  NAND2_X1 U5902 ( .A1(n9474), .A2(n9146), .ZN(n9440) );
  NAND2_X1 U5903 ( .A1(n9145), .A2(n9144), .ZN(n9476) );
  NAND2_X1 U5904 ( .A1(n4909), .A2(n4913), .ZN(n9173) );
  NAND2_X1 U5905 ( .A1(n7438), .A2(n4915), .ZN(n4909) );
  NAND2_X1 U5906 ( .A1(n4898), .A2(n8806), .ZN(n7106) );
  INV_X1 U5907 ( .A(n9847), .ZN(n9861) );
  INV_X1 U5908 ( .A(n9845), .ZN(n9644) );
  AND2_X1 U5909 ( .A1(n4700), .A2(n4699), .ZN(n9493) );
  OR2_X1 U5910 ( .A1(n9490), .A2(n9934), .ZN(n4700) );
  AND2_X1 U5911 ( .A1(n5098), .A2(n5097), .ZN(n5096) );
  INV_X1 U5912 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5097) );
  INV_X1 U5913 ( .A(n5129), .ZN(n7593) );
  INV_X1 U5914 ( .A(n8979), .ZN(n9023) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6563) );
  INV_X1 U5916 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10239) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10476) );
  OAI21_X1 U5918 ( .B1(n5319), .B2(n5342), .A(n4653), .ZN(n5366) );
  OR2_X1 U5919 ( .A1(n5322), .A2(n4751), .ZN(n6576) );
  INV_X1 U5920 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5921 ( .A(n7050), .ZN(n8084) );
  NOR2_X1 U5922 ( .A1(n6498), .A2(P1_U3084), .ZN(P1_U4006) );
  OAI21_X1 U5923 ( .B1(n9237), .B2(n8760), .A(n5939), .ZN(n5940) );
  NAND2_X1 U5924 ( .A1(n4643), .A2(n9068), .ZN(P1_U3240) );
  NAND2_X1 U5925 ( .A1(n4646), .A2(n4644), .ZN(n4643) );
  NOR2_X1 U5926 ( .A1(n9498), .A2(n9640), .ZN(n9232) );
  NAND2_X1 U5927 ( .A1(n9573), .A2(n9906), .ZN(n4781) );
  INV_X1 U5928 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4780) );
  NAND2_X4 U5929 ( .A1(n4787), .A2(n4786), .ZN(n6040) );
  AND4_X1 U5931 ( .A1(n4487), .A2(n4475), .A3(n6108), .A4(n4972), .ZN(n6025)
         );
  INV_X1 U5932 ( .A(n5105), .ZN(n4799) );
  OR2_X1 U5933 ( .A1(n8585), .A2(n8196), .ZN(n4485) );
  AND2_X1 U5934 ( .A1(n4548), .A2(n4791), .ZN(n4486) );
  AND2_X2 U5935 ( .A1(n5130), .A2(n5129), .ZN(n5217) );
  INV_X1 U5936 ( .A(n8238), .ZN(n8234) );
  AND2_X1 U5937 ( .A1(n4887), .A2(n7945), .ZN(n4488) );
  INV_X1 U5938 ( .A(n6964), .ZN(n9894) );
  AND2_X1 U5939 ( .A1(n4941), .A2(n9012), .ZN(n4489) );
  OR2_X1 U5940 ( .A1(n7648), .A2(n6915), .ZN(n4490) );
  OR2_X1 U5941 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4491) );
  INV_X1 U5942 ( .A(n4748), .ZN(n5762) );
  AND2_X1 U5943 ( .A1(n4779), .A2(n8198), .ZN(n4492) );
  INV_X1 U5944 ( .A(n8984), .ZN(n9195) );
  OR2_X1 U5945 ( .A1(n9511), .A2(n9279), .ZN(n8984) );
  INV_X1 U5946 ( .A(n4634), .ZN(n4633) );
  NAND2_X1 U5947 ( .A1(n8443), .A2(n4485), .ZN(n4634) );
  AND2_X1 U5948 ( .A1(n4988), .A2(n5472), .ZN(n4493) );
  NAND2_X1 U5949 ( .A1(n9221), .A2(n8958), .ZN(n9238) );
  INV_X1 U5950 ( .A(n9238), .ZN(n9235) );
  NAND2_X1 U5951 ( .A1(n8691), .A2(n8693), .ZN(n8692) );
  NAND2_X1 U5952 ( .A1(n6314), .A2(n6313), .ZN(n8585) );
  OR2_X1 U5953 ( .A1(n8577), .A2(n8445), .ZN(n7960) );
  AND3_X1 U5954 ( .A1(n6128), .A2(n6127), .A3(n6126), .ZN(n10030) );
  AND2_X1 U5955 ( .A1(n5802), .A2(n5801), .ZN(n9294) );
  AND2_X1 U5956 ( .A1(n5064), .A2(n9147), .ZN(n4495) );
  AND2_X1 U5957 ( .A1(n9287), .A2(n9294), .ZN(n4496) );
  AND2_X1 U5958 ( .A1(n4608), .A2(n7848), .ZN(n4497) );
  INV_X1 U5959 ( .A(n5582), .ZN(n4720) );
  NOR2_X1 U5960 ( .A1(n5025), .A2(n4728), .ZN(n4498) );
  NAND2_X1 U5961 ( .A1(n9147), .A2(n4792), .ZN(n4791) );
  NAND2_X1 U5962 ( .A1(n5434), .A2(n5433), .ZN(n9140) );
  INV_X1 U5963 ( .A(n9140), .ZN(n4789) );
  AND2_X1 U5964 ( .A1(n4772), .A2(n4771), .ZN(n4499) );
  AND2_X1 U5965 ( .A1(n4860), .A2(n8070), .ZN(n4500) );
  AND2_X1 U5966 ( .A1(n8488), .A2(n4515), .ZN(n4501) );
  OR2_X1 U5967 ( .A1(n4534), .A2(n4734), .ZN(n4502) );
  AND2_X1 U5968 ( .A1(n8040), .A2(n5049), .ZN(n4503) );
  AND2_X1 U5969 ( .A1(n6002), .A2(n4895), .ZN(n4504) );
  AND2_X1 U5970 ( .A1(n8209), .A2(n4565), .ZN(n4505) );
  OR2_X1 U5971 ( .A1(n8727), .A2(n5024), .ZN(n4506) );
  AND2_X1 U5972 ( .A1(n9251), .A2(n9167), .ZN(n4507) );
  OR2_X1 U5973 ( .A1(n4766), .A2(n4765), .ZN(n4508) );
  OR2_X1 U5974 ( .A1(n4691), .A2(n5819), .ZN(n4509) );
  AND2_X1 U5975 ( .A1(n4886), .A2(n7935), .ZN(n4510) );
  AND2_X1 U5976 ( .A1(n9144), .A2(n5064), .ZN(n4511) );
  INV_X1 U5977 ( .A(n7069), .ZN(n5909) );
  NAND2_X1 U5978 ( .A1(n8070), .A2(n8068), .ZN(n4512) );
  OR2_X1 U5979 ( .A1(n8198), .A2(n8435), .ZN(n4513) );
  OR2_X1 U5980 ( .A1(n10064), .A2(n7548), .ZN(n4514) );
  OR2_X1 U5981 ( .A1(n9616), .A2(n8492), .ZN(n4515) );
  AND2_X1 U5982 ( .A1(n4761), .A2(n4760), .ZN(n4516) );
  AND2_X1 U5983 ( .A1(n5168), .A2(n5096), .ZN(n5127) );
  AND2_X1 U5984 ( .A1(n5348), .A2(n5320), .ZN(n5292) );
  AND2_X1 U5985 ( .A1(n4930), .A2(n4928), .ZN(n4517) );
  NAND2_X1 U5986 ( .A1(n6759), .A2(n6914), .ZN(n6871) );
  AND2_X1 U5987 ( .A1(n4926), .A2(n4924), .ZN(n4518) );
  NAND2_X1 U5988 ( .A1(n5150), .A2(n5122), .ZN(n5144) );
  AND2_X1 U5989 ( .A1(n8271), .A2(n4499), .ZN(n4519) );
  OR2_X1 U5990 ( .A1(n8190), .A2(n7872), .ZN(n4520) );
  INV_X1 U5991 ( .A(n5033), .ZN(n5032) );
  INV_X1 U5992 ( .A(n5342), .ZN(n5343) );
  XNOR2_X1 U5993 ( .A(n5345), .B(SI_6_), .ZN(n5342) );
  NAND2_X1 U5994 ( .A1(n4521), .A2(n4806), .ZN(n4805) );
  OAI211_X1 U5995 ( .C1(n5347), .C2(n6480), .A(n5267), .B(n5266), .ZN(n6952)
         );
  INV_X1 U5996 ( .A(n8410), .ZN(n4872) );
  AND2_X1 U5997 ( .A1(n5263), .A2(n5111), .ZN(n5294) );
  AND2_X1 U5998 ( .A1(n5421), .A2(n5396), .ZN(n4521) );
  AND2_X1 U5999 ( .A1(n9933), .A2(n4789), .ZN(n4522) );
  OAI211_X1 U6000 ( .C1(n5347), .C2(n6472), .A(n5216), .B(n5215), .ZN(n6855)
         );
  OR2_X1 U6001 ( .A1(n4820), .A2(n4816), .ZN(n4523) );
  INV_X1 U6002 ( .A(n9668), .ZN(n9643) );
  AND3_X1 U6003 ( .A1(n7873), .A2(n4892), .A3(n4891), .ZN(n4524) );
  NAND2_X1 U6004 ( .A1(n9140), .A2(n9837), .ZN(n9171) );
  AND2_X1 U6005 ( .A1(n7226), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U6006 ( .A1(n5626), .A2(n5625), .ZN(n9555) );
  AND2_X1 U6007 ( .A1(n4599), .A2(n4598), .ZN(n4526) );
  AND2_X1 U6008 ( .A1(n5996), .A2(n4504), .ZN(n4527) );
  XNOR2_X1 U6009 ( .A(n4743), .B(n6815), .ZN(n5274) );
  AND2_X1 U6010 ( .A1(n8467), .A2(n7951), .ZN(n4528) );
  AND2_X1 U6011 ( .A1(n7629), .A2(n4595), .ZN(n4529) );
  NAND2_X1 U6012 ( .A1(n8942), .A2(n8941), .ZN(n9277) );
  INV_X1 U6013 ( .A(n5586), .ZN(n5004) );
  AND3_X1 U6014 ( .A1(n7767), .A2(n7824), .A3(n7768), .ZN(n4530) );
  NOR2_X1 U6015 ( .A1(n5838), .A2(n5837), .ZN(n4531) );
  AND2_X1 U6016 ( .A1(n4488), .A2(n4883), .ZN(n4532) );
  XNOR2_X1 U6017 ( .A(n5473), .B(SI_11_), .ZN(n5472) );
  NAND2_X1 U6018 ( .A1(n8719), .A2(n8718), .ZN(n4533) );
  AND2_X1 U6019 ( .A1(n4735), .A2(n7057), .ZN(n4534) );
  INV_X1 U6020 ( .A(n4940), .ZN(n4939) );
  NAND2_X1 U6021 ( .A1(n9012), .A2(n8984), .ZN(n4940) );
  OR2_X1 U6022 ( .A1(n8570), .A2(n8433), .ZN(n8387) );
  INV_X1 U6023 ( .A(n8895), .ZN(n4918) );
  OR2_X1 U6024 ( .A1(n9548), .A2(n8782), .ZN(n9187) );
  INV_X1 U6025 ( .A(n6902), .ZN(n5045) );
  AND3_X1 U6026 ( .A1(n7984), .A2(n7983), .A3(n8054), .ZN(n4535) );
  AND2_X1 U6027 ( .A1(n4616), .A2(n4505), .ZN(n4536) );
  NAND2_X1 U6028 ( .A1(n4746), .A2(n4745), .ZN(n4748) );
  INV_X1 U6029 ( .A(n4805), .ZN(n4804) );
  AND2_X1 U6030 ( .A1(n9495), .A2(n9169), .ZN(n4537) );
  AND2_X1 U6031 ( .A1(n5500), .A2(n5499), .ZN(n4538) );
  XNOR2_X1 U6032 ( .A(n7865), .B(n7864), .ZN(n8613) );
  NAND2_X1 U6033 ( .A1(n5394), .A2(n10469), .ZN(n5421) );
  INV_X1 U6034 ( .A(n5421), .ZN(n4990) );
  AND2_X1 U6035 ( .A1(n6988), .A2(n7041), .ZN(n4539) );
  INV_X1 U6036 ( .A(n7238), .ZN(n5053) );
  INV_X1 U6037 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U6038 ( .A1(n4882), .A2(n4880), .ZN(n4879) );
  AND2_X1 U6039 ( .A1(n5137), .A2(n5138), .ZN(n5040) );
  AND2_X1 U6040 ( .A1(n8283), .A2(n7991), .ZN(n4540) );
  OR2_X1 U6041 ( .A1(n9262), .A2(n9263), .ZN(n4541) );
  AND2_X1 U6042 ( .A1(n5345), .A2(SI_6_), .ZN(n4542) );
  INV_X1 U6043 ( .A(n5525), .ZN(n4722) );
  AND2_X1 U6044 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4543) );
  AND2_X1 U6045 ( .A1(n5094), .A2(n5294), .ZN(n5150) );
  NAND2_X1 U6046 ( .A1(n6029), .A2(n5990), .ZN(n4544) );
  AND2_X1 U6047 ( .A1(n4669), .A2(n4665), .ZN(n4545) );
  NAND2_X1 U6048 ( .A1(n5428), .A2(n5137), .ZN(n4546) );
  AND2_X1 U6049 ( .A1(n4641), .A2(n4637), .ZN(n4547) );
  NOR2_X1 U6050 ( .A1(n9151), .A2(n5090), .ZN(n4548) );
  OR2_X1 U6051 ( .A1(n9356), .A2(n4930), .ZN(n4929) );
  INV_X1 U6052 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U6053 ( .A1(n4938), .A2(n4936), .ZN(n4935) );
  OAI21_X1 U6054 ( .B1(n5005), .B2(n5004), .A(n5614), .ZN(n5003) );
  AND2_X1 U6055 ( .A1(n5474), .A2(SI_11_), .ZN(n4549) );
  OR2_X1 U6056 ( .A1(n7477), .A2(n4885), .ZN(n4550) );
  NAND2_X1 U6057 ( .A1(n7049), .A2(n10030), .ZN(n5051) );
  NAND2_X1 U6058 ( .A1(n7837), .A2(n4513), .ZN(n4551) );
  INV_X1 U6059 ( .A(n5061), .ZN(n5060) );
  NAND2_X1 U6060 ( .A1(n7475), .A2(n4514), .ZN(n5061) );
  NAND2_X1 U6061 ( .A1(n8343), .A2(n4626), .ZN(n4552) );
  AND2_X1 U6062 ( .A1(n7929), .A2(n7928), .ZN(n4553) );
  AND2_X1 U6063 ( .A1(n6084), .A2(n6083), .ZN(n4554) );
  AND2_X1 U6064 ( .A1(n9180), .A2(n4902), .ZN(n4555) );
  AND2_X1 U6065 ( .A1(n5007), .A2(n5586), .ZN(n4556) );
  NAND2_X1 U6066 ( .A1(n7946), .A2(n7945), .ZN(n8047) );
  INV_X1 U6067 ( .A(n8047), .ZN(n4880) );
  NAND2_X1 U6068 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4557) );
  AND2_X1 U6069 ( .A1(n4927), .A2(n8986), .ZN(n4558) );
  OR2_X1 U6070 ( .A1(n8004), .A2(n8005), .ZN(n4559) );
  NOR2_X1 U6071 ( .A1(n5054), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4560) );
  INV_X1 U6072 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4980) );
  OR2_X1 U6073 ( .A1(n4523), .A2(n4507), .ZN(n4561) );
  OR2_X1 U6074 ( .A1(n4805), .A2(n4799), .ZN(n4562) );
  NAND2_X1 U6075 ( .A1(n4506), .A2(n4744), .ZN(n4563) );
  INV_X1 U6076 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4895) );
  OR2_X1 U6077 ( .A1(n8249), .A2(n4859), .ZN(n4564) );
  OR2_X1 U6078 ( .A1(n8324), .A2(n8346), .ZN(n4565) );
  OR2_X1 U6079 ( .A1(n5840), .A2(n5014), .ZN(n4566) );
  INV_X1 U6080 ( .A(n5761), .ZN(n5024) );
  NOR2_X1 U6081 ( .A1(n8738), .A2(n8737), .ZN(n8646) );
  NAND2_X1 U6082 ( .A1(n4511), .A2(n9145), .ZN(n9474) );
  NAND2_X1 U6083 ( .A1(n4615), .A2(n4619), .ZN(n8328) );
  AND2_X1 U6084 ( .A1(n9441), .A2(n4905), .ZN(n4567) );
  NAND2_X1 U6085 ( .A1(n5540), .A2(n5539), .ZN(n9150) );
  NAND2_X1 U6086 ( .A1(n4718), .A2(n4721), .ZN(n8626) );
  NAND2_X1 U6087 ( .A1(n5093), .A2(n9154), .ZN(n9379) );
  NAND2_X1 U6088 ( .A1(n4723), .A2(n5031), .ZN(n8717) );
  INV_X1 U6089 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U6090 ( .A1(n6291), .A2(n6290), .ZN(n8580) );
  INV_X1 U6091 ( .A(n8375), .ZN(n4831) );
  INV_X1 U6092 ( .A(n8748), .ZN(n4728) );
  NAND2_X1 U6093 ( .A1(n8011), .A2(n8012), .ZN(n8221) );
  NAND2_X1 U6094 ( .A1(n7721), .A2(n7720), .ZN(n8517) );
  INV_X1 U6095 ( .A(n8517), .ZN(n4771) );
  AND2_X1 U6096 ( .A1(n8727), .A2(n5024), .ZN(n4568) );
  NAND2_X1 U6097 ( .A1(n5585), .A2(n5584), .ZN(n8682) );
  AND2_X1 U6098 ( .A1(n9339), .A2(n9324), .ZN(n4569) );
  OR2_X1 U6099 ( .A1(n9409), .A2(n4706), .ZN(n4570) );
  NAND2_X1 U6100 ( .A1(n7996), .A2(n7998), .ZN(n8264) );
  NAND2_X1 U6101 ( .A1(n5294), .A2(n10261), .ZN(n5349) );
  INV_X1 U6102 ( .A(n5349), .ZN(n4751) );
  NAND2_X1 U6103 ( .A1(n8961), .A2(n9198), .ZN(n9222) );
  NAND2_X1 U6104 ( .A1(n7726), .A2(n7671), .ZN(n4571) );
  AND2_X1 U6105 ( .A1(n4881), .A2(n4878), .ZN(n4572) );
  NOR3_X1 U6106 ( .A1(n9305), .A2(n4703), .A3(n9505), .ZN(n4705) );
  AND4_X1 U6107 ( .A1(n6433), .A2(n6432), .A3(n6431), .A4(n6430), .ZN(n8345)
         );
  AND2_X1 U6108 ( .A1(n8422), .A2(n8445), .ZN(n4573) );
  INV_X1 U6109 ( .A(n4950), .ZN(n4949) );
  OAI21_X1 U6110 ( .B1(n7811), .B2(n7659), .A(n7673), .ZN(n4950) );
  NAND2_X1 U6111 ( .A1(n7645), .A2(n7644), .ZN(n8529) );
  AND2_X1 U6112 ( .A1(n7609), .A2(n7608), .ZN(n8366) );
  INV_X1 U6113 ( .A(n8366), .ZN(n8555) );
  NAND2_X1 U6114 ( .A1(n6398), .A2(n6397), .ZN(n8570) );
  OR2_X1 U6115 ( .A1(n9352), .A2(n9157), .ZN(n4574) );
  OR2_X1 U6116 ( .A1(n8395), .A2(n8412), .ZN(n4575) );
  NAND2_X1 U6117 ( .A1(n7847), .A2(n7846), .ZN(n8183) );
  INV_X1 U6118 ( .A(n4701), .ZN(n9268) );
  NOR2_X1 U6119 ( .A1(n9305), .A2(n4703), .ZN(n4701) );
  AND2_X1 U6120 ( .A1(n8342), .A2(n7979), .ZN(n4576) );
  AND2_X1 U6121 ( .A1(n4499), .A2(n8511), .ZN(n4577) );
  INV_X1 U6122 ( .A(n4693), .ZN(n4691) );
  AND2_X1 U6123 ( .A1(n5771), .A2(n4694), .ZN(n4693) );
  NOR2_X1 U6124 ( .A1(n7731), .A2(n7730), .ZN(n4578) );
  INV_X1 U6125 ( .A(n4709), .ZN(n9381) );
  NOR2_X1 U6126 ( .A1(n9409), .A2(n4710), .ZN(n4709) );
  INV_X1 U6127 ( .A(n4773), .ZN(n8334) );
  NOR2_X1 U6128 ( .A1(n8393), .A2(n4775), .ZN(n4773) );
  OAI21_X1 U6129 ( .B1(n8459), .B2(n4634), .A(n4632), .ZN(n8418) );
  AND4_X1 U6130 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n7049)
         );
  AND2_X1 U6131 ( .A1(n9555), .A2(n9403), .ZN(n4579) );
  AND2_X1 U6132 ( .A1(n5670), .A2(SI_18_), .ZN(n4580) );
  NAND2_X1 U6133 ( .A1(n9505), .A2(n9265), .ZN(n5082) );
  NAND2_X1 U6134 ( .A1(n6328), .A2(n6327), .ZN(n8577) );
  INV_X1 U6135 ( .A(n9287), .ZN(n9517) );
  AND2_X1 U6136 ( .A1(n5792), .A2(n5791), .ZN(n9287) );
  AND2_X1 U6137 ( .A1(n5740), .A2(n5724), .ZN(n4581) );
  AND2_X1 U6138 ( .A1(n4678), .A2(n4677), .ZN(n4582) );
  NOR2_X1 U6139 ( .A1(n5666), .A2(n4730), .ZN(n4583) );
  AND2_X1 U6140 ( .A1(n4635), .A2(n4485), .ZN(n4584) );
  AND2_X1 U6141 ( .A1(n7515), .A2(n5471), .ZN(n4585) );
  AND4_X1 U6142 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n8490)
         );
  NAND2_X1 U6143 ( .A1(n7532), .A2(n8047), .ZN(n8194) );
  OR2_X1 U6144 ( .A1(n5999), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4586) );
  AND2_X1 U6145 ( .A1(n4696), .A2(n9668), .ZN(n4587) );
  AND2_X1 U6146 ( .A1(n5307), .A2(n5037), .ZN(n7058) );
  OAI22_X1 U6147 ( .A1(n7017), .A2(n5047), .B1(n7238), .B2(n4503), .ZN(n7298)
         );
  NAND2_X1 U6148 ( .A1(n7023), .A2(n7913), .ZN(n7242) );
  NAND2_X1 U6149 ( .A1(n4736), .A2(n7057), .ZN(n7082) );
  NAND2_X1 U6150 ( .A1(n4731), .A2(n4502), .ZN(n7335) );
  AND2_X1 U6151 ( .A1(n9443), .A2(n8992), .ZN(n9475) );
  INV_X1 U6152 ( .A(n9475), .ZN(n5064) );
  NAND2_X1 U6153 ( .A1(n5652), .A2(n5651), .ZN(n9548) );
  INV_X1 U6154 ( .A(n9548), .ZN(n4707) );
  OR2_X1 U6155 ( .A1(n9906), .A2(n4780), .ZN(n4588) );
  NAND2_X1 U6156 ( .A1(n5035), .A2(n5034), .ZN(n7416) );
  AND2_X1 U6157 ( .A1(n4737), .A2(n4738), .ZN(n4589) );
  INV_X1 U6158 ( .A(n4589), .ZN(n4724) );
  NAND2_X1 U6159 ( .A1(n5086), .A2(n7446), .ZN(n7447) );
  NAND2_X1 U6160 ( .A1(n4589), .A2(n5468), .ZN(n7515) );
  INV_X1 U6161 ( .A(n5788), .ZN(n5017) );
  INV_X1 U6162 ( .A(n4915), .ZN(n4914) );
  NOR2_X1 U6163 ( .A1(n8810), .A2(n8894), .ZN(n4915) );
  OR2_X1 U6164 ( .A1(n7483), .A2(n7548), .ZN(n7935) );
  AND2_X1 U6165 ( .A1(n7474), .A2(n5060), .ZN(n4590) );
  AND2_X1 U6166 ( .A1(n7589), .A2(n7588), .ZN(n4591) );
  AND2_X1 U6167 ( .A1(n7553), .A2(n6250), .ZN(n4592) );
  INV_X1 U6168 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10261) );
  AND2_X1 U6169 ( .A1(n7877), .A2(n7876), .ZN(n4593) );
  NAND2_X1 U6170 ( .A1(n8070), .A2(n4593), .ZN(n4594) );
  INV_X1 U6171 ( .A(n7189), .ZN(n4766) );
  INV_X1 U6172 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n4765) );
  INV_X1 U6173 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4784) );
  INV_X1 U6174 ( .A(n8469), .ZN(n8491) );
  INV_X2 U6175 ( .A(n9597), .ZN(n9595) );
  AOI21_X2 U6177 ( .B1(n7788), .B2(n7787), .A(n7620), .ZN(n7626) );
  NAND2_X2 U6178 ( .A1(n7800), .A2(n6415), .ZN(n7709) );
  NAND2_X1 U6179 ( .A1(n5116), .A2(n5115), .ZN(n5136) );
  OAI21_X1 U6180 ( .B1(n6438), .B2(n4977), .A(n4974), .ZN(n6175) );
  NOR2_X1 U6181 ( .A1(n9333), .A2(n4807), .ZN(n9159) );
  NAND2_X1 U6182 ( .A1(n6693), .A2(n6692), .ZN(n6691) );
  NAND2_X1 U6183 ( .A1(n4781), .A2(n4588), .ZN(P1_U3519) );
  OAI21_X2 U6184 ( .B1(n9624), .B2(n9668), .A(n9143), .ZN(n9145) );
  NOR2_X1 U6185 ( .A1(n9365), .A2(n4809), .ZN(n9348) );
  INV_X1 U6186 ( .A(n5065), .ZN(n9290) );
  NAND2_X1 U6187 ( .A1(n7284), .A2(n7283), .ZN(n7352) );
  NOR2_X1 U6188 ( .A1(n7330), .A2(n7329), .ZN(n7328) );
  NOR2_X1 U6189 ( .A1(n8120), .A2(n8119), .ZN(n8134) );
  XNOR2_X2 U6190 ( .A(n6068), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U6191 ( .A1(n8341), .A2(n5101), .ZN(n8314) );
  INV_X1 U6192 ( .A(n8357), .ZN(n4601) );
  NAND2_X1 U6193 ( .A1(n5422), .A2(n4493), .ZN(n4986) );
  INV_X1 U6194 ( .A(n8488), .ZN(n4887) );
  NAND2_X1 U6195 ( .A1(n5528), .A2(n5527), .ZN(n5556) );
  NAND2_X1 U6196 ( .A1(n4877), .A2(n4876), .ZN(n8487) );
  NAND2_X2 U6197 ( .A1(n5369), .A2(n5368), .ZN(n5392) );
  OR2_X1 U6198 ( .A1(n5058), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U6199 ( .A1(n5058), .A2(n5055), .ZN(n8233) );
  NAND3_X1 U6200 ( .A1(n4606), .A2(n4605), .A3(n4602), .ZN(n8510) );
  NAND2_X1 U6201 ( .A1(n4611), .A2(n4612), .ZN(n7017) );
  NAND3_X1 U6202 ( .A1(n8030), .A2(n4613), .A3(n5042), .ZN(n4611) );
  NAND2_X1 U6203 ( .A1(n8353), .A2(n4619), .ZN(n4617) );
  NAND2_X1 U6204 ( .A1(n5997), .A2(n4629), .ZN(n6038) );
  INV_X1 U6205 ( .A(n6038), .ZN(n6012) );
  NAND2_X1 U6206 ( .A1(n5997), .A2(n5996), .ZN(n5999) );
  NAND2_X1 U6207 ( .A1(n8459), .A2(n4632), .ZN(n4630) );
  NAND2_X1 U6208 ( .A1(n4630), .A2(n4631), .ZN(n8402) );
  NAND2_X1 U6209 ( .A1(n5237), .A2(n5236), .ZN(n5240) );
  NAND3_X1 U6210 ( .A1(n9056), .A2(n4648), .A3(n4647), .ZN(n4646) );
  NAND2_X1 U6211 ( .A1(n5319), .A2(n4653), .ZN(n4650) );
  NAND2_X1 U6212 ( .A1(n4650), .A2(n4651), .ZN(n5369) );
  NAND2_X1 U6213 ( .A1(n5503), .A2(n5501), .ZN(n4657) );
  NAND2_X1 U6214 ( .A1(n4656), .A2(n4655), .ZN(n5617) );
  NAND2_X1 U6215 ( .A1(n5503), .A2(n4658), .ZN(n4656) );
  NAND3_X1 U6216 ( .A1(n8942), .A2(n8984), .A3(n4667), .ZN(n4666) );
  NAND2_X1 U6217 ( .A1(n5647), .A2(n4582), .ZN(n4676) );
  OAI21_X1 U6218 ( .B1(n5647), .B2(n4682), .A(n5646), .ZN(n5669) );
  NAND2_X1 U6219 ( .A1(n5765), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6220 ( .A1(n5765), .A2(n5763), .ZN(n4688) );
  OR2_X1 U6221 ( .A1(n5765), .A2(n5764), .ZN(n4692) );
  NAND2_X1 U6222 ( .A1(n9894), .A2(n9900), .ZN(n4698) );
  NAND3_X1 U6223 ( .A1(n9888), .A2(n6801), .A3(n6852), .ZN(n6961) );
  INV_X1 U6224 ( .A(n4483), .ZN(n9888) );
  NAND2_X1 U6225 ( .A1(n5094), .A2(n4907), .ZN(n5169) );
  NAND2_X1 U6226 ( .A1(n5164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5165) );
  INV_X1 U6227 ( .A(n4705), .ZN(n9248) );
  NOR2_X1 U6228 ( .A1(n9409), .A2(n9561), .ZN(n9396) );
  AOI21_X2 U6229 ( .B1(n4484), .B2(n5032), .A(n4722), .ZN(n4721) );
  NAND2_X1 U6230 ( .A1(n4589), .A2(n4719), .ZN(n4715) );
  NAND2_X1 U6231 ( .A1(n4589), .A2(n4484), .ZN(n4718) );
  NAND3_X1 U6232 ( .A1(n4716), .A2(n4715), .A3(n5576), .ZN(n8761) );
  NAND2_X1 U6233 ( .A1(n4719), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U6234 ( .A1(n5210), .A2(n4725), .ZN(n5212) );
  NAND3_X1 U6235 ( .A1(n5210), .A2(n5110), .A3(n4725), .ZN(n5243) );
  NAND3_X1 U6236 ( .A1(n8701), .A2(n4729), .A3(n8636), .ZN(n4727) );
  NAND3_X1 U6237 ( .A1(n8701), .A2(n8636), .A3(n5030), .ZN(n5027) );
  NAND3_X1 U6238 ( .A1(n5037), .A2(n4732), .A3(n5307), .ZN(n4731) );
  NAND3_X1 U6239 ( .A1(n5037), .A2(n5307), .A3(n7056), .ZN(n4736) );
  NAND2_X1 U6240 ( .A1(n5035), .A2(n4740), .ZN(n4737) );
  OAI21_X1 U6241 ( .B1(n5951), .B2(n9870), .A(n5268), .ZN(n4743) );
  OAI21_X1 U6242 ( .B1(n8657), .B2(n4563), .A(n4747), .ZN(n5811) );
  INV_X1 U6243 ( .A(n5811), .ZN(n5813) );
  XNOR2_X2 U6244 ( .A(n4770), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7120) );
  INV_X1 U6245 ( .A(n4777), .ZN(n8320) );
  NAND2_X1 U6246 ( .A1(n5997), .A2(n4527), .ZN(n6033) );
  NAND3_X1 U6247 ( .A1(n9129), .A2(n4785), .A3(n4784), .ZN(n4787) );
  NAND3_X1 U6248 ( .A1(n4788), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4786) );
  INV_X1 U6249 ( .A(n9146), .ZN(n4792) );
  NAND2_X1 U6250 ( .A1(n5392), .A2(n4797), .ZN(n4793) );
  NAND2_X1 U6251 ( .A1(n5392), .A2(n5390), .ZN(n4800) );
  OR2_X1 U6252 ( .A1(n5392), .A2(n5391), .ZN(n4803) );
  AND2_X2 U6253 ( .A1(n4813), .A2(n4811), .ZN(n9236) );
  OR2_X2 U6254 ( .A1(n9290), .A2(n4561), .ZN(n4813) );
  NAND2_X1 U6255 ( .A1(n4828), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U6256 ( .A1(n4828), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U6257 ( .A1(n4828), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U6258 ( .A1(n4828), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U6259 ( .A1(n4828), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U6260 ( .A1(n4828), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U6261 ( .A1(n4828), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U6262 ( .A1(n4828), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U6263 ( .A1(n4828), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U6264 ( .A1(n4828), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U6265 ( .A1(n4828), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U6266 ( .A1(n4828), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U6267 ( .A1(n4828), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U6268 ( .A1(n7737), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n4828), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n7604) );
  AOI22_X1 U6269 ( .A1(n7737), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n4828), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n7639) );
  OR2_X1 U6270 ( .A1(n7050), .A2(n6904), .ZN(n7045) );
  NAND2_X1 U6271 ( .A1(n7930), .A2(n4553), .ZN(n7932) );
  INV_X1 U6272 ( .A(n4839), .ZN(n7957) );
  AOI211_X1 U6273 ( .C1(n7948), .C2(n4844), .A(n4843), .B(n4840), .ZN(n4839)
         );
  OAI22_X1 U6274 ( .A1(n4845), .A2(n4841), .B1(n7956), .B2(n8020), .ZN(n4840)
         );
  NAND2_X1 U6275 ( .A1(n4842), .A2(n8047), .ZN(n4841) );
  NOR2_X1 U6276 ( .A1(n4845), .A2(n4846), .ZN(n4844) );
  NAND2_X1 U6277 ( .A1(n4848), .A2(n4847), .ZN(n8006) );
  NAND2_X1 U6278 ( .A1(n4535), .A2(n4849), .ZN(n4847) );
  AOI21_X1 U6279 ( .B1(n4850), .B2(n4849), .A(n4559), .ZN(n4848) );
  NOR2_X1 U6280 ( .A1(n5999), .A2(n5054), .ZN(n6036) );
  NAND2_X1 U6281 ( .A1(n6038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U6282 ( .A1(n4858), .A2(n4854), .ZN(P2_U3244) );
  OAI21_X1 U6283 ( .B1(n4500), .B2(n4857), .A(n4856), .ZN(n4855) );
  NAND2_X1 U6284 ( .A1(n5104), .A2(n4512), .ZN(n4856) );
  NAND2_X1 U6285 ( .A1(n4512), .A2(n4594), .ZN(n4857) );
  NAND2_X1 U6286 ( .A1(n8064), .A2(n4512), .ZN(n4858) );
  OAI211_X2 U6287 ( .C1(n6149), .C2(n6489), .A(n6148), .B(n6147), .ZN(n10033)
         );
  MUX2_X1 U6288 ( .A(n7944), .B(n7943), .S(n8020), .Z(n7948) );
  NAND2_X1 U6289 ( .A1(n8025), .A2(n8024), .ZN(n8061) );
  NAND2_X1 U6290 ( .A1(n4984), .A2(n4982), .ZN(n8064) );
  INV_X1 U6291 ( .A(n7844), .ZN(n8266) );
  OAI21_X1 U6292 ( .B1(n7844), .B2(n4564), .A(n8001), .ZN(n8239) );
  INV_X1 U6293 ( .A(n7878), .ZN(n4860) );
  NAND2_X1 U6294 ( .A1(n6871), .A2(n6872), .ZN(n6876) );
  NAND2_X1 U6295 ( .A1(n6761), .A2(n7888), .ZN(n6872) );
  NAND2_X2 U6296 ( .A1(n6884), .A2(n6769), .ZN(n7888) );
  NAND2_X1 U6297 ( .A1(n7023), .A2(n4862), .ZN(n7243) );
  NAND2_X1 U6298 ( .A1(n6996), .A2(n8035), .ZN(n7023) );
  NOR2_X1 U6299 ( .A1(n4864), .A2(n4863), .ZN(n4862) );
  AND2_X2 U6300 ( .A1(n4867), .A2(n4865), .ZN(n8390) );
  OR2_X2 U6301 ( .A1(n8428), .A2(n4871), .ZN(n4867) );
  INV_X1 U6302 ( .A(n7960), .ZN(n4873) );
  INV_X1 U6303 ( .A(n5995), .ZN(n5997) );
  NAND4_X1 U6304 ( .A1(n4875), .A2(n5062), .A3(n4475), .A4(n4487), .ZN(n5995)
         );
  NAND2_X1 U6305 ( .A1(n7478), .A2(n4532), .ZN(n4877) );
  NAND2_X1 U6306 ( .A1(n7849), .A2(n4524), .ZN(n4888) );
  NAND2_X1 U6307 ( .A1(n4888), .A2(n4889), .ZN(n7875) );
  NAND2_X1 U6308 ( .A1(n4898), .A2(n4896), .ZN(n7258) );
  OAI21_X1 U6309 ( .B1(n9444), .B2(n4904), .A(n4555), .ZN(n9416) );
  AND2_X2 U6310 ( .A1(n5294), .A2(n4908), .ZN(n4907) );
  NAND3_X1 U6311 ( .A1(n9171), .A2(n4913), .A3(n4914), .ZN(n4911) );
  INV_X1 U6312 ( .A(n9190), .ZN(n4928) );
  OAI21_X1 U6313 ( .B1(n9356), .B2(n4921), .A(n4919), .ZN(n4923) );
  NOR2_X1 U6314 ( .A1(n4517), .A2(n4925), .ZN(n4922) );
  INV_X1 U6315 ( .A(n4923), .ZN(n9193) );
  INV_X1 U6316 ( .A(n4929), .ZN(n9353) );
  INV_X1 U6317 ( .A(n9276), .ZN(n4941) );
  NAND2_X1 U6318 ( .A1(n7812), .A2(n4945), .ZN(n4942) );
  NAND2_X1 U6319 ( .A1(n4942), .A2(n4943), .ZN(n7733) );
  NAND2_X1 U6320 ( .A1(n7812), .A2(n4949), .ZN(n4944) );
  AOI21_X1 U6321 ( .B1(n7812), .B2(n7659), .A(n7811), .ZN(n7674) );
  INV_X1 U6322 ( .A(n6713), .ZN(n4954) );
  AOI21_X1 U6323 ( .B1(n4951), .B2(n6746), .A(n4554), .ZN(n4955) );
  NAND3_X1 U6324 ( .A1(n4955), .A2(n4953), .A3(n4952), .ZN(n6097) );
  INV_X1 U6325 ( .A(n6072), .ZN(n4960) );
  OAI21_X2 U6326 ( .B1(n7544), .B2(n4964), .A(n4961), .ZN(n7697) );
  INV_X1 U6327 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4971) );
  NAND4_X1 U6328 ( .A1(n4487), .A2(n4475), .A3(n6108), .A4(n5989), .ZN(n6324)
         );
  NAND2_X2 U6329 ( .A1(n5187), .A2(n6057), .ZN(n5206) );
  OR2_X2 U6330 ( .A1(n6468), .A2(n4557), .ZN(n5187) );
  NAND2_X1 U6331 ( .A1(n5944), .A2(n5943), .ZN(n4993) );
  NAND2_X1 U6332 ( .A1(n4997), .A2(n4581), .ZN(n5743) );
  NAND2_X1 U6333 ( .A1(n5000), .A2(n7868), .ZN(n8502) );
  NAND2_X1 U6334 ( .A1(n5528), .A2(n5007), .ZN(n5001) );
  NAND2_X1 U6335 ( .A1(n5789), .A2(n5012), .ZN(n5011) );
  OAI211_X1 U6336 ( .C1(n5023), .C2(n5975), .A(n5021), .B(n5018), .ZN(P1_U3218) );
  OR2_X1 U6337 ( .A1(n5969), .A2(n5968), .ZN(n5019) );
  NAND3_X1 U6338 ( .A1(n5023), .A2(n5977), .A3(n5022), .ZN(n5021) );
  OAI21_X1 U6339 ( .B1(n5974), .B2(n5973), .A(n5972), .ZN(n5023) );
  NAND3_X1 U6340 ( .A1(n8701), .A2(n8636), .A3(n8700), .ZN(n8699) );
  AND2_X1 U6341 ( .A1(n5418), .A2(n5389), .ZN(n5034) );
  NOR2_X1 U6342 ( .A1(n5374), .A2(n5135), .ZN(n5428) );
  NAND2_X1 U6343 ( .A1(n6900), .A2(n5044), .ZN(n5042) );
  OAI21_X1 U6344 ( .B1(n6900), .B2(n4478), .A(n5043), .ZN(n6903) );
  AOI21_X1 U6345 ( .B1(n8031), .B2(n5046), .A(n5045), .ZN(n5043) );
  NOR2_X1 U6346 ( .A1(n5046), .A2(n5045), .ZN(n5044) );
  NAND3_X1 U6347 ( .A1(n6002), .A2(n4895), .A3(n6034), .ZN(n5054) );
  AOI21_X1 U6348 ( .B1(n8263), .B2(n8264), .A(n8215), .ZN(n8248) );
  NAND2_X1 U6349 ( .A1(n8263), .A2(n5059), .ZN(n5058) );
  NAND2_X1 U6350 ( .A1(n8194), .A2(n4501), .ZN(n8477) );
  NAND3_X1 U6351 ( .A1(n4487), .A2(n4475), .A3(n6108), .ZN(n6322) );
  NOR2_X1 U6352 ( .A1(n9159), .A2(n4569), .ZN(n9329) );
  INV_X1 U6353 ( .A(n4569), .ZN(n5072) );
  NAND2_X1 U6354 ( .A1(n5073), .A2(n5074), .ZN(n9170) );
  NAND2_X1 U6355 ( .A1(n9247), .A2(n5076), .ZN(n5073) );
  NAND2_X1 U6356 ( .A1(n5088), .A2(n5087), .ZN(n9153) );
  NAND2_X1 U6357 ( .A1(n9149), .A2(n9148), .ZN(n9435) );
  NAND2_X1 U6358 ( .A1(n9394), .A2(n9395), .ZN(n5093) );
  NAND2_X1 U6359 ( .A1(n5093), .A2(n5091), .ZN(n9156) );
  NAND3_X1 U6360 ( .A1(n5121), .A2(n5294), .A3(n10261), .ZN(n5887) );
  NAND2_X1 U6361 ( .A1(n5168), .A2(n5098), .ZN(n5166) );
  NAND2_X2 U6362 ( .A1(n8616), .A2(n6018), .ZN(n6086) );
  INV_X1 U6363 ( .A(n8314), .ZN(n8340) );
  AND2_X1 U6364 ( .A1(n7704), .A2(n7703), .ZN(n7777) );
  INV_X1 U6365 ( .A(n8088), .ZN(n6682) );
  XNOR2_X1 U6366 ( .A(n8239), .B(n8238), .ZN(n8245) );
  OR2_X1 U6367 ( .A1(n7648), .A2(n10234), .ZN(n6054) );
  NAND2_X1 U6368 ( .A1(n5278), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6369 ( .A1(n5278), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5133) );
  INV_X1 U6370 ( .A(n5278), .ZN(n5962) );
  INV_X1 U6371 ( .A(n5130), .ZN(n9593) );
  NOR2_X2 U6372 ( .A1(n8487), .A2(n7836), .ZN(n8468) );
  AND2_X1 U6373 ( .A1(n5738), .A2(n5737), .ZN(n5099) );
  OR2_X1 U6374 ( .A1(n9161), .A2(n9160), .ZN(n5100) );
  AND2_X1 U6375 ( .A1(n8332), .A2(n8342), .ZN(n5101) );
  INV_X1 U6376 ( .A(n9495), .ZN(n9219) );
  OR2_X1 U6377 ( .A1(n9301), .A2(n9280), .ZN(n5102) );
  NOR2_X1 U6378 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5103) );
  NAND2_X1 U6379 ( .A1(n8314), .A2(n5109), .ZN(n8300) );
  AND2_X1 U6380 ( .A1(n5935), .A2(n5934), .ZN(n9203) );
  AND2_X1 U6381 ( .A1(n5451), .A2(n5427), .ZN(n5105) );
  AND2_X1 U6382 ( .A1(n6454), .A2(n6449), .ZN(n8471) );
  INV_X1 U6383 ( .A(n8471), .ZN(n8434) );
  AND2_X1 U6384 ( .A1(n5527), .A2(n5507), .ZN(n5106) );
  OR2_X1 U6385 ( .A1(n9565), .A2(n9427), .ZN(n5107) );
  NOR2_X1 U6386 ( .A1(n8326), .A2(n8315), .ZN(n5109) );
  INV_X1 U6387 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5990) );
  INV_X1 U6388 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5114) );
  INV_X1 U6389 ( .A(n8059), .ZN(n7873) );
  INV_X1 U6390 ( .A(n8029), .ZN(n6873) );
  OR2_X1 U6391 ( .A1(n9251), .A2(n5951), .ZN(n5861) );
  INV_X1 U6392 ( .A(n5850), .ZN(n5848) );
  INV_X1 U6393 ( .A(n9203), .ZN(n9169) );
  INV_X1 U6394 ( .A(n6272), .ZN(n6271) );
  INV_X1 U6395 ( .A(n6425), .ZN(n6427) );
  INV_X1 U6396 ( .A(n6301), .ZN(n6293) );
  INV_X1 U6397 ( .A(n6372), .ZN(n6370) );
  OR2_X1 U6398 ( .A1(n7601), .A2(n10380), .ZN(n7635) );
  INV_X1 U6399 ( .A(n5778), .ZN(n5776) );
  NAND2_X1 U6400 ( .A1(n6858), .A2(n5953), .ZN(n5194) );
  INV_X1 U6401 ( .A(n5303), .ZN(n5301) );
  INV_X1 U6402 ( .A(n5953), .ZN(n5401) );
  INV_X1 U6403 ( .A(n5705), .ZN(n5704) );
  INV_X1 U6404 ( .A(n5542), .ZN(n5541) );
  NAND2_X1 U6405 ( .A1(n5848), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5928) );
  INV_X1 U6406 ( .A(n5136), .ZN(n5137) );
  INV_X1 U6407 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5530) );
  INV_X1 U6408 ( .A(SI_9_), .ZN(n10469) );
  INV_X1 U6409 ( .A(SI_8_), .ZN(n10442) );
  NAND2_X1 U6410 ( .A1(n6271), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U6411 ( .A1(n6427), .A2(n6426), .ZN(n6656) );
  AND2_X1 U6412 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6099) );
  OR2_X1 U6413 ( .A1(n6656), .A2(n10489), .ZN(n6663) );
  NAND2_X1 U6414 ( .A1(n6293), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6303) );
  AND2_X1 U6415 ( .A1(n6881), .A2(n6878), .ZN(n6359) );
  NAND2_X1 U6416 ( .A1(n6370), .A2(n6369), .ZN(n6407) );
  INV_X1 U6417 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10470) );
  INV_X1 U6418 ( .A(n8301), .ZN(n8209) );
  INV_X1 U6419 ( .A(n7841), .ZN(n8315) );
  OR2_X1 U6420 ( .A1(n6156), .A2(n7190), .ZN(n6179) );
  AND2_X1 U6421 ( .A1(n7923), .A2(n7922), .ZN(n8041) );
  NAND2_X1 U6422 ( .A1(n6896), .A2(n7893), .ZN(n6925) );
  OR2_X1 U6423 ( .A1(n7526), .A2(n6340), .ZN(n6341) );
  INV_X1 U6424 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U6425 ( .A1(n5776), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5795) );
  INV_X1 U6426 ( .A(n7419), .ZN(n5418) );
  XNOR2_X1 U6427 ( .A(n5836), .B(n6815), .ZN(n5838) );
  INV_X1 U6428 ( .A(n5655), .ZN(n5653) );
  NOR2_X1 U6429 ( .A1(n5863), .A2(n5862), .ZN(n8749) );
  NAND2_X1 U6430 ( .A1(n5704), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5727) );
  OR2_X1 U6431 ( .A1(n5403), .A2(n5402), .ZN(n5436) );
  OR2_X1 U6432 ( .A1(n9786), .A2(n9785), .ZN(n9782) );
  OAI22_X1 U6433 ( .A1(n9203), .A2(n9871), .B1(n9202), .B2(n9201), .ZN(n9204)
         );
  INV_X1 U6434 ( .A(n9532), .ZN(n9161) );
  OR2_X1 U6435 ( .A1(n5727), .A2(n8658), .ZN(n5752) );
  XNOR2_X1 U6436 ( .A(n9492), .B(n9227), .ZN(n9199) );
  NAND2_X1 U6437 ( .A1(n8982), .A2(n9863), .ZN(n8969) );
  AND2_X1 U6438 ( .A1(n5788), .A2(n5770), .ZN(n5771) );
  INV_X1 U6439 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6440 ( .A1(n5558), .A2(n10276), .ZN(n5586) );
  NAND2_X1 U6441 ( .A1(n5478), .A2(n5477), .ZN(n5501) );
  OR2_X1 U6442 ( .A1(n7646), .A2(n10460), .ZN(n7680) );
  NAND2_X1 U6443 ( .A1(n6099), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6118) );
  OR2_X1 U6444 ( .A1(n6303), .A2(n8128), .ZN(n6372) );
  INV_X1 U6445 ( .A(n7840), .ZN(n8346) );
  INV_X1 U6446 ( .A(n8183), .ZN(n8511) );
  INV_X1 U6447 ( .A(n8549), .ZN(n8339) );
  INV_X1 U6448 ( .A(n7540), .ZN(n9616) );
  AND2_X1 U6449 ( .A1(n7929), .A2(n7931), .ZN(n8043) );
  OR2_X1 U6450 ( .A1(n6447), .A2(n6354), .ZN(n6460) );
  OR2_X1 U6451 ( .A1(n5677), .A2(n8650), .ZN(n5705) );
  OR2_X1 U6452 ( .A1(n5826), .A2(n8676), .ZN(n5850) );
  AOI21_X1 U6453 ( .B1(n6803), .B2(n4477), .A(n5174), .ZN(n6673) );
  NAND2_X1 U6454 ( .A1(n5653), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5677) );
  INV_X1 U6455 ( .A(n5958), .ZN(n5852) );
  AND2_X1 U6456 ( .A1(n6582), .A2(n6555), .ZN(n6557) );
  AND2_X1 U6457 ( .A1(n9525), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U6458 ( .A1(n9142), .A2(n9141), .ZN(n9624) );
  AND2_X1 U6459 ( .A1(n8876), .A2(n8873), .ZN(n9865) );
  NAND2_X1 U6460 ( .A1(n5617), .A2(n5616), .ZN(n5647) );
  NOR2_X1 U6461 ( .A1(n5431), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5532) );
  INV_X1 U6462 ( .A(SI_4_), .ZN(n5261) );
  INV_X1 U6463 ( .A(n8200), .ZN(n8433) );
  AND4_X1 U6464 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n8445)
         );
  INV_X1 U6465 ( .A(n9962), .ZN(n9964) );
  INV_X1 U6466 ( .A(n9965), .ZN(n9602) );
  OR2_X1 U6467 ( .A1(n6660), .A2(n6659), .ZN(n8317) );
  INV_X1 U6468 ( .A(n9989), .ZN(n8499) );
  INV_X1 U6469 ( .A(n8486), .ZN(n10004) );
  INV_X1 U6470 ( .A(n9988), .ZN(n8455) );
  AND2_X1 U6471 ( .A1(n6343), .A2(n6342), .ZN(n6881) );
  AND2_X1 U6472 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  INV_X1 U6473 ( .A(n10069), .ZN(n10078) );
  INV_X1 U6474 ( .A(n6460), .ZN(n9996) );
  AND2_X1 U6475 ( .A1(n5850), .A2(n5827), .ZN(n9270) );
  AND2_X1 U6476 ( .A1(n9723), .A2(n9060), .ZN(n9811) );
  INV_X1 U6477 ( .A(n9823), .ZN(n9806) );
  NAND2_X1 U6478 ( .A1(n8984), .A2(n8983), .ZN(n9263) );
  NAND2_X1 U6479 ( .A1(n9939), .A2(n5910), .ZN(n9847) );
  AND2_X1 U6480 ( .A1(n6803), .A2(n7572), .ZN(n6804) );
  INV_X1 U6481 ( .A(n9856), .ZN(n9934) );
  AND2_X1 U6482 ( .A1(n9843), .A2(n7504), .ZN(n9660) );
  INV_X1 U6483 ( .A(n9660), .ZN(n9924) );
  INV_X1 U6484 ( .A(n7504), .ZN(n9939) );
  AND2_X1 U6485 ( .A1(n5624), .A2(n5648), .ZN(n9114) );
  XNOR2_X1 U6486 ( .A(n5367), .B(n5346), .ZN(n5365) );
  XNOR2_X1 U6487 ( .A(n5317), .B(n10357), .ZN(n5315) );
  AND2_X1 U6488 ( .A1(n7458), .A2(n6005), .ZN(n6447) );
  INV_X1 U6489 ( .A(n8570), .ZN(n8408) );
  INV_X1 U6490 ( .A(n7379), .ZN(n8079) );
  INV_X1 U6491 ( .A(n9993), .ZN(n8496) );
  NAND2_X1 U6492 ( .A1(n9993), .A2(n9986), .ZN(n8501) );
  INV_X1 U6493 ( .A(n10097), .ZN(n10095) );
  INV_X1 U6494 ( .A(n10083), .ZN(n10081) );
  AND2_X1 U6495 ( .A1(n6446), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10003) );
  INV_X1 U6496 ( .A(n5940), .ZN(n5941) );
  INV_X1 U6497 ( .A(n9511), .ZN(n9261) );
  INV_X1 U6498 ( .A(n9167), .ZN(n9265) );
  INV_X1 U6499 ( .A(n9294), .ZN(n9266) );
  OR2_X1 U6500 ( .A1(P1_U3083), .A2(n6499), .ZN(n9828) );
  OR2_X1 U6501 ( .A1(n6727), .A2(n6806), .ZN(n9957) );
  OR2_X1 U6502 ( .A1(n6727), .A2(n6721), .ZN(n9940) );
  INV_X1 U6503 ( .A(n9878), .ZN(n9877) );
  INV_X1 U6504 ( .A(n9063), .ZN(n8982) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10236) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6587) );
  AND2_X1 U6507 ( .A1(n6447), .A2(n10003), .ZN(P2_U3966) );
  NOR2_X1 U6508 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5119) );
  NOR2_X1 U6509 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5118) );
  NOR2_X1 U6510 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5117) );
  NAND4_X1 U6511 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n10454), .ZN(n5120)
         );
  INV_X1 U6512 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5122) );
  INV_X1 U6513 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6514 ( .A1(n5166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5125) );
  INV_X1 U6515 ( .A(n5126), .ZN(n5128) );
  NAND2_X1 U6516 ( .A1(n5217), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5134) );
  AND2_X4 U6517 ( .A1(n5129), .A2(n9593), .ZN(n5278) );
  NAND2_X1 U6518 ( .A1(n4482), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6519 ( .A1(n5282), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5131) );
  INV_X1 U6520 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U6521 ( .A1(n10454), .A2(n10339), .ZN(n5135) );
  INV_X1 U6522 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5138) );
  INV_X1 U6523 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5139) );
  XNOR2_X2 U6524 ( .A(n5140), .B(n5139), .ZN(n7069) );
  OR2_X1 U6525 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5141) );
  NOR2_X1 U6526 ( .A1(n5142), .A2(n5103), .ZN(n5155) );
  AND2_X2 U6527 ( .A1(n5155), .A2(n5143), .ZN(n8979) );
  NAND2_X1 U6528 ( .A1(n5144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5147) );
  INV_X1 U6529 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6530 ( .A1(n5147), .A2(n5146), .ZN(n5149) );
  NAND2_X1 U6531 ( .A1(n5149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6532 ( .A1(n5147), .A2(n5146), .ZN(n5148) );
  NAND2_X1 U6533 ( .A1(n5149), .A2(n5148), .ZN(n7561) );
  INV_X1 U6534 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6535 ( .A1(n5151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5152) );
  MUX2_X1 U6536 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5152), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5153) );
  NAND2_X1 U6537 ( .A1(n5153), .A2(n5144), .ZN(n7472) );
  NOR2_X1 U6538 ( .A1(n7561), .A2(n7472), .ZN(n5154) );
  NAND2_X1 U6539 ( .A1(n5155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6540 ( .A1(n4546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5157) );
  MUX2_X1 U6541 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5157), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5159) );
  AND2_X1 U6542 ( .A1(n7069), .A2(n9327), .ZN(n5914) );
  INV_X1 U6543 ( .A(n5914), .ZN(n5886) );
  AND2_X2 U6544 ( .A1(n5953), .A2(n5160), .ZN(n5713) );
  INV_X1 U6545 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U6546 ( .A1(n4479), .A2(SI_0_), .ZN(n5162) );
  INV_X1 U6547 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6548 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  AND2_X1 U6549 ( .A1(n5163), .A2(n5187), .ZN(n9601) );
  NAND2_X1 U6550 ( .A1(n5169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U6551 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5170), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5171) );
  NAND2_X2 U6552 ( .A1(n5923), .A2(n9688), .ZN(n5348) );
  MUX2_X1 U6553 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9601), .S(n5348), .Z(n7572) );
  AND2_X4 U6554 ( .A1(n5172), .A2(n5978), .ZN(n5634) );
  NAND2_X1 U6555 ( .A1(n7572), .A2(n5634), .ZN(n5173) );
  OAI21_X1 U6556 ( .B1(n6623), .B2(n5978), .A(n5173), .ZN(n5174) );
  NAND2_X1 U6557 ( .A1(n6803), .A2(n5634), .ZN(n5177) );
  INV_X1 U6558 ( .A(n5978), .ZN(n5175) );
  AOI22_X1 U6559 ( .A1(n7572), .A2(n5953), .B1(n5175), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6560 ( .A1(n5177), .A2(n5176), .ZN(n6671) );
  NAND2_X1 U6561 ( .A1(n6673), .A2(n6671), .ZN(n6672) );
  INV_X1 U6562 ( .A(n6671), .ZN(n5179) );
  INV_X1 U6563 ( .A(n5917), .ZN(n5178) );
  NAND2_X1 U6564 ( .A1(n5179), .A2(n6815), .ZN(n5180) );
  NAND2_X1 U6565 ( .A1(n6672), .A2(n5180), .ZN(n6705) );
  INV_X1 U6566 ( .A(n6705), .ZN(n5197) );
  NAND2_X1 U6567 ( .A1(n5235), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6568 ( .A1(n5217), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5181) );
  AND2_X1 U6569 ( .A1(n5182), .A2(n5181), .ZN(n5184) );
  NAND2_X1 U6570 ( .A1(n5282), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6571 ( .A1(n4480), .A2(n5634), .ZN(n5195) );
  AND2_X4 U6572 ( .A1(n5348), .A2(n4479), .ZN(n8848) );
  AND2_X1 U6573 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6574 ( .A1(n5320), .A2(n5186), .ZN(n6057) );
  INV_X1 U6575 ( .A(SI_1_), .ZN(n5188) );
  MUX2_X1 U6576 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6040), .Z(n5204) );
  XNOR2_X1 U6577 ( .A(n5205), .B(n5204), .ZN(n6482) );
  INV_X1 U6578 ( .A(n6482), .ZN(n5189) );
  NAND2_X1 U6579 ( .A1(n8848), .A2(n5189), .ZN(n5193) );
  NAND2_X1 U6580 ( .A1(n5292), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5192) );
  INV_X2 U6581 ( .A(n5348), .ZN(n5538) );
  NAND2_X1 U6582 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5190) );
  XNOR2_X1 U6583 ( .A(n5190), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U6584 ( .A1(n5538), .A2(n6630), .ZN(n5191) );
  NAND2_X1 U6585 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  XNOR2_X1 U6586 ( .A(n5196), .B(n5327), .ZN(n5198) );
  INV_X1 U6587 ( .A(n5198), .ZN(n6707) );
  NAND2_X1 U6588 ( .A1(n5197), .A2(n6707), .ZN(n5203) );
  NAND2_X1 U6589 ( .A1(n6705), .A2(n5198), .ZN(n5201) );
  NAND2_X1 U6590 ( .A1(n4480), .A2(n5713), .ZN(n5200) );
  OR2_X1 U6591 ( .A1(n6801), .A2(n5951), .ZN(n5199) );
  NAND2_X1 U6592 ( .A1(n5200), .A2(n5199), .ZN(n6704) );
  NAND2_X1 U6593 ( .A1(n5201), .A2(n6704), .ZN(n5202) );
  NAND2_X1 U6594 ( .A1(n5203), .A2(n5202), .ZN(n7577) );
  INV_X1 U6595 ( .A(n7577), .ZN(n5232) );
  NAND2_X1 U6596 ( .A1(n5205), .A2(n5204), .ZN(n5208) );
  NAND2_X1 U6597 ( .A1(n5206), .A2(SI_1_), .ZN(n5207) );
  NAND2_X1 U6598 ( .A1(n5208), .A2(n5207), .ZN(n5237) );
  XNOR2_X1 U6599 ( .A(n5237), .B(n5236), .ZN(n6472) );
  NAND2_X1 U6600 ( .A1(n5292), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5216) );
  NOR2_X1 U6601 ( .A1(n5210), .A2(n5453), .ZN(n5211) );
  MUX2_X1 U6602 ( .A(n5453), .B(n5211), .S(P1_IR_REG_2__SCAN_IN), .Z(n5214) );
  INV_X1 U6603 ( .A(n5212), .ZN(n5213) );
  NOR2_X1 U6604 ( .A1(n5214), .A2(n5213), .ZN(n6518) );
  NAND2_X1 U6605 ( .A1(n5538), .A2(n6518), .ZN(n5215) );
  NAND2_X1 U6606 ( .A1(n4483), .A2(n5953), .ZN(n5223) );
  NAND2_X1 U6607 ( .A1(n5278), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6608 ( .A1(n5217), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6609 ( .A1(n5282), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6610 ( .A1(n4482), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6611 ( .A1(n6850), .A2(n5634), .ZN(n5222) );
  NAND2_X1 U6612 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  XNOR2_X1 U6613 ( .A(n5224), .B(n5327), .ZN(n5229) );
  INV_X1 U6614 ( .A(n5229), .ZN(n5227) );
  AND2_X1 U6615 ( .A1(n4483), .A2(n5634), .ZN(n5225) );
  AOI21_X1 U6616 ( .B1(n6850), .B2(n5713), .A(n5225), .ZN(n5228) );
  INV_X1 U6617 ( .A(n5228), .ZN(n5226) );
  NAND2_X1 U6618 ( .A1(n5227), .A2(n5226), .ZN(n5230) );
  NAND2_X1 U6619 ( .A1(n5229), .A2(n5228), .ZN(n5233) );
  NAND2_X1 U6620 ( .A1(n5230), .A2(n5233), .ZN(n7576) );
  INV_X1 U6621 ( .A(n7576), .ZN(n5231) );
  NAND2_X1 U6622 ( .A1(n5232), .A2(n5231), .ZN(n7578) );
  NAND2_X1 U6623 ( .A1(n7578), .A2(n5233), .ZN(n6792) );
  NAND2_X1 U6624 ( .A1(n5278), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6840) );
  INV_X1 U6625 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6626 ( .A1(n5217), .A2(n5234), .ZN(n6839) );
  NAND2_X1 U6627 ( .A1(n5282), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U6628 ( .A1(n4482), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6837) );
  NAND4_X1 U6629 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n9077)
         );
  NAND2_X1 U6630 ( .A1(n9077), .A2(n5634), .ZN(n5248) );
  NAND2_X1 U6631 ( .A1(n5238), .A2(SI_2_), .ZN(n5239) );
  NAND2_X1 U6632 ( .A1(n5240), .A2(n5239), .ZN(n5257) );
  MUX2_X1 U6633 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6040), .Z(n5258) );
  XNOR2_X1 U6634 ( .A(n5257), .B(n5256), .ZN(n6478) );
  NAND2_X1 U6635 ( .A1(n5292), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6636 ( .A1(n5212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5242) );
  MUX2_X1 U6637 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5242), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5244) );
  AND2_X1 U6638 ( .A1(n5244), .A2(n5243), .ZN(n6546) );
  NAND2_X1 U6639 ( .A1(n5538), .A2(n6546), .ZN(n5245) );
  NAND2_X1 U6640 ( .A1(n6964), .A2(n5953), .ZN(n5247) );
  NAND2_X1 U6641 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  XNOR2_X1 U6642 ( .A(n5249), .B(n6815), .ZN(n5270) );
  AND2_X1 U6643 ( .A1(n6964), .A2(n5634), .ZN(n5250) );
  AOI21_X1 U6644 ( .B1(n9077), .B2(n5713), .A(n5250), .ZN(n5271) );
  XNOR2_X1 U6645 ( .A(n5270), .B(n5271), .ZN(n6793) );
  NAND2_X1 U6646 ( .A1(n6792), .A2(n6793), .ZN(n6791) );
  INV_X1 U6647 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5251) );
  XNOR2_X1 U6648 ( .A(n5251), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U6649 ( .A1(n5217), .A2(n6951), .ZN(n5255) );
  NAND2_X1 U6650 ( .A1(n5278), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6651 ( .A1(n5282), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6652 ( .A1(n4482), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5252) );
  NAND4_X1 U6653 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n9076)
         );
  NAND2_X1 U6654 ( .A1(n5257), .A2(n5256), .ZN(n5260) );
  NAND2_X1 U6655 ( .A1(n5258), .A2(SI_3_), .ZN(n5259) );
  NAND2_X1 U6656 ( .A1(n5260), .A2(n5259), .ZN(n5288) );
  MUX2_X1 U6657 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6040), .Z(n5289) );
  XNOR2_X1 U6658 ( .A(n5288), .B(n5287), .ZN(n6480) );
  NAND2_X1 U6659 ( .A1(n8838), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6660 ( .A1(n5243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5262) );
  MUX2_X1 U6661 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5262), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5265) );
  INV_X1 U6662 ( .A(n5263), .ZN(n5264) );
  AND2_X1 U6663 ( .A1(n5265), .A2(n5264), .ZN(n9703) );
  NAND2_X1 U6664 ( .A1(n5538), .A2(n9703), .ZN(n5266) );
  NAND2_X1 U6665 ( .A1(n6952), .A2(n5953), .ZN(n5268) );
  AND2_X1 U6666 ( .A1(n6952), .A2(n5634), .ZN(n5269) );
  AOI21_X1 U6667 ( .B1(n9076), .B2(n5713), .A(n5269), .ZN(n5275) );
  XNOR2_X1 U6668 ( .A(n5274), .B(n5275), .ZN(n6835) );
  INV_X1 U6669 ( .A(n5270), .ZN(n5272) );
  NAND2_X1 U6670 ( .A1(n5272), .A2(n5271), .ZN(n6833) );
  AND2_X1 U6671 ( .A1(n6835), .A2(n6833), .ZN(n5273) );
  NAND2_X1 U6672 ( .A1(n6791), .A2(n5273), .ZN(n6834) );
  INV_X1 U6673 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6674 ( .A1(n5274), .A2(n5276), .ZN(n5277) );
  NAND2_X1 U6675 ( .A1(n6834), .A2(n5277), .ZN(n5304) );
  INV_X1 U6676 ( .A(n5304), .ZN(n5302) );
  NAND2_X1 U6677 ( .A1(n5278), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5286) );
  NAND3_X1 U6678 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5309) );
  INV_X1 U6679 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6680 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5279) );
  NAND2_X1 U6681 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  AND2_X1 U6682 ( .A1(n5309), .A2(n5281), .ZN(n9860) );
  NAND2_X1 U6683 ( .A1(n5958), .A2(n9860), .ZN(n5285) );
  NAND2_X1 U6684 ( .A1(n8851), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6685 ( .A1(n4482), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5283) );
  NAND4_X1 U6686 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9075)
         );
  NAND2_X1 U6687 ( .A1(n9075), .A2(n5634), .ZN(n5299) );
  NAND2_X1 U6688 ( .A1(n5288), .A2(n5287), .ZN(n5291) );
  NAND2_X1 U6689 ( .A1(n5289), .A2(SI_4_), .ZN(n5290) );
  MUX2_X1 U6690 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4479), .Z(n5317) );
  NAND2_X1 U6691 ( .A1(n8838), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5297) );
  NOR2_X1 U6692 ( .A1(n5263), .A2(n5453), .ZN(n5293) );
  MUX2_X1 U6693 ( .A(n5453), .B(n5293), .S(P1_IR_REG_5__SCAN_IN), .Z(n5295) );
  OR2_X1 U6694 ( .A1(n5295), .A2(n5294), .ZN(n6593) );
  INV_X1 U6695 ( .A(n6593), .ZN(n6537) );
  NAND2_X1 U6696 ( .A1(n5538), .A2(n6537), .ZN(n5296) );
  OAI211_X1 U6697 ( .C1(n5347), .C2(n6476), .A(n5297), .B(n5296), .ZN(n9858)
         );
  NAND2_X1 U6698 ( .A1(n9858), .A2(n5953), .ZN(n5298) );
  NAND2_X1 U6699 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  XNOR2_X1 U6700 ( .A(n5300), .B(n6815), .ZN(n5303) );
  NAND2_X1 U6701 ( .A1(n5302), .A2(n5301), .ZN(n5307) );
  NAND2_X1 U6702 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  AND2_X1 U6703 ( .A1(n9858), .A2(n5634), .ZN(n5306) );
  AOI21_X1 U6704 ( .B1(n9075), .B2(n5713), .A(n5306), .ZN(n7006) );
  NAND2_X1 U6705 ( .A1(n5278), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5314) );
  INV_X1 U6706 ( .A(n5309), .ZN(n5308) );
  INV_X1 U6707 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U6708 ( .A1(n5309), .A2(n6575), .ZN(n5310) );
  AND2_X1 U6709 ( .A1(n5336), .A2(n5310), .ZN(n7313) );
  NAND2_X1 U6710 ( .A1(n5958), .A2(n7313), .ZN(n5313) );
  NAND2_X1 U6711 ( .A1(n8851), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6712 ( .A1(n8841), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5311) );
  NAND4_X1 U6713 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n9074)
         );
  NAND2_X1 U6714 ( .A1(n9074), .A2(n5634), .ZN(n5326) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U6716 ( .A1(n5317), .A2(SI_5_), .ZN(n5318) );
  MUX2_X1 U6717 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6040), .Z(n5345) );
  XNOR2_X1 U6718 ( .A(n5344), .B(n5342), .ZN(n6484) );
  NAND2_X1 U6719 ( .A1(n8848), .A2(n6484), .ZN(n5324) );
  NOR2_X1 U6720 ( .A1(n5294), .A2(n5453), .ZN(n5321) );
  MUX2_X1 U6721 ( .A(n5453), .B(n5321), .S(P1_IR_REG_6__SCAN_IN), .Z(n5322) );
  INV_X1 U6722 ( .A(n6576), .ZN(n6554) );
  NAND2_X1 U6723 ( .A1(n5538), .A2(n6554), .ZN(n5323) );
  NAND2_X1 U6724 ( .A1(n8882), .A2(n5953), .ZN(n5325) );
  NAND2_X1 U6725 ( .A1(n5326), .A2(n5325), .ZN(n5328) );
  XNOR2_X1 U6726 ( .A(n5328), .B(n5327), .ZN(n5330) );
  AND2_X1 U6727 ( .A1(n8882), .A2(n5634), .ZN(n5329) );
  AOI21_X1 U6728 ( .B1(n9074), .B2(n5713), .A(n5329), .ZN(n5331) );
  NAND2_X1 U6729 ( .A1(n5330), .A2(n5331), .ZN(n7056) );
  INV_X1 U6730 ( .A(n5330), .ZN(n5333) );
  INV_X1 U6731 ( .A(n5331), .ZN(n5332) );
  NAND2_X1 U6732 ( .A1(n5333), .A2(n5332), .ZN(n7057) );
  NAND2_X1 U6733 ( .A1(n5278), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5341) );
  INV_X1 U6734 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6735 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  AND2_X1 U6736 ( .A1(n5359), .A2(n5337), .ZN(n7111) );
  NAND2_X1 U6737 ( .A1(n5958), .A2(n7111), .ZN(n5340) );
  NAND2_X1 U6738 ( .A1(n8851), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6739 ( .A1(n8841), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6740 ( .A1(n9073), .A2(n5713), .ZN(n5354) );
  MUX2_X1 U6741 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4479), .Z(n5367) );
  XNOR2_X1 U6742 ( .A(n5366), .B(n5365), .ZN(n6489) );
  NOR2_X1 U6743 ( .A1(n6489), .A2(n5347), .ZN(n5352) );
  INV_X1 U6744 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U6745 ( .A1(n5349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5350) );
  XNOR2_X1 U6746 ( .A(n5350), .B(n4750), .ZN(n6610) );
  OAI22_X1 U6747 ( .A1(n5377), .A2(n10273), .B1(n5982), .B2(n6610), .ZN(n5351)
         );
  NAND2_X1 U6748 ( .A1(n8872), .A2(n5634), .ZN(n5353) );
  NAND2_X1 U6749 ( .A1(n5354), .A2(n5353), .ZN(n7084) );
  NAND2_X1 U6750 ( .A1(n9073), .A2(n5634), .ZN(n5356) );
  NAND2_X1 U6751 ( .A1(n8872), .A2(n5953), .ZN(n5355) );
  NAND2_X1 U6752 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  XNOR2_X1 U6753 ( .A(n5357), .B(n6815), .ZN(n7083) );
  INV_X1 U6754 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U6755 ( .A1(n5359), .A2(n7340), .ZN(n5360) );
  AND2_X1 U6756 ( .A1(n5403), .A2(n5360), .ZN(n7339) );
  NAND2_X1 U6757 ( .A1(n5958), .A2(n7339), .ZN(n5364) );
  NAND2_X1 U6758 ( .A1(n5278), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6759 ( .A1(n8851), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6760 ( .A1(n8841), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5361) );
  NAND4_X1 U6761 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), .ZN(n9072)
         );
  NAND2_X1 U6762 ( .A1(n9072), .A2(n5634), .ZN(n5382) );
  NAND2_X1 U6763 ( .A1(n5367), .A2(SI_7_), .ZN(n5368) );
  INV_X1 U6764 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6765 ( .A(n5370), .B(n10476), .S(n4479), .Z(n5371) );
  NAND2_X1 U6766 ( .A1(n5371), .A2(n10442), .ZN(n5390) );
  INV_X1 U6767 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6768 ( .A1(n5372), .A2(SI_8_), .ZN(n5373) );
  XNOR2_X1 U6769 ( .A(n5392), .B(n5391), .ZN(n6490) );
  NAND2_X1 U6770 ( .A1(n6490), .A2(n8848), .ZN(n5380) );
  NAND2_X1 U6771 ( .A1(n5374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6772 ( .A1(n5375), .A2(n10454), .ZN(n5397) );
  OR2_X1 U6773 ( .A1(n5375), .A2(n10454), .ZN(n5376) );
  NAND2_X1 U6774 ( .A1(n5397), .A2(n5376), .ZN(n9727) );
  OAI22_X1 U6775 ( .A1(n5377), .A2(n10476), .B1(n5982), .B2(n9727), .ZN(n5378)
         );
  INV_X1 U6776 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6777 ( .A1(n7440), .A2(n5953), .ZN(n5381) );
  NAND2_X1 U6778 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  XNOR2_X1 U6779 ( .A(n5383), .B(n5327), .ZN(n7337) );
  NAND2_X1 U6780 ( .A1(n9072), .A2(n5713), .ZN(n5385) );
  NAND2_X1 U6781 ( .A1(n7440), .A2(n5634), .ZN(n5384) );
  AND2_X1 U6782 ( .A1(n5385), .A2(n5384), .ZN(n5387) );
  NAND2_X1 U6783 ( .A1(n7337), .A2(n5387), .ZN(n5386) );
  INV_X1 U6784 ( .A(n7337), .ZN(n5388) );
  INV_X1 U6785 ( .A(n5387), .ZN(n7336) );
  NAND2_X1 U6786 ( .A1(n5388), .A2(n7336), .ZN(n5389) );
  INV_X1 U6787 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5393) );
  MUX2_X1 U6788 ( .A(n5393), .B(n10239), .S(n4479), .Z(n5394) );
  INV_X1 U6789 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6790 ( .A1(n5395), .A2(SI_9_), .ZN(n5396) );
  XNOR2_X1 U6791 ( .A(n5420), .B(n4521), .ZN(n6493) );
  NAND2_X1 U6792 ( .A1(n6493), .A2(n8848), .ZN(n5400) );
  NAND2_X1 U6793 ( .A1(n5397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5398) );
  XNOR2_X1 U6794 ( .A(n5398), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U6795 ( .A1(n8838), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5538), .B2(
        n6647), .ZN(n5399) );
  AND2_X2 U6796 ( .A1(n5400), .A2(n5399), .ZN(n9933) );
  NAND2_X1 U6797 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  AND2_X1 U6798 ( .A1(n5436), .A2(n5404), .ZN(n9846) );
  NAND2_X1 U6799 ( .A1(n5958), .A2(n9846), .ZN(n5408) );
  NAND2_X1 U6800 ( .A1(n5278), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6801 ( .A1(n8851), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6802 ( .A1(n8841), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5405) );
  NAND4_X1 U6803 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n9071)
         );
  NAND2_X1 U6804 ( .A1(n9071), .A2(n5634), .ZN(n5409) );
  OAI21_X1 U6805 ( .B1(n9933), .B2(n5401), .A(n5409), .ZN(n5410) );
  XNOR2_X1 U6806 ( .A(n5410), .B(n5327), .ZN(n5413) );
  OR2_X1 U6807 ( .A1(n9933), .A2(n5951), .ZN(n5412) );
  NAND2_X1 U6808 ( .A1(n9071), .A2(n5713), .ZN(n5411) );
  AND2_X1 U6809 ( .A1(n5412), .A2(n5411), .ZN(n5414) );
  NAND2_X1 U6810 ( .A1(n5413), .A2(n5414), .ZN(n5419) );
  INV_X1 U6811 ( .A(n5413), .ZN(n5416) );
  INV_X1 U6812 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6813 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  NAND2_X1 U6814 ( .A1(n5419), .A2(n5417), .ZN(n7419) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5423) );
  MUX2_X1 U6816 ( .A(n5423), .B(n6563), .S(n4479), .Z(n5425) );
  INV_X1 U6817 ( .A(SI_10_), .ZN(n5424) );
  INV_X1 U6818 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U6819 ( .A1(n5426), .A2(SI_10_), .ZN(n5427) );
  NAND2_X1 U6820 ( .A1(n6496), .A2(n8848), .ZN(n5434) );
  NAND2_X1 U6821 ( .A1(n5431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5429) );
  MUX2_X1 U6822 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5429), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5430) );
  INV_X1 U6823 ( .A(n5430), .ZN(n5432) );
  NOR2_X1 U6824 ( .A1(n5432), .A2(n5532), .ZN(n6735) );
  AOI22_X1 U6825 ( .A1(n8838), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5538), .B2(
        n6735), .ZN(n5433) );
  NAND2_X1 U6826 ( .A1(n9140), .A2(n5953), .ZN(n5443) );
  INV_X1 U6827 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6828 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  AND2_X1 U6829 ( .A1(n5459), .A2(n5437), .ZN(n7449) );
  NAND2_X1 U6830 ( .A1(n5958), .A2(n7449), .ZN(n5441) );
  NAND2_X1 U6831 ( .A1(n5278), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6832 ( .A1(n8851), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6833 ( .A1(n8841), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5438) );
  NAND4_X1 U6834 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n9633)
         );
  NAND2_X1 U6835 ( .A1(n9633), .A2(n5634), .ZN(n5442) );
  NAND2_X1 U6836 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  XNOR2_X1 U6837 ( .A(n5444), .B(n6815), .ZN(n5447) );
  NAND2_X1 U6838 ( .A1(n9140), .A2(n5634), .ZN(n5446) );
  NAND2_X1 U6839 ( .A1(n9633), .A2(n5713), .ZN(n5445) );
  NAND2_X1 U6840 ( .A1(n5446), .A2(n5445), .ZN(n5448) );
  NAND2_X1 U6841 ( .A1(n5447), .A2(n5448), .ZN(n7428) );
  INV_X1 U6842 ( .A(n5447), .ZN(n5450) );
  INV_X1 U6843 ( .A(n5448), .ZN(n5449) );
  NAND2_X1 U6844 ( .A1(n5450), .A2(n5449), .ZN(n7427) );
  INV_X1 U6845 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5452) );
  MUX2_X1 U6846 ( .A(n5452), .B(n6587), .S(n4479), .Z(n5473) );
  XNOR2_X1 U6847 ( .A(n5475), .B(n5472), .ZN(n6532) );
  NAND2_X1 U6848 ( .A1(n6532), .A2(n8848), .ZN(n5456) );
  OR2_X1 U6849 ( .A1(n5532), .A2(n5453), .ZN(n5454) );
  XNOR2_X1 U6850 ( .A(n5454), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6738) );
  AOI22_X1 U6851 ( .A1(n8838), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5538), .B2(
        n6738), .ZN(n5455) );
  NAND2_X1 U6852 ( .A1(n5278), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5464) );
  INV_X1 U6853 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6854 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  AND2_X1 U6855 ( .A1(n5488), .A2(n5460), .ZN(n9628) );
  NAND2_X1 U6856 ( .A1(n5958), .A2(n9628), .ZN(n5463) );
  NAND2_X1 U6857 ( .A1(n8851), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6858 ( .A1(n8841), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5461) );
  NAND4_X1 U6859 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n9462)
         );
  OAI22_X1 U6860 ( .A1(n9668), .A2(n5401), .B1(n9143), .B2(n5951), .ZN(n5465)
         );
  XNOR2_X1 U6861 ( .A(n5465), .B(n6815), .ZN(n5470) );
  OR2_X1 U6862 ( .A1(n9668), .A2(n5951), .ZN(n5467) );
  NAND2_X1 U6863 ( .A1(n9462), .A2(n5713), .ZN(n5466) );
  NAND2_X1 U6864 ( .A1(n5467), .A2(n5466), .ZN(n5469) );
  XNOR2_X1 U6865 ( .A(n5470), .B(n5469), .ZN(n7514) );
  INV_X1 U6866 ( .A(n7514), .ZN(n5468) );
  NAND2_X1 U6867 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  INV_X1 U6868 ( .A(n5473), .ZN(n5474) );
  INV_X1 U6869 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5476) );
  INV_X1 U6870 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6670) );
  MUX2_X1 U6871 ( .A(n5476), .B(n6670), .S(n4479), .Z(n5478) );
  INV_X1 U6872 ( .A(SI_12_), .ZN(n5477) );
  INV_X1 U6873 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U6874 ( .A1(n5479), .A2(SI_12_), .ZN(n5480) );
  NAND2_X1 U6875 ( .A1(n6637), .A2(n8848), .ZN(n5485) );
  INV_X1 U6876 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6877 ( .A1(n5532), .A2(n5529), .ZN(n5481) );
  NAND2_X1 U6878 ( .A1(n5481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6879 ( .A1(n5482), .A2(n10479), .ZN(n5508) );
  OR2_X1 U6880 ( .A1(n5482), .A2(n10479), .ZN(n5483) );
  AOI22_X1 U6881 ( .A1(n8838), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5538), .B2(
        n9094), .ZN(n5484) );
  NAND2_X1 U6882 ( .A1(n9471), .A2(n5953), .ZN(n5495) );
  NAND2_X1 U6883 ( .A1(n5278), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5493) );
  INV_X1 U6884 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6885 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  AND2_X1 U6886 ( .A1(n5513), .A2(n5489), .ZN(n9467) );
  NAND2_X1 U6887 ( .A1(n5958), .A2(n9467), .ZN(n5492) );
  NAND2_X1 U6888 ( .A1(n8851), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6889 ( .A1(n8841), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5490) );
  NAND4_X1 U6890 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n9634)
         );
  NAND2_X1 U6891 ( .A1(n9634), .A2(n5634), .ZN(n5494) );
  NAND2_X1 U6892 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  XNOR2_X1 U6893 ( .A(n5496), .B(n6815), .ZN(n5498) );
  AND2_X1 U6894 ( .A1(n9634), .A2(n5713), .ZN(n5497) );
  AOI21_X1 U6895 ( .B1(n9471), .B2(n5634), .A(n5497), .ZN(n5499) );
  XNOR2_X1 U6896 ( .A(n5498), .B(n5499), .ZN(n8665) );
  INV_X1 U6897 ( .A(n5498), .ZN(n5500) );
  INV_X1 U6898 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5504) );
  MUX2_X1 U6899 ( .A(n5504), .B(n10236), .S(n4479), .Z(n5505) );
  INV_X1 U6900 ( .A(SI_13_), .ZN(n10296) );
  NAND2_X1 U6901 ( .A1(n5505), .A2(n10296), .ZN(n5527) );
  INV_X1 U6902 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U6903 ( .A1(n5506), .A2(SI_13_), .ZN(n5507) );
  XNOR2_X1 U6904 ( .A(n5526), .B(n5106), .ZN(n6680) );
  NAND2_X1 U6905 ( .A1(n6680), .A2(n8848), .ZN(n5511) );
  NAND2_X1 U6906 ( .A1(n5508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5509) );
  XNOR2_X1 U6907 ( .A(n5509), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U6908 ( .A1(n8838), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5538), .B2(
        n9746), .ZN(n5510) );
  NAND2_X1 U6909 ( .A1(n9452), .A2(n5953), .ZN(n5520) );
  INV_X1 U6910 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6911 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  AND2_X1 U6912 ( .A1(n5542), .A2(n5514), .ZN(n9451) );
  NAND2_X1 U6913 ( .A1(n5958), .A2(n9451), .ZN(n5518) );
  NAND2_X1 U6914 ( .A1(n5278), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6915 ( .A1(n8851), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6916 ( .A1(n8841), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5515) );
  NAND4_X1 U6917 ( .A1(n5518), .A2(n5517), .A3(n5516), .A4(n5515), .ZN(n9461)
         );
  NAND2_X1 U6918 ( .A1(n9461), .A2(n5634), .ZN(n5519) );
  NAND2_X1 U6919 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  XNOR2_X1 U6920 ( .A(n5521), .B(n5327), .ZN(n8719) );
  AND2_X1 U6921 ( .A1(n9461), .A2(n5713), .ZN(n5522) );
  AOI21_X1 U6922 ( .B1(n9452), .B2(n5634), .A(n5522), .ZN(n8718) );
  INV_X1 U6923 ( .A(n8719), .ZN(n5524) );
  INV_X1 U6924 ( .A(n8718), .ZN(n5523) );
  NAND2_X1 U6925 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  MUX2_X1 U6926 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4479), .Z(n5553) );
  INV_X1 U6927 ( .A(SI_14_), .ZN(n10248) );
  NAND2_X1 U6928 ( .A1(n6700), .A2(n8848), .ZN(n5540) );
  AND3_X1 U6929 ( .A1(n10479), .A2(n5530), .A3(n5529), .ZN(n5531) );
  AND2_X1 U6930 ( .A1(n5532), .A2(n5531), .ZN(n5535) );
  NOR2_X1 U6931 ( .A1(n5535), .A2(n5453), .ZN(n5533) );
  MUX2_X1 U6932 ( .A(n5453), .B(n5533), .S(P1_IR_REG_14__SCAN_IN), .Z(n5534)
         );
  INV_X1 U6933 ( .A(n5534), .ZN(n5536) );
  NAND2_X1 U6934 ( .A1(n5535), .A2(n10247), .ZN(n5593) );
  NAND2_X1 U6935 ( .A1(n5536), .A2(n5593), .ZN(n9761) );
  INV_X1 U6936 ( .A(n9761), .ZN(n5537) );
  AOI22_X1 U6937 ( .A1(n8838), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5538), .B2(
        n5537), .ZN(n5539) );
  NAND2_X1 U6938 ( .A1(n9150), .A2(n5953), .ZN(n5549) );
  NAND2_X1 U6939 ( .A1(n5278), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5547) );
  INV_X1 U6940 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U6941 ( .A1(n5542), .A2(n8630), .ZN(n5543) );
  AND2_X1 U6942 ( .A1(n5565), .A2(n5543), .ZN(n9430) );
  NAND2_X1 U6943 ( .A1(n5958), .A2(n9430), .ZN(n5546) );
  NAND2_X1 U6944 ( .A1(n8851), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6945 ( .A1(n8841), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5544) );
  NAND4_X1 U6946 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n9418)
         );
  NAND2_X1 U6947 ( .A1(n9418), .A2(n5634), .ZN(n5548) );
  NAND2_X1 U6948 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  XNOR2_X1 U6949 ( .A(n5550), .B(n5327), .ZN(n8628) );
  AND2_X1 U6950 ( .A1(n9418), .A2(n5713), .ZN(n5551) );
  AOI21_X1 U6951 ( .B1(n9150), .B2(n5634), .A(n5551), .ZN(n5574) );
  NAND2_X1 U6952 ( .A1(n8628), .A2(n5574), .ZN(n5582) );
  NAND2_X1 U6953 ( .A1(n5553), .A2(SI_14_), .ZN(n5554) );
  INV_X1 U6954 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5557) );
  INV_X1 U6955 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6790) );
  MUX2_X1 U6956 ( .A(n5557), .B(n6790), .S(n4479), .Z(n5558) );
  INV_X1 U6957 ( .A(SI_15_), .ZN(n10276) );
  INV_X1 U6958 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U6959 ( .A1(n5559), .A2(SI_15_), .ZN(n5560) );
  XNOR2_X1 U6960 ( .A(n5588), .B(n5587), .ZN(n6751) );
  NAND2_X1 U6961 ( .A1(n6751), .A2(n8848), .ZN(n5563) );
  NAND2_X1 U6962 ( .A1(n5593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5561) );
  XNOR2_X1 U6963 ( .A(n5561), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9775) );
  AOI22_X1 U6964 ( .A1(n8838), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5538), .B2(
        n9775), .ZN(n5562) );
  NAND2_X1 U6965 ( .A1(n9565), .A2(n5953), .ZN(n5572) );
  INV_X1 U6966 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U6967 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  AND2_X1 U6968 ( .A1(n5598), .A2(n5566), .ZN(n9411) );
  NAND2_X1 U6969 ( .A1(n5958), .A2(n9411), .ZN(n5570) );
  NAND2_X1 U6970 ( .A1(n5278), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6971 ( .A1(n8851), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6972 ( .A1(n8841), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5567) );
  NAND4_X1 U6973 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n9427)
         );
  NAND2_X1 U6974 ( .A1(n9427), .A2(n5634), .ZN(n5571) );
  NAND2_X1 U6975 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  XNOR2_X1 U6976 ( .A(n5573), .B(n5327), .ZN(n5581) );
  INV_X1 U6977 ( .A(n8628), .ZN(n5575) );
  INV_X1 U6978 ( .A(n5574), .ZN(n8627) );
  NAND2_X1 U6979 ( .A1(n5575), .A2(n8627), .ZN(n5579) );
  AND2_X1 U6980 ( .A1(n5581), .A2(n5579), .ZN(n5576) );
  NAND2_X1 U6981 ( .A1(n9565), .A2(n5634), .ZN(n5578) );
  NAND2_X1 U6982 ( .A1(n9427), .A2(n5713), .ZN(n5577) );
  NAND2_X1 U6983 ( .A1(n5578), .A2(n5577), .ZN(n8763) );
  NAND2_X1 U6984 ( .A1(n8761), .A2(n8763), .ZN(n8684) );
  INV_X1 U6985 ( .A(n8626), .ZN(n5580) );
  NAND2_X1 U6986 ( .A1(n5580), .A2(n5579), .ZN(n5585) );
  INV_X1 U6987 ( .A(n5581), .ZN(n5583) );
  AND2_X1 U6988 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  INV_X1 U6989 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5589) );
  INV_X1 U6990 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10445) );
  MUX2_X1 U6991 ( .A(n5589), .B(n10445), .S(n4479), .Z(n5590) );
  INV_X1 U6992 ( .A(SI_16_), .ZN(n10444) );
  NAND2_X1 U6993 ( .A1(n5590), .A2(n10444), .ZN(n5616) );
  INV_X1 U6994 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U6995 ( .A1(n5591), .A2(SI_16_), .ZN(n5592) );
  XNOR2_X1 U6996 ( .A(n5615), .B(n5614), .ZN(n6776) );
  NAND2_X1 U6997 ( .A1(n6776), .A2(n8848), .ZN(n5596) );
  OR2_X1 U6998 ( .A1(n5593), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6999 ( .A1(n5594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U7000 ( .A(n5620), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9789) );
  AOI22_X1 U7001 ( .A1(n8838), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5538), .B2(
        n9789), .ZN(n5595) );
  NAND2_X1 U7002 ( .A1(n9561), .A2(n5953), .ZN(n5605) );
  NAND2_X1 U7003 ( .A1(n5278), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5603) );
  INV_X1 U7004 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U7005 ( .A1(n5598), .A2(n9781), .ZN(n5599) );
  AND2_X1 U7006 ( .A1(n5628), .A2(n5599), .ZN(n9397) );
  NAND2_X1 U7007 ( .A1(n5958), .A2(n9397), .ZN(n5602) );
  NAND2_X1 U7008 ( .A1(n8851), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7009 ( .A1(n8841), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5600) );
  NAND4_X1 U7010 ( .A1(n5603), .A2(n5602), .A3(n5601), .A4(n5600), .ZN(n9419)
         );
  NAND2_X1 U7011 ( .A1(n9419), .A2(n5634), .ZN(n5604) );
  NAND2_X1 U7012 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  XNOR2_X1 U7013 ( .A(n5606), .B(n5327), .ZN(n5608) );
  AND2_X1 U7014 ( .A1(n9419), .A2(n5713), .ZN(n5607) );
  AOI21_X1 U7015 ( .B1(n9561), .B2(n5634), .A(n5607), .ZN(n5609) );
  NAND2_X1 U7016 ( .A1(n5608), .A2(n5609), .ZN(n5613) );
  INV_X1 U7017 ( .A(n5608), .ZN(n5611) );
  INV_X1 U7018 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7019 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  AND2_X1 U7020 ( .A1(n5613), .A2(n5612), .ZN(n8683) );
  NAND3_X1 U7021 ( .A1(n8684), .A2(n8682), .A3(n8683), .ZN(n8681) );
  NAND2_X1 U7022 ( .A1(n8681), .A2(n5613), .ZN(n8691) );
  INV_X1 U7023 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5618) );
  INV_X1 U7024 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6847) );
  MUX2_X1 U7025 ( .A(n5618), .B(n6847), .S(n4479), .Z(n5644) );
  XNOR2_X1 U7026 ( .A(n5644), .B(SI_17_), .ZN(n5643) );
  XNOR2_X1 U7027 ( .A(n5647), .B(n5643), .ZN(n6831) );
  NAND2_X1 U7028 ( .A1(n6831), .A2(n8848), .ZN(n5626) );
  AOI21_X1 U7029 ( .B1(n5620), .B2(n5619), .A(n5453), .ZN(n5621) );
  NAND2_X1 U7030 ( .A1(n5621), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5624) );
  INV_X1 U7031 ( .A(n5621), .ZN(n5623) );
  NAND2_X1 U7032 ( .A1(n5623), .A2(n5622), .ZN(n5648) );
  AOI22_X1 U7033 ( .A1(n9114), .A2(n5538), .B1(n8838), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7034 ( .A1(n9555), .A2(n5953), .ZN(n5636) );
  INV_X1 U7035 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7036 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  AND2_X1 U7037 ( .A1(n5655), .A2(n5629), .ZN(n9383) );
  NAND2_X1 U7038 ( .A1(n5958), .A2(n9383), .ZN(n5633) );
  NAND2_X1 U7039 ( .A1(n5278), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7040 ( .A1(n8851), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7041 ( .A1(n8841), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5630) );
  NAND4_X1 U7042 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5630), .ZN(n9403)
         );
  NAND2_X1 U7043 ( .A1(n9403), .A2(n5634), .ZN(n5635) );
  NAND2_X1 U7044 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  XNOR2_X1 U7045 ( .A(n5637), .B(n6815), .ZN(n5639) );
  AND2_X1 U7046 ( .A1(n9403), .A2(n5713), .ZN(n5638) );
  AOI21_X1 U7047 ( .B1(n9555), .B2(n5634), .A(n5638), .ZN(n5640) );
  XNOR2_X1 U7048 ( .A(n5639), .B(n5640), .ZN(n8693) );
  INV_X1 U7049 ( .A(n5639), .ZN(n5641) );
  NAND2_X1 U7050 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  INV_X1 U7051 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7052 ( .A1(n5645), .A2(SI_17_), .ZN(n5646) );
  MUX2_X1 U7053 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4479), .Z(n5670) );
  XNOR2_X1 U7054 ( .A(n5670), .B(SI_18_), .ZN(n5668) );
  XNOR2_X1 U7055 ( .A(n5669), .B(n5668), .ZN(n6958) );
  NAND2_X1 U7056 ( .A1(n6958), .A2(n8848), .ZN(n5652) );
  NAND2_X1 U7057 ( .A1(n5648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5649) );
  XNOR2_X1 U7058 ( .A(n5649), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9104) );
  INV_X1 U7059 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10326) );
  NOR2_X1 U7060 ( .A1(n5377), .A2(n10326), .ZN(n5650) );
  AOI21_X1 U7061 ( .B1(n9104), .B2(n5538), .A(n5650), .ZN(n5651) );
  NAND2_X1 U7062 ( .A1(n9548), .A2(n5953), .ZN(n5662) );
  NAND2_X1 U7063 ( .A1(n5278), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5660) );
  INV_X1 U7064 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7065 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  AND2_X1 U7066 ( .A1(n5677), .A2(n5656), .ZN(n9373) );
  NAND2_X1 U7067 ( .A1(n5958), .A2(n9373), .ZN(n5659) );
  NAND2_X1 U7068 ( .A1(n8851), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7069 ( .A1(n8841), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5657) );
  NAND4_X1 U7070 ( .A1(n5660), .A2(n5659), .A3(n5658), .A4(n5657), .ZN(n9389)
         );
  NAND2_X1 U7071 ( .A1(n9389), .A2(n5634), .ZN(n5661) );
  NAND2_X1 U7072 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  XNOR2_X1 U7073 ( .A(n5663), .B(n5327), .ZN(n5666) );
  NAND2_X1 U7074 ( .A1(n9548), .A2(n5634), .ZN(n5665) );
  NAND2_X1 U7075 ( .A1(n9389), .A2(n5713), .ZN(n5664) );
  NAND2_X1 U7076 ( .A1(n5665), .A2(n5664), .ZN(n8737) );
  INV_X1 U7077 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5671) );
  INV_X1 U7078 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10330) );
  MUX2_X1 U7079 ( .A(n5671), .B(n10330), .S(n4479), .Z(n5672) );
  INV_X1 U7080 ( .A(SI_19_), .ZN(n10355) );
  NAND2_X1 U7081 ( .A1(n5672), .A2(n10355), .ZN(n5692) );
  INV_X1 U7082 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7083 ( .A1(n5673), .A2(SI_19_), .ZN(n5674) );
  NAND2_X1 U7084 ( .A1(n5692), .A2(n5674), .ZN(n5693) );
  XNOR2_X1 U7085 ( .A(n5694), .B(n5693), .ZN(n7002) );
  NAND2_X1 U7086 ( .A1(n7002), .A2(n8848), .ZN(n5676) );
  AOI22_X1 U7087 ( .A1(n8838), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9863), .B2(
        n5538), .ZN(n5675) );
  NAND2_X1 U7088 ( .A1(n9542), .A2(n5953), .ZN(n5684) );
  NAND2_X1 U7089 ( .A1(n5278), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5682) );
  INV_X1 U7090 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U7091 ( .A1(n5677), .A2(n8650), .ZN(n5678) );
  AND2_X1 U7092 ( .A1(n5705), .A2(n5678), .ZN(n9350) );
  NAND2_X1 U7093 ( .A1(n5958), .A2(n9350), .ZN(n5681) );
  NAND2_X1 U7094 ( .A1(n8851), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7095 ( .A1(n8841), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5679) );
  NAND4_X1 U7096 ( .A1(n5682), .A2(n5681), .A3(n5680), .A4(n5679), .ZN(n9369)
         );
  NAND2_X1 U7097 ( .A1(n9369), .A2(n5634), .ZN(n5683) );
  NAND2_X1 U7098 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  XNOR2_X1 U7099 ( .A(n5685), .B(n5327), .ZN(n5687) );
  AND2_X1 U7100 ( .A1(n9369), .A2(n5713), .ZN(n5686) );
  AOI21_X1 U7101 ( .B1(n9542), .B2(n5634), .A(n5686), .ZN(n5688) );
  NAND2_X1 U7102 ( .A1(n5687), .A2(n5688), .ZN(n8710) );
  INV_X1 U7103 ( .A(n5687), .ZN(n5690) );
  INV_X1 U7104 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U7105 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  OAI21_X1 U7106 ( .B1(n8646), .B2(n8740), .A(n8647), .ZN(n8645) );
  INV_X1 U7107 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5695) );
  INV_X1 U7108 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7068) );
  MUX2_X1 U7109 ( .A(n5695), .B(n7068), .S(n4479), .Z(n5697) );
  INV_X1 U7110 ( .A(SI_20_), .ZN(n5696) );
  NAND2_X1 U7111 ( .A1(n5697), .A2(n5696), .ZN(n5724) );
  INV_X1 U7112 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7113 ( .A1(n5698), .A2(SI_20_), .ZN(n5699) );
  XNOR2_X1 U7114 ( .A(n5723), .B(n5722), .ZN(n7066) );
  NAND2_X1 U7115 ( .A1(n7066), .A2(n8848), .ZN(n5701) );
  NAND2_X1 U7116 ( .A1(n8838), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7117 ( .A1(n9537), .A2(n5953), .ZN(n5711) );
  INV_X1 U7118 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7119 ( .A1(n8851), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7120 ( .A1(n8841), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5702) );
  AND2_X1 U7121 ( .A1(n5703), .A2(n5702), .ZN(n5708) );
  INV_X1 U7122 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U7123 ( .A1(n5705), .A2(n8712), .ZN(n5706) );
  NAND2_X1 U7124 ( .A1(n5727), .A2(n5706), .ZN(n9336) );
  OR2_X1 U7125 ( .A1(n5852), .A2(n9336), .ZN(n5707) );
  OAI211_X1 U7126 ( .C1(n5962), .C2(n5709), .A(n5708), .B(n5707), .ZN(n9358)
         );
  NAND2_X1 U7127 ( .A1(n9358), .A2(n5634), .ZN(n5710) );
  NAND2_X1 U7128 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  XNOR2_X1 U7129 ( .A(n5712), .B(n5327), .ZN(n5715) );
  AND2_X1 U7130 ( .A1(n9358), .A2(n5713), .ZN(n5714) );
  AOI21_X1 U7131 ( .B1(n9537), .B2(n5634), .A(n5714), .ZN(n5716) );
  NAND2_X1 U7132 ( .A1(n5715), .A2(n5716), .ZN(n5720) );
  INV_X1 U7133 ( .A(n5715), .ZN(n5718) );
  INV_X1 U7134 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7135 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  NAND2_X1 U7136 ( .A1(n5720), .A2(n5719), .ZN(n8709) );
  AOI21_X1 U7137 ( .B1(n8645), .B2(n8710), .A(n8709), .ZN(n8708) );
  INV_X1 U7138 ( .A(n5720), .ZN(n5721) );
  MUX2_X1 U7139 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4479), .Z(n5741) );
  INV_X1 U7140 ( .A(SI_21_), .ZN(n10486) );
  XNOR2_X1 U7141 ( .A(n5741), .B(n10486), .ZN(n5740) );
  XNOR2_X1 U7142 ( .A(n5739), .B(n5740), .ZN(n7607) );
  NAND2_X1 U7143 ( .A1(n7607), .A2(n8848), .ZN(n5726) );
  NAND2_X1 U7144 ( .A1(n8838), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7145 ( .A1(n9532), .A2(n5953), .ZN(n5733) );
  INV_X1 U7146 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U7147 ( .A1(n5727), .A2(n8658), .ZN(n5728) );
  NAND2_X1 U7148 ( .A1(n5752), .A2(n5728), .ZN(n9321) );
  OR2_X1 U7149 ( .A1(n9321), .A2(n5852), .ZN(n5731) );
  AOI22_X1 U7150 ( .A1(n5278), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n8851), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7151 ( .A1(n8841), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5729) );
  INV_X1 U7152 ( .A(n9160), .ZN(n9343) );
  NAND2_X1 U7153 ( .A1(n9343), .A2(n5634), .ZN(n5732) );
  NAND2_X1 U7154 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  XNOR2_X1 U7155 ( .A(n5734), .B(n6815), .ZN(n5735) );
  INV_X1 U7156 ( .A(n5713), .ZN(n5882) );
  OAI22_X1 U7157 ( .A1(n9161), .A2(n5951), .B1(n9160), .B2(n5882), .ZN(n5736)
         );
  XNOR2_X1 U7158 ( .A(n5735), .B(n5736), .ZN(n8656) );
  INV_X1 U7159 ( .A(n5735), .ZN(n5738) );
  INV_X1 U7160 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7161 ( .A1(n5741), .A2(SI_21_), .ZN(n5742) );
  INV_X1 U7162 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5745) );
  INV_X1 U7163 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5744) );
  MUX2_X1 U7164 ( .A(n5745), .B(n5744), .S(n4479), .Z(n5747) );
  INV_X1 U7165 ( .A(SI_22_), .ZN(n5746) );
  NAND2_X1 U7166 ( .A1(n5747), .A2(n5746), .ZN(n5763) );
  INV_X1 U7167 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7168 ( .A1(n5748), .A2(SI_22_), .ZN(n5749) );
  NAND2_X1 U7169 ( .A1(n5763), .A2(n5749), .ZN(n5764) );
  XNOR2_X1 U7170 ( .A(n5765), .B(n5764), .ZN(n7614) );
  NAND2_X1 U7171 ( .A1(n7614), .A2(n8848), .ZN(n5751) );
  NAND2_X1 U7172 ( .A1(n8838), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5750) );
  INV_X1 U7173 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U7174 ( .A1(n5752), .A2(n8729), .ZN(n5753) );
  NAND2_X1 U7175 ( .A1(n5778), .A2(n5753), .ZN(n8732) );
  INV_X1 U7176 ( .A(n8732), .ZN(n9307) );
  NAND2_X1 U7177 ( .A1(n9307), .A2(n5958), .ZN(n5759) );
  INV_X1 U7178 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7179 ( .A1(n8841), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7180 ( .A1(n8851), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U7181 ( .C1(n5962), .C2(n5756), .A(n5755), .B(n5754), .ZN(n5757)
         );
  INV_X1 U7182 ( .A(n5757), .ZN(n5758) );
  OAI22_X1 U7183 ( .A1(n9309), .A2(n5951), .B1(n9325), .B2(n5882), .ZN(n5761)
         );
  OAI22_X1 U7184 ( .A1(n9309), .A2(n5401), .B1(n9325), .B2(n5951), .ZN(n5760)
         );
  XOR2_X1 U7185 ( .A(n6815), .B(n5760), .Z(n8727) );
  INV_X1 U7186 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5767) );
  INV_X1 U7187 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5766) );
  MUX2_X1 U7188 ( .A(n5767), .B(n5766), .S(n4479), .Z(n5768) );
  INV_X1 U7189 ( .A(SI_23_), .ZN(n10345) );
  NAND2_X1 U7190 ( .A1(n5768), .A2(n10345), .ZN(n5788) );
  INV_X1 U7191 ( .A(n5768), .ZN(n5769) );
  NAND2_X1 U7192 ( .A1(n5769), .A2(SI_23_), .ZN(n5770) );
  OR2_X1 U7193 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U7194 ( .A1(n5789), .A2(n5773), .ZN(n7621) );
  NAND2_X1 U7195 ( .A1(n7621), .A2(n8848), .ZN(n5775) );
  NAND2_X1 U7196 ( .A1(n8838), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5774) );
  INV_X1 U7197 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7198 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  NAND2_X1 U7199 ( .A1(n5795), .A2(n5779), .ZN(n9297) );
  OR2_X1 U7200 ( .A1(n9297), .A2(n5852), .ZN(n5785) );
  INV_X1 U7201 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7202 ( .A1(n8841), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7203 ( .A1(n8851), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5780) );
  OAI211_X1 U7204 ( .C1(n5962), .C2(n5782), .A(n5781), .B(n5780), .ZN(n5783)
         );
  INV_X1 U7205 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U7206 ( .A1(n5785), .A2(n5784), .ZN(n9313) );
  OAI22_X1 U7207 ( .A1(n9301), .A2(n5401), .B1(n9280), .B2(n5951), .ZN(n5786)
         );
  XNOR2_X1 U7208 ( .A(n5786), .B(n6815), .ZN(n5812) );
  INV_X1 U7209 ( .A(n5812), .ZN(n5787) );
  OAI22_X1 U7210 ( .A1(n9301), .A2(n5951), .B1(n9280), .B2(n5882), .ZN(n8639)
         );
  NAND2_X1 U7211 ( .A1(n8637), .A2(n8639), .ZN(n8701) );
  INV_X1 U7212 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5790) );
  INV_X1 U7213 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10294) );
  MUX2_X1 U7214 ( .A(n5790), .B(n10294), .S(n4479), .Z(n5816) );
  XNOR2_X1 U7215 ( .A(n5816), .B(SI_24_), .ZN(n5815) );
  NAND2_X1 U7216 ( .A1(n7598), .A2(n8848), .ZN(n5792) );
  NAND2_X1 U7217 ( .A1(n8838), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5791) );
  INV_X1 U7218 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7219 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7220 ( .A1(n5826), .A2(n5796), .ZN(n9283) );
  OR2_X1 U7221 ( .A1(n9283), .A2(n5852), .ZN(n5802) );
  INV_X1 U7222 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7223 ( .A1(n8851), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7224 ( .A1(n8841), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5797) );
  OAI211_X1 U7225 ( .C1(n5962), .C2(n5799), .A(n5798), .B(n5797), .ZN(n5800)
         );
  INV_X1 U7226 ( .A(n5800), .ZN(n5801) );
  OAI22_X1 U7227 ( .A1(n9287), .A2(n5401), .B1(n9294), .B2(n5951), .ZN(n5803)
         );
  XNOR2_X1 U7228 ( .A(n5803), .B(n5327), .ZN(n5806) );
  NAND2_X1 U7229 ( .A1(n9266), .A2(n5713), .ZN(n5804) );
  NAND2_X1 U7230 ( .A1(n5806), .A2(n5807), .ZN(n5814) );
  INV_X1 U7231 ( .A(n5806), .ZN(n5809) );
  INV_X1 U7232 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7233 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U7234 ( .A1(n5813), .A2(n5812), .ZN(n8636) );
  INV_X1 U7235 ( .A(n5815), .ZN(n5819) );
  INV_X1 U7236 ( .A(n5816), .ZN(n5817) );
  NAND2_X1 U7237 ( .A1(n5817), .A2(SI_24_), .ZN(n5818) );
  INV_X1 U7238 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5820) );
  INV_X1 U7239 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7563) );
  MUX2_X1 U7240 ( .A(n5820), .B(n7563), .S(n6040), .Z(n5821) );
  INV_X1 U7241 ( .A(SI_25_), .ZN(n10429) );
  NAND2_X1 U7242 ( .A1(n5821), .A2(n10429), .ZN(n5839) );
  INV_X1 U7243 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7244 ( .A1(n5822), .A2(SI_25_), .ZN(n5823) );
  NAND2_X1 U7245 ( .A1(n5839), .A2(n5823), .ZN(n5840) );
  NAND2_X1 U7246 ( .A1(n7631), .A2(n8848), .ZN(n5825) );
  NAND2_X1 U7247 ( .A1(n8838), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5824) );
  INV_X1 U7248 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U7249 ( .A1(n5826), .A2(n8676), .ZN(n5827) );
  NAND2_X1 U7250 ( .A1(n9270), .A2(n5958), .ZN(n5833) );
  INV_X1 U7251 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7252 ( .A1(n8851), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7253 ( .A1(n8841), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5828) );
  OAI211_X1 U7254 ( .C1(n5830), .C2(n5962), .A(n5829), .B(n5828), .ZN(n5831)
         );
  INV_X1 U7255 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U7256 ( .A1(n9511), .A2(n5953), .ZN(n5835) );
  NAND2_X1 U7257 ( .A1(n9254), .A2(n5634), .ZN(n5834) );
  NAND2_X1 U7258 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XOR2_X1 U7259 ( .A(n5837), .B(n5838), .Z(n8674) );
  INV_X1 U7260 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5842) );
  INV_X1 U7261 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U7262 ( .A(n5842), .B(n7564), .S(n6040), .Z(n5843) );
  INV_X1 U7263 ( .A(SI_26_), .ZN(n10324) );
  NAND2_X1 U7264 ( .A1(n5843), .A2(n10324), .ZN(n5866) );
  INV_X1 U7265 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7266 ( .A1(n5844), .A2(SI_26_), .ZN(n5845) );
  AND2_X1 U7267 ( .A1(n5866), .A2(n5845), .ZN(n5864) );
  NAND2_X1 U7268 ( .A1(n7643), .A2(n8848), .ZN(n5847) );
  NAND2_X1 U7269 ( .A1(n8838), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5846) );
  INV_X1 U7270 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7271 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  NAND2_X1 U7272 ( .A1(n5928), .A2(n5851), .ZN(n8753) );
  INV_X1 U7273 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7274 ( .A1(n8841), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7275 ( .A1(n8851), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5853) );
  OAI211_X1 U7276 ( .C1(n5962), .C2(n5855), .A(n5854), .B(n5853), .ZN(n5856)
         );
  INV_X1 U7277 ( .A(n5856), .ZN(n5857) );
  OAI22_X1 U7278 ( .A1(n9251), .A2(n5401), .B1(n9167), .B2(n5951), .ZN(n5859)
         );
  XNOR2_X1 U7279 ( .A(n5859), .B(n6815), .ZN(n5863) );
  NAND2_X1 U7280 ( .A1(n9265), .A2(n5713), .ZN(n5860) );
  NAND2_X1 U7281 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7282 ( .A1(n5863), .A2(n5862), .ZN(n8748) );
  INV_X1 U7283 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5869) );
  INV_X1 U7284 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5868) );
  MUX2_X1 U7285 ( .A(n5869), .B(n5868), .S(n6040), .Z(n5870) );
  INV_X1 U7286 ( .A(SI_27_), .ZN(n10352) );
  NAND2_X1 U7287 ( .A1(n5870), .A2(n10352), .ZN(n5945) );
  INV_X1 U7288 ( .A(n5870), .ZN(n5871) );
  NAND2_X1 U7289 ( .A1(n5871), .A2(SI_27_), .ZN(n5872) );
  AND2_X1 U7290 ( .A1(n5945), .A2(n5872), .ZN(n5943) );
  NAND2_X1 U7291 ( .A1(n7595), .A2(n8848), .ZN(n5874) );
  NAND2_X1 U7292 ( .A1(n8838), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U7293 ( .A(n5928), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U7294 ( .A1(n9242), .A2(n5958), .ZN(n5880) );
  INV_X1 U7295 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7296 ( .A1(n8851), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7297 ( .A1(n8841), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5875) );
  OAI211_X1 U7298 ( .C1(n5962), .C2(n5877), .A(n5876), .B(n5875), .ZN(n5878)
         );
  INV_X1 U7299 ( .A(n5878), .ZN(n5879) );
  OAI22_X1 U7300 ( .A1(n9237), .A2(n5401), .B1(n9168), .B2(n5951), .ZN(n5881)
         );
  XNOR2_X1 U7301 ( .A(n5881), .B(n6815), .ZN(n5973) );
  INV_X1 U7302 ( .A(n5973), .ZN(n5884) );
  NOR2_X1 U7303 ( .A1(n9168), .A2(n5882), .ZN(n5883) );
  AOI21_X1 U7304 ( .B1(n9501), .B2(n5634), .A(n5883), .ZN(n5971) );
  XNOR2_X1 U7305 ( .A(n5884), .B(n5971), .ZN(n5885) );
  XNOR2_X1 U7306 ( .A(n5974), .B(n5885), .ZN(n5908) );
  AND2_X1 U7307 ( .A1(n8982), .A2(n9023), .ZN(n6813) );
  NAND2_X1 U7308 ( .A1(n9063), .A2(n8979), .ZN(n5980) );
  INV_X1 U7309 ( .A(n5980), .ZN(n6817) );
  OR2_X1 U7310 ( .A1(n9647), .A2(n6817), .ZN(n5912) );
  NAND2_X1 U7311 ( .A1(n5887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  INV_X1 U7312 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5888) );
  XNOR2_X1 U7313 ( .A(n5889), .B(n5888), .ZN(n7392) );
  AND2_X1 U7314 ( .A1(n7392), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7315 ( .A1(n5978), .A2(n5890), .ZN(n9881) );
  NOR2_X1 U7316 ( .A1(n5912), .A2(n9881), .ZN(n5907) );
  NAND2_X1 U7317 ( .A1(n7561), .A2(P1_B_REG_SCAN_IN), .ZN(n5891) );
  MUX2_X1 U7318 ( .A(P1_B_REG_SCAN_IN), .B(n5891), .S(n7472), .Z(n5892) );
  NAND2_X1 U7319 ( .A1(n5892), .A2(n5905), .ZN(n5906) );
  INV_X1 U7320 ( .A(n7561), .ZN(n5893) );
  OAI22_X1 U7321 ( .A1(n5906), .A2(P1_D_REG_1__SCAN_IN), .B1(n5905), .B2(n5893), .ZN(n6719) );
  INV_X1 U7322 ( .A(n6719), .ZN(n5904) );
  NOR4_X1 U7323 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5897) );
  NOR4_X1 U7324 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5896) );
  NOR4_X1 U7325 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5895) );
  NOR4_X1 U7326 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5894) );
  NAND4_X1 U7327 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n5903)
         );
  NOR2_X1 U7328 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5901) );
  NOR4_X1 U7329 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5900) );
  NOR4_X1 U7330 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5899) );
  NOR4_X1 U7331 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5898) );
  NAND4_X1 U7332 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5902)
         );
  INV_X1 U7333 ( .A(n5906), .ZN(n9587) );
  OAI21_X1 U7334 ( .B1(n5903), .B2(n5902), .A(n9587), .ZN(n6718) );
  AND2_X1 U7335 ( .A1(n5904), .A2(n6718), .ZN(n6808) );
  INV_X1 U7336 ( .A(n5905), .ZN(n7565) );
  NAND2_X1 U7337 ( .A1(n7565), .A2(n7472), .ZN(n9588) );
  OAI21_X1 U7338 ( .B1(n5906), .B2(P1_D_REG_0__SCAN_IN), .A(n9588), .ZN(n6806)
         );
  INV_X1 U7339 ( .A(n6806), .ZN(n6721) );
  NAND2_X1 U7340 ( .A1(n5908), .A2(n8751), .ZN(n5942) );
  NAND2_X1 U7341 ( .A1(n6813), .A2(n5909), .ZN(n6827) );
  NOR2_X1 U7342 ( .A1(n6827), .A2(n9881), .ZN(n5918) );
  NAND2_X1 U7343 ( .A1(n6676), .A2(n5918), .ZN(n5911) );
  NOR2_X1 U7344 ( .A1(n9881), .A2(n8979), .ZN(n5910) );
  INV_X1 U7345 ( .A(n5912), .ZN(n5913) );
  INV_X1 U7346 ( .A(n6676), .ZN(n5921) );
  NAND2_X1 U7347 ( .A1(n5913), .A2(n5921), .ZN(n5915) );
  OR2_X1 U7348 ( .A1(n5980), .A2(n5914), .ZN(n6809) );
  NAND4_X1 U7349 ( .A1(n5915), .A2(n5978), .A3(n7392), .A4(n6809), .ZN(n5916)
         );
  NAND2_X1 U7350 ( .A1(n5916), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7351 ( .A1(n5917), .A2(n5172), .ZN(n6816) );
  OR2_X1 U7352 ( .A1(n6816), .A2(n9881), .ZN(n9067) );
  INV_X1 U7353 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U7354 ( .A1(n9067), .A2(n5919), .ZN(n5920) );
  NAND2_X1 U7355 ( .A1(n5921), .A2(n5920), .ZN(n6674) );
  NAND2_X1 U7356 ( .A1(n5922), .A2(n6674), .ZN(n8764) );
  NOR2_X1 U7357 ( .A1(n9067), .A2(n5923), .ZN(n5924) );
  NAND2_X1 U7358 ( .A1(n6676), .A2(n5924), .ZN(n8755) );
  INV_X1 U7359 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5926) );
  OAI22_X1 U7360 ( .A1(n9167), .A2(n8755), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5926), .ZN(n5938) );
  INV_X1 U7361 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U7362 ( .B1(n5928), .B2(n5926), .A(n5925), .ZN(n5929) );
  NAND2_X1 U7363 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5927) );
  NAND2_X1 U7364 ( .A1(n9217), .A2(n5958), .ZN(n5935) );
  INV_X1 U7365 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7366 ( .A1(n8851), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7367 ( .A1(n8841), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U7368 ( .C1(n5962), .C2(n5932), .A(n5931), .B(n5930), .ZN(n5933)
         );
  INV_X1 U7369 ( .A(n5933), .ZN(n5934) );
  INV_X1 U7370 ( .A(n5923), .ZN(n9060) );
  NOR2_X1 U7371 ( .A1(n9067), .A2(n9060), .ZN(n5936) );
  INV_X1 U7372 ( .A(n8757), .ZN(n8768) );
  NOR2_X1 U7373 ( .A1(n9203), .A2(n8768), .ZN(n5937) );
  AOI211_X1 U7374 ( .C1(n9242), .C2(n8764), .A(n5938), .B(n5937), .ZN(n5939)
         );
  NAND2_X1 U7375 ( .A1(n5942), .A2(n5941), .ZN(P1_U3212) );
  MUX2_X1 U7376 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6040), .Z(n7587) );
  INV_X1 U7377 ( .A(SI_28_), .ZN(n7588) );
  XNOR2_X1 U7378 ( .A(n7587), .B(n7588), .ZN(n7585) );
  NAND2_X1 U7379 ( .A1(n7719), .A2(n8848), .ZN(n5947) );
  NAND2_X1 U7380 ( .A1(n8838), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7381 ( .A1(n9495), .A2(n5634), .ZN(n5949) );
  NAND2_X1 U7382 ( .A1(n9169), .A2(n5713), .ZN(n5948) );
  NAND2_X1 U7383 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  XNOR2_X1 U7384 ( .A(n5950), .B(n6815), .ZN(n5955) );
  NOR2_X1 U7385 ( .A1(n9203), .A2(n5951), .ZN(n5952) );
  AOI21_X1 U7386 ( .B1(n9495), .B2(n5953), .A(n5952), .ZN(n5954) );
  XNOR2_X1 U7387 ( .A(n5955), .B(n5954), .ZN(n5976) );
  INV_X1 U7388 ( .A(n5976), .ZN(n5956) );
  NAND2_X1 U7389 ( .A1(n5956), .A2(n8751), .ZN(n5975) );
  INV_X1 U7390 ( .A(n5975), .ZN(n5970) );
  NOR2_X1 U7391 ( .A1(n9219), .A2(n8760), .ZN(n5969) );
  AOI22_X1 U7392 ( .A1(n9217), .A2(n8764), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5967) );
  INV_X1 U7393 ( .A(n5957), .ZN(n9207) );
  NAND2_X1 U7394 ( .A1(n9207), .A2(n5958), .ZN(n5965) );
  INV_X1 U7395 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7396 ( .A1(n8851), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7397 ( .A1(n8841), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5959) );
  OAI211_X1 U7398 ( .C1(n5962), .C2(n5961), .A(n5960), .B(n5959), .ZN(n5963)
         );
  INV_X1 U7399 ( .A(n5963), .ZN(n5964) );
  NAND2_X1 U7400 ( .A1(n5965), .A2(n5964), .ZN(n9227) );
  NAND2_X1 U7401 ( .A1(n9227), .A2(n8757), .ZN(n5966) );
  OAI211_X1 U7402 ( .C1(n9168), .C2(n8755), .A(n5967), .B(n5966), .ZN(n5968)
         );
  INV_X1 U7403 ( .A(n5971), .ZN(n5972) );
  INV_X1 U7404 ( .A(n7392), .ZN(n5979) );
  OR2_X1 U7405 ( .A1(n5978), .A2(n5979), .ZN(n6498) );
  OR2_X1 U7406 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  AND2_X1 U7407 ( .A1(n5981), .A2(n6498), .ZN(n6508) );
  NAND2_X1 U7408 ( .A1(n6508), .A2(n5982), .ZN(n6567) );
  NAND2_X1 U7409 ( .A1(n6567), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U7410 ( .A1(n5995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6024) );
  INV_X1 U7411 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7412 ( .A1(n6024), .A2(n6023), .ZN(n5992) );
  NAND2_X1 U7413 ( .A1(n5992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  INV_X1 U7414 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7415 ( .A1(n6007), .A2(n6006), .ZN(n6009) );
  NAND2_X1 U7416 ( .A1(n6009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5994) );
  INV_X1 U7417 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U7418 ( .A(n5994), .B(n5993), .ZN(n6339) );
  INV_X1 U7419 ( .A(n6339), .ZN(n7458) );
  NOR3_X1 U7420 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7421 ( .A1(n5999), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5998) );
  MUX2_X1 U7422 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5998), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6000) );
  AND2_X1 U7423 ( .A1(n6000), .A2(n4586), .ZN(n7526) );
  INV_X1 U7424 ( .A(n7526), .ZN(n6004) );
  NAND2_X1 U7425 ( .A1(n4586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  MUX2_X1 U7426 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6001), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6003) );
  INV_X1 U7427 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7428 ( .A1(n6003), .A2(n6033), .ZN(n6337) );
  NOR2_X1 U7429 ( .A1(n6004), .A2(n6337), .ZN(n6005) );
  OR2_X1 U7430 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U7431 ( .A1(n6009), .A2(n6008), .ZN(n6446) );
  INV_X1 U7432 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U7433 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7434 ( .A1(n6012), .A2(n6011), .ZN(n6014) );
  XNOR2_X2 U7435 ( .A(n6015), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6017) );
  INV_X1 U7436 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6915) );
  INV_X2 U7437 ( .A(n6017), .ZN(n6020) );
  INV_X1 U7438 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7439 ( .A1(n6085), .A2(n6016), .ZN(n6022) );
  INV_X1 U7440 ( .A(n6086), .ZN(n6019) );
  NAND2_X1 U7441 ( .A1(n6019), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7442 ( .A(n6024), .B(n6023), .ZN(n7880) );
  NAND2_X1 U7443 ( .A1(n7880), .A2(n8062), .ZN(n10008) );
  NAND2_X1 U7444 ( .A1(n4544), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6026) );
  MUX2_X1 U7445 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6026), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6028) );
  NAND2_X1 U7446 ( .A1(n6028), .A2(n6027), .ZN(n8024) );
  INV_X1 U7447 ( .A(n6029), .ZN(n6030) );
  NAND2_X1 U7448 ( .A1(n6030), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  INV_X1 U7449 ( .A(n8066), .ZN(n6032) );
  INV_X2 U7450 ( .A(n7877), .ZN(n7722) );
  NOR2_X1 U7451 ( .A1(n6884), .A2(n7722), .ZN(n6044) );
  INV_X1 U7452 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6034) );
  OR2_X1 U7453 ( .A1(n6036), .A2(n6195), .ZN(n6037) );
  NAND2_X1 U7454 ( .A1(n6039), .A2(n6038), .ZN(n6368) );
  NAND2_X2 U7455 ( .A1(n7567), .A2(n6368), .ZN(n6059) );
  NAND2_X1 U7456 ( .A1(n6326), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7457 ( .A1(n6404), .A2(n7120), .ZN(n6041) );
  INV_X1 U7458 ( .A(n7880), .ZN(n8069) );
  NAND2_X1 U7459 ( .A1(n8069), .A2(n9980), .ZN(n8027) );
  NAND3_X1 U7460 ( .A1(n10008), .A2(n8027), .A3(n8062), .ZN(n6043) );
  NAND2_X1 U7461 ( .A1(n7890), .A2(n8024), .ZN(n6883) );
  NAND2_X2 U7462 ( .A1(n6043), .A2(n6883), .ZN(n7660) );
  XNOR2_X1 U7463 ( .A(n6769), .B(n7660), .ZN(n6045) );
  NAND2_X1 U7464 ( .A1(n6044), .A2(n6045), .ZN(n6048) );
  INV_X1 U7465 ( .A(n6044), .ZN(n6047) );
  INV_X1 U7466 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7467 ( .A1(n6047), .A2(n6046), .ZN(n6061) );
  AND2_X1 U7468 ( .A1(n6048), .A2(n6061), .ZN(n6693) );
  INV_X1 U7469 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10234) );
  INV_X1 U7470 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6049) );
  INV_X1 U7471 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7472 ( .A1(n6085), .A2(n6050), .ZN(n6052) );
  NAND2_X1 U7473 ( .A1(n7637), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7474 ( .A1(n8088), .A2(n7877), .ZN(n6060) );
  NAND2_X1 U7475 ( .A1(n6468), .A2(SI_0_), .ZN(n6056) );
  INV_X1 U7476 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7477 ( .A1(n6056), .A2(n6055), .ZN(n6058) );
  AND2_X1 U7478 ( .A1(n6058), .A2(n6057), .ZN(n8625) );
  MUX2_X1 U7479 ( .A(n9960), .B(n8625), .S(n6059), .Z(n6768) );
  MUX2_X1 U7480 ( .A(n7660), .B(n6060), .S(n6768), .Z(n6692) );
  NAND2_X1 U7481 ( .A1(n6691), .A2(n6061), .ZN(n6713) );
  INV_X1 U7482 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10285) );
  OR2_X1 U7483 ( .A1(n7648), .A2(n10285), .ZN(n6066) );
  NAND2_X1 U7484 ( .A1(n6115), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6065) );
  INV_X1 U7485 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7134) );
  OR2_X1 U7486 ( .A1(n6274), .A2(n7134), .ZN(n6064) );
  INV_X1 U7487 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6062) );
  OR2_X1 U7488 ( .A1(n6085), .A2(n6062), .ZN(n6063) );
  OR2_X1 U7489 ( .A1(n6870), .A2(n7722), .ZN(n6071) );
  NAND2_X1 U7490 ( .A1(n6326), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7491 ( .A1(n6067), .A2(n6195), .ZN(n6068) );
  NAND2_X1 U7492 ( .A1(n6404), .A2(n9607), .ZN(n6069) );
  XNOR2_X1 U7493 ( .A(n6869), .B(n7723), .ZN(n6072) );
  XNOR2_X1 U7494 ( .A(n6071), .B(n6072), .ZN(n6712) );
  NAND2_X1 U7495 ( .A1(n6115), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6077) );
  OR2_X1 U7496 ( .A1(n7648), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6076) );
  INV_X1 U7497 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7129) );
  OR2_X1 U7498 ( .A1(n6274), .A2(n7129), .ZN(n6075) );
  INV_X1 U7499 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7500 ( .A1(n6085), .A2(n6073), .ZN(n6074) );
  OR2_X1 U7501 ( .A1(n6901), .A2(n7722), .ZN(n6082) );
  NAND2_X1 U7502 ( .A1(n6326), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7503 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6078), .ZN(n6079) );
  XNOR2_X1 U7504 ( .A(n6079), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U7505 ( .A1(n6404), .A2(n7149), .ZN(n6080) );
  OAI211_X1 U7506 ( .C1(n6149), .C2(n6478), .A(n6081), .B(n6080), .ZN(n6935)
         );
  XNOR2_X1 U7507 ( .A(n6935), .B(n7660), .ZN(n6083) );
  XNOR2_X1 U7508 ( .A(n6082), .B(n6083), .ZN(n6746) );
  INV_X1 U7509 ( .A(n6082), .ZN(n6084) );
  XNOR2_X1 U7510 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6907) );
  OR2_X1 U7511 ( .A1(n7648), .A2(n6907), .ZN(n6090) );
  INV_X1 U7512 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7128) );
  OR2_X1 U7513 ( .A1(n6274), .A2(n7128), .ZN(n6089) );
  INV_X1 U7514 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7515 ( .A1(n6086), .A2(n6087), .ZN(n6088) );
  OR2_X1 U7516 ( .A1(n7050), .A2(n7722), .ZN(n6096) );
  NAND2_X1 U7517 ( .A1(n7867), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6094) );
  INV_X1 U7518 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7519 ( .A1(n6108), .A2(n6195), .ZN(n6092) );
  XNOR2_X1 U7520 ( .A(n6092), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7226) );
  NAND2_X1 U7521 ( .A1(n6404), .A2(n7226), .ZN(n6093) );
  OAI211_X1 U7522 ( .C1(n6149), .C2(n6480), .A(n6094), .B(n6093), .ZN(n6904)
         );
  XNOR2_X1 U7523 ( .A(n6904), .B(n7723), .ZN(n6095) );
  NOR2_X1 U7524 ( .A1(n6096), .A2(n6095), .ZN(n6780) );
  NAND2_X1 U7525 ( .A1(n6096), .A2(n6095), .ZN(n6778) );
  NAND2_X1 U7526 ( .A1(n6097), .A2(n6778), .ZN(n6439) );
  NAND2_X1 U7527 ( .A1(n7737), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6106) );
  INV_X1 U7528 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6098) );
  OR2_X1 U7529 ( .A1(n6085), .A2(n6098), .ZN(n6105) );
  INV_X1 U7530 ( .A(n6099), .ZN(n6101) );
  INV_X1 U7531 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7532 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7533 ( .A1(n6118), .A2(n6102), .ZN(n9973) );
  OR2_X1 U7534 ( .A1(n7648), .A2(n9973), .ZN(n6104) );
  INV_X1 U7535 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7138) );
  OR2_X1 U7536 ( .A1(n6274), .A2(n7138), .ZN(n6103) );
  NOR2_X1 U7537 ( .A1(n6988), .A2(n7722), .ZN(n6111) );
  NAND2_X1 U7538 ( .A1(n7867), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6110) );
  INV_X1 U7539 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7540 ( .A1(n6108), .A2(n6107), .ZN(n6166) );
  NAND2_X1 U7541 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7542 ( .A(n6124), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7173) );
  NAND2_X1 U7543 ( .A1(n6404), .A2(n7173), .ZN(n6109) );
  XNOR2_X1 U7544 ( .A(n9975), .B(n7660), .ZN(n6979) );
  NAND2_X1 U7545 ( .A1(n6111), .A2(n6979), .ZN(n6129) );
  INV_X1 U7546 ( .A(n6111), .ZN(n6113) );
  INV_X1 U7547 ( .A(n6979), .ZN(n6112) );
  NAND2_X1 U7548 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7549 ( .A1(n6129), .A2(n6114), .ZN(n6440) );
  OR2_X1 U7550 ( .A1(n6439), .A2(n6440), .ZN(n6438) );
  NAND2_X1 U7551 ( .A1(n7737), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6123) );
  INV_X1 U7552 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6116) );
  OR2_X1 U7553 ( .A1(n6085), .A2(n6116), .ZN(n6122) );
  INV_X1 U7554 ( .A(n6118), .ZN(n6117) );
  NAND2_X1 U7555 ( .A1(n6117), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6138) );
  INV_X1 U7556 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U7557 ( .A1(n6118), .A2(n10341), .ZN(n6119) );
  NAND2_X1 U7558 ( .A1(n6138), .A2(n6119), .ZN(n6990) );
  OR2_X1 U7559 ( .A1(n7648), .A2(n6990), .ZN(n6121) );
  INV_X1 U7560 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7172) );
  OR2_X1 U7561 ( .A1(n6274), .A2(n7172), .ZN(n6120) );
  OR2_X1 U7562 ( .A1(n7049), .A2(n7722), .ZN(n6133) );
  NAND2_X1 U7563 ( .A1(n6185), .A2(n6484), .ZN(n6128) );
  NAND2_X1 U7564 ( .A1(n7867), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7565 ( .A1(n6124), .A2(n6163), .ZN(n6125) );
  NAND2_X1 U7566 ( .A1(n6125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7567 ( .A(n6144), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U7568 ( .A1(n6404), .A2(n7171), .ZN(n6126) );
  XNOR2_X1 U7569 ( .A(n10030), .B(n7660), .ZN(n6132) );
  XNOR2_X1 U7570 ( .A(n6133), .B(n6132), .ZN(n6980) );
  INV_X1 U7571 ( .A(n6129), .ZN(n6130) );
  NOR2_X1 U7572 ( .A1(n6980), .A2(n6130), .ZN(n6131) );
  NAND2_X1 U7573 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  NAND2_X1 U7574 ( .A1(n7737), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6143) );
  INV_X1 U7575 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7576 ( .A1(n6085), .A2(n6135), .ZN(n6142) );
  INV_X1 U7577 ( .A(n6138), .ZN(n6136) );
  NAND2_X1 U7578 ( .A1(n6136), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6156) );
  INV_X1 U7579 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7580 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U7581 ( .A1(n6156), .A2(n6139), .ZN(n7033) );
  OR2_X1 U7582 ( .A1(n7648), .A2(n7033), .ZN(n6141) );
  INV_X1 U7583 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7170) );
  OR2_X1 U7584 ( .A1(n6274), .A2(n7170), .ZN(n6140) );
  NOR2_X1 U7585 ( .A1(n7077), .A2(n7722), .ZN(n6150) );
  NAND2_X1 U7586 ( .A1(n6326), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6148) );
  INV_X1 U7587 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7588 ( .A1(n6144), .A2(n6164), .ZN(n6145) );
  NAND2_X1 U7589 ( .A1(n6145), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U7590 ( .A(n6146), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U7591 ( .A1(n6404), .A2(n7213), .ZN(n6147) );
  XNOR2_X1 U7592 ( .A(n10033), .B(n7660), .ZN(n6151) );
  NAND2_X1 U7593 ( .A1(n6150), .A2(n6151), .ZN(n6154) );
  INV_X1 U7594 ( .A(n6150), .ZN(n6152) );
  INV_X1 U7595 ( .A(n6151), .ZN(n7074) );
  NAND2_X1 U7596 ( .A1(n6152), .A2(n7074), .ZN(n6153) );
  NAND2_X1 U7597 ( .A1(n6154), .A2(n6153), .ZN(n7030) );
  NAND2_X1 U7598 ( .A1(n7737), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6161) );
  INV_X1 U7599 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6155) );
  OR2_X1 U7600 ( .A1(n6085), .A2(n6155), .ZN(n6160) );
  NAND2_X1 U7601 ( .A1(n6156), .A2(n7190), .ZN(n6157) );
  NAND2_X1 U7602 ( .A1(n6179), .A2(n6157), .ZN(n7250) );
  OR2_X1 U7603 ( .A1(n7648), .A2(n7250), .ZN(n6159) );
  INV_X1 U7604 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7169) );
  OR2_X1 U7605 ( .A1(n6274), .A2(n7169), .ZN(n6158) );
  NOR2_X1 U7606 ( .A1(n7295), .A2(n7722), .ZN(n6171) );
  NAND2_X1 U7607 ( .A1(n6185), .A2(n6490), .ZN(n6170) );
  NAND2_X1 U7608 ( .A1(n6326), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6169) );
  INV_X1 U7609 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6162) );
  NAND3_X1 U7610 ( .A1(n6164), .A2(n6163), .A3(n6162), .ZN(n6165) );
  NAND2_X1 U7611 ( .A1(n6186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U7612 ( .A(n6167), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7189) );
  NAND2_X1 U7613 ( .A1(n6404), .A2(n7189), .ZN(n6168) );
  XNOR2_X1 U7614 ( .A(n10041), .B(n7723), .ZN(n7362) );
  NAND2_X1 U7615 ( .A1(n6171), .A2(n7362), .ZN(n6189) );
  INV_X1 U7616 ( .A(n6171), .ZN(n6173) );
  INV_X1 U7617 ( .A(n7362), .ZN(n6172) );
  NAND2_X1 U7618 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  AND2_X1 U7619 ( .A1(n6189), .A2(n6174), .ZN(n7071) );
  NAND2_X1 U7620 ( .A1(n6175), .A2(n7071), .ZN(n7364) );
  NAND2_X1 U7621 ( .A1(n7737), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6184) );
  INV_X1 U7622 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6176) );
  OR2_X1 U7623 ( .A1(n6085), .A2(n6176), .ZN(n6183) );
  INV_X1 U7624 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7625 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NAND2_X1 U7626 ( .A1(n6202), .A2(n6180), .ZN(n7366) );
  OR2_X1 U7627 ( .A1(n7648), .A2(n7366), .ZN(n6182) );
  INV_X1 U7628 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7168) );
  OR2_X1 U7629 ( .A1(n6274), .A2(n7168), .ZN(n6181) );
  OR2_X1 U7630 ( .A1(n7379), .A2(n7722), .ZN(n6193) );
  NAND2_X1 U7631 ( .A1(n6493), .A2(n6185), .ZN(n6188) );
  NOR2_X1 U7632 ( .A1(n6186), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7633 ( .A1(n6235), .A2(n6195), .ZN(n6196) );
  XNOR2_X1 U7634 ( .A(n6196), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8093) );
  AOI22_X1 U7635 ( .A1(n7867), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6404), .B2(
        n8093), .ZN(n6187) );
  NAND2_X1 U7636 ( .A1(n6188), .A2(n6187), .ZN(n10047) );
  XNOR2_X1 U7637 ( .A(n10047), .B(n7723), .ZN(n6192) );
  XNOR2_X1 U7638 ( .A(n6193), .B(n6192), .ZN(n7375) );
  INV_X1 U7639 ( .A(n6189), .ZN(n6190) );
  NOR2_X1 U7640 ( .A1(n7375), .A2(n6190), .ZN(n6191) );
  NAND2_X1 U7641 ( .A1(n7364), .A2(n6191), .ZN(n7371) );
  NAND2_X1 U7642 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  NAND2_X1 U7643 ( .A1(n7371), .A2(n6194), .ZN(n7407) );
  NAND2_X1 U7644 ( .A1(n6496), .A2(n6185), .ZN(n6201) );
  INV_X1 U7645 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6233) );
  AOI21_X1 U7646 ( .B1(n6196), .B2(n6233), .A(n6195), .ZN(n6197) );
  NAND2_X1 U7647 ( .A1(n6197), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6199) );
  INV_X1 U7648 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7649 ( .A1(n6198), .A2(n6232), .ZN(n6214) );
  AND2_X1 U7650 ( .A1(n6199), .A2(n6214), .ZN(n7280) );
  AOI22_X1 U7651 ( .A1(n6326), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6404), .B2(
        n7280), .ZN(n6200) );
  XNOR2_X1 U7652 ( .A(n10055), .B(n7723), .ZN(n6209) );
  NAND2_X1 U7653 ( .A1(n7637), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7654 ( .A1(n6202), .A2(n10470), .ZN(n6203) );
  NAND2_X1 U7655 ( .A1(n6220), .A2(n6203), .ZN(n7410) );
  OR2_X1 U7656 ( .A1(n7648), .A2(n7410), .ZN(n6207) );
  INV_X1 U7657 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7383) );
  OR2_X1 U7658 ( .A1(n6086), .A2(n7383), .ZN(n6206) );
  INV_X1 U7659 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6204) );
  OR2_X1 U7660 ( .A1(n6085), .A2(n6204), .ZN(n6205) );
  NAND4_X1 U7661 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(n8078)
         );
  AND2_X1 U7662 ( .A1(n8078), .A2(n7877), .ZN(n6210) );
  NAND2_X1 U7663 ( .A1(n6209), .A2(n6210), .ZN(n6213) );
  INV_X1 U7664 ( .A(n6209), .ZN(n7464) );
  INV_X1 U7665 ( .A(n6210), .ZN(n6211) );
  NAND2_X1 U7666 ( .A1(n7464), .A2(n6211), .ZN(n6212) );
  NAND2_X1 U7667 ( .A1(n6213), .A2(n6212), .ZN(n7408) );
  NAND2_X1 U7668 ( .A1(n7462), .A2(n6213), .ZN(n6230) );
  NAND2_X1 U7669 ( .A1(n6532), .A2(n6185), .ZN(n6217) );
  NAND2_X1 U7670 ( .A1(n6214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7671 ( .A(n6215), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8106) );
  AOI22_X1 U7672 ( .A1(n6326), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6404), .B2(
        n8106), .ZN(n6216) );
  XNOR2_X1 U7673 ( .A(n7483), .B(n7660), .ZN(n6226) );
  INV_X1 U7674 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7401) );
  OR2_X1 U7675 ( .A1(n6086), .A2(n7401), .ZN(n6224) );
  INV_X1 U7676 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7677 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U7678 ( .A1(n6239), .A2(n6221), .ZN(n7467) );
  OR2_X1 U7679 ( .A1(n7648), .A2(n7467), .ZN(n6223) );
  INV_X1 U7680 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7271) );
  OR2_X1 U7681 ( .A1(n6274), .A2(n7271), .ZN(n6222) );
  NOR2_X1 U7682 ( .A1(n7548), .A2(n7722), .ZN(n6227) );
  NAND2_X1 U7683 ( .A1(n6226), .A2(n6227), .ZN(n6245) );
  INV_X1 U7684 ( .A(n6226), .ZN(n7545) );
  INV_X1 U7685 ( .A(n6227), .ZN(n6228) );
  NAND2_X1 U7686 ( .A1(n7545), .A2(n6228), .ZN(n6229) );
  AND2_X1 U7687 ( .A1(n6245), .A2(n6229), .ZN(n7460) );
  NAND2_X1 U7688 ( .A1(n6637), .A2(n6185), .ZN(n6238) );
  INV_X1 U7689 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6231) );
  AND3_X1 U7690 ( .A1(n6233), .A2(n6232), .A3(n6231), .ZN(n6234) );
  AND2_X1 U7691 ( .A1(n6235), .A2(n6234), .ZN(n6252) );
  OR2_X1 U7692 ( .A1(n6252), .A2(n6195), .ZN(n6236) );
  XNOR2_X1 U7693 ( .A(n6236), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U7694 ( .A1(n6326), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6404), .B2(
        n7333), .ZN(n6237) );
  XNOR2_X1 U7695 ( .A(n10072), .B(n7723), .ZN(n6249) );
  INV_X1 U7696 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7481) );
  OR2_X1 U7697 ( .A1(n6086), .A2(n7481), .ZN(n6243) );
  INV_X1 U7698 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U7699 ( .A1(n6239), .A2(n10485), .ZN(n6240) );
  NAND2_X1 U7700 ( .A1(n6255), .A2(n6240), .ZN(n7552) );
  OR2_X1 U7701 ( .A1(n7648), .A2(n7552), .ZN(n6242) );
  INV_X1 U7702 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7275) );
  OR2_X1 U7703 ( .A1(n6274), .A2(n7275), .ZN(n6241) );
  NOR2_X1 U7704 ( .A1(n8075), .A2(n7722), .ZN(n6247) );
  XNOR2_X1 U7705 ( .A(n6249), .B(n6247), .ZN(n7557) );
  AND2_X1 U7706 ( .A1(n7557), .A2(n6245), .ZN(n6246) );
  INV_X1 U7707 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7708 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U7709 ( .A1(n6680), .A2(n6185), .ZN(n6254) );
  INV_X1 U7710 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7711 ( .A1(n6252), .A2(n6251), .ZN(n6288) );
  NAND2_X1 U7712 ( .A1(n6288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6266) );
  XNOR2_X1 U7713 ( .A(n6266), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7353) );
  AOI22_X1 U7714 ( .A1(n6326), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6404), .B2(
        n7353), .ZN(n6253) );
  XNOR2_X1 U7715 ( .A(n7540), .B(n7660), .ZN(n6262) );
  INV_X1 U7716 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7286) );
  NAND2_X1 U7717 ( .A1(n6255), .A2(n7286), .ZN(n6256) );
  NAND2_X1 U7718 ( .A1(n6272), .A2(n6256), .ZN(n7534) );
  OR2_X1 U7719 ( .A1(n7648), .A2(n7534), .ZN(n6260) );
  INV_X1 U7720 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6257) );
  OR2_X1 U7721 ( .A1(n6274), .A2(n6257), .ZN(n6259) );
  INV_X1 U7722 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7535) );
  OR2_X1 U7723 ( .A1(n6086), .A2(n7535), .ZN(n6258) );
  NOR2_X1 U7724 ( .A1(n8492), .A2(n7722), .ZN(n6263) );
  NAND2_X1 U7725 ( .A1(n6262), .A2(n6263), .ZN(n6279) );
  INV_X1 U7726 ( .A(n6262), .ZN(n7691) );
  INV_X1 U7727 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7728 ( .A1(n7691), .A2(n6264), .ZN(n6265) );
  AND2_X1 U7729 ( .A1(n6279), .A2(n6265), .ZN(n7521) );
  NAND2_X1 U7730 ( .A1(n6700), .A2(n6185), .ZN(n6269) );
  NAND2_X1 U7731 ( .A1(n6266), .A2(n6286), .ZN(n6267) );
  NAND2_X1 U7732 ( .A1(n6267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6310) );
  XNOR2_X1 U7733 ( .A(n6310), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7492) );
  AOI22_X1 U7734 ( .A1(n7867), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6404), .B2(
        n7492), .ZN(n6268) );
  NAND2_X2 U7735 ( .A1(n6269), .A2(n6268), .ZN(n8590) );
  XNOR2_X1 U7736 ( .A(n8590), .B(n7723), .ZN(n6283) );
  INV_X1 U7737 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6270) );
  OR2_X1 U7738 ( .A1(n6086), .A2(n6270), .ZN(n6277) );
  INV_X1 U7739 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U7740 ( .A1(n6272), .A2(n10478), .ZN(n6273) );
  NAND2_X1 U7741 ( .A1(n6301), .A2(n6273), .ZN(n8482) );
  OR2_X1 U7742 ( .A1(n7648), .A2(n8482), .ZN(n6276) );
  INV_X1 U7743 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7495) );
  OR2_X1 U7744 ( .A1(n6274), .A2(n7495), .ZN(n6275) );
  NOR2_X1 U7745 ( .A1(n8073), .A2(n7722), .ZN(n6281) );
  XNOR2_X1 U7746 ( .A(n6283), .B(n6281), .ZN(n7701) );
  AND2_X1 U7747 ( .A1(n7701), .A2(n6279), .ZN(n6280) );
  INV_X1 U7748 ( .A(n6281), .ZN(n6282) );
  NAND2_X1 U7749 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U7750 ( .A1(n7697), .A2(n6284), .ZN(n7766) );
  NAND2_X1 U7751 ( .A1(n6776), .A2(n6185), .ZN(n6291) );
  INV_X1 U7752 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6309) );
  INV_X1 U7753 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6285) );
  NAND3_X1 U7754 ( .A1(n6309), .A2(n6286), .A3(n6285), .ZN(n6287) );
  OAI21_X1 U7755 ( .B1(n6288), .B2(n6287), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6289) );
  XNOR2_X1 U7756 ( .A(n6289), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8135) );
  AOI22_X1 U7757 ( .A1(n6326), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6404), .B2(
        n8135), .ZN(n6290) );
  XNOR2_X1 U7758 ( .A(n8580), .B(n7660), .ZN(n7769) );
  NAND2_X1 U7759 ( .A1(n7737), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6298) );
  INV_X1 U7760 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6292) );
  OR2_X1 U7761 ( .A1(n6085), .A2(n6292), .ZN(n6297) );
  INV_X1 U7762 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U7763 ( .A1(n6303), .A2(n8128), .ZN(n6294) );
  NAND2_X1 U7764 ( .A1(n6372), .A2(n6294), .ZN(n8452) );
  OR2_X1 U7765 ( .A1(n7648), .A2(n8452), .ZN(n6296) );
  INV_X1 U7766 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8142) );
  OR2_X1 U7767 ( .A1(n4481), .A2(n8142), .ZN(n6295) );
  NOR2_X1 U7768 ( .A1(n8435), .A2(n7722), .ZN(n6317) );
  INV_X1 U7769 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6299) );
  OR2_X1 U7770 ( .A1(n6086), .A2(n6299), .ZN(n6307) );
  INV_X1 U7771 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7772 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7773 ( .A1(n6303), .A2(n6302), .ZN(n8463) );
  OR2_X1 U7774 ( .A1(n7648), .A2(n8463), .ZN(n6306) );
  INV_X1 U7775 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6304) );
  OR2_X1 U7776 ( .A1(n6274), .A2(n6304), .ZN(n6305) );
  NOR2_X1 U7777 ( .A1(n8490), .A2(n7722), .ZN(n6316) );
  NAND2_X1 U7778 ( .A1(n6751), .A2(n6185), .ZN(n6314) );
  NAND2_X1 U7779 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  NAND2_X1 U7780 ( .A1(n6311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6312) );
  XNOR2_X1 U7781 ( .A(n6312), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8122) );
  AOI22_X1 U7782 ( .A1(n6326), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6404), .B2(
        n8122), .ZN(n6313) );
  XNOR2_X1 U7783 ( .A(n8585), .B(n7660), .ZN(n7765) );
  AOI22_X1 U7784 ( .A1(n7769), .A2(n6317), .B1(n6316), .B2(n7765), .ZN(n6315)
         );
  NAND2_X1 U7785 ( .A1(n7766), .A2(n6315), .ZN(n6321) );
  INV_X1 U7786 ( .A(n7769), .ZN(n6319) );
  OAI21_X1 U7787 ( .B1(n7765), .B2(n6316), .A(n6317), .ZN(n6318) );
  INV_X1 U7788 ( .A(n7765), .ZN(n7767) );
  INV_X1 U7789 ( .A(n6316), .ZN(n7824) );
  INV_X1 U7790 ( .A(n6317), .ZN(n7768) );
  AOI21_X1 U7791 ( .B1(n6319), .B2(n6318), .A(n4530), .ZN(n6320) );
  NAND2_X1 U7792 ( .A1(n6321), .A2(n6320), .ZN(n6358) );
  NAND2_X1 U7793 ( .A1(n6831), .A2(n6185), .ZN(n6328) );
  NAND2_X1 U7794 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U7795 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6323), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6325) );
  AND2_X1 U7796 ( .A1(n6325), .A2(n6324), .ZN(n8156) );
  AOI22_X1 U7797 ( .A1(n6326), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6404), .B2(
        n8156), .ZN(n6327) );
  XNOR2_X1 U7798 ( .A(n8577), .B(n7660), .ZN(n6333) );
  INV_X1 U7799 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8424) );
  OR2_X1 U7800 ( .A1(n6086), .A2(n8424), .ZN(n6331) );
  INV_X1 U7801 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8139) );
  XNOR2_X1 U7802 ( .A(n6372), .B(n8139), .ZN(n8423) );
  OR2_X1 U7803 ( .A1(n7648), .A2(n8423), .ZN(n6330) );
  INV_X1 U7804 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8152) );
  OR2_X1 U7805 ( .A1(n6274), .A2(n8152), .ZN(n6329) );
  NOR2_X1 U7806 ( .A1(n8445), .A2(n7722), .ZN(n6334) );
  NAND2_X1 U7807 ( .A1(n6333), .A2(n6334), .ZN(n6395) );
  INV_X1 U7808 ( .A(n6333), .ZN(n7799) );
  INV_X1 U7809 ( .A(n6334), .ZN(n6335) );
  NAND2_X1 U7810 ( .A1(n7799), .A2(n6335), .ZN(n6336) );
  NAND2_X1 U7811 ( .A1(n6395), .A2(n6336), .ZN(n6357) );
  AND2_X1 U7812 ( .A1(n6339), .A2(n6337), .ZN(n9998) );
  INV_X1 U7813 ( .A(n9998), .ZN(n6343) );
  INV_X1 U7814 ( .A(n6337), .ZN(n7559) );
  INV_X1 U7815 ( .A(P2_B_REG_SCAN_IN), .ZN(n6338) );
  XNOR2_X1 U7816 ( .A(n6339), .B(n6338), .ZN(n6340) );
  INV_X1 U7817 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U7818 ( .A1(n9995), .A2(n9999), .ZN(n6342) );
  INV_X1 U7819 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10001) );
  NOR2_X1 U7820 ( .A1(n7526), .A2(n7559), .ZN(n10002) );
  AOI21_X1 U7821 ( .B1(n9995), .B2(n10001), .A(n10002), .ZN(n6755) );
  NOR4_X1 U7822 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6347) );
  NOR4_X1 U7823 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6346) );
  NOR4_X1 U7824 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6345) );
  NOR4_X1 U7825 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6344) );
  NAND4_X1 U7826 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6353)
         );
  NOR2_X1 U7827 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6351) );
  NOR4_X1 U7828 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6350) );
  NOR4_X1 U7829 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6349) );
  NOR4_X1 U7830 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6348) );
  NAND4_X1 U7831 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n6352)
         );
  OAI21_X1 U7832 ( .B1(n6353), .B2(n6352), .A(n9995), .ZN(n6754) );
  AND2_X1 U7833 ( .A1(n6755), .A2(n6754), .ZN(n6878) );
  INV_X1 U7834 ( .A(n6359), .ZN(n6363) );
  INV_X1 U7835 ( .A(n10003), .ZN(n6354) );
  NOR2_X1 U7836 ( .A1(n6363), .A2(n6460), .ZN(n6367) );
  OR2_X1 U7837 ( .A1(n10008), .A2(n8066), .ZN(n10063) );
  NAND2_X1 U7838 ( .A1(n8069), .A2(n7890), .ZN(n6461) );
  AND2_X1 U7839 ( .A1(n10063), .A2(n6461), .ZN(n6355) );
  OR2_X2 U7840 ( .A1(n6358), .A2(n6357), .ZN(n7798) );
  INV_X1 U7841 ( .A(n7798), .ZN(n6356) );
  INV_X1 U7843 ( .A(n8577), .ZN(n8422) );
  NOR2_X1 U7844 ( .A1(n10008), .A2(n8024), .ZN(n9974) );
  NAND3_X1 U7845 ( .A1(n6359), .A2(n9996), .A3(n9974), .ZN(n6362) );
  AND2_X1 U7846 ( .A1(n8024), .A2(n9980), .ZN(n6360) );
  NAND2_X1 U7847 ( .A1(n7880), .A2(n6360), .ZN(n10056) );
  OR2_X1 U7848 ( .A1(n10056), .A2(n7890), .ZN(n6753) );
  INV_X1 U7849 ( .A(n6753), .ZN(n6361) );
  NAND2_X1 U7850 ( .A1(n6362), .A2(n8451), .ZN(n7793) );
  INV_X1 U7851 ( .A(n7793), .ZN(n7835) );
  NOR2_X1 U7852 ( .A1(n8422), .A2(n7835), .ZN(n6381) );
  NAND2_X1 U7853 ( .A1(n6363), .A2(n6753), .ZN(n6366) );
  OR2_X1 U7854 ( .A1(n6461), .A2(n8066), .ZN(n6879) );
  NAND2_X1 U7855 ( .A1(n6879), .A2(n6446), .ZN(n6364) );
  NOR2_X1 U7856 ( .A1(n6447), .A2(n6364), .ZN(n6365) );
  NAND2_X1 U7857 ( .A1(n6366), .A2(n6365), .ZN(n6685) );
  OAI22_X1 U7858 ( .A1(n7828), .A2(n8423), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8139), .ZN(n6380) );
  NAND2_X1 U7859 ( .A1(n6367), .A2(n8066), .ZN(n6697) );
  INV_X1 U7860 ( .A(n6697), .ZN(n7819) );
  NOR2_X1 U7861 ( .A1(n6454), .A2(n6461), .ZN(n8469) );
  AND2_X1 U7862 ( .A1(n7819), .A2(n8469), .ZN(n7745) );
  AND2_X1 U7863 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6369) );
  INV_X1 U7864 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6371) );
  OAI21_X1 U7865 ( .B1(n6372), .B2(n8139), .A(n6371), .ZN(n6373) );
  NAND2_X1 U7866 ( .A1(n6407), .A2(n6373), .ZN(n7803) );
  OR2_X1 U7867 ( .A1(n7648), .A2(n7803), .ZN(n6377) );
  INV_X1 U7868 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8170) );
  OR2_X1 U7869 ( .A1(n6274), .A2(n8170), .ZN(n6376) );
  INV_X1 U7870 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6374) );
  OR2_X1 U7871 ( .A1(n6086), .A2(n6374), .ZN(n6375) );
  NAND4_X1 U7872 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n8200)
         );
  INV_X1 U7873 ( .A(n6461), .ZN(n6449) );
  OAI22_X1 U7874 ( .A1(n7830), .A2(n8435), .B1(n8433), .B2(n7829), .ZN(n6379)
         );
  OR4_X1 U7875 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(P2_U3230)
         );
  NAND2_X1 U7876 ( .A1(n7066), .A2(n6185), .ZN(n6384) );
  NAND2_X1 U7877 ( .A1(n7867), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6383) );
  XNOR2_X1 U7878 ( .A(n8560), .B(n7660), .ZN(n6391) );
  NAND2_X1 U7879 ( .A1(n7737), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6390) );
  INV_X1 U7880 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6385) );
  OR2_X1 U7881 ( .A1(n6085), .A2(n6385), .ZN(n6389) );
  INV_X1 U7882 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10426) );
  INV_X1 U7883 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6424) );
  XNOR2_X1 U7884 ( .A(n6425), .B(n6424), .ZN(n8371) );
  OR2_X1 U7885 ( .A1(n8371), .A2(n7648), .ZN(n6388) );
  INV_X1 U7886 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6386) );
  OR2_X1 U7887 ( .A1(n6274), .A2(n6386), .ZN(n6387) );
  NOR2_X1 U7888 ( .A1(n8392), .A2(n7722), .ZN(n6392) );
  NAND2_X1 U7889 ( .A1(n6391), .A2(n6392), .ZN(n7606) );
  INV_X1 U7890 ( .A(n6391), .ZN(n7751) );
  INV_X1 U7891 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U7892 ( .A1(n7751), .A2(n6393), .ZN(n6394) );
  NAND2_X1 U7893 ( .A1(n7606), .A2(n6394), .ZN(n6422) );
  NAND2_X1 U7894 ( .A1(n7798), .A2(n6395), .ZN(n6403) );
  NAND2_X1 U7895 ( .A1(n6958), .A2(n6185), .ZN(n6398) );
  NAND2_X1 U7896 ( .A1(n6324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6396) );
  XNOR2_X1 U7897 ( .A(n6396), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8157) );
  AOI22_X1 U7898 ( .A1(n7867), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6404), .B2(
        n8157), .ZN(n6397) );
  XNOR2_X1 U7899 ( .A(n8570), .B(n7660), .ZN(n6399) );
  AND2_X1 U7900 ( .A1(n8200), .A2(n7877), .ZN(n6400) );
  NAND2_X1 U7901 ( .A1(n6399), .A2(n6400), .ZN(n6414) );
  INV_X1 U7902 ( .A(n6399), .ZN(n7713) );
  INV_X1 U7903 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U7904 ( .A1(n7713), .A2(n6401), .ZN(n6402) );
  AND2_X1 U7905 ( .A1(n6414), .A2(n6402), .ZN(n7796) );
  NAND2_X1 U7906 ( .A1(n7002), .A2(n6185), .ZN(n6406) );
  AOI22_X1 U7907 ( .A1(n7867), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6404), .B2(
        n9980), .ZN(n6405) );
  XNOR2_X1 U7908 ( .A(n8567), .B(n7660), .ZN(n6416) );
  NAND2_X1 U7909 ( .A1(n7637), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7910 ( .A1(n6407), .A2(n10426), .ZN(n6408) );
  NAND2_X1 U7911 ( .A1(n6425), .A2(n6408), .ZN(n8396) );
  OR2_X1 U7912 ( .A1(n7648), .A2(n8396), .ZN(n6412) );
  INV_X1 U7913 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7914 ( .A1(n6086), .A2(n8397), .ZN(n6411) );
  INV_X1 U7915 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6409) );
  OR2_X1 U7916 ( .A1(n6085), .A2(n6409), .ZN(n6410) );
  NAND4_X1 U7917 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .ZN(n8378)
         );
  NAND2_X1 U7918 ( .A1(n8378), .A2(n7877), .ZN(n6417) );
  XNOR2_X1 U7919 ( .A(n6416), .B(n6417), .ZN(n7714) );
  AND2_X1 U7920 ( .A1(n7714), .A2(n6414), .ZN(n6415) );
  INV_X1 U7921 ( .A(n6416), .ZN(n6418) );
  NAND2_X1 U7922 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  INV_X1 U7923 ( .A(n7750), .ZN(n6420) );
  AOI211_X1 U7924 ( .C1(n6422), .C2(n6421), .A(n7810), .B(n6420), .ZN(n6437)
         );
  INV_X1 U7925 ( .A(n8560), .ZN(n8374) );
  NOR2_X1 U7926 ( .A1(n8374), .A2(n7835), .ZN(n6436) );
  OAI22_X1 U7927 ( .A1(n7828), .A2(n8371), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6424), .ZN(n6435) );
  NAND2_X1 U7928 ( .A1(n7737), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6433) );
  INV_X1 U7929 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6423) );
  OR2_X1 U7930 ( .A1(n6085), .A2(n6423), .ZN(n6432) );
  INV_X1 U7931 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10455) );
  OAI21_X1 U7932 ( .B1(n6425), .B2(n6424), .A(n10455), .ZN(n6428) );
  AND2_X1 U7933 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n6426) );
  NAND2_X1 U7934 ( .A1(n6428), .A2(n6656), .ZN(n8362) );
  OR2_X1 U7935 ( .A1(n7648), .A2(n8362), .ZN(n6431) );
  INV_X1 U7936 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6429) );
  OR2_X1 U7937 ( .A1(n4481), .A2(n6429), .ZN(n6430) );
  OAI22_X1 U7938 ( .A1(n7830), .A2(n8412), .B1(n8345), .B2(n7829), .ZN(n6434)
         );
  OR4_X1 U7939 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(P2_U3235)
         );
  INV_X1 U7940 ( .A(n6438), .ZN(n6976) );
  AOI211_X1 U7941 ( .C1(n6440), .C2(n6439), .A(n7810), .B(n6976), .ZN(n6444)
         );
  NOR2_X1 U7942 ( .A1(n7828), .A2(n9973), .ZN(n6443) );
  OAI22_X1 U7943 ( .A1(n7835), .A2(n7041), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6100), .ZN(n6442) );
  OAI22_X1 U7944 ( .A1(n7830), .A2(n7050), .B1(n7049), .B2(n7829), .ZN(n6441)
         );
  OR4_X1 U7945 ( .A1(n6444), .A2(n6443), .A3(n6442), .A4(n6441), .ZN(P2_U3229)
         );
  NAND2_X1 U7946 ( .A1(n9960), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6453) );
  INV_X1 U7947 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6445) );
  INV_X1 U7948 ( .A(n9960), .ZN(n9968) );
  NOR2_X1 U7949 ( .A1(n6454), .A2(P2_U3152), .ZN(n8622) );
  NOR2_X1 U7950 ( .A1(n6446), .A2(P2_U3152), .ZN(n8065) );
  AOI21_X1 U7951 ( .B1(n8622), .B2(n6447), .A(n8065), .ZN(n6448) );
  OAI21_X1 U7952 ( .B1(n6460), .B2(n6449), .A(n6448), .ZN(n6457) );
  NAND2_X1 U7953 ( .A1(n6457), .A2(n6059), .ZN(n6450) );
  INV_X2 U7954 ( .A(P2_U3966), .ZN(n8087) );
  NAND2_X1 U7955 ( .A1(n6450), .A2(n8087), .ZN(n6455) );
  INV_X1 U7956 ( .A(n6455), .ZN(n6451) );
  NOR3_X2 U7957 ( .A1(n6451), .A2(n6454), .A3(n7567), .ZN(n9965) );
  AOI211_X1 U7958 ( .C1(n6453), .C2(n6452), .A(n7119), .B(n9602), .ZN(n6467)
         );
  NAND2_X1 U7959 ( .A1(n6455), .A2(n6454), .ZN(n9961) );
  INV_X1 U7960 ( .A(n7120), .ZN(n7132) );
  NOR2_X1 U7961 ( .A1(n9961), .A2(n7132), .ZN(n6466) );
  INV_X1 U7962 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10084) );
  OR2_X1 U7963 ( .A1(n9968), .A2(n10084), .ZN(n6459) );
  INV_X1 U7964 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7133) );
  MUX2_X1 U7965 ( .A(n7133), .B(P2_REG1_REG_1__SCAN_IN), .S(n7120), .Z(n6458)
         );
  NOR3_X1 U7966 ( .A1(n6458), .A2(n10084), .A3(n9968), .ZN(n7130) );
  AND2_X1 U7967 ( .A1(n6059), .A2(n7567), .ZN(n6456) );
  NAND2_X1 U7968 ( .A1(n6457), .A2(n6456), .ZN(n9962) );
  AOI211_X1 U7969 ( .C1(n6459), .C2(n6458), .A(n7130), .B(n9962), .ZN(n6465)
         );
  INV_X1 U7970 ( .A(n8065), .ZN(n8068) );
  OAI21_X1 U7971 ( .B1(n6059), .B2(n8068), .A(n6460), .ZN(n6463) );
  NAND2_X1 U7972 ( .A1(n6059), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U7973 ( .A1(n6463), .A2(n6462), .ZN(n8181) );
  INV_X1 U7974 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10101) );
  OAI22_X1 U7975 ( .A1(n8181), .A2(n10101), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6915), .ZN(n6464) );
  OR4_X1 U7976 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(P2_U3246)
         );
  NOR2_X1 U7977 ( .A1(n5320), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8623) );
  AOI22_X1 U7978 ( .A1(n8623), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n7120), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6469) );
  OAI21_X1 U7979 ( .B1(n6482), .B2(n6488), .A(n6469), .ZN(P2_U3357) );
  AOI22_X1 U7980 ( .A1(n8623), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9607), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6470) );
  OAI21_X1 U7981 ( .B1(n6472), .B2(n6488), .A(n6470), .ZN(P2_U3356) );
  AOI22_X1 U7982 ( .A1(n8623), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7149), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6471) );
  OAI21_X1 U7983 ( .B1(n6478), .B2(n6488), .A(n6471), .ZN(P2_U3355) );
  NOR2_X1 U7984 ( .A1(n6040), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9597) );
  INV_X1 U7985 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7986 ( .A1(n6040), .A2(P1_U3084), .ZN(n9599) );
  INV_X1 U7987 ( .A(n6518), .ZN(n9687) );
  OAI222_X1 U7988 ( .A1(n9595), .A2(n6473), .B1(n9599), .B2(n6472), .C1(
        P1_U3084), .C2(n9687), .ZN(P1_U3351) );
  AOI22_X1 U7989 ( .A1(n8623), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7226), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6474) );
  OAI21_X1 U7990 ( .B1(n6480), .B2(n6488), .A(n6474), .ZN(P2_U3354) );
  AOI22_X1 U7991 ( .A1(n7173), .A2(P2_STATE_REG_SCAN_IN), .B1(n8623), .B2(
        P1_DATAO_REG_5__SCAN_IN), .ZN(n6475) );
  OAI21_X1 U7992 ( .B1(n6476), .B2(n6488), .A(n6475), .ZN(P2_U3353) );
  INV_X1 U7993 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6477) );
  OAI222_X1 U7994 ( .A1(n9595), .A2(n6477), .B1(n9599), .B2(n6476), .C1(
        P1_U3084), .C2(n6593), .ZN(P1_U3348) );
  INV_X1 U7995 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6479) );
  CLKBUF_X1 U7996 ( .A(n9599), .Z(n7594) );
  INV_X1 U7997 ( .A(n6546), .ZN(n6513) );
  OAI222_X1 U7998 ( .A1(n9595), .A2(n6479), .B1(n7594), .B2(n6478), .C1(
        P1_U3084), .C2(n6513), .ZN(P1_U3350) );
  INV_X1 U7999 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6481) );
  INV_X1 U8000 ( .A(n9703), .ZN(n6550) );
  OAI222_X1 U8001 ( .A1(n9595), .A2(n6481), .B1(n7594), .B2(n6480), .C1(
        P1_U3084), .C2(n6550), .ZN(P1_U3349) );
  INV_X1 U8002 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6483) );
  INV_X1 U8003 ( .A(n6630), .ZN(n6628) );
  OAI222_X1 U8004 ( .A1(n9595), .A2(n6483), .B1(n7594), .B2(n6482), .C1(
        P1_U3084), .C2(n6628), .ZN(P1_U3352) );
  INV_X1 U8005 ( .A(n6484), .ZN(n6486) );
  CLKBUF_X1 U8006 ( .A(n8623), .Z(n8618) );
  AOI22_X1 U8007 ( .A1(n7171), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8618), .ZN(n6485) );
  OAI21_X1 U8008 ( .B1(n6486), .B2(n6488), .A(n6485), .ZN(P2_U3352) );
  OAI222_X1 U8009 ( .A1(n9595), .A2(n10323), .B1(n7594), .B2(n6486), .C1(
        P1_U3084), .C2(n6576), .ZN(P1_U3347) );
  AOI22_X1 U8010 ( .A1(n7213), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8618), .ZN(n6487) );
  OAI21_X1 U8011 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(P2_U3351) );
  INV_X1 U8012 ( .A(n8181), .ZN(n9966) );
  NOR2_X1 U8013 ( .A1(n9966), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8014 ( .A(n6490), .ZN(n6492) );
  AOI22_X1 U8015 ( .A1(n7189), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8618), .ZN(n6491) );
  OAI21_X1 U8016 ( .B1(n6492), .B2(n6488), .A(n6491), .ZN(P2_U3350) );
  OAI222_X1 U8017 ( .A1(n9595), .A2(n10476), .B1(n7594), .B2(n6492), .C1(
        P1_U3084), .C2(n9727), .ZN(P1_U3345) );
  INV_X1 U8018 ( .A(n6493), .ZN(n6495) );
  AOI22_X1 U8019 ( .A1(n8093), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8618), .ZN(n6494) );
  OAI21_X1 U8020 ( .B1(n6495), .B2(n6488), .A(n6494), .ZN(P2_U3349) );
  INV_X1 U8021 ( .A(n6647), .ZN(n6613) );
  OAI222_X1 U8022 ( .A1(n7594), .A2(n6495), .B1(n6613), .B2(P1_U3084), .C1(
        n10239), .C2(n9595), .ZN(P1_U3344) );
  INV_X1 U8023 ( .A(n6496), .ZN(n6562) );
  AOI22_X1 U8024 ( .A1(n7280), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8618), .ZN(n6497) );
  OAI21_X1 U8025 ( .B1(n6562), .B2(n6488), .A(n6497), .ZN(P2_U3348) );
  INV_X1 U8026 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6527) );
  INV_X1 U8027 ( .A(n6498), .ZN(n6499) );
  NOR2_X1 U8028 ( .A1(n9688), .A2(P1_U3084), .ZN(n7569) );
  AND2_X1 U8029 ( .A1(n6508), .A2(n7569), .ZN(n9723) );
  NAND2_X1 U8030 ( .A1(n9723), .A2(n5923), .ZN(n9817) );
  NOR2_X1 U8031 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5234), .ZN(n6796) );
  INV_X1 U8032 ( .A(n6796), .ZN(n6512) );
  INV_X1 U8033 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U8034 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6500), .S(n6546), .Z(n6510)
         );
  INV_X1 U8035 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9943) );
  XNOR2_X1 U8036 ( .A(n6518), .B(n9943), .ZN(n9697) );
  INV_X1 U8037 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6501) );
  MUX2_X1 U8038 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6501), .S(n6630), .Z(n6503)
         );
  AND2_X1 U8039 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6502) );
  NAND2_X1 U8040 ( .A1(n6503), .A2(n6502), .ZN(n6625) );
  NAND2_X1 U8041 ( .A1(n6630), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8042 ( .A1(n6625), .A2(n6504), .ZN(n9698) );
  NAND2_X1 U8043 ( .A1(n9697), .A2(n9698), .ZN(n6506) );
  NAND2_X1 U8044 ( .A1(n6518), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U8045 ( .A1(n6506), .A2(n6505), .ZN(n6509) );
  NOR2_X1 U8046 ( .A1(n5923), .A2(P1_U3084), .ZN(n9596) );
  AND2_X1 U8047 ( .A1(n9596), .A2(n9688), .ZN(n6507) );
  NAND2_X1 U8048 ( .A1(n6508), .A2(n6507), .ZN(n9823) );
  NAND2_X1 U8049 ( .A1(n6509), .A2(n6510), .ZN(n6535) );
  OAI211_X1 U8050 ( .C1(n6510), .C2(n6509), .A(n9806), .B(n6535), .ZN(n6511)
         );
  OAI211_X1 U8051 ( .C1(n9817), .C2(n6513), .A(n6512), .B(n6511), .ZN(n6514)
         );
  INV_X1 U8052 ( .A(n6514), .ZN(n6526) );
  INV_X1 U8053 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6515) );
  MUX2_X1 U8054 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6515), .S(n6518), .Z(n9685)
         );
  INV_X1 U8055 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6826) );
  MUX2_X1 U8056 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6826), .S(n6630), .Z(n6516)
         );
  AND2_X1 U8057 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6629) );
  NAND2_X1 U8058 ( .A1(n6516), .A2(n6629), .ZN(n6631) );
  NAND2_X1 U8059 ( .A1(n6630), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8060 ( .A1(n6631), .A2(n6517), .ZN(n9684) );
  NAND2_X1 U8061 ( .A1(n9685), .A2(n9684), .ZN(n9683) );
  NAND2_X1 U8062 ( .A1(n6518), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8063 ( .A1(n9683), .A2(n6523), .ZN(n6520) );
  INV_X1 U8064 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6521) );
  MUX2_X1 U8065 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6521), .S(n6546), .Z(n6519)
         );
  NAND2_X1 U8066 ( .A1(n6520), .A2(n6519), .ZN(n6548) );
  MUX2_X1 U8067 ( .A(n6521), .B(P1_REG2_REG_3__SCAN_IN), .S(n6546), .Z(n6522)
         );
  NAND3_X1 U8068 ( .A1(n9683), .A2(n6523), .A3(n6522), .ZN(n6524) );
  NAND3_X1 U8069 ( .A1(n9811), .A2(n6548), .A3(n6524), .ZN(n6525) );
  OAI211_X1 U8070 ( .C1(n6527), .C2(n9828), .A(n6526), .B(n6525), .ZN(P1_U3244) );
  INV_X1 U8071 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10458) );
  INV_X1 U8072 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8073 ( .A1(n7637), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6529) );
  INV_X1 U8074 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8184) );
  OR2_X1 U8075 ( .A1(n6086), .A2(n8184), .ZN(n6528) );
  OAI211_X1 U8076 ( .C1(n6085), .C2(n6530), .A(n6529), .B(n6528), .ZN(n8186)
         );
  NAND2_X1 U8077 ( .A1(n8186), .A2(P2_U3966), .ZN(n6531) );
  OAI21_X1 U8078 ( .B1(n10458), .B2(P2_U3966), .A(n6531), .ZN(P2_U3583) );
  INV_X1 U8079 ( .A(n6532), .ZN(n6586) );
  AOI22_X1 U8080 ( .A1(n8106), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8618), .ZN(n6533) );
  OAI21_X1 U8081 ( .B1(n6586), .B2(n6488), .A(n6533), .ZN(P2_U3347) );
  INV_X1 U8082 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6561) );
  INV_X1 U8083 ( .A(n9817), .ZN(n9790) );
  INV_X1 U8084 ( .A(n6610), .ZN(n6545) );
  AND2_X1 U8085 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7086) );
  NAND2_X1 U8086 ( .A1(n6546), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6534) );
  AND2_X1 U8087 ( .A1(n6535), .A2(n6534), .ZN(n9713) );
  INV_X1 U8088 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U8089 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9946), .S(n9703), .Z(n9714)
         );
  NAND2_X1 U8090 ( .A1(n9713), .A2(n9714), .ZN(n9712) );
  NAND2_X1 U8091 ( .A1(n6550), .A2(n9946), .ZN(n6536) );
  NAND2_X1 U8092 ( .A1(n9712), .A2(n6536), .ZN(n6589) );
  INV_X1 U8093 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U8094 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9949), .S(n6593), .Z(n6588)
         );
  OR2_X1 U8095 ( .A1(n6589), .A2(n6588), .ZN(n6591) );
  NAND2_X1 U8096 ( .A1(n6537), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6538) );
  AND2_X1 U8097 ( .A1(n6591), .A2(n6538), .ZN(n6574) );
  INV_X1 U8098 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9951) );
  MUX2_X1 U8099 ( .A(n9951), .B(P1_REG1_REG_6__SCAN_IN), .S(n6576), .Z(n6573)
         );
  NAND2_X1 U8100 ( .A1(n6574), .A2(n6573), .ZN(n6572) );
  NAND2_X1 U8101 ( .A1(n6576), .A2(n9951), .ZN(n6541) );
  NAND2_X1 U8102 ( .A1(n6572), .A2(n6541), .ZN(n6539) );
  INV_X1 U8103 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U8104 ( .A(n9953), .B(P1_REG1_REG_7__SCAN_IN), .S(n6610), .Z(n6540)
         );
  NAND2_X1 U8105 ( .A1(n6539), .A2(n6540), .ZN(n6612) );
  INV_X1 U8106 ( .A(n6540), .ZN(n6542) );
  NAND3_X1 U8107 ( .A1(n6572), .A2(n6542), .A3(n6541), .ZN(n6543) );
  AOI21_X1 U8108 ( .B1(n6612), .B2(n6543), .A(n9823), .ZN(n6544) );
  AOI211_X1 U8109 ( .C1(n9790), .C2(n6545), .A(n7086), .B(n6544), .ZN(n6560)
         );
  NAND2_X1 U8110 ( .A1(n6546), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6547) );
  AND2_X1 U8111 ( .A1(n6548), .A2(n6547), .ZN(n9706) );
  INV_X1 U8112 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U8113 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6549), .S(n9703), .Z(n9705)
         );
  NAND2_X1 U8114 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  NAND2_X1 U8115 ( .A1(n6550), .A2(n6549), .ZN(n6595) );
  NAND2_X1 U8116 ( .A1(n9704), .A2(n6595), .ZN(n6551) );
  INV_X1 U8117 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U8118 ( .A(n9876), .B(P1_REG2_REG_5__SCAN_IN), .S(n6593), .Z(n6594)
         );
  NAND2_X1 U8119 ( .A1(n6551), .A2(n6594), .ZN(n6598) );
  NAND2_X1 U8120 ( .A1(n6593), .A2(n9876), .ZN(n6552) );
  NAND2_X1 U8121 ( .A1(n6598), .A2(n6552), .ZN(n6580) );
  INV_X1 U8122 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8123 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6553), .S(n6576), .Z(n6579)
         );
  NAND2_X1 U8124 ( .A1(n6554), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6555) );
  INV_X1 U8125 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7113) );
  MUX2_X1 U8126 ( .A(n7113), .B(P1_REG2_REG_7__SCAN_IN), .S(n6610), .Z(n6556)
         );
  NAND2_X1 U8127 ( .A1(n6557), .A2(n6556), .ZN(n6604) );
  OAI21_X1 U8128 ( .B1(n6557), .B2(n6556), .A(n6604), .ZN(n6558) );
  NAND2_X1 U8129 ( .A1(n9811), .A2(n6558), .ZN(n6559) );
  OAI211_X1 U8130 ( .C1(n6561), .C2(n9828), .A(n6560), .B(n6559), .ZN(P1_U3248) );
  INV_X1 U8131 ( .A(n6735), .ZN(n6731) );
  OAI222_X1 U8132 ( .A1(n9595), .A2(n6563), .B1(n6731), .B2(P1_U3084), .C1(
        n7594), .C2(n6562), .ZN(P1_U3343) );
  INV_X1 U8133 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6571) );
  INV_X1 U8134 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6730) );
  OAI22_X1 U8135 ( .A1(n9688), .A2(n6629), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6730), .ZN(n6565) );
  NOR2_X1 U8136 ( .A1(n9688), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6564) );
  OAI21_X1 U8137 ( .B1(n5923), .B2(n6564), .A(n6623), .ZN(n9691) );
  OAI211_X1 U8138 ( .C1(n5923), .C2(n6565), .A(n9691), .B(P1_STATE_REG_SCAN_IN), .ZN(n6566) );
  NOR2_X1 U8139 ( .A1(n6567), .A2(n6566), .ZN(n6569) );
  AND3_X1 U8140 ( .A1(n9806), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6730), .ZN(n6568) );
  AOI211_X1 U8141 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6569), .B(
        n6568), .ZN(n6570) );
  OAI21_X1 U8142 ( .B1(n9828), .B2(n6571), .A(n6570), .ZN(P1_U3241) );
  INV_X1 U8143 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6585) );
  OAI21_X1 U8144 ( .B1(n6574), .B2(n6573), .A(n6572), .ZN(n6578) );
  NOR2_X1 U8145 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6575), .ZN(n7060) );
  NOR2_X1 U8146 ( .A1(n9817), .A2(n6576), .ZN(n6577) );
  AOI211_X1 U8147 ( .C1(n9806), .C2(n6578), .A(n7060), .B(n6577), .ZN(n6584)
         );
  NAND2_X1 U8148 ( .A1(n6580), .A2(n6579), .ZN(n6581) );
  NAND3_X1 U8149 ( .A1(n9811), .A2(n6582), .A3(n6581), .ZN(n6583) );
  OAI211_X1 U8150 ( .C1(n6585), .C2(n9828), .A(n6584), .B(n6583), .ZN(P1_U3247) );
  INV_X1 U8151 ( .A(n6738), .ZN(n9082) );
  OAI222_X1 U8152 ( .A1(n9595), .A2(n6587), .B1(n9082), .B2(P1_U3084), .C1(
        n9599), .C2(n6586), .ZN(P1_U3342) );
  INV_X1 U8153 ( .A(n9828), .ZN(n9696) );
  NAND2_X1 U8154 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U8155 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  NAND3_X1 U8156 ( .A1(n9806), .A2(n6591), .A3(n6590), .ZN(n6592) );
  OAI211_X1 U8157 ( .C1(n9817), .C2(n6593), .A(n7008), .B(n6592), .ZN(n6600)
         );
  INV_X1 U8158 ( .A(n6594), .ZN(n6596) );
  NAND3_X1 U8159 ( .A1(n9704), .A2(n6596), .A3(n6595), .ZN(n6597) );
  INV_X1 U8160 ( .A(n9811), .ZN(n9784) );
  AOI21_X1 U8161 ( .B1(n6598), .B2(n6597), .A(n9784), .ZN(n6599) );
  AOI211_X1 U8162 ( .C1(P1_ADDR_REG_5__SCAN_IN), .C2(n9696), .A(n6600), .B(
        n6599), .ZN(n6601) );
  INV_X1 U8163 ( .A(n6601), .ZN(P1_U3246) );
  NAND2_X1 U8164 ( .A1(n6647), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6602) );
  OAI21_X1 U8165 ( .B1(n6647), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6602), .ZN(
        n6609) );
  NAND2_X1 U8166 ( .A1(n6610), .A2(n7113), .ZN(n6603) );
  AND2_X1 U8167 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  NAND2_X1 U8168 ( .A1(n6605), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U8169 ( .A1(n9720), .A2(n9727), .ZN(n6608) );
  INV_X1 U8170 ( .A(n6605), .ZN(n9728) );
  INV_X1 U8171 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8172 ( .A1(n9728), .A2(n6606), .ZN(n6607) );
  NAND2_X1 U8173 ( .A1(n6608), .A2(n6607), .ZN(n9730) );
  NOR2_X1 U8174 ( .A1(n9730), .A2(n6609), .ZN(n6646) );
  AOI211_X1 U8175 ( .C1(n6609), .C2(n9730), .A(n6646), .B(n9784), .ZN(n6621)
         );
  NAND2_X1 U8176 ( .A1(n6610), .A2(n9953), .ZN(n6611) );
  NAND2_X1 U8177 ( .A1(n6612), .A2(n6611), .ZN(n9732) );
  INV_X1 U8178 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9955) );
  MUX2_X1 U8179 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9955), .S(n9727), .Z(n9731)
         );
  OR2_X1 U8180 ( .A1(n9732), .A2(n9731), .ZN(n9734) );
  OAI21_X1 U8181 ( .B1(n9727), .B2(n9955), .A(n9734), .ZN(n6615) );
  INV_X1 U8182 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U8183 ( .A1(n6647), .A2(n9958), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6613), .ZN(n6614) );
  NOR2_X1 U8184 ( .A1(n6615), .A2(n6614), .ZN(n6639) );
  AOI21_X1 U8185 ( .B1(n6615), .B2(n6614), .A(n6639), .ZN(n6616) );
  NOR2_X1 U8186 ( .A1(n6616), .A2(n9823), .ZN(n6620) );
  INV_X1 U8187 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8188 ( .A1(n9790), .A2(n6647), .ZN(n6617) );
  NAND2_X1 U8189 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7420) );
  OAI211_X1 U8190 ( .C1(n6618), .C2(n9828), .A(n6617), .B(n7420), .ZN(n6619)
         );
  OR3_X1 U8191 ( .A1(n6621), .A2(n6620), .A3(n6619), .ZN(P1_U3250) );
  NAND2_X1 U8192 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6627) );
  MUX2_X1 U8193 ( .A(n6501), .B(P1_REG1_REG_1__SCAN_IN), .S(n6630), .Z(n6622)
         );
  OAI21_X1 U8194 ( .B1(n6730), .B2(n6623), .A(n6622), .ZN(n6624) );
  NAND3_X1 U8195 ( .A1(n9806), .A2(n6625), .A3(n6624), .ZN(n6626) );
  OAI211_X1 U8196 ( .C1(n9817), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6635)
         );
  INV_X1 U8197 ( .A(n6629), .ZN(n9690) );
  MUX2_X1 U8198 ( .A(n6826), .B(P1_REG2_REG_1__SCAN_IN), .S(n6630), .Z(n6633)
         );
  INV_X1 U8199 ( .A(n6631), .ZN(n6632) );
  AOI211_X1 U8200 ( .C1(n9690), .C2(n6633), .A(n6632), .B(n9784), .ZN(n6634)
         );
  AOI211_X1 U8201 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9696), .A(n6635), .B(
        n6634), .ZN(n6636) );
  INV_X1 U8202 ( .A(n6636), .ZN(P1_U3242) );
  INV_X1 U8203 ( .A(n6637), .ZN(n6669) );
  AOI22_X1 U8204 ( .A1(n7333), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8618), .ZN(n6638) );
  OAI21_X1 U8205 ( .B1(n6669), .B2(n6488), .A(n6638), .ZN(P2_U3346) );
  NOR2_X1 U8206 ( .A1(n6647), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6640) );
  NOR2_X1 U8207 ( .A1(n6640), .A2(n6639), .ZN(n6645) );
  INV_X1 U8208 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7513) );
  MUX2_X1 U8209 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7513), .S(n6735), .Z(n6641)
         );
  INV_X1 U8210 ( .A(n6641), .ZN(n6644) );
  INV_X1 U8211 ( .A(n6645), .ZN(n6642) );
  NAND2_X1 U8212 ( .A1(n6642), .A2(n6641), .ZN(n9087) );
  INV_X1 U8213 ( .A(n9087), .ZN(n6643) );
  AOI21_X1 U8214 ( .B1(n6645), .B2(n6644), .A(n6643), .ZN(n6653) );
  NAND2_X1 U8215 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7431) );
  OAI21_X1 U8216 ( .B1(n9817), .B2(n6731), .A(n7431), .ZN(n6651) );
  AOI21_X1 U8217 ( .B1(n6647), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6646), .ZN(
        n6649) );
  XNOR2_X1 U8218 ( .A(n6735), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6648) );
  NOR2_X1 U8219 ( .A1(n6649), .A2(n6648), .ZN(n6734) );
  AOI211_X1 U8220 ( .C1(n6649), .C2(n6648), .A(n9784), .B(n6734), .ZN(n6650)
         );
  AOI211_X1 U8221 ( .C1(n9696), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6651), .B(
        n6650), .ZN(n6652) );
  OAI21_X1 U8222 ( .B1(n6653), .B2(n9823), .A(n6652), .ZN(P1_U3251) );
  INV_X1 U8223 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8224 ( .A1(n7737), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U8225 ( .B1(n6085), .B2(n6655), .A(n6654), .ZN(n6660) );
  INV_X1 U8226 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U8227 ( .A1(n6656), .A2(n10489), .ZN(n6657) );
  NAND2_X1 U8228 ( .A1(n6663), .A2(n6657), .ZN(n8336) );
  NAND2_X1 U8229 ( .A1(n7637), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U8230 ( .B1(n8336), .B2(n7648), .A(n6658), .ZN(n6659) );
  NAND2_X1 U8231 ( .A1(n8317), .A2(P2_U3966), .ZN(n6661) );
  OAI21_X1 U8232 ( .B1(n5744), .B2(P2_U3966), .A(n6661), .ZN(P2_U3574) );
  INV_X1 U8233 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6667) );
  INV_X1 U8234 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U8235 ( .A1(n6663), .A2(n10461), .ZN(n6664) );
  NAND2_X1 U8236 ( .A1(n7601), .A2(n6664), .ZN(n8321) );
  OR2_X1 U8237 ( .A1(n8321), .A2(n7648), .ZN(n6666) );
  OAI211_X1 U8238 ( .C1(n4481), .C2(n6667), .A(n6666), .B(n6665), .ZN(n7840)
         );
  NAND2_X1 U8239 ( .A1(n7840), .A2(P2_U3966), .ZN(n6668) );
  OAI21_X1 U8240 ( .B1(n5766), .B2(P2_U3966), .A(n6668), .ZN(P2_U3575) );
  INV_X1 U8241 ( .A(n9094), .ZN(n9108) );
  OAI222_X1 U8242 ( .A1(n9595), .A2(n6670), .B1(n7594), .B2(n6669), .C1(
        P1_U3084), .C2(n9108), .ZN(P1_U3341) );
  OAI21_X1 U8243 ( .B1(n6673), .B2(n6671), .A(n6672), .ZN(n9689) );
  INV_X1 U8244 ( .A(n9689), .ZN(n6679) );
  INV_X1 U8245 ( .A(n8751), .ZN(n8772) );
  INV_X1 U8246 ( .A(n9881), .ZN(n6805) );
  AND2_X1 U8247 ( .A1(n6809), .A2(n6805), .ZN(n6675) );
  OAI211_X1 U8248 ( .C1(n6676), .C2(n9647), .A(n6675), .B(n6674), .ZN(n7582)
         );
  INV_X1 U8249 ( .A(n4480), .ZN(n6859) );
  INV_X1 U8250 ( .A(n7572), .ZN(n6852) );
  OAI22_X1 U8251 ( .A1(n6859), .A2(n8768), .B1(n8760), .B2(n6852), .ZN(n6677)
         );
  AOI21_X1 U8252 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7582), .A(n6677), .ZN(
        n6678) );
  OAI21_X1 U8253 ( .B1(n6679), .B2(n8772), .A(n6678), .ZN(P1_U3230) );
  INV_X1 U8254 ( .A(n6680), .ZN(n6703) );
  AOI22_X1 U8255 ( .A1(n7353), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8618), .ZN(n6681) );
  OAI21_X1 U8256 ( .B1(n6703), .B2(n6488), .A(n6681), .ZN(P2_U3345) );
  NAND2_X1 U8257 ( .A1(n6682), .A2(n6768), .ZN(n6761) );
  INV_X1 U8258 ( .A(n6761), .ZN(n6765) );
  AOI21_X1 U8259 ( .B1(n6768), .B2(n7722), .A(n6765), .ZN(n6688) );
  OR2_X1 U8260 ( .A1(n6884), .A2(n8434), .ZN(n10005) );
  INV_X1 U8261 ( .A(n10005), .ZN(n6684) );
  OR2_X1 U8262 ( .A1(n7810), .A2(n7722), .ZN(n7808) );
  INV_X1 U8263 ( .A(n7808), .ZN(n7822) );
  INV_X1 U8264 ( .A(n6768), .ZN(n10007) );
  NAND2_X1 U8265 ( .A1(n8088), .A2(n10007), .ZN(n9985) );
  INV_X1 U8266 ( .A(n9985), .ZN(n6683) );
  AOI22_X1 U8267 ( .A1(n6684), .A2(n7819), .B1(n7822), .B2(n6683), .ZN(n6687)
         );
  OR2_X1 U8268 ( .A1(n6685), .A2(P2_U3152), .ZN(n6714) );
  AOI22_X1 U8269 ( .A1(n6714), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n7793), .B2(
        n6768), .ZN(n6686) );
  OAI211_X1 U8270 ( .C1(n6688), .C2(n7810), .A(n6687), .B(n6686), .ZN(P2_U3234) );
  OR2_X1 U8271 ( .A1(n6870), .A2(n8434), .ZN(n6690) );
  NAND2_X1 U8272 ( .A1(n8088), .A2(n8469), .ZN(n6689) );
  NAND2_X1 U8273 ( .A1(n6690), .A2(n6689), .ZN(n6766) );
  INV_X1 U8274 ( .A(n6766), .ZN(n6698) );
  OAI21_X1 U8275 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6694) );
  INV_X1 U8276 ( .A(n7810), .ZN(n7823) );
  NAND2_X1 U8277 ( .A1(n6694), .A2(n7823), .ZN(n6696) );
  AOI22_X1 U8278 ( .A1(n6714), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n7793), .B2(
        n6769), .ZN(n6695) );
  OAI211_X1 U8279 ( .C1(n6698), .C2(n6697), .A(n6696), .B(n6695), .ZN(P2_U3224) );
  CLKBUF_X2 U8280 ( .A(P1_U4006), .Z(n9692) );
  NAND2_X1 U8281 ( .A1(n9313), .A2(n9692), .ZN(n6699) );
  OAI21_X1 U8282 ( .B1(n9692), .B2(n5767), .A(n6699), .ZN(P1_U3578) );
  INV_X1 U8283 ( .A(n6700), .ZN(n6702) );
  AOI22_X1 U8284 ( .A1(n7492), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n8618), .ZN(n6701) );
  OAI21_X1 U8285 ( .B1(n6702), .B2(n6488), .A(n6701), .ZN(P2_U3344) );
  INV_X1 U8286 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10245) );
  OAI222_X1 U8287 ( .A1(n7594), .A2(n6702), .B1(n9761), .B2(P1_U3084), .C1(
        n10245), .C2(n9595), .ZN(P1_U3339) );
  INV_X1 U8288 ( .A(n9746), .ZN(n9109) );
  OAI222_X1 U8289 ( .A1(n9595), .A2(n10236), .B1(n9109), .B2(P1_U3084), .C1(
        n9599), .C2(n6703), .ZN(P1_U3340) );
  XNOR2_X1 U8290 ( .A(n6705), .B(n6704), .ZN(n6706) );
  XNOR2_X1 U8291 ( .A(n6707), .B(n6706), .ZN(n6711) );
  INV_X1 U8292 ( .A(n8755), .ZN(n8765) );
  AOI22_X1 U8293 ( .A1(n8765), .A2(n6803), .B1(n8757), .B2(n6850), .ZN(n6708)
         );
  OAI21_X1 U8294 ( .B1(n6801), .B2(n8760), .A(n6708), .ZN(n6709) );
  AOI21_X1 U8295 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7582), .A(n6709), .ZN(
        n6710) );
  OAI21_X1 U8296 ( .B1(n6711), .B2(n8772), .A(n6710), .ZN(P1_U3220) );
  XNOR2_X1 U8297 ( .A(n6713), .B(n6712), .ZN(n6717) );
  AOI22_X1 U8298 ( .A1(n6714), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n7793), .B2(
        n6869), .ZN(n6716) );
  INV_X1 U8299 ( .A(n7829), .ZN(n7694) );
  INV_X1 U8300 ( .A(n6901), .ZN(n8085) );
  AOI22_X1 U8301 ( .A1(n7745), .A2(n6759), .B1(n7694), .B2(n8085), .ZN(n6715)
         );
  OAI211_X1 U8302 ( .C1(n6717), .C2(n7810), .A(n6716), .B(n6715), .ZN(P2_U3239) );
  AND2_X1 U8303 ( .A1(n6809), .A2(n6718), .ZN(n6720) );
  AND2_X1 U8304 ( .A1(n6719), .A2(n6805), .ZN(n9879) );
  OAI211_X1 U8305 ( .C1(n7504), .C2(n8979), .A(n6720), .B(n9879), .ZN(n6727)
         );
  INV_X2 U8306 ( .A(n9940), .ZN(n9906) );
  INV_X1 U8307 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6726) );
  INV_X1 U8308 ( .A(n6813), .ZN(n6724) );
  AND2_X1 U8309 ( .A1(n6803), .A2(n6852), .ZN(n8795) );
  NOR2_X1 U8310 ( .A1(n6819), .A2(n8795), .ZN(n8996) );
  INV_X1 U8311 ( .A(n6816), .ZN(n6722) );
  NOR3_X1 U8312 ( .A1(n8996), .A2(n6722), .A3(n6813), .ZN(n6723) );
  AOI21_X1 U8313 ( .B1(n9635), .B2(n4480), .A(n6723), .ZN(n7575) );
  OAI21_X1 U8314 ( .B1(n6852), .B2(n6724), .A(n7575), .ZN(n6728) );
  NAND2_X1 U8315 ( .A1(n6728), .A2(n9906), .ZN(n6725) );
  OAI21_X1 U8316 ( .B1(n9906), .B2(n6726), .A(n6725), .ZN(P1_U3454) );
  INV_X2 U8317 ( .A(n9957), .ZN(n9948) );
  NAND2_X1 U8318 ( .A1(n6728), .A2(n9948), .ZN(n6729) );
  OAI21_X1 U8319 ( .B1(n9948), .B2(n6730), .A(n6729), .ZN(P1_U3523) );
  INV_X1 U8320 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U8321 ( .A1(n6731), .A2(n7513), .ZN(n9085) );
  MUX2_X1 U8322 ( .A(n9674), .B(P1_REG1_REG_11__SCAN_IN), .S(n6738), .Z(n9086)
         );
  AOI21_X1 U8323 ( .B1(n9087), .B2(n9085), .A(n9086), .ZN(n9089) );
  AOI21_X1 U8324 ( .B1(n9674), .B2(n9082), .A(n9089), .ZN(n6733) );
  INV_X1 U8325 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U8326 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9108), .B1(n9094), .B2(
        n9667), .ZN(n6732) );
  NOR2_X1 U8327 ( .A1(n6733), .A2(n6732), .ZN(n9107) );
  AOI21_X1 U8328 ( .B1(n6733), .B2(n6732), .A(n9107), .ZN(n6745) );
  NAND2_X1 U8329 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8667) );
  OAI21_X1 U8330 ( .B1(n9817), .B2(n9108), .A(n8667), .ZN(n6743) );
  AOI21_X1 U8331 ( .B1(n6735), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6734), .ZN(
        n9080) );
  INV_X1 U8332 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8333 ( .A(n6736), .B(P1_REG2_REG_11__SCAN_IN), .S(n6738), .Z(n6737)
         );
  INV_X1 U8334 ( .A(n6737), .ZN(n9079) );
  NAND2_X1 U8335 ( .A1(n9080), .A2(n9079), .ZN(n9078) );
  OAI21_X1 U8336 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6738), .A(n9078), .ZN(
        n6741) );
  NAND2_X1 U8337 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9094), .ZN(n6739) );
  OAI21_X1 U8338 ( .B1(n9094), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6739), .ZN(
        n6740) );
  NOR2_X1 U8339 ( .A1(n6741), .A2(n6740), .ZN(n9093) );
  AOI211_X1 U8340 ( .C1(n6741), .C2(n6740), .A(n9784), .B(n9093), .ZN(n6742)
         );
  AOI211_X1 U8341 ( .C1(n9696), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6743), .B(
        n6742), .ZN(n6744) );
  OAI21_X1 U8342 ( .B1(n6745), .B2(n9823), .A(n6744), .ZN(P1_U3253) );
  XNOR2_X1 U8343 ( .A(n6747), .B(n6746), .ZN(n6750) );
  OAI22_X1 U8344 ( .A1(n6870), .A2(n8491), .B1(n7050), .B2(n8434), .ZN(n6926)
         );
  AOI22_X1 U8345 ( .A1(n6926), .A2(n7819), .B1(n6935), .B2(n7793), .ZN(n6749)
         );
  MUX2_X1 U8346 ( .A(n7828), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6748) );
  OAI211_X1 U8347 ( .C1(n6750), .C2(n7810), .A(n6749), .B(n6748), .ZN(P2_U3220) );
  INV_X1 U8348 ( .A(n6751), .ZN(n6789) );
  AOI22_X1 U8349 ( .A1(n8122), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8618), .ZN(n6752) );
  OAI21_X1 U8350 ( .B1(n6789), .B2(n6488), .A(n6752), .ZN(P2_U3343) );
  NAND4_X1 U8351 ( .A1(n6754), .A2(n9996), .A3(n6753), .A4(n6879), .ZN(n6756)
         );
  NOR2_X1 U8352 ( .A1(n6756), .A2(n6755), .ZN(n6773) );
  INV_X1 U8353 ( .A(n6881), .ZN(n6757) );
  AND2_X2 U8354 ( .A1(n6773), .A2(n6757), .ZN(n10083) );
  XNOR2_X1 U8355 ( .A(n8069), .B(n6883), .ZN(n6758) );
  NAND2_X1 U8356 ( .A1(n6758), .A2(n8275), .ZN(n7241) );
  NAND2_X1 U8357 ( .A1(n7241), .A2(n10056), .ZN(n10069) );
  INV_X1 U8358 ( .A(n6769), .ZN(n6914) );
  NAND2_X1 U8359 ( .A1(n8088), .A2(n6768), .ZN(n6760) );
  OAI21_X1 U8360 ( .B1(n6764), .B2(n6760), .A(n6886), .ZN(n6919) );
  INV_X1 U8361 ( .A(n6919), .ZN(n6771) );
  INV_X1 U8362 ( .A(n8024), .ZN(n8033) );
  NAND2_X1 U8363 ( .A1(n7890), .A2(n8033), .ZN(n7876) );
  INV_X1 U8364 ( .A(n6871), .ZN(n6762) );
  NOR2_X1 U8365 ( .A1(n6872), .A2(n6762), .ZN(n6763) );
  AOI211_X1 U8366 ( .C1(n6765), .C2(n6764), .A(n8486), .B(n6763), .ZN(n6767)
         );
  NOR2_X1 U8367 ( .A1(n6767), .A2(n6766), .ZN(n6922) );
  AOI211_X1 U8368 ( .C1(n6768), .C2(n6769), .A(n10065), .B(n6889), .ZN(n6918)
         );
  AOI21_X1 U8369 ( .B1(n10073), .B2(n6769), .A(n6918), .ZN(n6770) );
  OAI211_X1 U8370 ( .C1(n10078), .C2(n6771), .A(n6922), .B(n6770), .ZN(n6774)
         );
  NAND2_X1 U8371 ( .A1(n6774), .A2(n10083), .ZN(n6772) );
  OAI21_X1 U8372 ( .B1(n10083), .B2(n6016), .A(n6772), .ZN(P2_U3454) );
  AND2_X2 U8373 ( .A1(n6773), .A2(n6881), .ZN(n10097) );
  NAND2_X1 U8374 ( .A1(n6774), .A2(n10097), .ZN(n6775) );
  OAI21_X1 U8375 ( .B1(n10097), .B2(n7133), .A(n6775), .ZN(P2_U3521) );
  INV_X1 U8376 ( .A(n6776), .ZN(n6799) );
  AOI22_X1 U8377 ( .A1(n8135), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8618), .ZN(n6777) );
  OAI21_X1 U8378 ( .B1(n6799), .B2(n6488), .A(n6777), .ZN(P2_U3342) );
  INV_X1 U8379 ( .A(n6778), .ZN(n6779) );
  NOR2_X1 U8380 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  XNOR2_X1 U8381 ( .A(n6782), .B(n6781), .ZN(n6788) );
  INV_X1 U8382 ( .A(n6907), .ZN(n6786) );
  INV_X1 U8383 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U8384 ( .A1(n10356), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7227) );
  INV_X1 U8385 ( .A(n7227), .ZN(n6783) );
  OAI21_X1 U8386 ( .B1(n7835), .B2(n10023), .A(n6783), .ZN(n6785) );
  OAI22_X1 U8387 ( .A1(n7830), .A2(n6901), .B1(n6988), .B2(n7829), .ZN(n6784)
         );
  AOI211_X1 U8388 ( .C1(n6786), .C2(n7805), .A(n6785), .B(n6784), .ZN(n6787)
         );
  OAI21_X1 U8389 ( .B1(n6788), .B2(n7810), .A(n6787), .ZN(P2_U3232) );
  INV_X1 U8390 ( .A(n9775), .ZN(n9111) );
  OAI222_X1 U8391 ( .A1(n9595), .A2(n6790), .B1(n7594), .B2(n6789), .C1(
        P1_U3084), .C2(n9111), .ZN(P1_U3338) );
  INV_X1 U8392 ( .A(n8764), .ZN(n8733) );
  OAI21_X1 U8393 ( .B1(n6793), .B2(n6792), .A(n6791), .ZN(n6794) );
  NAND2_X1 U8394 ( .A1(n6794), .A2(n8751), .ZN(n6798) );
  OAI22_X1 U8395 ( .A1(n8760), .A2(n9894), .B1(n6939), .B2(n8755), .ZN(n6795)
         );
  AOI211_X1 U8396 ( .C1(n8757), .C2(n9076), .A(n6796), .B(n6795), .ZN(n6797)
         );
  OAI211_X1 U8397 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8733), .A(n6798), .B(
        n6797), .ZN(P1_U3216) );
  INV_X1 U8398 ( .A(n9789), .ZN(n6800) );
  OAI222_X1 U8399 ( .A1(n9595), .A2(n10445), .B1(n6800), .B2(P1_U3084), .C1(
        n9599), .C2(n6799), .ZN(P1_U3337) );
  NAND2_X1 U8400 ( .A1(n6804), .A2(n6818), .ZN(n6849) );
  OAI21_X1 U8401 ( .B1(n6818), .B2(n6804), .A(n6849), .ZN(n9882) );
  AND2_X1 U8402 ( .A1(n6806), .A2(n6805), .ZN(n6807) );
  AND2_X1 U8403 ( .A1(n6808), .A2(n6807), .ZN(n7110) );
  NAND2_X1 U8404 ( .A1(n7110), .A2(n6809), .ZN(n6810) );
  NOR2_X1 U8405 ( .A1(n6811), .A2(n9327), .ZN(n6812) );
  AND2_X1 U8406 ( .A1(n9874), .A2(n6812), .ZN(n9834) );
  INV_X1 U8407 ( .A(n9834), .ZN(n6830) );
  XNOR2_X1 U8408 ( .A(n6801), .B(n7572), .ZN(n6814) );
  NAND2_X1 U8409 ( .A1(n6814), .A2(n9856), .ZN(n9883) );
  NOR2_X1 U8410 ( .A1(n9883), .A2(n9863), .ZN(n6824) );
  NAND2_X1 U8411 ( .A1(n6816), .A2(n6815), .ZN(n7101) );
  OR2_X1 U8412 ( .A1(n7101), .A2(n9863), .ZN(n9843) );
  AOI22_X1 U8413 ( .A1(n9632), .A2(n6803), .B1(n6850), .B2(n9635), .ZN(n6823)
         );
  NAND2_X1 U8414 ( .A1(n8995), .A2(n6819), .ZN(n6861) );
  OAI21_X1 U8415 ( .B1(n8995), .B2(n6819), .A(n6861), .ZN(n6821) );
  NAND2_X1 U8416 ( .A1(n9063), .A2(n9863), .ZN(n8980) );
  NAND2_X1 U8417 ( .A1(n8979), .A2(n5909), .ZN(n6820) );
  NAND2_X1 U8418 ( .A1(n8980), .A2(n6820), .ZN(n9840) );
  NAND2_X1 U8419 ( .A1(n6821), .A2(n9840), .ZN(n6822) );
  OAI211_X1 U8420 ( .C1(n9882), .C2(n9843), .A(n6823), .B(n6822), .ZN(n9884)
         );
  AOI211_X1 U8421 ( .C1(n9861), .C2(P1_REG3_REG_1__SCAN_IN), .A(n6824), .B(
        n9884), .ZN(n6825) );
  MUX2_X1 U8422 ( .A(n6826), .B(n6825), .S(n9874), .Z(n6829) );
  INV_X1 U8423 ( .A(n6827), .ZN(n9859) );
  NAND2_X1 U8424 ( .A1(n9874), .A2(n9859), .ZN(n9845) );
  INV_X1 U8425 ( .A(n6801), .ZN(n6858) );
  NAND2_X1 U8426 ( .A1(n9644), .A2(n6858), .ZN(n6828) );
  OAI211_X1 U8427 ( .C1(n9882), .C2(n6830), .A(n6829), .B(n6828), .ZN(P1_U3290) );
  INV_X1 U8428 ( .A(n6831), .ZN(n6846) );
  AOI22_X1 U8429 ( .A1(n8156), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8623), .ZN(n6832) );
  OAI21_X1 U8430 ( .B1(n6846), .B2(n6488), .A(n6832), .ZN(P2_U3341) );
  INV_X1 U8431 ( .A(n6951), .ZN(n6845) );
  AND2_X1 U8432 ( .A1(n6791), .A2(n6833), .ZN(n6836) );
  OAI211_X1 U8433 ( .C1(n6836), .C2(n6835), .A(n8751), .B(n6834), .ZN(n6844)
         );
  NAND2_X1 U8434 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9718) );
  INV_X1 U8435 ( .A(n9718), .ZN(n6842) );
  OAI22_X1 U8436 ( .A1(n8760), .A2(n9900), .B1(n6945), .B2(n8755), .ZN(n6841)
         );
  AOI211_X1 U8437 ( .C1(n8757), .C2(n9075), .A(n6842), .B(n6841), .ZN(n6843)
         );
  OAI211_X1 U8438 ( .C1(n8733), .C2(n6845), .A(n6844), .B(n6843), .ZN(P1_U3228) );
  INV_X1 U8439 ( .A(n9114), .ZN(n9802) );
  OAI222_X1 U8440 ( .A1(n9595), .A2(n6847), .B1(n9802), .B2(P1_U3084), .C1(
        n7594), .C2(n6846), .ZN(P1_U3336) );
  NAND2_X1 U8441 ( .A1(n4480), .A2(n6858), .ZN(n6848) );
  AND2_X1 U8442 ( .A1(n6849), .A2(n6848), .ZN(n6851) );
  NAND2_X1 U8443 ( .A1(n6939), .A2(n4483), .ZN(n8799) );
  NAND2_X1 U8444 ( .A1(n6850), .A2(n9888), .ZN(n8800) );
  NAND2_X1 U8445 ( .A1(n6851), .A2(n6857), .ZN(n6941) );
  OAI21_X1 U8446 ( .B1(n6851), .B2(n6857), .A(n6941), .ZN(n9892) );
  NAND2_X1 U8447 ( .A1(n9874), .A2(n9327), .ZN(n9376) );
  NAND2_X1 U8448 ( .A1(n6801), .A2(n6852), .ZN(n6853) );
  NAND2_X1 U8449 ( .A1(n6853), .A2(n4483), .ZN(n6854) );
  NAND2_X1 U8450 ( .A1(n6961), .A2(n6854), .ZN(n9889) );
  AOI22_X1 U8451 ( .A1(n9644), .A2(n4483), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9861), .ZN(n6856) );
  OAI21_X1 U8452 ( .B1(n9455), .B2(n9889), .A(n6856), .ZN(n6867) );
  INV_X1 U8453 ( .A(n9843), .ZN(n9639) );
  NAND2_X1 U8454 ( .A1(n9892), .A2(n9639), .ZN(n6865) );
  AOI22_X1 U8455 ( .A1(n9632), .A2(n4480), .B1(n9077), .B2(n9635), .ZN(n6864)
         );
  INV_X1 U8456 ( .A(n6857), .ZN(n8997) );
  NAND2_X1 U8457 ( .A1(n6859), .A2(n6858), .ZN(n6860) );
  NAND2_X1 U8458 ( .A1(n8802), .A2(n8997), .ZN(n6944) );
  OAI21_X1 U8459 ( .B1(n8997), .B2(n8802), .A(n6944), .ZN(n6862) );
  NAND2_X1 U8460 ( .A1(n6862), .A2(n9840), .ZN(n6863) );
  NAND3_X1 U8461 ( .A1(n6865), .A2(n6864), .A3(n6863), .ZN(n9890) );
  MUX2_X1 U8462 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9890), .S(n9874), .Z(n6866)
         );
  AOI211_X1 U8463 ( .C1(n9834), .C2(n9892), .A(n6867), .B(n6866), .ZN(n6868)
         );
  INV_X1 U8464 ( .A(n6868), .ZN(P1_U3289) );
  INV_X1 U8465 ( .A(n6870), .ZN(n8086) );
  NAND2_X1 U8466 ( .A1(n8086), .A2(n10011), .ZN(n7891) );
  NAND2_X1 U8467 ( .A1(n6870), .A2(n6869), .ZN(n7893) );
  NAND2_X1 U8468 ( .A1(n7891), .A2(n7893), .ZN(n8029) );
  INV_X1 U8469 ( .A(n6876), .ZN(n6874) );
  NAND2_X1 U8470 ( .A1(n6874), .A2(n6873), .ZN(n6896) );
  INV_X1 U8471 ( .A(n6896), .ZN(n6875) );
  AOI21_X1 U8472 ( .B1(n8029), .B2(n6876), .A(n6875), .ZN(n6877) );
  OAI222_X1 U8473 ( .A1(n8434), .A2(n6901), .B1(n8491), .B2(n6884), .C1(n8486), 
        .C2(n6877), .ZN(n10013) );
  INV_X1 U8474 ( .A(n10013), .ZN(n6895) );
  NAND2_X1 U8475 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  NOR2_X1 U8476 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  NAND2_X1 U8477 ( .A1(n6882), .A2(n9996), .ZN(n6888) );
  INV_X1 U8478 ( .A(n9993), .ZN(n8289) );
  OR2_X1 U8479 ( .A1(n6883), .A2(n8275), .ZN(n8449) );
  NAND2_X1 U8480 ( .A1(n7241), .A2(n8449), .ZN(n9986) );
  INV_X1 U8481 ( .A(n8501), .ZN(n8329) );
  NAND2_X1 U8482 ( .A1(n6884), .A2(n6914), .ZN(n6885) );
  OAI21_X1 U8483 ( .B1(n6887), .B2(n8029), .A(n6900), .ZN(n10015) );
  OR2_X1 U8484 ( .A1(n6888), .A2(n9980), .ZN(n7385) );
  NAND2_X1 U8485 ( .A1(n8427), .A2(n10074), .ZN(n9989) );
  NAND2_X1 U8486 ( .A1(n6889), .A2(n10011), .ZN(n6930) );
  OAI21_X1 U8487 ( .B1(n6889), .B2(n10011), .A(n6930), .ZN(n10012) );
  NOR2_X1 U8488 ( .A1(n8451), .A2(n10285), .ZN(n6891) );
  NOR2_X1 U8489 ( .A1(n9988), .A2(n10011), .ZN(n6890) );
  AOI211_X1 U8490 ( .C1(n8289), .C2(P2_REG2_REG_2__SCAN_IN), .A(n6891), .B(
        n6890), .ZN(n6892) );
  OAI21_X1 U8491 ( .B1(n9989), .B2(n10012), .A(n6892), .ZN(n6893) );
  AOI21_X1 U8492 ( .B1(n8329), .B2(n10015), .A(n6893), .ZN(n6894) );
  OAI21_X1 U8493 ( .B1(n6895), .B2(n8289), .A(n6894), .ZN(P2_U3294) );
  NAND2_X1 U8494 ( .A1(n6901), .A2(n6935), .ZN(n6993) );
  INV_X1 U8495 ( .A(n6935), .ZN(n10018) );
  NAND2_X1 U8496 ( .A1(n8085), .A2(n10018), .ZN(n7903) );
  NAND2_X1 U8497 ( .A1(n6993), .A2(n7903), .ZN(n8031) );
  NAND2_X1 U8498 ( .A1(n6925), .A2(n4478), .ZN(n6994) );
  NAND2_X1 U8499 ( .A1(n6994), .A2(n6993), .ZN(n6897) );
  NAND2_X1 U8500 ( .A1(n7050), .A2(n6904), .ZN(n7881) );
  NAND2_X1 U8501 ( .A1(n7881), .A2(n7045), .ZN(n8032) );
  XNOR2_X1 U8502 ( .A(n6897), .B(n8032), .ZN(n6898) );
  OAI222_X1 U8503 ( .A1(n8434), .A2(n6988), .B1(n8491), .B2(n6901), .C1(n6898), 
        .C2(n8486), .ZN(n10024) );
  INV_X1 U8504 ( .A(n10024), .ZN(n6913) );
  NAND2_X1 U8505 ( .A1(n6870), .A2(n10011), .ZN(n6899) );
  NAND2_X1 U8506 ( .A1(n6901), .A2(n10018), .ZN(n6902) );
  OAI21_X1 U8507 ( .B1(n6903), .B2(n8032), .A(n6987), .ZN(n10026) );
  OR2_X1 U8508 ( .A1(n6930), .A2(n6935), .ZN(n6931) );
  INV_X1 U8509 ( .A(n6931), .ZN(n6906) );
  INV_X1 U8510 ( .A(n7042), .ZN(n6905) );
  OAI211_X1 U8511 ( .C1(n10023), .C2(n6906), .A(n6905), .B(n10074), .ZN(n10022) );
  NOR2_X1 U8512 ( .A1(n8451), .A2(n6907), .ZN(n6909) );
  NOR2_X1 U8513 ( .A1(n9988), .A2(n10023), .ZN(n6908) );
  AOI211_X1 U8514 ( .C1(n8289), .C2(P2_REG2_REG_4__SCAN_IN), .A(n6909), .B(
        n6908), .ZN(n6910) );
  OAI21_X1 U8515 ( .B1(n10022), .B2(n7385), .A(n6910), .ZN(n6911) );
  AOI21_X1 U8516 ( .B1(n10026), .B2(n8329), .A(n6911), .ZN(n6912) );
  OAI21_X1 U8517 ( .B1(n6913), .B2(n8289), .A(n6912), .ZN(P2_U3292) );
  NOR2_X1 U8518 ( .A1(n9988), .A2(n6914), .ZN(n6917) );
  OAI22_X1 U8519 ( .A1(n9993), .A2(n6445), .B1(n6915), .B2(n8451), .ZN(n6916)
         );
  AOI211_X1 U8520 ( .C1(n6918), .C2(n8427), .A(n6917), .B(n6916), .ZN(n6921)
         );
  NAND2_X1 U8521 ( .A1(n6919), .A2(n8329), .ZN(n6920) );
  OAI211_X1 U8522 ( .C1(n6922), .C2(n8289), .A(n6921), .B(n6920), .ZN(P2_U3295) );
  OAI21_X1 U8523 ( .B1(n6924), .B2(n8031), .A(n6923), .ZN(n10021) );
  INV_X1 U8524 ( .A(n10021), .ZN(n6938) );
  XNOR2_X1 U8525 ( .A(n8031), .B(n6925), .ZN(n6928) );
  INV_X1 U8526 ( .A(n6926), .ZN(n6927) );
  OAI21_X1 U8527 ( .B1(n6928), .B2(n8486), .A(n6927), .ZN(n10020) );
  NAND2_X1 U8528 ( .A1(n10020), .A2(n9993), .ZN(n6937) );
  INV_X1 U8529 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6929) );
  OAI22_X1 U8530 ( .A1(n9993), .A2(n6929), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8451), .ZN(n6934) );
  INV_X1 U8531 ( .A(n6930), .ZN(n6932) );
  OAI211_X1 U8532 ( .C1(n6932), .C2(n10018), .A(n10074), .B(n6931), .ZN(n10016) );
  NOR2_X1 U8533 ( .A1(n10016), .A2(n7385), .ZN(n6933) );
  AOI211_X1 U8534 ( .C1(n8455), .C2(n6935), .A(n6934), .B(n6933), .ZN(n6936)
         );
  OAI211_X1 U8535 ( .C1(n6938), .C2(n8501), .A(n6937), .B(n6936), .ZN(P2_U3293) );
  NAND2_X1 U8536 ( .A1(n6939), .A2(n9888), .ZN(n6940) );
  NAND2_X1 U8537 ( .A1(n6941), .A2(n6940), .ZN(n6960) );
  NAND2_X1 U8538 ( .A1(n6945), .A2(n6964), .ZN(n9026) );
  NAND2_X1 U8539 ( .A1(n9077), .A2(n9894), .ZN(n8804) );
  NAND2_X1 U8540 ( .A1(n9026), .A2(n8804), .ZN(n8994) );
  NAND2_X1 U8541 ( .A1(n6960), .A2(n8994), .ZN(n6943) );
  NAND2_X1 U8542 ( .A1(n6945), .A2(n9894), .ZN(n6942) );
  NAND2_X1 U8543 ( .A1(n6943), .A2(n6942), .ZN(n7093) );
  INV_X1 U8544 ( .A(n9076), .ZN(n9870) );
  NAND2_X1 U8545 ( .A1(n9870), .A2(n6952), .ZN(n9025) );
  NAND2_X1 U8546 ( .A1(n9076), .A2(n9900), .ZN(n9028) );
  NAND2_X1 U8547 ( .A1(n9025), .A2(n9028), .ZN(n8993) );
  XOR2_X1 U8548 ( .A(n7093), .B(n8993), .Z(n6949) );
  NAND2_X1 U8549 ( .A1(n6944), .A2(n8799), .ZN(n6966) );
  NAND2_X1 U8550 ( .A1(n6966), .A2(n8804), .ZN(n9027) );
  NAND2_X1 U8551 ( .A1(n9027), .A2(n9026), .ZN(n8875) );
  XOR2_X1 U8552 ( .A(n8875), .B(n8993), .Z(n6947) );
  INV_X1 U8553 ( .A(n9075), .ZN(n7096) );
  INV_X1 U8554 ( .A(n9635), .ZN(n9869) );
  OAI22_X1 U8555 ( .A1(n7096), .A2(n9869), .B1(n6945), .B2(n9871), .ZN(n6946)
         );
  AOI21_X1 U8556 ( .B1(n6947), .B2(n9840), .A(n6946), .ZN(n6948) );
  OAI21_X1 U8557 ( .B1(n6949), .B2(n9843), .A(n6948), .ZN(n9902) );
  INV_X1 U8558 ( .A(n9902), .ZN(n6957) );
  INV_X2 U8559 ( .A(n9874), .ZN(n9640) );
  INV_X1 U8560 ( .A(n6949), .ZN(n9904) );
  AND2_X1 U8561 ( .A1(n6963), .A2(n6952), .ZN(n6950) );
  OR2_X1 U8562 ( .A1(n6950), .A2(n9857), .ZN(n9901) );
  AOI22_X1 U8563 ( .A1(n9640), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6951), .B2(
        n9861), .ZN(n6954) );
  NAND2_X1 U8564 ( .A1(n9644), .A2(n6952), .ZN(n6953) );
  OAI211_X1 U8565 ( .C1(n9901), .C2(n9455), .A(n6954), .B(n6953), .ZN(n6955)
         );
  AOI21_X1 U8566 ( .B1(n9904), .B2(n9834), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8567 ( .B1(n6957), .B2(n9640), .A(n6956), .ZN(P1_U3287) );
  INV_X1 U8568 ( .A(n6958), .ZN(n6973) );
  AOI22_X1 U8569 ( .A1(n8157), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8618), .ZN(n6959) );
  OAI21_X1 U8570 ( .B1(n6973), .B2(n6488), .A(n6959), .ZN(P2_U3340) );
  XNOR2_X1 U8571 ( .A(n6960), .B(n8994), .ZN(n9898) );
  NAND2_X1 U8572 ( .A1(n6961), .A2(n6964), .ZN(n6962) );
  NAND2_X1 U8573 ( .A1(n6963), .A2(n6962), .ZN(n9895) );
  AOI22_X1 U8574 ( .A1(n9644), .A2(n6964), .B1(n5234), .B2(n9861), .ZN(n6965)
         );
  OAI21_X1 U8575 ( .B1(n9455), .B2(n9895), .A(n6965), .ZN(n6971) );
  INV_X1 U8576 ( .A(n9840), .ZN(n9866) );
  XNOR2_X1 U8577 ( .A(n6966), .B(n8994), .ZN(n6969) );
  NAND2_X1 U8578 ( .A1(n9898), .A2(n9639), .ZN(n6968) );
  AOI22_X1 U8579 ( .A1(n9635), .A2(n9076), .B1(n6850), .B2(n9632), .ZN(n6967)
         );
  OAI211_X1 U8580 ( .C1(n9866), .C2(n6969), .A(n6968), .B(n6967), .ZN(n9896)
         );
  MUX2_X1 U8581 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9896), .S(n9874), .Z(n6970)
         );
  AOI211_X1 U8582 ( .C1(n9834), .C2(n9898), .A(n6971), .B(n6970), .ZN(n6972)
         );
  INV_X1 U8583 ( .A(n6972), .ZN(P1_U3288) );
  INV_X1 U8584 ( .A(n9104), .ZN(n9818) );
  OAI222_X1 U8585 ( .A1(n9595), .A2(n10326), .B1(n7594), .B2(n6973), .C1(
        P1_U3084), .C2(n9818), .ZN(P1_U3335) );
  INV_X1 U8586 ( .A(n6974), .ZN(n6975) );
  AOI21_X1 U8587 ( .B1(n6980), .B2(n6976), .A(n6975), .ZN(n6985) );
  INV_X1 U8588 ( .A(n10030), .ZN(n6989) );
  NAND2_X1 U8589 ( .A1(n7694), .A2(n8081), .ZN(n6978) );
  NOR2_X1 U8590 ( .A1(n10341), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7201) );
  INV_X1 U8591 ( .A(n7201), .ZN(n6977) );
  OAI211_X1 U8592 ( .C1(n7828), .C2(n6990), .A(n6978), .B(n6977), .ZN(n6983)
         );
  NAND3_X1 U8593 ( .A1(n6980), .A2(n7822), .A3(n6979), .ZN(n6981) );
  AOI21_X1 U8594 ( .B1(n6981), .B2(n7830), .A(n6988), .ZN(n6982) );
  AOI211_X1 U8595 ( .C1(n6989), .C2(n7793), .A(n6983), .B(n6982), .ZN(n6984)
         );
  OAI21_X1 U8596 ( .B1(n6985), .B2(n7810), .A(n6984), .ZN(P2_U3241) );
  NAND2_X1 U8597 ( .A1(n7050), .A2(n10023), .ZN(n6986) );
  NAND2_X1 U8598 ( .A1(n6988), .A2(n9975), .ZN(n7884) );
  NAND2_X1 U8599 ( .A1(n7884), .A2(n7902), .ZN(n8030) );
  NAND2_X1 U8600 ( .A1(n7049), .A2(n6989), .ZN(n7913) );
  INV_X1 U8601 ( .A(n7049), .ZN(n8082) );
  NAND2_X1 U8602 ( .A1(n8082), .A2(n10030), .ZN(n7908) );
  XOR2_X1 U8603 ( .A(n7017), .B(n8035), .Z(n10032) );
  INV_X1 U8604 ( .A(n10032), .ZN(n7001) );
  NAND2_X1 U8605 ( .A1(n7043), .A2(n10030), .ZN(n7018) );
  OAI211_X1 U8606 ( .C1(n7043), .C2(n10030), .A(n10074), .B(n7018), .ZN(n10028) );
  INV_X1 U8607 ( .A(n10028), .ZN(n6992) );
  OAI22_X1 U8608 ( .A1(n10030), .A2(n9988), .B1(n8451), .B2(n6990), .ZN(n6991)
         );
  AOI21_X1 U8609 ( .B1(n6992), .B2(n8427), .A(n6991), .ZN(n7000) );
  INV_X1 U8610 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6998) );
  AND2_X1 U8611 ( .A1(n7881), .A2(n6993), .ZN(n7885) );
  NAND2_X1 U8612 ( .A1(n6994), .A2(n7885), .ZN(n7046) );
  NAND2_X1 U8613 ( .A1(n7046), .A2(n7904), .ZN(n6995) );
  NAND2_X1 U8614 ( .A1(n6995), .A2(n7884), .ZN(n6996) );
  OAI21_X1 U8615 ( .B1(n8035), .B2(n6996), .A(n7023), .ZN(n6997) );
  AOI222_X1 U8616 ( .A1(n10004), .A2(n6997), .B1(n8081), .B2(n8471), .C1(n8083), .C2(n8469), .ZN(n10029) );
  MUX2_X1 U8617 ( .A(n6998), .B(n10029), .S(n9993), .Z(n6999) );
  OAI211_X1 U8618 ( .C1(n7001), .C2(n8501), .A(n7000), .B(n6999), .ZN(P2_U3290) );
  INV_X1 U8619 ( .A(n7002), .ZN(n7016) );
  AOI22_X1 U8620 ( .A1(n9980), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n8623), .ZN(n7003) );
  OAI21_X1 U8621 ( .B1(n7016), .B2(n6488), .A(n7003), .ZN(P2_U3339) );
  INV_X1 U8622 ( .A(n9860), .ZN(n7015) );
  OAI21_X1 U8623 ( .B1(n7006), .B2(n7005), .A(n7004), .ZN(n7007) );
  NAND2_X1 U8624 ( .A1(n7007), .A2(n8751), .ZN(n7014) );
  INV_X1 U8625 ( .A(n9858), .ZN(n9908) );
  INV_X1 U8626 ( .A(n7008), .ZN(n7009) );
  AOI21_X1 U8627 ( .B1(n8757), .B2(n9074), .A(n7009), .ZN(n7011) );
  NAND2_X1 U8628 ( .A1(n8765), .A2(n9076), .ZN(n7010) );
  OAI211_X1 U8629 ( .C1(n8760), .C2(n9908), .A(n7011), .B(n7010), .ZN(n7012)
         );
  INV_X1 U8630 ( .A(n7012), .ZN(n7013) );
  OAI211_X1 U8631 ( .C1(n8733), .C2(n7015), .A(n7014), .B(n7013), .ZN(P1_U3225) );
  OAI222_X1 U8632 ( .A1(n9595), .A2(n10330), .B1(n7594), .B2(n7016), .C1(
        P1_U3084), .C2(n9327), .ZN(P1_U3334) );
  NAND2_X1 U8633 ( .A1(n7077), .A2(n10033), .ZN(n7917) );
  INV_X1 U8634 ( .A(n10033), .ZN(n7038) );
  NAND2_X1 U8635 ( .A1(n8081), .A2(n7038), .ZN(n7918) );
  XNOR2_X1 U8636 ( .A(n7239), .B(n8040), .ZN(n10038) );
  NAND2_X1 U8637 ( .A1(n7018), .A2(n10033), .ZN(n7019) );
  NAND2_X1 U8638 ( .A1(n7236), .A2(n7019), .ZN(n10036) );
  INV_X1 U8639 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7020) );
  OAI22_X1 U8640 ( .A1(n9993), .A2(n7020), .B1(n7033), .B2(n8451), .ZN(n7021)
         );
  AOI21_X1 U8641 ( .B1(n8455), .B2(n10033), .A(n7021), .ZN(n7022) );
  OAI21_X1 U8642 ( .B1(n10036), .B2(n9989), .A(n7022), .ZN(n7028) );
  INV_X1 U8643 ( .A(n8040), .ZN(n7024) );
  XNOR2_X1 U8644 ( .A(n7242), .B(n7024), .ZN(n7026) );
  OAI22_X1 U8645 ( .A1(n7049), .A2(n8491), .B1(n7295), .B2(n8434), .ZN(n7025)
         );
  AOI21_X1 U8646 ( .B1(n7026), .B2(n10004), .A(n7025), .ZN(n10035) );
  NOR2_X1 U8647 ( .A1(n10035), .A2(n8289), .ZN(n7027) );
  AOI211_X1 U8648 ( .C1(n8329), .C2(n10038), .A(n7028), .B(n7027), .ZN(n7029)
         );
  INV_X1 U8649 ( .A(n7029), .ZN(P2_U3289) );
  AOI21_X1 U8650 ( .B1(n7031), .B2(n7030), .A(n7810), .ZN(n7032) );
  NAND2_X1 U8651 ( .A1(n7032), .A2(n7073), .ZN(n7037) );
  NOR2_X1 U8652 ( .A1(n7829), .A2(n7295), .ZN(n7035) );
  OAI22_X1 U8653 ( .A1(n7828), .A2(n7033), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6137), .ZN(n7034) );
  AOI211_X1 U8654 ( .C1(n7745), .C2(n8082), .A(n7035), .B(n7034), .ZN(n7036)
         );
  OAI211_X1 U8655 ( .C1(n7038), .C2(n7835), .A(n7037), .B(n7036), .ZN(P2_U3215) );
  OAI21_X1 U8656 ( .B1(n7040), .B2(n8030), .A(n7039), .ZN(n9982) );
  INV_X1 U8657 ( .A(n9982), .ZN(n7052) );
  OAI21_X1 U8658 ( .B1(n7042), .B2(n7041), .A(n10074), .ZN(n7044) );
  NOR2_X1 U8659 ( .A1(n7044), .A2(n7043), .ZN(n9971) );
  NAND2_X1 U8660 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  XOR2_X1 U8661 ( .A(n8030), .B(n7047), .Z(n7048) );
  OAI222_X1 U8662 ( .A1(n8491), .A2(n7050), .B1(n8434), .B2(n7049), .C1(n8486), 
        .C2(n7048), .ZN(n9972) );
  AOI211_X1 U8663 ( .C1(n10073), .C2(n9975), .A(n9971), .B(n9972), .ZN(n7051)
         );
  OAI21_X1 U8664 ( .B1(n10078), .B2(n7052), .A(n7051), .ZN(n7054) );
  NAND2_X1 U8665 ( .A1(n7054), .A2(n10097), .ZN(n7053) );
  OAI21_X1 U8666 ( .B1(n10097), .B2(n7138), .A(n7053), .ZN(P2_U3525) );
  NAND2_X1 U8667 ( .A1(n7054), .A2(n10083), .ZN(n7055) );
  OAI21_X1 U8668 ( .B1(n10083), .B2(n6098), .A(n7055), .ZN(P2_U3466) );
  NAND2_X1 U8669 ( .A1(n7057), .A2(n7056), .ZN(n7059) );
  XOR2_X1 U8670 ( .A(n7059), .B(n7058), .Z(n7065) );
  NAND2_X1 U8671 ( .A1(n8764), .A2(n7313), .ZN(n7062) );
  AOI21_X1 U8672 ( .B1(n8765), .B2(n9075), .A(n7060), .ZN(n7061) );
  OAI211_X1 U8673 ( .C1(n8868), .C2(n8768), .A(n7062), .B(n7061), .ZN(n7063)
         );
  AOI21_X1 U8674 ( .B1(n8882), .B2(n8770), .A(n7063), .ZN(n7064) );
  OAI21_X1 U8675 ( .B1(n7065), .B2(n8772), .A(n7064), .ZN(P1_U3237) );
  INV_X1 U8676 ( .A(n7066), .ZN(n7070) );
  AOI22_X1 U8677 ( .A1(n8033), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n8623), .ZN(n7067) );
  OAI21_X1 U8678 ( .B1(n7070), .B2(n6488), .A(n7067), .ZN(P2_U3338) );
  OAI222_X1 U8679 ( .A1(n7594), .A2(n7070), .B1(n7069), .B2(P1_U3084), .C1(
        n7068), .C2(n9595), .ZN(P1_U3333) );
  INV_X1 U8680 ( .A(n7071), .ZN(n7072) );
  AOI21_X1 U8681 ( .B1(n7073), .B2(n7072), .A(n7810), .ZN(n7076) );
  NOR3_X1 U8682 ( .A1(n7074), .A2(n7808), .A3(n7077), .ZN(n7075) );
  OAI21_X1 U8683 ( .B1(n7076), .B2(n7075), .A(n7364), .ZN(n7081) );
  OR2_X1 U8684 ( .A1(n7077), .A2(n8491), .ZN(n7078) );
  OAI21_X1 U8685 ( .B1(n7379), .B2(n8434), .A(n7078), .ZN(n7244) );
  OAI22_X1 U8686 ( .A1(n7828), .A2(n7250), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7190), .ZN(n7079) );
  AOI21_X1 U8687 ( .B1(n7819), .B2(n7244), .A(n7079), .ZN(n7080) );
  OAI211_X1 U8688 ( .C1(n10041), .C2(n7835), .A(n7081), .B(n7080), .ZN(
        P2_U3223) );
  XOR2_X1 U8689 ( .A(n7084), .B(n7083), .Z(n7085) );
  XNOR2_X1 U8690 ( .A(n7082), .B(n7085), .ZN(n7091) );
  INV_X1 U8691 ( .A(n9072), .ZN(n9838) );
  NAND2_X1 U8692 ( .A1(n8764), .A2(n7111), .ZN(n7088) );
  AOI21_X1 U8693 ( .B1(n8765), .B2(n9074), .A(n7086), .ZN(n7087) );
  OAI211_X1 U8694 ( .C1(n9838), .C2(n8768), .A(n7088), .B(n7087), .ZN(n7089)
         );
  AOI21_X1 U8695 ( .B1(n8872), .B2(n8770), .A(n7089), .ZN(n7090) );
  OAI21_X1 U8696 ( .B1(n7091), .B2(n8772), .A(n7090), .ZN(P1_U3211) );
  INV_X1 U8697 ( .A(n7607), .ZN(n7307) );
  AOI22_X1 U8698 ( .A1(n7890), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n8618), .ZN(n7092) );
  OAI21_X1 U8699 ( .B1(n7307), .B2(n6488), .A(n7092), .ZN(P2_U3337) );
  NAND2_X1 U8700 ( .A1(n7093), .A2(n8993), .ZN(n7095) );
  NAND2_X1 U8701 ( .A1(n9870), .A2(n9900), .ZN(n7094) );
  NAND2_X1 U8702 ( .A1(n7095), .A2(n7094), .ZN(n9854) );
  NAND2_X1 U8703 ( .A1(n7096), .A2(n9858), .ZN(n8876) );
  NAND2_X1 U8704 ( .A1(n9075), .A2(n9908), .ZN(n8873) );
  NAND2_X1 U8705 ( .A1(n9075), .A2(n9858), .ZN(n7097) );
  INV_X1 U8706 ( .A(n7309), .ZN(n7099) );
  NAND2_X1 U8707 ( .A1(n9868), .A2(n8882), .ZN(n8878) );
  INV_X1 U8708 ( .A(n8882), .ZN(n9913) );
  NAND2_X1 U8709 ( .A1(n9074), .A2(n9913), .ZN(n8863) );
  NAND2_X1 U8710 ( .A1(n7099), .A2(n7098), .ZN(n7308) );
  NAND2_X1 U8711 ( .A1(n9868), .A2(n9913), .ZN(n7100) );
  NAND2_X1 U8712 ( .A1(n7308), .A2(n7100), .ZN(n7255) );
  NAND2_X1 U8713 ( .A1(n8868), .A2(n8872), .ZN(n8877) );
  INV_X1 U8714 ( .A(n8872), .ZN(n9920) );
  NAND2_X1 U8715 ( .A1(n9073), .A2(n9920), .ZN(n8864) );
  NAND2_X1 U8716 ( .A1(n8877), .A2(n8864), .ZN(n8999) );
  XNOR2_X1 U8717 ( .A(n7255), .B(n8999), .ZN(n9923) );
  INV_X1 U8718 ( .A(n9923), .ZN(n7118) );
  INV_X1 U8719 ( .A(n7101), .ZN(n9873) );
  NAND2_X1 U8720 ( .A1(n9874), .A2(n9873), .ZN(n9477) );
  NAND2_X1 U8721 ( .A1(n8875), .A2(n9028), .ZN(n7102) );
  NAND2_X2 U8722 ( .A1(n7102), .A2(n9025), .ZN(n9864) );
  INV_X1 U8723 ( .A(n9864), .ZN(n7104) );
  NAND2_X1 U8724 ( .A1(n8878), .A2(n8876), .ZN(n9030) );
  INV_X1 U8725 ( .A(n9030), .ZN(n7103) );
  NAND2_X1 U8726 ( .A1(n8873), .A2(n8863), .ZN(n9000) );
  NAND2_X1 U8727 ( .A1(n9000), .A2(n8878), .ZN(n8806) );
  INV_X1 U8728 ( .A(n7258), .ZN(n7105) );
  AOI21_X1 U8729 ( .B1(n8999), .B2(n7106), .A(n7105), .ZN(n7107) );
  OAI222_X1 U8730 ( .A1(n9869), .A2(n9838), .B1(n9871), .B2(n9868), .C1(n9866), 
        .C2(n7107), .ZN(n9921) );
  NAND2_X1 U8731 ( .A1(n9857), .A2(n9908), .ZN(n9855) );
  INV_X1 U8732 ( .A(n7312), .ZN(n7109) );
  INV_X1 U8733 ( .A(n7265), .ZN(n7108) );
  OAI211_X1 U8734 ( .C1(n9920), .C2(n7109), .A(n7108), .B(n9856), .ZN(n9919)
         );
  AND2_X1 U8735 ( .A1(n7110), .A2(n9327), .ZN(n9433) );
  INV_X1 U8736 ( .A(n9433), .ZN(n9473) );
  INV_X1 U8737 ( .A(n7111), .ZN(n7112) );
  OAI22_X1 U8738 ( .A1(n9874), .A2(n7113), .B1(n7112), .B2(n9847), .ZN(n7114)
         );
  AOI21_X1 U8739 ( .B1(n9644), .B2(n8872), .A(n7114), .ZN(n7115) );
  OAI21_X1 U8740 ( .B1(n9919), .B2(n9473), .A(n7115), .ZN(n7116) );
  AOI21_X1 U8741 ( .B1(n9921), .B2(n9874), .A(n7116), .ZN(n7117) );
  OAI21_X1 U8742 ( .B1(n7118), .B2(n9477), .A(n7117), .ZN(P1_U3284) );
  AOI21_X1 U8743 ( .B1(n7120), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7119), .ZN(
        n9605) );
  NAND2_X1 U8744 ( .A1(n9607), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7121) );
  OAI21_X1 U8745 ( .B1(n9607), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7121), .ZN(
        n9604) );
  NOR2_X1 U8746 ( .A1(n9605), .A2(n9604), .ZN(n9603) );
  NAND2_X1 U8747 ( .A1(n7149), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7122) );
  OAI21_X1 U8748 ( .B1(n7149), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7122), .ZN(
        n7147) );
  NOR2_X1 U8749 ( .A1(n7148), .A2(n7147), .ZN(n7146) );
  NAND2_X1 U8750 ( .A1(n7226), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7123) );
  OAI21_X1 U8751 ( .B1(n7226), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7123), .ZN(
        n7224) );
  NAND2_X1 U8752 ( .A1(n7173), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7124) );
  OAI21_X1 U8753 ( .B1(n7173), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7124), .ZN(
        n7125) );
  AOI211_X1 U8754 ( .C1(n7126), .C2(n7125), .A(n7159), .B(n9602), .ZN(n7145)
         );
  INV_X1 U8755 ( .A(n7173), .ZN(n7143) );
  NOR2_X1 U8756 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6100), .ZN(n7127) );
  AOI21_X1 U8757 ( .B1(n9966), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7127), .ZN(
        n7142) );
  NAND2_X1 U8758 ( .A1(n7226), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7137) );
  MUX2_X1 U8759 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7128), .S(n7226), .Z(n7229)
         );
  NAND2_X1 U8760 ( .A1(n7149), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7136) );
  MUX2_X1 U8761 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7129), .S(n7149), .Z(n7152)
         );
  INV_X1 U8762 ( .A(n7130), .ZN(n7131) );
  OAI21_X1 U8763 ( .B1(n7133), .B2(n7132), .A(n7131), .ZN(n9611) );
  MUX2_X1 U8764 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7134), .S(n9607), .Z(n9610)
         );
  NAND2_X1 U8765 ( .A1(n9611), .A2(n9610), .ZN(n9609) );
  NAND2_X1 U8766 ( .A1(n9607), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U8767 ( .A1(n9609), .A2(n7135), .ZN(n7153) );
  NAND2_X1 U8768 ( .A1(n7152), .A2(n7153), .ZN(n7151) );
  NAND2_X1 U8769 ( .A1(n7136), .A2(n7151), .ZN(n7230) );
  NAND2_X1 U8770 ( .A1(n7229), .A2(n7230), .ZN(n7228) );
  NAND2_X1 U8771 ( .A1(n7137), .A2(n7228), .ZN(n7140) );
  MUX2_X1 U8772 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7138), .S(n7173), .Z(n7139)
         );
  NAND2_X1 U8773 ( .A1(n7139), .A2(n7140), .ZN(n7174) );
  OAI211_X1 U8774 ( .C1(n7140), .C2(n7139), .A(n9964), .B(n7174), .ZN(n7141)
         );
  OAI211_X1 U8775 ( .C1(n9961), .C2(n7143), .A(n7142), .B(n7141), .ZN(n7144)
         );
  OR2_X1 U8776 ( .A1(n7145), .A2(n7144), .ZN(P2_U3250) );
  AOI211_X1 U8777 ( .C1(n7148), .C2(n7147), .A(n7146), .B(n9602), .ZN(n7158)
         );
  INV_X1 U8778 ( .A(n7149), .ZN(n7156) );
  INV_X1 U8779 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10457) );
  NOR2_X1 U8780 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10457), .ZN(n7150) );
  AOI21_X1 U8781 ( .B1(n9966), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7150), .ZN(
        n7155) );
  OAI211_X1 U8782 ( .C1(n7153), .C2(n7152), .A(n9964), .B(n7151), .ZN(n7154)
         );
  OAI211_X1 U8783 ( .C1(n9961), .C2(n7156), .A(n7155), .B(n7154), .ZN(n7157)
         );
  OR2_X1 U8784 ( .A1(n7158), .A2(n7157), .ZN(P2_U3248) );
  MUX2_X1 U8785 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6998), .S(n7171), .Z(n7160)
         );
  INV_X1 U8786 ( .A(n7160), .ZN(n7200) );
  NOR2_X1 U8787 ( .A1(n4526), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U8788 ( .A1(n7213), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7161) );
  OAI21_X1 U8789 ( .B1(n7213), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7161), .ZN(
        n7211) );
  NOR2_X1 U8790 ( .A1(n7212), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U8791 ( .A1(n7189), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7162) );
  OAI21_X1 U8792 ( .B1(n7189), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7162), .ZN(
        n7187) );
  NAND2_X1 U8793 ( .A1(n8093), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7163) );
  OAI21_X1 U8794 ( .B1(n8093), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7163), .ZN(
        n8090) );
  NAND2_X1 U8795 ( .A1(n7280), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7164) );
  OAI21_X1 U8796 ( .B1(n7280), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7164), .ZN(
        n7165) );
  AOI211_X1 U8797 ( .C1(n7166), .C2(n7165), .A(n4516), .B(n9602), .ZN(n7185)
         );
  INV_X1 U8798 ( .A(n7280), .ZN(n7273) );
  NOR2_X1 U8799 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10470), .ZN(n7167) );
  AOI21_X1 U8800 ( .B1(n9966), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7167), .ZN(
        n7183) );
  INV_X1 U8801 ( .A(n8093), .ZN(n7178) );
  MUX2_X1 U8802 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7168), .S(n8093), .Z(n8096)
         );
  NAND2_X1 U8803 ( .A1(n7189), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7177) );
  MUX2_X1 U8804 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7169), .S(n7189), .Z(n7193)
         );
  NAND2_X1 U8805 ( .A1(n7213), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7176) );
  MUX2_X1 U8806 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7170), .S(n7213), .Z(n7216)
         );
  INV_X1 U8807 ( .A(n7171), .ZN(n7207) );
  MUX2_X1 U8808 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7172), .S(n7171), .Z(n7203)
         );
  NAND2_X1 U8809 ( .A1(n7173), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8810 ( .A1(n7175), .A2(n7174), .ZN(n7204) );
  NAND2_X1 U8811 ( .A1(n7203), .A2(n7204), .ZN(n7202) );
  OAI21_X1 U8812 ( .B1(n7207), .B2(n7172), .A(n7202), .ZN(n7217) );
  NAND2_X1 U8813 ( .A1(n7216), .A2(n7217), .ZN(n7215) );
  NAND2_X1 U8814 ( .A1(n7176), .A2(n7215), .ZN(n7194) );
  NAND2_X1 U8815 ( .A1(n7193), .A2(n7194), .ZN(n7192) );
  NAND2_X1 U8816 ( .A1(n7177), .A2(n7192), .ZN(n8097) );
  NAND2_X1 U8817 ( .A1(n8096), .A2(n8097), .ZN(n8095) );
  OAI21_X1 U8818 ( .B1(n7178), .B2(n7168), .A(n8095), .ZN(n7181) );
  INV_X1 U8819 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7179) );
  MUX2_X1 U8820 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7179), .S(n7280), .Z(n7180)
         );
  NAND2_X1 U8821 ( .A1(n7180), .A2(n7181), .ZN(n7272) );
  OAI211_X1 U8822 ( .C1(n7181), .C2(n7180), .A(n9964), .B(n7272), .ZN(n7182)
         );
  OAI211_X1 U8823 ( .C1(n9961), .C2(n7273), .A(n7183), .B(n7182), .ZN(n7184)
         );
  OR2_X1 U8824 ( .A1(n7185), .A2(n7184), .ZN(P2_U3255) );
  AOI211_X1 U8825 ( .C1(n7188), .C2(n7187), .A(n7186), .B(n9602), .ZN(n7198)
         );
  NOR2_X1 U8826 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7190), .ZN(n7191) );
  AOI21_X1 U8827 ( .B1(n9966), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7191), .ZN(
        n7196) );
  OAI211_X1 U8828 ( .C1(n7194), .C2(n7193), .A(n9964), .B(n7192), .ZN(n7195)
         );
  OAI211_X1 U8829 ( .C1(n9961), .C2(n4766), .A(n7196), .B(n7195), .ZN(n7197)
         );
  OR2_X1 U8830 ( .A1(n7198), .A2(n7197), .ZN(P2_U3253) );
  AOI211_X1 U8831 ( .C1(n4526), .C2(n7200), .A(n7199), .B(n9602), .ZN(n7209)
         );
  AOI21_X1 U8832 ( .B1(n9966), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7201), .ZN(
        n7206) );
  OAI211_X1 U8833 ( .C1(n7204), .C2(n7203), .A(n9964), .B(n7202), .ZN(n7205)
         );
  OAI211_X1 U8834 ( .C1(n9961), .C2(n7207), .A(n7206), .B(n7205), .ZN(n7208)
         );
  OR2_X1 U8835 ( .A1(n7209), .A2(n7208), .ZN(P2_U3251) );
  AOI211_X1 U8836 ( .C1(n7212), .C2(n7211), .A(n7210), .B(n9602), .ZN(n7222)
         );
  INV_X1 U8837 ( .A(n7213), .ZN(n7220) );
  NOR2_X1 U8838 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6137), .ZN(n7214) );
  AOI21_X1 U8839 ( .B1(n9966), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7214), .ZN(
        n7219) );
  OAI211_X1 U8840 ( .C1(n7217), .C2(n7216), .A(n9964), .B(n7215), .ZN(n7218)
         );
  OAI211_X1 U8841 ( .C1(n9961), .C2(n7220), .A(n7219), .B(n7218), .ZN(n7221)
         );
  OR2_X1 U8842 ( .A1(n7222), .A2(n7221), .ZN(P2_U3252) );
  AOI211_X1 U8843 ( .C1(n7225), .C2(n7224), .A(n7223), .B(n9602), .ZN(n7235)
         );
  INV_X1 U8844 ( .A(n7226), .ZN(n7233) );
  AOI21_X1 U8845 ( .B1(n9966), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7227), .ZN(
        n7232) );
  OAI211_X1 U8846 ( .C1(n7230), .C2(n7229), .A(n9964), .B(n7228), .ZN(n7231)
         );
  OAI211_X1 U8847 ( .C1(n9961), .C2(n7233), .A(n7232), .B(n7231), .ZN(n7234)
         );
  OR2_X1 U8848 ( .A1(n7235), .A2(n7234), .ZN(P2_U3249) );
  AND2_X1 U8849 ( .A1(n7236), .A2(n7924), .ZN(n7237) );
  OR2_X1 U8850 ( .A1(n7237), .A2(n7300), .ZN(n10042) );
  NOR2_X1 U8851 ( .A1(n8081), .A2(n10033), .ZN(n7238) );
  NAND2_X1 U8852 ( .A1(n7295), .A2(n10041), .ZN(n7923) );
  NAND2_X1 U8853 ( .A1(n8080), .A2(n7924), .ZN(n7922) );
  INV_X1 U8854 ( .A(n8041), .ZN(n7240) );
  XNOR2_X1 U8855 ( .A(n7298), .B(n7240), .ZN(n10040) );
  INV_X1 U8856 ( .A(n7241), .ZN(n10061) );
  NAND2_X1 U8857 ( .A1(n10040), .A2(n10061), .ZN(n7247) );
  XNOR2_X1 U8858 ( .A(n7293), .B(n8041), .ZN(n7245) );
  AOI21_X1 U8859 ( .B1(n7245), .B2(n10004), .A(n7244), .ZN(n7246) );
  NAND2_X1 U8860 ( .A1(n7247), .A2(n7246), .ZN(n10045) );
  INV_X1 U8861 ( .A(n10040), .ZN(n7248) );
  NOR2_X1 U8862 ( .A1(n7248), .A2(n8449), .ZN(n7249) );
  OAI21_X1 U8863 ( .B1(n10045), .B2(n7249), .A(n9993), .ZN(n7253) );
  OAI22_X1 U8864 ( .A1(n9993), .A2(n4765), .B1(n7250), .B2(n8451), .ZN(n7251)
         );
  AOI21_X1 U8865 ( .B1(n8455), .B2(n7924), .A(n7251), .ZN(n7252) );
  OAI211_X1 U8866 ( .C1(n9989), .C2(n10042), .A(n7253), .B(n7252), .ZN(
        P2_U3288) );
  NOR2_X1 U8867 ( .A1(n9073), .A2(n8872), .ZN(n7254) );
  NAND2_X1 U8868 ( .A1(n9838), .A2(n7440), .ZN(n8895) );
  NAND2_X1 U8869 ( .A1(n9072), .A2(n9927), .ZN(n8809) );
  NAND2_X1 U8870 ( .A1(n8895), .A2(n8809), .ZN(n7259) );
  NAND2_X1 U8871 ( .A1(n7256), .A2(n7259), .ZN(n7442) );
  OR2_X1 U8872 ( .A1(n7256), .A2(n7259), .ZN(n7257) );
  NAND2_X1 U8873 ( .A1(n7442), .A2(n7257), .ZN(n7263) );
  NAND2_X1 U8874 ( .A1(n7258), .A2(n8877), .ZN(n7438) );
  INV_X1 U8875 ( .A(n7259), .ZN(n8890) );
  XNOR2_X1 U8876 ( .A(n7438), .B(n8890), .ZN(n7261) );
  INV_X1 U8877 ( .A(n9071), .ZN(n7443) );
  OAI22_X1 U8878 ( .A1(n8868), .A2(n9871), .B1(n7443), .B2(n9869), .ZN(n7260)
         );
  AOI21_X1 U8879 ( .B1(n7261), .B2(n9840), .A(n7260), .ZN(n7262) );
  OAI21_X1 U8880 ( .B1(n7263), .B2(n9843), .A(n7262), .ZN(n9928) );
  INV_X1 U8881 ( .A(n9928), .ZN(n7270) );
  INV_X1 U8882 ( .A(n7263), .ZN(n9930) );
  AND2_X2 U8883 ( .A1(n7265), .A2(n9927), .ZN(n9831) );
  INV_X1 U8884 ( .A(n9831), .ZN(n7264) );
  OAI211_X1 U8885 ( .C1(n9927), .C2(n7265), .A(n7264), .B(n9856), .ZN(n9926)
         );
  AOI22_X1 U8886 ( .A1(n9640), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7339), .B2(
        n9861), .ZN(n7267) );
  NAND2_X1 U8887 ( .A1(n9644), .A2(n7440), .ZN(n7266) );
  OAI211_X1 U8888 ( .C1(n9926), .C2(n9376), .A(n7267), .B(n7266), .ZN(n7268)
         );
  AOI21_X1 U8889 ( .B1(n9930), .B2(n9834), .A(n7268), .ZN(n7269) );
  OAI21_X1 U8890 ( .B1(n7270), .B2(n9640), .A(n7269), .ZN(P1_U3283) );
  INV_X1 U8891 ( .A(n7333), .ZN(n7276) );
  INV_X1 U8892 ( .A(n8106), .ZN(n7274) );
  MUX2_X1 U8893 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7271), .S(n8106), .Z(n8108)
         );
  OAI21_X1 U8894 ( .B1(n7273), .B2(n7179), .A(n7272), .ZN(n8109) );
  NAND2_X1 U8895 ( .A1(n8108), .A2(n8109), .ZN(n8107) );
  OAI21_X1 U8896 ( .B1(n7274), .B2(n7271), .A(n8107), .ZN(n7325) );
  MUX2_X1 U8897 ( .A(n7275), .B(P2_REG1_REG_12__SCAN_IN), .S(n7333), .Z(n7324)
         );
  NOR2_X1 U8898 ( .A1(n7325), .A2(n7324), .ZN(n7323) );
  AOI21_X1 U8899 ( .B1(n7276), .B2(n7275), .A(n7323), .ZN(n7278) );
  INV_X1 U8900 ( .A(n7353), .ZN(n7349) );
  AOI22_X1 U8901 ( .A1(n7353), .A2(n6257), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7349), .ZN(n7277) );
  NOR2_X1 U8902 ( .A1(n7278), .A2(n7277), .ZN(n7348) );
  AOI21_X1 U8903 ( .B1(n7278), .B2(n7277), .A(n7348), .ZN(n7291) );
  NAND2_X1 U8904 ( .A1(n7333), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U8905 ( .B1(n7333), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7279), .ZN(
        n7329) );
  MUX2_X1 U8906 ( .A(n7401), .B(P2_REG2_REG_11__SCAN_IN), .S(n8106), .Z(n7281)
         );
  INV_X1 U8907 ( .A(n7281), .ZN(n8103) );
  NAND2_X1 U8908 ( .A1(n8102), .A2(n8103), .ZN(n8101) );
  OAI21_X1 U8909 ( .B1(n8106), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8101), .ZN(
        n7330) );
  NOR2_X1 U8910 ( .A1(n7353), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7282) );
  AOI21_X1 U8911 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7353), .A(n7282), .ZN(
        n7283) );
  OAI21_X1 U8912 ( .B1(n7284), .B2(n7283), .A(n7352), .ZN(n7285) );
  NAND2_X1 U8913 ( .A1(n7285), .A2(n9965), .ZN(n7290) );
  INV_X1 U8914 ( .A(n9961), .ZN(n9608) );
  INV_X1 U8915 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7287) );
  OAI22_X1 U8916 ( .A1(n8181), .A2(n7287), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7286), .ZN(n7288) );
  AOI21_X1 U8917 ( .B1(n9608), .B2(n7353), .A(n7288), .ZN(n7289) );
  OAI211_X1 U8918 ( .C1(n7291), .C2(n9962), .A(n7290), .B(n7289), .ZN(P2_U3258) );
  NAND2_X1 U8919 ( .A1(n7295), .A2(n7924), .ZN(n7292) );
  NAND2_X1 U8920 ( .A1(n7379), .A2(n10047), .ZN(n7926) );
  INV_X1 U8921 ( .A(n10047), .ZN(n7370) );
  NAND2_X1 U8922 ( .A1(n8079), .A2(n7370), .ZN(n7928) );
  NAND2_X1 U8923 ( .A1(n7926), .A2(n7928), .ZN(n8039) );
  INV_X1 U8924 ( .A(n8039), .ZN(n7921) );
  XNOR2_X1 U8925 ( .A(n7377), .B(n7921), .ZN(n7296) );
  NAND2_X1 U8926 ( .A1(n8078), .A2(n8471), .ZN(n7294) );
  OAI21_X1 U8927 ( .B1(n7295), .B2(n8491), .A(n7294), .ZN(n7365) );
  AOI21_X1 U8928 ( .B1(n7296), .B2(n10004), .A(n7365), .ZN(n10049) );
  INV_X1 U8929 ( .A(n7922), .ZN(n7297) );
  NAND2_X1 U8930 ( .A1(n7299), .A2(n8039), .ZN(n7382) );
  OAI21_X1 U8931 ( .B1(n7299), .B2(n8039), .A(n7382), .ZN(n10052) );
  NAND2_X1 U8932 ( .A1(n10052), .A2(n8329), .ZN(n7306) );
  INV_X1 U8933 ( .A(n7300), .ZN(n7301) );
  AOI211_X1 U8934 ( .C1(n10047), .C2(n7301), .A(n10065), .B(n7384), .ZN(n10046) );
  NOR2_X1 U8935 ( .A1(n9988), .A2(n7370), .ZN(n7304) );
  INV_X1 U8936 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7302) );
  OAI22_X1 U8937 ( .A1(n9993), .A2(n7302), .B1(n7366), .B2(n8451), .ZN(n7303)
         );
  AOI211_X1 U8938 ( .C1(n10046), .C2(n8427), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI211_X1 U8939 ( .C1(n8289), .C2(n10049), .A(n7306), .B(n7305), .ZN(
        P2_U3287) );
  INV_X1 U8940 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10490) );
  OAI222_X1 U8941 ( .A1(n7594), .A2(n7307), .B1(n9023), .B2(P1_U3084), .C1(
        n10490), .C2(n9595), .ZN(P1_U3332) );
  NAND2_X1 U8942 ( .A1(n7309), .A2(n7315), .ZN(n7310) );
  NAND2_X1 U8943 ( .A1(n7308), .A2(n7310), .ZN(n9917) );
  NAND2_X1 U8944 ( .A1(n9855), .A2(n8882), .ZN(n7311) );
  NAND2_X1 U8945 ( .A1(n7312), .A2(n7311), .ZN(n9914) );
  AOI22_X1 U8946 ( .A1(n9644), .A2(n8882), .B1(n7313), .B2(n9861), .ZN(n7314)
         );
  OAI21_X1 U8947 ( .B1(n9914), .B2(n9455), .A(n7314), .ZN(n7321) );
  INV_X1 U8948 ( .A(n8876), .ZN(n8866) );
  AOI21_X1 U8949 ( .B1(n9864), .B2(n9865), .A(n8866), .ZN(n7316) );
  XNOR2_X1 U8950 ( .A(n7316), .B(n7315), .ZN(n7319) );
  NAND2_X1 U8951 ( .A1(n9917), .A2(n9639), .ZN(n7318) );
  AOI22_X1 U8952 ( .A1(n9635), .A2(n9073), .B1(n9075), .B2(n9632), .ZN(n7317)
         );
  OAI211_X1 U8953 ( .C1(n7319), .C2(n9866), .A(n7318), .B(n7317), .ZN(n9915)
         );
  MUX2_X1 U8954 ( .A(n9915), .B(P1_REG2_REG_6__SCAN_IN), .S(n9640), .Z(n7320)
         );
  AOI211_X1 U8955 ( .C1(n9834), .C2(n9917), .A(n7321), .B(n7320), .ZN(n7322)
         );
  INV_X1 U8956 ( .A(n7322), .ZN(P1_U3285) );
  AOI21_X1 U8957 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n7327) );
  NOR2_X1 U8958 ( .A1(n10485), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7549) );
  AOI21_X1 U8959 ( .B1(n9966), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7549), .ZN(
        n7326) );
  OAI21_X1 U8960 ( .B1(n7327), .B2(n9962), .A(n7326), .ZN(n7332) );
  AOI211_X1 U8961 ( .C1(n7330), .C2(n7329), .A(n7328), .B(n9602), .ZN(n7331)
         );
  AOI211_X1 U8962 ( .C1(n9608), .C2(n7333), .A(n7332), .B(n7331), .ZN(n7334)
         );
  INV_X1 U8963 ( .A(n7334), .ZN(P2_U3257) );
  XNOR2_X1 U8964 ( .A(n7337), .B(n7336), .ZN(n7338) );
  XNOR2_X1 U8965 ( .A(n7335), .B(n7338), .ZN(n7345) );
  NAND2_X1 U8966 ( .A1(n8764), .A2(n7339), .ZN(n7342) );
  NOR2_X1 U8967 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7340), .ZN(n9724) );
  AOI21_X1 U8968 ( .B1(n8757), .B2(n9071), .A(n9724), .ZN(n7341) );
  OAI211_X1 U8969 ( .C1(n8868), .C2(n8755), .A(n7342), .B(n7341), .ZN(n7343)
         );
  AOI21_X1 U8970 ( .B1(n7440), .B2(n8770), .A(n7343), .ZN(n7344) );
  OAI21_X1 U8971 ( .B1(n7345), .B2(n8772), .A(n7344), .ZN(P1_U3219) );
  INV_X1 U8972 ( .A(n7614), .ZN(n7347) );
  AOI22_X1 U8973 ( .A1(n8069), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8623), .ZN(n7346) );
  OAI21_X1 U8974 ( .B1(n7347), .B2(n6488), .A(n7346), .ZN(P2_U3336) );
  OAI222_X1 U8975 ( .A1(n8982), .A2(P1_U3084), .B1(n7594), .B2(n7347), .C1(
        n9595), .C2(n5744), .ZN(P1_U3331) );
  AOI21_X1 U8976 ( .B1(n7349), .B2(n6257), .A(n7348), .ZN(n7351) );
  INV_X1 U8977 ( .A(n7492), .ZN(n7496) );
  AOI22_X1 U8978 ( .A1(n7492), .A2(n7495), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7496), .ZN(n7350) );
  NOR2_X1 U8979 ( .A1(n7351), .A2(n7350), .ZN(n7494) );
  AOI21_X1 U8980 ( .B1(n7351), .B2(n7350), .A(n7494), .ZN(n7361) );
  AOI22_X1 U8981 ( .A1(n7492), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6270), .B2(
        n7496), .ZN(n7355) );
  NAND2_X1 U8982 ( .A1(n7355), .A2(n7354), .ZN(n7491) );
  OAI21_X1 U8983 ( .B1(n7355), .B2(n7354), .A(n7491), .ZN(n7356) );
  NAND2_X1 U8984 ( .A1(n7356), .A2(n9965), .ZN(n7360) );
  INV_X1 U8985 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8986 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7695) );
  OAI21_X1 U8987 ( .B1(n8181), .B2(n7357), .A(n7695), .ZN(n7358) );
  AOI21_X1 U8988 ( .B1(n9608), .B2(n7492), .A(n7358), .ZN(n7359) );
  OAI211_X1 U8989 ( .C1(n7361), .C2(n9962), .A(n7360), .B(n7359), .ZN(P2_U3259) );
  NAND3_X1 U8990 ( .A1(n7822), .A2(n8080), .A3(n7362), .ZN(n7363) );
  OAI21_X1 U8991 ( .B1(n7364), .B2(n7810), .A(n7363), .ZN(n7374) );
  NAND2_X1 U8992 ( .A1(n7365), .A2(n7819), .ZN(n7369) );
  INV_X1 U8993 ( .A(n7366), .ZN(n7367) );
  AOI22_X1 U8994 ( .A1(n7805), .A2(n7367), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n7368) );
  OAI211_X1 U8995 ( .C1(n7370), .C2(n7835), .A(n7369), .B(n7368), .ZN(n7373)
         );
  NOR2_X1 U8996 ( .A1(n7371), .A2(n7810), .ZN(n7372) );
  AOI211_X1 U8997 ( .C1(n7375), .C2(n7374), .A(n7373), .B(n7372), .ZN(n7376)
         );
  INV_X1 U8998 ( .A(n7376), .ZN(P2_U3233) );
  NAND2_X1 U8999 ( .A1(n7377), .A2(n7921), .ZN(n7378) );
  NAND2_X1 U9000 ( .A1(n7378), .A2(n7926), .ZN(n7398) );
  NAND2_X1 U9001 ( .A1(n10055), .A2(n8078), .ZN(n7929) );
  INV_X1 U9002 ( .A(n10055), .ZN(n7388) );
  NAND2_X1 U9003 ( .A1(n7388), .A2(n7463), .ZN(n7931) );
  XNOR2_X1 U9004 ( .A(n7398), .B(n8043), .ZN(n7381) );
  OR2_X1 U9005 ( .A1(n7379), .A2(n8491), .ZN(n7380) );
  OAI21_X1 U9006 ( .B1(n7548), .B2(n8434), .A(n7380), .ZN(n7409) );
  AOI21_X1 U9007 ( .B1(n7381), .B2(n10004), .A(n7409), .ZN(n10054) );
  OAI21_X1 U9008 ( .B1(n10047), .B2(n8079), .A(n7382), .ZN(n7395) );
  XOR2_X1 U9009 ( .A(n8043), .B(n7395), .Z(n10060) );
  NAND2_X1 U9010 ( .A1(n10060), .A2(n8329), .ZN(n7390) );
  OAI22_X1 U9011 ( .A1(n9993), .A2(n7383), .B1(n7410), .B2(n8451), .ZN(n7387)
         );
  NAND2_X1 U9012 ( .A1(n7384), .A2(n10055), .ZN(n7484) );
  OAI211_X1 U9013 ( .C1(n7384), .C2(n10055), .A(n10074), .B(n7484), .ZN(n10053) );
  NOR2_X1 U9014 ( .A1(n10053), .A2(n7385), .ZN(n7386) );
  AOI211_X1 U9015 ( .C1(n8455), .C2(n7388), .A(n7387), .B(n7386), .ZN(n7389)
         );
  OAI211_X1 U9016 ( .C1(n8496), .C2(n10054), .A(n7390), .B(n7389), .ZN(
        P2_U3286) );
  INV_X1 U9017 ( .A(n7621), .ZN(n7394) );
  AOI21_X1 U9018 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8618), .A(n8065), .ZN(
        n7391) );
  OAI21_X1 U9019 ( .B1(n7394), .B2(n6488), .A(n7391), .ZN(P2_U3335) );
  NOR2_X1 U9020 ( .A1(n7392), .A2(P1_U3084), .ZN(n9061) );
  AOI21_X1 U9021 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9597), .A(n9061), .ZN(
        n7393) );
  OAI21_X1 U9022 ( .B1(n7394), .B2(n9599), .A(n7393), .ZN(P1_U3330) );
  NAND2_X1 U9023 ( .A1(n7483), .A2(n7548), .ZN(n7938) );
  NAND2_X1 U9024 ( .A1(n7935), .A2(n7938), .ZN(n7399) );
  OAI21_X1 U9025 ( .B1(n7396), .B2(n7399), .A(n7474), .ZN(n10062) );
  INV_X1 U9026 ( .A(n7931), .ZN(n7397) );
  AOI21_X2 U9027 ( .B1(n7398), .B2(n7929), .A(n7397), .ZN(n7478) );
  INV_X1 U9028 ( .A(n7399), .ZN(n8044) );
  XNOR2_X1 U9029 ( .A(n7478), .B(n8044), .ZN(n7400) );
  OAI222_X1 U9030 ( .A1(n8434), .A2(n8075), .B1(n8491), .B2(n7463), .C1(n7400), 
        .C2(n8486), .ZN(n10068) );
  XNOR2_X1 U9031 ( .A(n7484), .B(n7483), .ZN(n10066) );
  OAI22_X1 U9032 ( .A1(n9993), .A2(n7401), .B1(n7467), .B2(n8451), .ZN(n7402)
         );
  AOI21_X1 U9033 ( .B1(n7483), .B2(n8455), .A(n7402), .ZN(n7403) );
  OAI21_X1 U9034 ( .B1(n10066), .B2(n9989), .A(n7403), .ZN(n7404) );
  AOI21_X1 U9035 ( .B1(n10068), .B2(n9993), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9036 ( .B1(n10062), .B2(n8501), .A(n7405), .ZN(P2_U3285) );
  INV_X1 U9037 ( .A(n7462), .ZN(n7406) );
  AOI211_X1 U9038 ( .C1(n7408), .C2(n7407), .A(n7810), .B(n7406), .ZN(n7415)
         );
  NAND2_X1 U9039 ( .A1(n7409), .A2(n7819), .ZN(n7413) );
  INV_X1 U9040 ( .A(n7410), .ZN(n7411) );
  AOI22_X1 U9041 ( .A1(n7805), .A2(n7411), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7412) );
  OAI211_X1 U9042 ( .C1(n10055), .C2(n7835), .A(n7413), .B(n7412), .ZN(n7414)
         );
  OR2_X1 U9043 ( .A1(n7415), .A2(n7414), .ZN(P2_U3219) );
  INV_X1 U9044 ( .A(n7416), .ZN(n7417) );
  AOI21_X1 U9045 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n7426) );
  INV_X1 U9046 ( .A(n9933), .ZN(n7445) );
  NAND2_X1 U9047 ( .A1(n8764), .A2(n9846), .ZN(n7423) );
  INV_X1 U9048 ( .A(n7420), .ZN(n7421) );
  AOI21_X1 U9049 ( .B1(n8757), .B2(n9633), .A(n7421), .ZN(n7422) );
  OAI211_X1 U9050 ( .C1(n9838), .C2(n8755), .A(n7423), .B(n7422), .ZN(n7424)
         );
  AOI21_X1 U9051 ( .B1(n7445), .B2(n8770), .A(n7424), .ZN(n7425) );
  OAI21_X1 U9052 ( .B1(n7426), .B2(n8772), .A(n7425), .ZN(P1_U3229) );
  NAND2_X1 U9053 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  XNOR2_X1 U9054 ( .A(n7430), .B(n7429), .ZN(n7437) );
  NAND2_X1 U9055 ( .A1(n8764), .A2(n7449), .ZN(n7434) );
  INV_X1 U9056 ( .A(n7431), .ZN(n7432) );
  AOI21_X1 U9057 ( .B1(n8757), .B2(n9462), .A(n7432), .ZN(n7433) );
  OAI211_X1 U9058 ( .C1(n7443), .C2(n8755), .A(n7434), .B(n7433), .ZN(n7435)
         );
  AOI21_X1 U9059 ( .B1(n9140), .B2(n8770), .A(n7435), .ZN(n7436) );
  OAI21_X1 U9060 ( .B1(n7437), .B2(n8772), .A(n7436), .ZN(P1_U3215) );
  AND2_X1 U9061 ( .A1(n9933), .A2(n9071), .ZN(n8894) );
  NAND2_X1 U9062 ( .A1(n7443), .A2(n7445), .ZN(n8896) );
  INV_X1 U9063 ( .A(n9633), .ZN(n9837) );
  XNOR2_X1 U9064 ( .A(n9173), .B(n4494), .ZN(n7439) );
  AOI222_X1 U9065 ( .A1(n9840), .A2(n7439), .B1(n9462), .B2(n9635), .C1(n9071), 
        .C2(n9632), .ZN(n7507) );
  NAND2_X1 U9066 ( .A1(n9072), .A2(n7440), .ZN(n7441) );
  NAND2_X1 U9067 ( .A1(n7442), .A2(n7441), .ZN(n9829) );
  NAND2_X1 U9068 ( .A1(n9933), .A2(n7443), .ZN(n7444) );
  NAND2_X1 U9069 ( .A1(n7445), .A2(n9071), .ZN(n7446) );
  INV_X1 U9070 ( .A(n9142), .ZN(n7448) );
  AOI21_X1 U9071 ( .B1(n4494), .B2(n7447), .A(n7448), .ZN(n7508) );
  INV_X1 U9072 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7451) );
  INV_X1 U9073 ( .A(n7449), .ZN(n7450) );
  OAI22_X1 U9074 ( .A1(n9874), .A2(n7451), .B1(n7450), .B2(n9847), .ZN(n7452)
         );
  AOI21_X1 U9075 ( .B1(n9644), .B2(n9140), .A(n7452), .ZN(n7455) );
  AOI21_X1 U9076 ( .B1(n9830), .B2(n9140), .A(n9934), .ZN(n7453) );
  AND2_X1 U9077 ( .A1(n7453), .A2(n9625), .ZN(n7505) );
  NAND2_X1 U9078 ( .A1(n7505), .A2(n9433), .ZN(n7454) );
  OAI211_X1 U9079 ( .C1(n7508), .C2(n9477), .A(n7455), .B(n7454), .ZN(n7456)
         );
  INV_X1 U9080 ( .A(n7456), .ZN(n7457) );
  OAI21_X1 U9081 ( .B1(n9640), .B2(n7507), .A(n7457), .ZN(P1_U3281) );
  INV_X1 U9082 ( .A(n7598), .ZN(n7473) );
  AOI22_X1 U9083 ( .A1(n7458), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n8618), .ZN(n7459) );
  OAI21_X1 U9084 ( .B1(n7473), .B2(n6488), .A(n7459), .ZN(P2_U3334) );
  INV_X1 U9085 ( .A(n7483), .ZN(n10064) );
  INV_X1 U9086 ( .A(n7460), .ZN(n7461) );
  AOI21_X1 U9087 ( .B1(n7462), .B2(n7461), .A(n7810), .ZN(n7466) );
  NOR3_X1 U9088 ( .A1(n7464), .A2(n7463), .A3(n7808), .ZN(n7465) );
  OAI21_X1 U9089 ( .B1(n7466), .B2(n7465), .A(n7544), .ZN(n7471) );
  NOR2_X1 U9090 ( .A1(n7829), .A2(n8075), .ZN(n7469) );
  OAI22_X1 U9091 ( .A1(n7828), .A2(n7467), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6219), .ZN(n7468) );
  AOI211_X1 U9092 ( .C1(n7745), .C2(n8078), .A(n7469), .B(n7468), .ZN(n7470)
         );
  OAI211_X1 U9093 ( .C1(n10064), .C2(n7835), .A(n7471), .B(n7470), .ZN(
        P2_U3238) );
  OAI222_X1 U9094 ( .A1(n7594), .A2(n7473), .B1(P1_U3084), .B2(n7472), .C1(
        n10294), .C2(n9595), .ZN(P1_U3329) );
  NAND2_X1 U9095 ( .A1(n10072), .A2(n8075), .ZN(n7936) );
  AOI21_X1 U9096 ( .B1(n8045), .B2(n7476), .A(n4590), .ZN(n10079) );
  INV_X1 U9097 ( .A(n7935), .ZN(n7477) );
  XNOR2_X1 U9098 ( .A(n4510), .B(n8045), .ZN(n7480) );
  OAI22_X1 U9099 ( .A1(n7548), .A2(n8491), .B1(n8492), .B2(n8434), .ZN(n7479)
         );
  AOI21_X1 U9100 ( .B1(n7480), .B2(n10004), .A(n7479), .ZN(n10077) );
  OAI22_X1 U9101 ( .A1(n9993), .A2(n7481), .B1(n7552), .B2(n8451), .ZN(n7482)
         );
  AOI21_X1 U9102 ( .B1(n10072), .B2(n8455), .A(n7482), .ZN(n7488) );
  AND2_X1 U9103 ( .A1(n7485), .A2(n10072), .ZN(n7486) );
  NOR2_X1 U9104 ( .A1(n7537), .A2(n7486), .ZN(n10075) );
  NAND2_X1 U9105 ( .A1(n10075), .A2(n8499), .ZN(n7487) );
  OAI211_X1 U9106 ( .C1(n10077), .C2(n8496), .A(n7488), .B(n7487), .ZN(n7489)
         );
  INV_X1 U9107 ( .A(n7489), .ZN(n7490) );
  OAI21_X1 U9108 ( .B1(n10079), .B2(n8501), .A(n7490), .ZN(P2_U3284) );
  OAI21_X1 U9109 ( .B1(n7492), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7491), .ZN(
        n8114) );
  XNOR2_X1 U9110 ( .A(n8114), .B(n8122), .ZN(n7493) );
  NAND2_X1 U9111 ( .A1(n7493), .A2(n6299), .ZN(n8116) );
  OAI21_X1 U9112 ( .B1(n7493), .B2(n6299), .A(n8116), .ZN(n7502) );
  INV_X1 U9113 ( .A(n8122), .ZN(n8115) );
  AOI21_X1 U9114 ( .B1(n7496), .B2(n7495), .A(n7494), .ZN(n8121) );
  XNOR2_X1 U9115 ( .A(n8121), .B(n8115), .ZN(n7497) );
  NAND2_X1 U9116 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7497), .ZN(n8123) );
  OAI211_X1 U9117 ( .C1(n7497), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9964), .B(
        n8123), .ZN(n7500) );
  AND2_X1 U9118 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7498) );
  AOI21_X1 U9119 ( .B1(n9966), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7498), .ZN(
        n7499) );
  OAI211_X1 U9120 ( .C1(n9961), .C2(n8115), .A(n7500), .B(n7499), .ZN(n7501)
         );
  AOI21_X1 U9121 ( .B1(n9965), .B2(n7502), .A(n7501), .ZN(n7503) );
  INV_X1 U9122 ( .A(n7503), .ZN(P2_U3260) );
  INV_X1 U9123 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7510) );
  AOI21_X1 U9124 ( .B1(n9647), .B2(n9140), .A(n7505), .ZN(n7506) );
  OAI211_X1 U9125 ( .C1(n7508), .C2(n9660), .A(n7507), .B(n7506), .ZN(n7511)
         );
  NAND2_X1 U9126 ( .A1(n7511), .A2(n9906), .ZN(n7509) );
  OAI21_X1 U9127 ( .B1(n9906), .B2(n7510), .A(n7509), .ZN(P1_U3484) );
  NAND2_X1 U9128 ( .A1(n7511), .A2(n9948), .ZN(n7512) );
  OAI21_X1 U9129 ( .B1(n9948), .B2(n7513), .A(n7512), .ZN(P1_U3533) );
  AOI21_X1 U9130 ( .B1(n4724), .B2(n7514), .A(n8772), .ZN(n7516) );
  NAND2_X1 U9131 ( .A1(n7516), .A2(n7515), .ZN(n7520) );
  AND2_X1 U9132 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9084) );
  AOI21_X1 U9133 ( .B1(n8765), .B2(n9633), .A(n9084), .ZN(n7517) );
  OAI21_X1 U9134 ( .B1(n9448), .B2(n8768), .A(n7517), .ZN(n7518) );
  AOI21_X1 U9135 ( .B1(n9628), .B2(n8764), .A(n7518), .ZN(n7519) );
  OAI211_X1 U9136 ( .C1(n9668), .C2(n8760), .A(n7520), .B(n7519), .ZN(P1_U3234) );
  OAI211_X1 U9137 ( .C1(n7521), .C2(n4592), .A(n7690), .B(n7823), .ZN(n7525)
         );
  OAI22_X1 U9138 ( .A1(n7828), .A2(n7534), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7286), .ZN(n7523) );
  OAI22_X1 U9139 ( .A1(n7830), .A2(n8075), .B1(n8073), .B2(n7829), .ZN(n7522)
         );
  AOI211_X1 U9140 ( .C1(n7540), .C2(n7793), .A(n7523), .B(n7522), .ZN(n7524)
         );
  NAND2_X1 U9141 ( .A1(n7525), .A2(n7524), .ZN(P2_U3236) );
  INV_X1 U9142 ( .A(n7631), .ZN(n7562) );
  AOI22_X1 U9143 ( .A1(n7526), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8618), .ZN(n7527) );
  OAI21_X1 U9144 ( .B1(n7562), .B2(n6488), .A(n7527), .ZN(P2_U3333) );
  INV_X1 U9145 ( .A(n7936), .ZN(n7940) );
  OR2_X1 U9146 ( .A1(n7540), .A2(n8492), .ZN(n7946) );
  NAND2_X1 U9147 ( .A1(n7540), .A2(n8492), .ZN(n7945) );
  AOI21_X1 U9148 ( .B1(n7528), .B2(n8047), .A(n4572), .ZN(n7529) );
  OAI222_X1 U9149 ( .A1(n8434), .A2(n8073), .B1(n8491), .B2(n8075), .C1(n8486), 
        .C2(n7529), .ZN(n9619) );
  INV_X1 U9150 ( .A(n9619), .ZN(n7543) );
  INV_X1 U9151 ( .A(n10072), .ZN(n7530) );
  NAND2_X1 U9152 ( .A1(n7530), .A2(n8075), .ZN(n7531) );
  NOR2_X1 U9153 ( .A1(n7532), .A2(n8047), .ZN(n9615) );
  INV_X1 U9154 ( .A(n9615), .ZN(n7533) );
  NAND3_X1 U9155 ( .A1(n7533), .A2(n8329), .A3(n8194), .ZN(n7542) );
  OAI22_X1 U9156 ( .A1(n9993), .A2(n7535), .B1(n7534), .B2(n8451), .ZN(n7539)
         );
  AND2_X2 U9157 ( .A1(n7537), .A2(n9616), .ZN(n8481) );
  INV_X1 U9158 ( .A(n8481), .ZN(n7536) );
  OAI21_X1 U9159 ( .B1(n9616), .B2(n7537), .A(n7536), .ZN(n9617) );
  NOR2_X1 U9160 ( .A1(n9617), .A2(n9989), .ZN(n7538) );
  AOI211_X1 U9161 ( .C1(n8455), .C2(n7540), .A(n7539), .B(n7538), .ZN(n7541)
         );
  OAI211_X1 U9162 ( .C1(n8289), .C2(n7543), .A(n7542), .B(n7541), .ZN(P2_U3283) );
  INV_X1 U9163 ( .A(n7544), .ZN(n7547) );
  NOR3_X1 U9164 ( .A1(n7545), .A2(n7548), .A3(n7808), .ZN(n7546) );
  AOI21_X1 U9165 ( .B1(n7547), .B2(n7823), .A(n7546), .ZN(n7558) );
  INV_X1 U9166 ( .A(n7548), .ZN(n8077) );
  INV_X1 U9167 ( .A(n8492), .ZN(n8074) );
  AOI22_X1 U9168 ( .A1(n7745), .A2(n8077), .B1(n7694), .B2(n8074), .ZN(n7551)
         );
  INV_X1 U9169 ( .A(n7549), .ZN(n7550) );
  OAI211_X1 U9170 ( .C1(n7552), .C2(n7828), .A(n7551), .B(n7550), .ZN(n7555)
         );
  NOR2_X1 U9171 ( .A1(n7553), .A2(n7810), .ZN(n7554) );
  AOI211_X1 U9172 ( .C1(n10072), .C2(n7793), .A(n7555), .B(n7554), .ZN(n7556)
         );
  OAI21_X1 U9173 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(P2_U3226) );
  INV_X1 U9174 ( .A(n7643), .ZN(n7566) );
  AOI22_X1 U9175 ( .A1(n7559), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8618), .ZN(n7560) );
  OAI21_X1 U9176 ( .B1(n7566), .B2(n6488), .A(n7560), .ZN(P2_U3332) );
  OAI222_X1 U9177 ( .A1(n9595), .A2(n7563), .B1(n7594), .B2(n7562), .C1(n7561), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9178 ( .A1(n9599), .A2(n7566), .B1(P1_U3084), .B2(n7565), .C1(
        n7564), .C2(n9595), .ZN(P1_U3327) );
  INV_X1 U9179 ( .A(n7595), .ZN(n7571) );
  INV_X1 U9180 ( .A(n7567), .ZN(n8185) );
  AOI22_X1 U9181 ( .A1(n8185), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8618), .ZN(n7568) );
  OAI21_X1 U9182 ( .B1(n7571), .B2(n6488), .A(n7568), .ZN(P2_U3331) );
  AOI21_X1 U9183 ( .B1(n9597), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7569), .ZN(
        n7570) );
  OAI21_X1 U9184 ( .B1(n7571), .B2(n9599), .A(n7570), .ZN(P1_U3326) );
  AOI22_X1 U9185 ( .A1(n9640), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9861), .ZN(n7574) );
  OAI21_X1 U9186 ( .B1(n9833), .B2(n9644), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9187 ( .C1(n7575), .C2(n9640), .A(n7574), .B(n7573), .ZN(P1_U3291) );
  INV_X1 U9188 ( .A(n7578), .ZN(n7579) );
  AOI21_X1 U9189 ( .B1(n7576), .B2(n7577), .A(n7579), .ZN(n7584) );
  AOI22_X1 U9190 ( .A1(n8765), .A2(n4480), .B1(n8757), .B2(n9077), .ZN(n7580)
         );
  OAI21_X1 U9191 ( .B1(n9888), .B2(n8760), .A(n7580), .ZN(n7581) );
  AOI21_X1 U9192 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7582), .A(n7581), .ZN(
        n7583) );
  OAI21_X1 U9193 ( .B1(n7584), .B2(n8772), .A(n7583), .ZN(P1_U3235) );
  INV_X1 U9194 ( .A(n7587), .ZN(n7589) );
  MUX2_X1 U9195 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6040), .Z(n7850) );
  INV_X1 U9196 ( .A(SI_29_), .ZN(n7590) );
  XNOR2_X1 U9197 ( .A(n7850), .B(n7590), .ZN(n7591) );
  INV_X1 U9198 ( .A(n8774), .ZN(n8621) );
  INV_X1 U9199 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7592) );
  OAI222_X1 U9200 ( .A1(n7594), .A2(n8621), .B1(n7593), .B2(P1_U3084), .C1(
        n7592), .C2(n9595), .ZN(P1_U3324) );
  NAND2_X1 U9201 ( .A1(n7595), .A2(n6185), .ZN(n7597) );
  NAND2_X1 U9202 ( .A1(n7867), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7596) );
  INV_X1 U9203 ( .A(n8523), .ZN(n8254) );
  NAND2_X1 U9204 ( .A1(n7598), .A2(n6185), .ZN(n7600) );
  NAND2_X1 U9205 ( .A1(n7867), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7599) );
  XNOR2_X1 U9206 ( .A(n8540), .B(n7660), .ZN(n7627) );
  INV_X1 U9207 ( .A(n7627), .ZN(n7778) );
  INV_X1 U9208 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U9209 ( .A1(n7601), .A2(n10380), .ZN(n7602) );
  AND2_X1 U9210 ( .A1(n7635), .A2(n7602), .ZN(n8308) );
  INV_X1 U9211 ( .A(n7648), .ZN(n7742) );
  NAND2_X1 U9212 ( .A1(n8308), .A2(n7742), .ZN(n7605) );
  NAND2_X1 U9213 ( .A1(n7637), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7603) );
  NOR2_X1 U9214 ( .A1(n8285), .A2(n7722), .ZN(n7628) );
  INV_X1 U9215 ( .A(n7628), .ZN(n7781) );
  INV_X1 U9216 ( .A(n8285), .ZN(n8318) );
  NAND2_X1 U9217 ( .A1(n7607), .A2(n6185), .ZN(n7609) );
  NAND2_X1 U9218 ( .A1(n7867), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7608) );
  XNOR2_X1 U9219 ( .A(n8366), .B(n7660), .ZN(n7610) );
  NOR2_X1 U9220 ( .A1(n8345), .A2(n7722), .ZN(n7611) );
  XNOR2_X1 U9221 ( .A(n7610), .B(n7611), .ZN(n7748) );
  INV_X1 U9222 ( .A(n7610), .ZN(n7612) );
  NAND2_X1 U9223 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  NAND2_X1 U9224 ( .A1(n7614), .A2(n6185), .ZN(n7616) );
  NAND2_X1 U9225 ( .A1(n7867), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7615) );
  XNOR2_X1 U9226 ( .A(n8549), .B(n7723), .ZN(n7617) );
  NAND2_X1 U9227 ( .A1(n8317), .A2(n7877), .ZN(n7787) );
  INV_X1 U9228 ( .A(n7617), .ZN(n7618) );
  NOR2_X1 U9229 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  NAND2_X1 U9230 ( .A1(n7621), .A2(n6185), .ZN(n7623) );
  NAND2_X1 U9231 ( .A1(n7867), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7622) );
  XNOR2_X1 U9232 ( .A(n8324), .B(n7660), .ZN(n7624) );
  AND2_X1 U9233 ( .A1(n7840), .A2(n7877), .ZN(n7703) );
  OAI211_X1 U9234 ( .C1(n8318), .C2(n7627), .A(n7704), .B(n7703), .ZN(n7630)
         );
  INV_X1 U9235 ( .A(n7624), .ZN(n7625) );
  AND2_X1 U9236 ( .A1(n7626), .A2(n7625), .ZN(n7776) );
  OAI21_X1 U9237 ( .B1(n7628), .B2(n7627), .A(n7776), .ZN(n7629) );
  NAND2_X1 U9238 ( .A1(n7631), .A2(n6185), .ZN(n7633) );
  NAND2_X1 U9239 ( .A1(n7867), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7632) );
  XNOR2_X1 U9240 ( .A(n8535), .B(n7723), .ZN(n7809) );
  INV_X1 U9241 ( .A(n7635), .ZN(n7634) );
  NAND2_X1 U9242 ( .A1(n7634), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7646) );
  INV_X1 U9243 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U9244 ( .A1(n7635), .A2(n10473), .ZN(n7636) );
  NAND2_X1 U9245 ( .A1(n7646), .A2(n7636), .ZN(n8288) );
  OR2_X1 U9246 ( .A1(n8288), .A2(n7648), .ZN(n7640) );
  NAND2_X1 U9247 ( .A1(n7637), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7638) );
  INV_X1 U9248 ( .A(n8212), .ZN(n8072) );
  NAND2_X1 U9249 ( .A1(n8072), .A2(n7877), .ZN(n7641) );
  NOR2_X1 U9250 ( .A1(n7809), .A2(n7641), .ZN(n7642) );
  AOI21_X1 U9251 ( .B1(n7809), .B2(n7641), .A(n7642), .ZN(n7759) );
  INV_X1 U9252 ( .A(n7642), .ZN(n7659) );
  NAND2_X1 U9253 ( .A1(n7643), .A2(n6185), .ZN(n7645) );
  NAND2_X1 U9254 ( .A1(n7867), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7644) );
  XNOR2_X1 U9255 ( .A(n8529), .B(n7660), .ZN(n7655) );
  INV_X1 U9256 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U9257 ( .A1(n7646), .A2(n10460), .ZN(n7647) );
  NAND2_X1 U9258 ( .A1(n7680), .A2(n7647), .ZN(n8277) );
  OR2_X1 U9259 ( .A1(n8277), .A2(n7648), .ZN(n7654) );
  INV_X1 U9260 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9261 ( .A1(n7737), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7650) );
  OAI211_X1 U9262 ( .C1(n7651), .C2(n6274), .A(n7650), .B(n7649), .ZN(n7652)
         );
  INV_X1 U9263 ( .A(n7652), .ZN(n7653) );
  NOR2_X1 U9264 ( .A1(n8286), .A2(n7722), .ZN(n7656) );
  NAND2_X1 U9265 ( .A1(n7655), .A2(n7656), .ZN(n7673) );
  INV_X1 U9266 ( .A(n7655), .ZN(n7672) );
  INV_X1 U9267 ( .A(n7656), .ZN(n7657) );
  NAND2_X1 U9268 ( .A1(n7672), .A2(n7657), .ZN(n7658) );
  NAND2_X1 U9269 ( .A1(n7673), .A2(n7658), .ZN(n7811) );
  INV_X1 U9270 ( .A(n7674), .ZN(n7813) );
  XNOR2_X1 U9271 ( .A(n8523), .B(n7660), .ZN(n7667) );
  XNOR2_X1 U9272 ( .A(n7680), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9273 ( .A1(n8252), .A2(n7742), .ZN(n7666) );
  INV_X1 U9274 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U9275 ( .A1(n7737), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7661) );
  OAI211_X1 U9276 ( .C1(n4481), .C2(n7663), .A(n7662), .B(n7661), .ZN(n7664)
         );
  INV_X1 U9277 ( .A(n7664), .ZN(n7665) );
  AND2_X1 U9278 ( .A1(n8241), .A2(n7877), .ZN(n7668) );
  NAND2_X1 U9279 ( .A1(n7667), .A2(n7668), .ZN(n7726) );
  INV_X1 U9280 ( .A(n7667), .ZN(n7670) );
  INV_X1 U9281 ( .A(n7668), .ZN(n7669) );
  NAND2_X1 U9282 ( .A1(n7670), .A2(n7669), .ZN(n7671) );
  AOI21_X1 U9283 ( .B1(n7813), .B2(n4571), .A(n7810), .ZN(n7676) );
  NOR3_X1 U9284 ( .A1(n7672), .A2(n8286), .A3(n7808), .ZN(n7675) );
  OAI21_X1 U9285 ( .B1(n7676), .B2(n7675), .A(n7727), .ZN(n7689) );
  INV_X1 U9286 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7679) );
  OAI22_X1 U9287 ( .A1(n8286), .A2(n7830), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7679), .ZN(n7687) );
  NAND2_X1 U9288 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n7677) );
  INV_X1 U9289 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7678) );
  OAI21_X1 U9290 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  INV_X1 U9291 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U9292 ( .A1(n7737), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7683) );
  OAI211_X1 U9293 ( .C1(n7684), .C2(n4481), .A(n7683), .B(n7682), .ZN(n7685)
         );
  NOR2_X1 U9294 ( .A1(n8218), .A2(n7829), .ZN(n7686) );
  AOI211_X1 U9295 ( .C1(n7805), .C2(n8252), .A(n7687), .B(n7686), .ZN(n7688)
         );
  OAI211_X1 U9296 ( .C1(n8254), .C2(n7835), .A(n7689), .B(n7688), .ZN(P2_U3216) );
  INV_X1 U9297 ( .A(n7690), .ZN(n7693) );
  NOR3_X1 U9298 ( .A1(n7691), .A2(n8492), .A3(n7808), .ZN(n7692) );
  AOI21_X1 U9299 ( .B1(n7693), .B2(n7823), .A(n7692), .ZN(n7702) );
  AOI22_X1 U9300 ( .A1(n7745), .A2(n8074), .B1(n7694), .B2(n8196), .ZN(n7696)
         );
  OAI211_X1 U9301 ( .C1(n8482), .C2(n7828), .A(n7696), .B(n7695), .ZN(n7699)
         );
  NOR2_X1 U9302 ( .A1(n7697), .A2(n7810), .ZN(n7698) );
  AOI211_X1 U9303 ( .C1(n8590), .C2(n7793), .A(n7699), .B(n7698), .ZN(n7700)
         );
  OAI21_X1 U9304 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(P2_U3217) );
  AOI22_X1 U9305 ( .A1(n7704), .A2(n7823), .B1(n7822), .B2(n7840), .ZN(n7708)
         );
  OAI22_X1 U9306 ( .A1(n7828), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10461), .ZN(n7706) );
  OAI22_X1 U9307 ( .A1(n8285), .A2(n7829), .B1(n7830), .B2(n8359), .ZN(n7705)
         );
  AOI211_X1 U9308 ( .C1(n8543), .C2(n7793), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OAI21_X1 U9309 ( .B1(n7708), .B2(n7777), .A(n7707), .ZN(P2_U3218) );
  OAI21_X1 U9310 ( .B1(n7714), .B2(n7800), .A(n7709), .ZN(n7710) );
  NAND2_X1 U9311 ( .A1(n7710), .A2(n7823), .ZN(n7718) );
  NOR2_X1 U9312 ( .A1(n7829), .A2(n8392), .ZN(n7712) );
  OAI22_X1 U9313 ( .A1(n7828), .A2(n8396), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10426), .ZN(n7711) );
  AOI211_X1 U9314 ( .C1(n8567), .C2(n7793), .A(n7712), .B(n7711), .ZN(n7717)
         );
  NOR3_X1 U9315 ( .A1(n7714), .A2(n7713), .A3(n7808), .ZN(n7715) );
  OAI21_X1 U9316 ( .B1(n7715), .B2(n7745), .A(n8200), .ZN(n7716) );
  NAND3_X1 U9317 ( .A1(n7718), .A2(n7717), .A3(n7716), .ZN(P2_U3221) );
  NAND2_X1 U9318 ( .A1(n7719), .A2(n6185), .ZN(n7721) );
  NAND2_X1 U9319 ( .A1(n7867), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7720) );
  OR2_X1 U9320 ( .A1(n8218), .A2(n7722), .ZN(n7724) );
  XNOR2_X1 U9321 ( .A(n7724), .B(n7723), .ZN(n7728) );
  INV_X1 U9322 ( .A(n7728), .ZN(n7729) );
  NOR3_X1 U9323 ( .A1(n4771), .A2(n7729), .A3(n7793), .ZN(n7725) );
  AOI21_X1 U9324 ( .B1(n4771), .B2(n7729), .A(n7725), .ZN(n7735) );
  NOR3_X1 U9325 ( .A1(n4771), .A2(n7728), .A3(n7793), .ZN(n7731) );
  NOR2_X1 U9326 ( .A1(n8517), .A2(n7729), .ZN(n7730) );
  OAI21_X1 U9327 ( .B1(n4771), .B2(n7835), .A(n7810), .ZN(n7732) );
  OAI211_X1 U9328 ( .C1(n7735), .C2(n7734), .A(n7733), .B(n7732), .ZN(n7747)
         );
  INV_X1 U9329 ( .A(n7736), .ZN(n8227) );
  INV_X1 U9330 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U9331 ( .A1(n7737), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7738) );
  OAI211_X1 U9332 ( .C1(n6274), .C2(n7740), .A(n7739), .B(n7738), .ZN(n7741)
         );
  AOI21_X1 U9333 ( .B1(n8227), .B2(n7742), .A(n7741), .ZN(n8071) );
  AOI22_X1 U9334 ( .A1(n8235), .A2(n7805), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7743) );
  OAI21_X1 U9335 ( .B1(n8071), .B2(n7829), .A(n7743), .ZN(n7744) );
  AOI21_X1 U9336 ( .B1(n7745), .B2(n8241), .A(n7744), .ZN(n7746) );
  NAND2_X1 U9337 ( .A1(n7747), .A2(n7746), .ZN(P2_U3222) );
  INV_X1 U9338 ( .A(n7748), .ZN(n7749) );
  AOI21_X1 U9339 ( .B1(n7750), .B2(n7749), .A(n7810), .ZN(n7754) );
  NOR3_X1 U9340 ( .A1(n7751), .A2(n8392), .A3(n7808), .ZN(n7753) );
  OAI21_X1 U9341 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n7758) );
  OAI22_X1 U9342 ( .A1(n7828), .A2(n8362), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10455), .ZN(n7756) );
  OAI22_X1 U9343 ( .A1(n7830), .A2(n8392), .B1(n8359), .B2(n7829), .ZN(n7755)
         );
  AOI211_X1 U9344 ( .C1(n8555), .C2(n7793), .A(n7756), .B(n7755), .ZN(n7757)
         );
  NAND2_X1 U9345 ( .A1(n7758), .A2(n7757), .ZN(P2_U3225) );
  OAI211_X1 U9346 ( .C1(n7760), .C2(n7759), .A(n7812), .B(n7823), .ZN(n7764)
         );
  OAI22_X1 U9347 ( .A1(n8288), .A2(n7828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10473), .ZN(n7762) );
  OAI22_X1 U9348 ( .A1(n8286), .A2(n7829), .B1(n8285), .B2(n7830), .ZN(n7761)
         );
  AOI211_X1 U9349 ( .C1(n8535), .C2(n7793), .A(n7762), .B(n7761), .ZN(n7763)
         );
  NAND2_X1 U9350 ( .A1(n7764), .A2(n7763), .ZN(P2_U3227) );
  XNOR2_X1 U9351 ( .A(n7766), .B(n7765), .ZN(n7825) );
  AOI22_X1 U9352 ( .A1(n7825), .A2(n7824), .B1(n7767), .B2(n7766), .ZN(n7771)
         );
  XNOR2_X1 U9353 ( .A(n7769), .B(n7768), .ZN(n7770) );
  XNOR2_X1 U9354 ( .A(n7771), .B(n7770), .ZN(n7775) );
  OAI22_X1 U9355 ( .A1(n7828), .A2(n8452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8128), .ZN(n7773) );
  OAI22_X1 U9356 ( .A1(n7830), .A2(n8490), .B1(n8445), .B2(n7829), .ZN(n7772)
         );
  AOI211_X1 U9357 ( .C1(n8580), .C2(n7793), .A(n7773), .B(n7772), .ZN(n7774)
         );
  OAI21_X1 U9358 ( .B1(n7775), .B2(n7810), .A(n7774), .ZN(P2_U3228) );
  INV_X1 U9359 ( .A(n8540), .ZN(n8311) );
  NOR2_X1 U9360 ( .A1(n7777), .A2(n7776), .ZN(n7779) );
  XNOR2_X1 U9361 ( .A(n7779), .B(n7778), .ZN(n7782) );
  OAI22_X1 U9362 ( .A1(n7782), .A2(n7810), .B1(n8285), .B2(n7808), .ZN(n7780)
         );
  OAI21_X1 U9363 ( .B1(n7782), .B2(n7781), .A(n7780), .ZN(n7786) );
  OAI22_X1 U9364 ( .A1(n8212), .A2(n8434), .B1(n8346), .B2(n8491), .ZN(n8303)
         );
  INV_X1 U9365 ( .A(n8308), .ZN(n7783) );
  OAI22_X1 U9366 ( .A1(n7783), .A2(n7828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10380), .ZN(n7784) );
  AOI21_X1 U9367 ( .B1(n8303), .B2(n7819), .A(n7784), .ZN(n7785) );
  OAI211_X1 U9368 ( .C1(n8311), .C2(n7835), .A(n7786), .B(n7785), .ZN(P2_U3231) );
  NAND2_X1 U9369 ( .A1(n7822), .A2(n8317), .ZN(n7790) );
  NAND2_X1 U9370 ( .A1(n7787), .A2(n7823), .ZN(n7789) );
  MUX2_X1 U9371 ( .A(n7790), .B(n7789), .S(n7788), .Z(n7795) );
  OAI22_X1 U9372 ( .A1(n7828), .A2(n8336), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10489), .ZN(n7792) );
  OAI22_X1 U9373 ( .A1(n7830), .A2(n8345), .B1(n8346), .B2(n7829), .ZN(n7791)
         );
  AOI211_X1 U9374 ( .C1(n8549), .C2(n7793), .A(n7792), .B(n7791), .ZN(n7794)
         );
  NAND2_X1 U9375 ( .A1(n7795), .A2(n7794), .ZN(P2_U3237) );
  INV_X1 U9376 ( .A(n7796), .ZN(n7797) );
  AOI21_X1 U9377 ( .B1(n7798), .B2(n7797), .A(n7810), .ZN(n7802) );
  NOR3_X1 U9378 ( .A1(n7799), .A2(n8445), .A3(n7808), .ZN(n7801) );
  OAI21_X1 U9379 ( .B1(n7802), .B2(n7801), .A(n7800), .ZN(n7807) );
  INV_X1 U9380 ( .A(n7803), .ZN(n8406) );
  AND2_X1 U9381 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8161) );
  OAI22_X1 U9382 ( .A1(n7830), .A2(n8445), .B1(n8412), .B2(n7829), .ZN(n7804)
         );
  AOI211_X1 U9383 ( .C1(n7805), .C2(n8406), .A(n8161), .B(n7804), .ZN(n7806)
         );
  OAI211_X1 U9384 ( .C1(n8408), .C2(n7835), .A(n7807), .B(n7806), .ZN(P2_U3240) );
  INV_X1 U9385 ( .A(n8529), .ZN(n8182) );
  NOR3_X1 U9386 ( .A1(n7809), .A2(n8212), .A3(n7808), .ZN(n7815) );
  AOI21_X1 U9387 ( .B1(n7812), .B2(n7811), .A(n7810), .ZN(n7814) );
  OAI21_X1 U9388 ( .B1(n7815), .B2(n7814), .A(n7813), .ZN(n7821) );
  NAND2_X1 U9389 ( .A1(n8241), .A2(n8471), .ZN(n7817) );
  NAND2_X1 U9390 ( .A1(n8072), .A2(n8469), .ZN(n7816) );
  NAND2_X1 U9391 ( .A1(n7817), .A2(n7816), .ZN(n8269) );
  OAI22_X1 U9392 ( .A1(n8277), .A2(n7828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10460), .ZN(n7818) );
  AOI21_X1 U9393 ( .B1(n8269), .B2(n7819), .A(n7818), .ZN(n7820) );
  OAI211_X1 U9394 ( .C1(n8182), .C2(n7835), .A(n7821), .B(n7820), .ZN(P2_U3242) );
  INV_X1 U9395 ( .A(n8585), .ZN(n8466) );
  NAND2_X1 U9396 ( .A1(n7822), .A2(n8196), .ZN(n7827) );
  NAND2_X1 U9397 ( .A1(n7824), .A2(n7823), .ZN(n7826) );
  MUX2_X1 U9398 ( .A(n7827), .B(n7826), .S(n7825), .Z(n7834) );
  NOR2_X1 U9399 ( .A1(n7828), .A2(n8463), .ZN(n7832) );
  OAI22_X1 U9400 ( .A1(n7830), .A2(n8073), .B1(n8435), .B2(n7829), .ZN(n7831)
         );
  AOI211_X1 U9401 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(P2_U3152), .A(n7832), 
        .B(n7831), .ZN(n7833) );
  OAI211_X1 U9402 ( .C1(n8466), .C2(n7835), .A(n7834), .B(n7833), .ZN(P2_U3243) );
  INV_X1 U9403 ( .A(n7945), .ZN(n8489) );
  NAND2_X1 U9404 ( .A1(n8590), .A2(n8073), .ZN(n7950) );
  NAND2_X1 U9405 ( .A1(n7949), .A2(n7950), .ZN(n8488) );
  INV_X1 U9406 ( .A(n7949), .ZN(n7836) );
  NAND2_X1 U9407 ( .A1(n8585), .A2(n8490), .ZN(n7952) );
  NAND2_X1 U9408 ( .A1(n7953), .A2(n7952), .ZN(n8197) );
  OAI21_X2 U9409 ( .B1(n8468), .B2(n8197), .A(n7953), .ZN(n8442) );
  NAND2_X1 U9410 ( .A1(n8580), .A2(n8435), .ZN(n7956) );
  NOR2_X1 U9411 ( .A1(n8442), .A2(n8443), .ZN(n8428) );
  INV_X1 U9412 ( .A(n7956), .ZN(n8429) );
  NAND2_X1 U9413 ( .A1(n8577), .A2(n8445), .ZN(n7962) );
  INV_X1 U9414 ( .A(n8430), .ZN(n7837) );
  NAND2_X1 U9415 ( .A1(n8570), .A2(n8433), .ZN(n7969) );
  NAND2_X1 U9416 ( .A1(n8387), .A2(n7969), .ZN(n8410) );
  OR2_X1 U9417 ( .A1(n8567), .A2(n8412), .ZN(n7977) );
  NAND2_X1 U9418 ( .A1(n8567), .A2(n8412), .ZN(n8375) );
  NAND2_X1 U9419 ( .A1(n7977), .A2(n8375), .ZN(n8384) );
  NAND2_X1 U9420 ( .A1(n8560), .A2(n8392), .ZN(n7979) );
  INV_X1 U9421 ( .A(n8376), .ZN(n7838) );
  NAND2_X1 U9422 ( .A1(n7838), .A2(n8375), .ZN(n7839) );
  NAND2_X1 U9423 ( .A1(n8555), .A2(n8345), .ZN(n8342) );
  NAND2_X1 U9424 ( .A1(n7980), .A2(n8342), .ZN(n8356) );
  NAND2_X1 U9425 ( .A1(n8549), .A2(n8359), .ZN(n7974) );
  INV_X1 U9426 ( .A(n8343), .ZN(n8332) );
  NAND2_X1 U9427 ( .A1(n8324), .A2(n7840), .ZN(n7985) );
  NAND2_X1 U9428 ( .A1(n8540), .A2(n8285), .ZN(n7989) );
  NAND2_X1 U9429 ( .A1(n8300), .A2(n7842), .ZN(n8299) );
  NAND2_X1 U9430 ( .A1(n8299), .A2(n7990), .ZN(n8282) );
  NAND2_X1 U9431 ( .A1(n8535), .A2(n8212), .ZN(n7993) );
  NAND2_X1 U9432 ( .A1(n8282), .A2(n8283), .ZN(n7843) );
  NAND2_X1 U9433 ( .A1(n7843), .A2(n7995), .ZN(n8265) );
  INV_X1 U9434 ( .A(n8241), .ZN(n8216) );
  OR2_X1 U9435 ( .A1(n8523), .A2(n8216), .ZN(n8001) );
  NAND2_X1 U9436 ( .A1(n8517), .A2(n8218), .ZN(n8007) );
  NAND2_X1 U9437 ( .A1(n7845), .A2(n8007), .ZN(n8238) );
  INV_X1 U9438 ( .A(n7845), .ZN(n8005) );
  NAND2_X1 U9439 ( .A1(n8774), .A2(n6185), .ZN(n7847) );
  NAND2_X1 U9440 ( .A1(n7867), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U9441 ( .A1(n8183), .A2(n8071), .ZN(n8012) );
  INV_X1 U9442 ( .A(n8221), .ZN(n7848) );
  NAND2_X1 U9443 ( .A1(n8220), .A2(n7848), .ZN(n7849) );
  NOR2_X1 U9444 ( .A1(n7850), .A2(SI_29_), .ZN(n7852) );
  NAND2_X1 U9445 ( .A1(n7850), .A2(SI_29_), .ZN(n7851) );
  MUX2_X1 U9446 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6040), .Z(n7859) );
  XNOR2_X1 U9447 ( .A(n7857), .B(SI_30_), .ZN(n8837) );
  NAND2_X1 U9448 ( .A1(n8837), .A2(n6185), .ZN(n7855) );
  NAND2_X1 U9449 ( .A1(n7867), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7854) );
  NOR2_X1 U9450 ( .A1(n8186), .A2(n8062), .ZN(n7856) );
  INV_X1 U9451 ( .A(n7857), .ZN(n7858) );
  NAND2_X1 U9452 ( .A1(n7858), .A2(SI_30_), .ZN(n7862) );
  NAND2_X1 U9453 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  NAND2_X1 U9454 ( .A1(n7862), .A2(n7861), .ZN(n7865) );
  MUX2_X1 U9455 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6040), .Z(n7863) );
  XNOR2_X1 U9456 ( .A(n7863), .B(SI_31_), .ZN(n7864) );
  NAND2_X1 U9457 ( .A1(n7867), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7868) );
  INV_X1 U9458 ( .A(n8186), .ZN(n7874) );
  INV_X1 U9459 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U9460 ( .A1(n7737), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7869) );
  OAI211_X1 U9461 ( .C1(n4481), .C2(n7871), .A(n7870), .B(n7869), .ZN(n8222)
         );
  INV_X1 U9462 ( .A(n8222), .ZN(n7872) );
  NAND2_X1 U9463 ( .A1(n8190), .A2(n7872), .ZN(n8013) );
  NAND2_X1 U9464 ( .A1(n8502), .A2(n7874), .ZN(n8022) );
  XNOR2_X1 U9465 ( .A(n7875), .B(n9980), .ZN(n7878) );
  AND2_X1 U9466 ( .A1(n7890), .A2(n9980), .ZN(n7879) );
  AND2_X1 U9467 ( .A1(n7880), .A2(n7879), .ZN(n8017) );
  INV_X1 U9468 ( .A(n8017), .ZN(n8020) );
  NAND2_X1 U9469 ( .A1(n7884), .A2(n7881), .ZN(n7882) );
  NAND2_X1 U9470 ( .A1(n7886), .A2(n8020), .ZN(n7900) );
  NAND2_X1 U9471 ( .A1(n6871), .A2(n9985), .ZN(n7887) );
  NAND3_X1 U9472 ( .A1(n7893), .A2(n7888), .A3(n7887), .ZN(n7889) );
  NAND2_X1 U9473 ( .A1(n7889), .A2(n7891), .ZN(n7896) );
  AND2_X1 U9474 ( .A1(n9985), .A2(n7890), .ZN(n7892) );
  OAI211_X1 U9475 ( .C1(n6872), .C2(n7892), .A(n7891), .B(n6871), .ZN(n7894)
         );
  NAND2_X1 U9476 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  MUX2_X1 U9477 ( .A(n7896), .B(n7895), .S(n8020), .Z(n7898) );
  INV_X1 U9478 ( .A(n7897), .ZN(n7907) );
  NAND3_X1 U9479 ( .A1(n7898), .A2(n4478), .A3(n7907), .ZN(n7899) );
  NAND2_X1 U9480 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U9481 ( .A1(n7901), .A2(n7908), .ZN(n7912) );
  INV_X1 U9482 ( .A(n7902), .ZN(n7906) );
  NAND2_X1 U9483 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  NAND2_X1 U9484 ( .A1(n7909), .A2(n7908), .ZN(n7910) );
  NAND2_X1 U9485 ( .A1(n7910), .A2(n8017), .ZN(n7911) );
  NAND2_X1 U9486 ( .A1(n7912), .A2(n7911), .ZN(n7916) );
  NOR2_X1 U9487 ( .A1(n7913), .A2(n8020), .ZN(n7914) );
  NOR2_X1 U9488 ( .A1(n7914), .A2(n8040), .ZN(n7915) );
  NAND2_X1 U9489 ( .A1(n7916), .A2(n7915), .ZN(n7920) );
  MUX2_X1 U9490 ( .A(n7918), .B(n7917), .S(n8020), .Z(n7919) );
  MUX2_X1 U9491 ( .A(n8080), .B(n7924), .S(n8020), .Z(n7925) );
  NAND3_X1 U9492 ( .A1(n7930), .A2(n7931), .A3(n7926), .ZN(n7927) );
  NAND3_X1 U9493 ( .A1(n7927), .A2(n7935), .A3(n7929), .ZN(n7934) );
  NAND3_X1 U9494 ( .A1(n7932), .A2(n7938), .A3(n7931), .ZN(n7933) );
  NAND3_X1 U9495 ( .A1(n7939), .A2(n7941), .A3(n7935), .ZN(n7937) );
  NAND2_X1 U9496 ( .A1(n7937), .A2(n7936), .ZN(n7944) );
  NAND2_X1 U9497 ( .A1(n7939), .A2(n7938), .ZN(n7942) );
  AOI21_X1 U9498 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7943) );
  INV_X1 U9499 ( .A(n8488), .ZN(n8480) );
  MUX2_X1 U9500 ( .A(n7946), .B(n7945), .S(n8020), .Z(n7947) );
  INV_X1 U9501 ( .A(n8197), .ZN(n8467) );
  MUX2_X1 U9502 ( .A(n7950), .B(n7949), .S(n8020), .Z(n7951) );
  INV_X1 U9503 ( .A(n8443), .ZN(n7955) );
  MUX2_X1 U9504 ( .A(n7953), .B(n7952), .S(n8020), .Z(n7954) );
  NAND2_X1 U9505 ( .A1(n7957), .A2(n8430), .ZN(n7968) );
  INV_X1 U9506 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9507 ( .A1(n8430), .A2(n7959), .ZN(n7961) );
  NAND3_X1 U9508 ( .A1(n7961), .A2(n7960), .A3(n8387), .ZN(n7964) );
  INV_X1 U9509 ( .A(n7962), .ZN(n7963) );
  MUX2_X1 U9510 ( .A(n7964), .B(n7963), .S(n8017), .Z(n7966) );
  INV_X1 U9511 ( .A(n7969), .ZN(n7965) );
  NOR2_X1 U9512 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  NAND2_X1 U9513 ( .A1(n7968), .A2(n7967), .ZN(n7976) );
  NAND3_X1 U9514 ( .A1(n7976), .A2(n7969), .A3(n8375), .ZN(n7970) );
  NAND2_X1 U9515 ( .A1(n7970), .A2(n7977), .ZN(n7971) );
  NAND2_X1 U9516 ( .A1(n7971), .A2(n7979), .ZN(n7972) );
  NAND3_X1 U9517 ( .A1(n7972), .A2(n7978), .A3(n7980), .ZN(n7973) );
  NAND3_X1 U9518 ( .A1(n7973), .A2(n8342), .A3(n8020), .ZN(n7975) );
  MUX2_X1 U9519 ( .A(n8020), .B(n7975), .S(n7974), .Z(n7984) );
  NAND3_X1 U9520 ( .A1(n7981), .A2(n8017), .A3(n7980), .ZN(n7982) );
  MUX2_X1 U9521 ( .A(n7982), .B(n8017), .S(n8315), .Z(n7983) );
  INV_X1 U9522 ( .A(n8326), .ZN(n8054) );
  NAND2_X1 U9523 ( .A1(n7989), .A2(n8302), .ZN(n7987) );
  NAND2_X1 U9524 ( .A1(n8301), .A2(n7985), .ZN(n7986) );
  MUX2_X1 U9525 ( .A(n7987), .B(n7986), .S(n8017), .Z(n7988) );
  INV_X1 U9526 ( .A(n7988), .ZN(n7992) );
  MUX2_X1 U9527 ( .A(n7990), .B(n7989), .S(n8017), .Z(n7991) );
  INV_X1 U9528 ( .A(n8264), .ZN(n8267) );
  AOI21_X1 U9529 ( .B1(n8267), .B2(n7993), .A(n8017), .ZN(n7994) );
  NAND2_X1 U9530 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  NAND2_X1 U9531 ( .A1(n7997), .A2(n8017), .ZN(n8000) );
  OAI21_X1 U9532 ( .B1(n7998), .B2(n8020), .A(n8256), .ZN(n7999) );
  INV_X1 U9533 ( .A(n8001), .ZN(n8003) );
  OAI21_X1 U9534 ( .B1(n8254), .B2(n8241), .A(n8007), .ZN(n8002) );
  MUX2_X1 U9535 ( .A(n8003), .B(n8002), .S(n8020), .Z(n8004) );
  AOI21_X1 U9536 ( .B1(n8006), .B2(n8218), .A(n8221), .ZN(n8010) );
  AND2_X1 U9537 ( .A1(n8011), .A2(n8017), .ZN(n8009) );
  OAI211_X1 U9538 ( .C1(n8017), .C2(n8517), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI21_X1 U9539 ( .B1(n8010), .B2(n8009), .A(n8008), .ZN(n8016) );
  MUX2_X1 U9540 ( .A(n8012), .B(n8011), .S(n8020), .Z(n8015) );
  NAND2_X1 U9541 ( .A1(n4520), .A2(n8013), .ZN(n8014) );
  AOI21_X1 U9542 ( .B1(n8016), .B2(n8015), .A(n8014), .ZN(n8019) );
  NAND2_X1 U9543 ( .A1(n8022), .A2(n4520), .ZN(n8058) );
  MUX2_X1 U9544 ( .A(n8058), .B(n8059), .S(n8017), .Z(n8018) );
  MUX2_X1 U9545 ( .A(n8022), .B(n8021), .S(n8020), .Z(n8023) );
  INV_X1 U9546 ( .A(n10008), .ZN(n8026) );
  NOR2_X1 U9547 ( .A1(n8061), .A2(n8026), .ZN(n8028) );
  INV_X1 U9548 ( .A(n8384), .ZN(n8386) );
  NOR2_X1 U9549 ( .A1(n8030), .A2(n8029), .ZN(n8038) );
  NOR2_X1 U9550 ( .A1(n8032), .A2(n8031), .ZN(n8037) );
  NAND3_X1 U9551 ( .A1(n6871), .A2(n9985), .A3(n8033), .ZN(n8034) );
  NOR2_X1 U9552 ( .A1(n6872), .A2(n8034), .ZN(n8036) );
  NAND4_X1 U9553 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8042)
         );
  NOR4_X1 U9554 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n8046)
         );
  NAND4_X1 U9555 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(n8048)
         );
  NOR2_X1 U9556 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  NAND3_X1 U9557 ( .A1(n8467), .A2(n8480), .A3(n8049), .ZN(n8050) );
  NOR2_X1 U9558 ( .A1(n8443), .A2(n8050), .ZN(n8051) );
  NAND4_X1 U9559 ( .A1(n8386), .A2(n8430), .A3(n4872), .A4(n8051), .ZN(n8052)
         );
  NOR3_X1 U9560 ( .A1(n8356), .A2(n8376), .A3(n8052), .ZN(n8053) );
  NAND4_X1 U9561 ( .A1(n8301), .A2(n8054), .A3(n8332), .A4(n8053), .ZN(n8055)
         );
  NOR4_X1 U9562 ( .A1(n8238), .A2(n8264), .A3(n8211), .A4(n8055), .ZN(n8056)
         );
  NAND2_X1 U9563 ( .A1(n8056), .A2(n8256), .ZN(n8057) );
  NOR4_X1 U9564 ( .A1(n8059), .A2(n8058), .A3(n8221), .A4(n8057), .ZN(n8060)
         );
  XNOR2_X1 U9565 ( .A(n8060), .B(n8275), .ZN(n8063) );
  NAND4_X1 U9566 ( .A1(n9996), .A2(n8185), .A3(n8469), .A4(n8066), .ZN(n8067)
         );
  OAI211_X1 U9567 ( .C1(n8069), .C2(n8068), .A(n8067), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8070) );
  MUX2_X1 U9568 ( .A(n8222), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8087), .Z(
        P2_U3582) );
  INV_X1 U9569 ( .A(n8071), .ZN(n8240) );
  MUX2_X1 U9570 ( .A(n8240), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8087), .Z(
        P2_U3581) );
  INV_X1 U9571 ( .A(n8218), .ZN(n8258) );
  MUX2_X1 U9572 ( .A(n8258), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8087), .Z(
        P2_U3580) );
  MUX2_X1 U9573 ( .A(n8241), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8087), .Z(
        P2_U3579) );
  INV_X1 U9574 ( .A(n8286), .ZN(n8257) );
  MUX2_X1 U9575 ( .A(n8257), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8087), .Z(
        P2_U3578) );
  MUX2_X1 U9576 ( .A(n8072), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8087), .Z(
        P2_U3577) );
  MUX2_X1 U9577 ( .A(n8318), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8087), .Z(
        P2_U3576) );
  INV_X1 U9578 ( .A(n8345), .ZN(n8379) );
  MUX2_X1 U9579 ( .A(n8379), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8087), .Z(
        P2_U3573) );
  INV_X1 U9580 ( .A(n8392), .ZN(n8205) );
  MUX2_X1 U9581 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8205), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9582 ( .A(n8378), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8087), .Z(
        P2_U3571) );
  MUX2_X1 U9583 ( .A(n8200), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8087), .Z(
        P2_U3570) );
  INV_X1 U9584 ( .A(n8445), .ZN(n8199) );
  MUX2_X1 U9585 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8199), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U9586 ( .A(n8435), .ZN(n8472) );
  MUX2_X1 U9587 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8472), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9588 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8196), .S(P2_U3966), .Z(
        P2_U3567) );
  INV_X1 U9589 ( .A(n8073), .ZN(n8470) );
  MUX2_X1 U9590 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8470), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9591 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8074), .S(P2_U3966), .Z(
        P2_U3565) );
  INV_X1 U9592 ( .A(n8075), .ZN(n8076) );
  MUX2_X1 U9593 ( .A(n8076), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8087), .Z(
        P2_U3564) );
  MUX2_X1 U9594 ( .A(n8077), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8087), .Z(
        P2_U3563) );
  MUX2_X1 U9595 ( .A(n8078), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8087), .Z(
        P2_U3562) );
  MUX2_X1 U9596 ( .A(n8079), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8087), .Z(
        P2_U3561) );
  MUX2_X1 U9597 ( .A(n8080), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8087), .Z(
        P2_U3560) );
  MUX2_X1 U9598 ( .A(n8081), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8087), .Z(
        P2_U3559) );
  MUX2_X1 U9599 ( .A(n8082), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8087), .Z(
        P2_U3558) );
  MUX2_X1 U9600 ( .A(n8083), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8087), .Z(
        P2_U3557) );
  MUX2_X1 U9601 ( .A(n8084), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8087), .Z(
        P2_U3556) );
  MUX2_X1 U9602 ( .A(n8085), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8087), .Z(
        P2_U3555) );
  MUX2_X1 U9603 ( .A(n8086), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8087), .Z(
        P2_U3554) );
  MUX2_X1 U9604 ( .A(n6759), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8087), .Z(
        P2_U3553) );
  MUX2_X1 U9605 ( .A(n8088), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8087), .Z(
        P2_U3552) );
  AOI211_X1 U9606 ( .C1(n8091), .C2(n8090), .A(n8089), .B(n9602), .ZN(n8092)
         );
  AOI21_X1 U9607 ( .B1(n9608), .B2(n8093), .A(n8092), .ZN(n8100) );
  NOR2_X1 U9608 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6178), .ZN(n8094) );
  AOI21_X1 U9609 ( .B1(n9966), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8094), .ZN(
        n8099) );
  OAI211_X1 U9610 ( .C1(n8097), .C2(n8096), .A(n9964), .B(n8095), .ZN(n8098)
         );
  NAND3_X1 U9611 ( .A1(n8100), .A2(n8099), .A3(n8098), .ZN(P2_U3254) );
  OAI21_X1 U9612 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8104) );
  NAND2_X1 U9613 ( .A1(n9965), .A2(n8104), .ZN(n8113) );
  NOR2_X1 U9614 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6219), .ZN(n8105) );
  AOI21_X1 U9615 ( .B1(n9966), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8105), .ZN(
        n8112) );
  NAND2_X1 U9616 ( .A1(n9608), .A2(n8106), .ZN(n8111) );
  OAI211_X1 U9617 ( .C1(n8109), .C2(n8108), .A(n9964), .B(n8107), .ZN(n8110)
         );
  NAND4_X1 U9618 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(
        P2_U3256) );
  NAND2_X1 U9619 ( .A1(n8115), .A2(n8114), .ZN(n8117) );
  NAND2_X1 U9620 ( .A1(n8117), .A2(n8116), .ZN(n8120) );
  NAND2_X1 U9621 ( .A1(n8135), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8118) );
  OAI21_X1 U9622 ( .B1(n8135), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8118), .ZN(
        n8119) );
  AOI211_X1 U9623 ( .C1(n8120), .C2(n8119), .A(n8134), .B(n9602), .ZN(n8133)
         );
  NAND2_X1 U9624 ( .A1(n8122), .A2(n8121), .ZN(n8124) );
  NAND2_X1 U9625 ( .A1(n8124), .A2(n8123), .ZN(n8126) );
  XNOR2_X1 U9626 ( .A(n8135), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8125) );
  NOR2_X1 U9627 ( .A1(n8125), .A2(n8126), .ZN(n8141) );
  AOI21_X1 U9628 ( .B1(n8126), .B2(n8125), .A(n8141), .ZN(n8127) );
  NOR2_X1 U9629 ( .A1(n8127), .A2(n9962), .ZN(n8132) );
  INV_X1 U9630 ( .A(n8135), .ZN(n8143) );
  NOR2_X1 U9631 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8128), .ZN(n8129) );
  AOI21_X1 U9632 ( .B1(n9966), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8129), .ZN(
        n8130) );
  OAI21_X1 U9633 ( .B1(n9961), .B2(n8143), .A(n8130), .ZN(n8131) );
  OR3_X1 U9634 ( .A1(n8133), .A2(n8132), .A3(n8131), .ZN(P2_U3261) );
  NAND2_X1 U9635 ( .A1(n8156), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8136) );
  OAI21_X1 U9636 ( .B1(n8156), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8136), .ZN(
        n8137) );
  AOI211_X1 U9637 ( .C1(n8138), .C2(n8137), .A(n8155), .B(n9602), .ZN(n8149)
         );
  INV_X1 U9638 ( .A(n8156), .ZN(n8151) );
  NOR2_X1 U9639 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8139), .ZN(n8140) );
  AOI21_X1 U9640 ( .B1(n9966), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8140), .ZN(
        n8147) );
  XNOR2_X1 U9641 ( .A(n8151), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8145) );
  AOI21_X1 U9642 ( .B1(n8143), .B2(n8142), .A(n8141), .ZN(n8144) );
  NAND2_X1 U9643 ( .A1(n8145), .A2(n8144), .ZN(n8150) );
  OAI211_X1 U9644 ( .C1(n8145), .C2(n8144), .A(n9964), .B(n8150), .ZN(n8146)
         );
  OAI211_X1 U9645 ( .C1(n9961), .C2(n8151), .A(n8147), .B(n8146), .ZN(n8148)
         );
  OR2_X1 U9646 ( .A1(n8149), .A2(n8148), .ZN(P2_U3262) );
  OAI21_X1 U9647 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8154) );
  INV_X1 U9648 ( .A(n8157), .ZN(n8171) );
  AOI22_X1 U9649 ( .A1(n8157), .A2(n8170), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8171), .ZN(n8153) );
  NOR2_X1 U9650 ( .A1(n8154), .A2(n8153), .ZN(n8169) );
  AOI21_X1 U9651 ( .B1(n8154), .B2(n8153), .A(n8169), .ZN(n8164) );
  XNOR2_X1 U9652 ( .A(n8165), .B(n8157), .ZN(n8158) );
  NAND2_X1 U9653 ( .A1(n8158), .A2(n6374), .ZN(n8167) );
  OAI21_X1 U9654 ( .B1(n8158), .B2(n6374), .A(n8167), .ZN(n8159) );
  NAND2_X1 U9655 ( .A1(n8159), .A2(n9965), .ZN(n8163) );
  NOR2_X1 U9656 ( .A1(n9961), .A2(n8171), .ZN(n8160) );
  AOI211_X1 U9657 ( .C1(n9966), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8161), .B(
        n8160), .ZN(n8162) );
  OAI211_X1 U9658 ( .C1(n8164), .C2(n9962), .A(n8163), .B(n8162), .ZN(P2_U3263) );
  NAND2_X1 U9659 ( .A1(n8165), .A2(n8171), .ZN(n8166) );
  NAND2_X1 U9660 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  XNOR2_X1 U9661 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8168), .ZN(n8176) );
  INV_X1 U9662 ( .A(n8176), .ZN(n8174) );
  AOI21_X1 U9663 ( .B1(n8171), .B2(n8170), .A(n8169), .ZN(n8172) );
  XOR2_X1 U9664 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8172), .Z(n8175) );
  OAI21_X1 U9665 ( .B1(n8175), .B2(n9962), .A(n9961), .ZN(n8173) );
  AOI21_X1 U9666 ( .B1(n8174), .B2(n9965), .A(n8173), .ZN(n8178) );
  AOI22_X1 U9667 ( .A1(n8176), .A2(n9965), .B1(n9964), .B2(n8175), .ZN(n8177)
         );
  MUX2_X1 U9668 ( .A(n8178), .B(n8177), .S(n8275), .Z(n8180) );
  NAND2_X1 U9669 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8179) );
  OAI211_X1 U9670 ( .C1(n4784), .C2(n8181), .A(n8180), .B(n8179), .ZN(P2_U3264) );
  INV_X1 U9671 ( .A(n8590), .ZN(n8485) );
  NAND2_X1 U9672 ( .A1(n8421), .A2(n8408), .ZN(n8403) );
  XOR2_X1 U9673 ( .A(n8502), .B(n8189), .Z(n8504) );
  NOR2_X1 U9674 ( .A1(n9993), .A2(n8184), .ZN(n8187) );
  AOI21_X1 U9675 ( .B1(n8185), .B2(P2_B_REG_SCAN_IN), .A(n8434), .ZN(n8223) );
  NAND2_X1 U9676 ( .A1(n8186), .A2(n8223), .ZN(n8507) );
  NOR2_X1 U9677 ( .A1(n8507), .A2(n8289), .ZN(n8191) );
  AOI211_X1 U9678 ( .C1(n8502), .C2(n8455), .A(n8187), .B(n8191), .ZN(n8188)
         );
  OAI21_X1 U9679 ( .B1(n8504), .B2(n9989), .A(n8188), .ZN(P2_U3265) );
  INV_X1 U9680 ( .A(n8190), .ZN(n8509) );
  INV_X1 U9681 ( .A(n8189), .ZN(n8506) );
  NAND2_X1 U9682 ( .A1(n8190), .A2(n8226), .ZN(n8505) );
  NAND3_X1 U9683 ( .A1(n8506), .A2(n8499), .A3(n8505), .ZN(n8193) );
  AOI21_X1 U9684 ( .B1(n8496), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8191), .ZN(
        n8192) );
  OAI211_X1 U9685 ( .C1(n8509), .C2(n9988), .A(n8193), .B(n8192), .ZN(P2_U3266) );
  NAND2_X1 U9686 ( .A1(n8477), .A2(n8195), .ZN(n8459) );
  INV_X1 U9687 ( .A(n8490), .ZN(n8196) );
  INV_X1 U9688 ( .A(n8580), .ZN(n8198) );
  NAND2_X1 U9689 ( .A1(n8570), .A2(n8200), .ZN(n8202) );
  NAND2_X1 U9690 ( .A1(n8385), .A2(n8203), .ZN(n8204) );
  INV_X1 U9691 ( .A(n8567), .ZN(n8395) );
  NAND2_X1 U9692 ( .A1(n8204), .A2(n4575), .ZN(n8369) );
  NAND2_X1 U9693 ( .A1(n8369), .A2(n8376), .ZN(n8207) );
  NAND2_X1 U9694 ( .A1(n8560), .A2(n8205), .ZN(n8206) );
  NAND2_X1 U9695 ( .A1(n8207), .A2(n8206), .ZN(n8353) );
  NAND2_X1 U9696 ( .A1(n8311), .A2(n8285), .ZN(n8210) );
  NAND2_X1 U9697 ( .A1(n8281), .A2(n8211), .ZN(n8214) );
  NAND2_X1 U9698 ( .A1(n8293), .A2(n8212), .ZN(n8213) );
  NAND2_X1 U9699 ( .A1(n8214), .A2(n8213), .ZN(n8263) );
  NOR2_X1 U9700 ( .A1(n8529), .A2(n8257), .ZN(n8215) );
  NAND2_X1 U9701 ( .A1(n8254), .A2(n8216), .ZN(n8217) );
  NAND2_X1 U9702 ( .A1(n4771), .A2(n8218), .ZN(n8219) );
  INV_X1 U9703 ( .A(n8510), .ZN(n8232) );
  XNOR2_X1 U9704 ( .A(n8220), .B(n8221), .ZN(n8225) );
  AOI22_X1 U9705 ( .A1(n8258), .A2(n8469), .B1(n8223), .B2(n8222), .ZN(n8224)
         );
  OAI21_X1 U9706 ( .B1(n8225), .B2(n8486), .A(n8224), .ZN(n8514) );
  OAI21_X1 U9707 ( .B1(n4519), .B2(n8511), .A(n8226), .ZN(n8512) );
  NOR2_X1 U9708 ( .A1(n8512), .A2(n9989), .ZN(n8230) );
  INV_X1 U9709 ( .A(n8451), .ZN(n9991) );
  AOI22_X1 U9710 ( .A1(n8227), .A2(n9991), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8289), .ZN(n8228) );
  OAI21_X1 U9711 ( .B1(n8511), .B2(n9988), .A(n8228), .ZN(n8229) );
  AOI211_X1 U9712 ( .C1(n8514), .C2(n9993), .A(n8230), .B(n8229), .ZN(n8231)
         );
  OAI21_X1 U9713 ( .B1(n8232), .B2(n8501), .A(n8231), .ZN(P2_U3267) );
  AOI21_X1 U9714 ( .B1(n8517), .B2(n8250), .A(n4519), .ZN(n8518) );
  AOI22_X1 U9715 ( .A1(n8235), .A2(n9991), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8289), .ZN(n8236) );
  OAI21_X1 U9716 ( .B1(n4771), .B2(n9988), .A(n8236), .ZN(n8237) );
  AOI21_X1 U9717 ( .B1(n8518), .B2(n8499), .A(n8237), .ZN(n8247) );
  NAND2_X1 U9718 ( .A1(n8240), .A2(n8471), .ZN(n8243) );
  NAND2_X1 U9719 ( .A1(n8241), .A2(n8469), .ZN(n8242) );
  OR2_X1 U9720 ( .A1(n8520), .A2(n8496), .ZN(n8246) );
  OAI211_X1 U9721 ( .C1(n8522), .C2(n8501), .A(n8247), .B(n8246), .ZN(P2_U3268) );
  XNOR2_X1 U9722 ( .A(n8248), .B(n8249), .ZN(n8527) );
  INV_X1 U9723 ( .A(n8250), .ZN(n8251) );
  AOI21_X1 U9724 ( .B1(n8523), .B2(n8272), .A(n8251), .ZN(n8524) );
  AOI22_X1 U9725 ( .A1(n8252), .A2(n9991), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8289), .ZN(n8253) );
  OAI21_X1 U9726 ( .B1(n8254), .B2(n9988), .A(n8253), .ZN(n8261) );
  XNOR2_X1 U9727 ( .A(n8255), .B(n8256), .ZN(n8259) );
  AOI222_X1 U9728 ( .A1(n10004), .A2(n8259), .B1(n8258), .B2(n8471), .C1(n8257), .C2(n8469), .ZN(n8526) );
  NOR2_X1 U9729 ( .A1(n8526), .A2(n8289), .ZN(n8260) );
  OAI21_X1 U9730 ( .B1(n8527), .B2(n8501), .A(n8262), .ZN(P2_U3269) );
  XOR2_X1 U9731 ( .A(n8264), .B(n8263), .Z(n8532) );
  AOI22_X1 U9732 ( .A1(n8529), .A2(n8455), .B1(n8496), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8280) );
  INV_X1 U9733 ( .A(n8265), .ZN(n8268) );
  OAI21_X1 U9734 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8270) );
  AOI21_X1 U9735 ( .B1(n8270), .B2(n10004), .A(n8269), .ZN(n8531) );
  INV_X1 U9736 ( .A(n8271), .ZN(n8274) );
  INV_X1 U9737 ( .A(n8272), .ZN(n8273) );
  AOI211_X1 U9738 ( .C1(n8529), .C2(n8274), .A(n10065), .B(n8273), .ZN(n8528)
         );
  NAND2_X1 U9739 ( .A1(n8528), .A2(n8275), .ZN(n8276) );
  OAI211_X1 U9740 ( .C1(n8451), .C2(n8277), .A(n8531), .B(n8276), .ZN(n8278)
         );
  NAND2_X1 U9741 ( .A1(n8278), .A2(n9993), .ZN(n8279) );
  OAI211_X1 U9742 ( .C1(n8532), .C2(n8501), .A(n8280), .B(n8279), .ZN(P2_U3270) );
  XNOR2_X1 U9743 ( .A(n8281), .B(n8283), .ZN(n8537) );
  XNOR2_X1 U9744 ( .A(n8282), .B(n8283), .ZN(n8284) );
  OAI222_X1 U9745 ( .A1(n8434), .A2(n8286), .B1(n8491), .B2(n8285), .C1(n8486), 
        .C2(n8284), .ZN(n8533) );
  XNOR2_X1 U9746 ( .A(n8307), .B(n8293), .ZN(n8287) );
  NOR2_X1 U9747 ( .A1(n8287), .A2(n10065), .ZN(n8534) );
  NAND2_X1 U9748 ( .A1(n8534), .A2(n8427), .ZN(n8292) );
  INV_X1 U9749 ( .A(n8288), .ZN(n8290) );
  AOI22_X1 U9750 ( .A1(n8290), .A2(n9991), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8289), .ZN(n8291) );
  OAI211_X1 U9751 ( .C1(n8293), .C2(n9988), .A(n8292), .B(n8291), .ZN(n8294)
         );
  AOI21_X1 U9752 ( .B1(n8533), .B2(n9993), .A(n8294), .ZN(n8295) );
  OAI21_X1 U9753 ( .B1(n8537), .B2(n8501), .A(n8295), .ZN(P2_U3271) );
  INV_X1 U9754 ( .A(n8296), .ZN(n8297) );
  AOI21_X1 U9755 ( .B1(n8301), .B2(n8298), .A(n8297), .ZN(n8542) );
  NAND2_X1 U9756 ( .A1(n8299), .A2(n10004), .ZN(n8306) );
  AOI21_X1 U9757 ( .B1(n8300), .B2(n8302), .A(n8301), .ZN(n8305) );
  INV_X1 U9758 ( .A(n8303), .ZN(n8304) );
  OAI21_X1 U9759 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(n8538) );
  AOI211_X1 U9760 ( .C1(n8540), .C2(n8320), .A(n10065), .B(n8307), .ZN(n8539)
         );
  NAND2_X1 U9761 ( .A1(n8539), .A2(n8427), .ZN(n8310) );
  AOI22_X1 U9762 ( .A1(n8308), .A2(n9991), .B1(n8496), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8309) );
  OAI211_X1 U9763 ( .C1(n8311), .C2(n9988), .A(n8310), .B(n8309), .ZN(n8312)
         );
  AOI21_X1 U9764 ( .B1(n8538), .B2(n9993), .A(n8312), .ZN(n8313) );
  OAI21_X1 U9765 ( .B1(n8542), .B2(n8501), .A(n8313), .ZN(P2_U3272) );
  OAI21_X1 U9766 ( .B1(n8340), .B2(n8315), .A(n8326), .ZN(n8316) );
  NAND2_X1 U9767 ( .A1(n8316), .A2(n8300), .ZN(n8319) );
  AOI222_X1 U9768 ( .A1(n10004), .A2(n8319), .B1(n8318), .B2(n8471), .C1(n8317), .C2(n8469), .ZN(n8548) );
  AOI21_X1 U9769 ( .B1(n8543), .B2(n8334), .A(n4777), .ZN(n8544) );
  INV_X1 U9770 ( .A(n8321), .ZN(n8322) );
  AOI22_X1 U9771 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n8496), .B1(n8322), .B2(
        n9991), .ZN(n8323) );
  OAI21_X1 U9772 ( .B1(n8324), .B2(n9988), .A(n8323), .ZN(n8325) );
  AOI21_X1 U9773 ( .B1(n8544), .B2(n8499), .A(n8325), .ZN(n8331) );
  OR2_X1 U9774 ( .A1(n8327), .A2(n8326), .ZN(n8545) );
  NAND3_X1 U9775 ( .A1(n8545), .A2(n8328), .A3(n8329), .ZN(n8330) );
  OAI211_X1 U9776 ( .C1(n8548), .C2(n8496), .A(n8331), .B(n8330), .ZN(P2_U3273) );
  XNOR2_X1 U9777 ( .A(n8333), .B(n8332), .ZN(n8553) );
  INV_X1 U9778 ( .A(n8360), .ZN(n8335) );
  AOI21_X1 U9779 ( .B1(n8549), .B2(n8335), .A(n4773), .ZN(n8550) );
  INV_X1 U9780 ( .A(n8336), .ZN(n8337) );
  AOI22_X1 U9781 ( .A1(n8496), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8337), .B2(
        n9991), .ZN(n8338) );
  OAI21_X1 U9782 ( .B1(n8339), .B2(n9988), .A(n8338), .ZN(n8351) );
  NOR2_X1 U9783 ( .A1(n8340), .A2(n8486), .ZN(n8349) );
  INV_X1 U9784 ( .A(n8341), .ZN(n8355) );
  INV_X1 U9785 ( .A(n8342), .ZN(n8344) );
  OAI21_X1 U9786 ( .B1(n8355), .B2(n8344), .A(n8343), .ZN(n8348) );
  OAI22_X1 U9787 ( .A1(n8346), .A2(n8434), .B1(n8345), .B2(n8491), .ZN(n8347)
         );
  AOI21_X1 U9788 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8552) );
  NOR2_X1 U9789 ( .A1(n8552), .A2(n8496), .ZN(n8350) );
  AOI211_X1 U9790 ( .C1(n8550), .C2(n8499), .A(n8351), .B(n8350), .ZN(n8352)
         );
  OAI21_X1 U9791 ( .B1(n8553), .B2(n8501), .A(n8352), .ZN(P2_U3274) );
  INV_X1 U9792 ( .A(n8353), .ZN(n8354) );
  XOR2_X1 U9793 ( .A(n8356), .B(n8354), .Z(n8559) );
  AOI21_X1 U9794 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8358) );
  OAI222_X1 U9795 ( .A1(n8434), .A2(n8359), .B1(n8491), .B2(n8392), .C1(n8486), 
        .C2(n8358), .ZN(n8554) );
  INV_X1 U9796 ( .A(n8370), .ZN(n8361) );
  AOI21_X1 U9797 ( .B1(n8555), .B2(n8361), .A(n8360), .ZN(n8556) );
  NAND2_X1 U9798 ( .A1(n8556), .A2(n8499), .ZN(n8365) );
  INV_X1 U9799 ( .A(n8362), .ZN(n8363) );
  AOI22_X1 U9800 ( .A1(n8496), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8363), .B2(
        n9991), .ZN(n8364) );
  OAI211_X1 U9801 ( .C1(n8366), .C2(n9988), .A(n8365), .B(n8364), .ZN(n8367)
         );
  AOI21_X1 U9802 ( .B1(n8554), .B2(n9993), .A(n8367), .ZN(n8368) );
  OAI21_X1 U9803 ( .B1(n8501), .B2(n8559), .A(n8368), .ZN(P2_U3275) );
  XNOR2_X1 U9804 ( .A(n8369), .B(n8376), .ZN(n8564) );
  AOI21_X1 U9805 ( .B1(n8560), .B2(n8393), .A(n8370), .ZN(n8561) );
  INV_X1 U9806 ( .A(n8371), .ZN(n8372) );
  AOI22_X1 U9807 ( .A1(n8496), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8372), .B2(
        n9991), .ZN(n8373) );
  OAI21_X1 U9808 ( .B1(n8374), .B2(n9988), .A(n8373), .ZN(n8382) );
  NOR2_X1 U9809 ( .A1(n8390), .A2(n4831), .ZN(n8377) );
  XNOR2_X1 U9810 ( .A(n8377), .B(n8376), .ZN(n8380) );
  AOI222_X1 U9811 ( .A1(n10004), .A2(n8380), .B1(n8379), .B2(n8471), .C1(n8378), .C2(n8469), .ZN(n8563) );
  NOR2_X1 U9812 ( .A1(n8563), .A2(n8496), .ZN(n8381) );
  AOI211_X1 U9813 ( .C1(n8561), .C2(n8499), .A(n8382), .B(n8381), .ZN(n8383)
         );
  OAI21_X1 U9814 ( .B1(n8501), .B2(n8564), .A(n8383), .ZN(P2_U3276) );
  XNOR2_X1 U9815 ( .A(n8385), .B(n8384), .ZN(n8569) );
  INV_X1 U9816 ( .A(n8409), .ZN(n8388) );
  AOI21_X1 U9817 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8389) );
  NOR2_X1 U9818 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  OAI222_X1 U9819 ( .A1(n8434), .A2(n8392), .B1(n8491), .B2(n8433), .C1(n8486), 
        .C2(n8391), .ZN(n8565) );
  NAND2_X1 U9820 ( .A1(n8565), .A2(n9993), .ZN(n8401) );
  INV_X1 U9821 ( .A(n8393), .ZN(n8394) );
  AOI211_X1 U9822 ( .C1(n8567), .C2(n8403), .A(n10065), .B(n8394), .ZN(n8566)
         );
  NOR2_X1 U9823 ( .A1(n8395), .A2(n9988), .ZN(n8399) );
  OAI22_X1 U9824 ( .A1(n9993), .A2(n8397), .B1(n8396), .B2(n8451), .ZN(n8398)
         );
  AOI211_X1 U9825 ( .C1(n8566), .C2(n8427), .A(n8399), .B(n8398), .ZN(n8400)
         );
  OAI211_X1 U9826 ( .C1(n8569), .C2(n8501), .A(n8401), .B(n8400), .ZN(P2_U3277) );
  XNOR2_X1 U9827 ( .A(n8402), .B(n4872), .ZN(n8574) );
  INV_X1 U9828 ( .A(n8421), .ZN(n8405) );
  INV_X1 U9829 ( .A(n8403), .ZN(n8404) );
  AOI21_X1 U9830 ( .B1(n8570), .B2(n8405), .A(n8404), .ZN(n8571) );
  AOI22_X1 U9831 ( .A1(n8496), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8406), .B2(
        n9991), .ZN(n8407) );
  OAI21_X1 U9832 ( .B1(n8408), .B2(n9988), .A(n8407), .ZN(n8416) );
  AOI211_X1 U9833 ( .C1(n8411), .C2(n8410), .A(n8486), .B(n8409), .ZN(n8414)
         );
  OAI22_X1 U9834 ( .A1(n8412), .A2(n8434), .B1(n8445), .B2(n8491), .ZN(n8413)
         );
  NOR2_X1 U9835 ( .A1(n8414), .A2(n8413), .ZN(n8573) );
  NOR2_X1 U9836 ( .A1(n8573), .A2(n8496), .ZN(n8415) );
  AOI211_X1 U9837 ( .C1(n8571), .C2(n8499), .A(n8416), .B(n8415), .ZN(n8417)
         );
  OAI21_X1 U9838 ( .B1(n8574), .B2(n8501), .A(n8417), .ZN(P2_U3278) );
  INV_X1 U9839 ( .A(n8418), .ZN(n8419) );
  AOI21_X1 U9840 ( .B1(n8430), .B2(n8420), .A(n8419), .ZN(n8579) );
  AOI211_X1 U9841 ( .C1(n8577), .C2(n8438), .A(n10065), .B(n8421), .ZN(n8576)
         );
  NOR2_X1 U9842 ( .A1(n8422), .A2(n9988), .ZN(n8426) );
  OAI22_X1 U9843 ( .A1(n9993), .A2(n8424), .B1(n8423), .B2(n8451), .ZN(n8425)
         );
  AOI211_X1 U9844 ( .C1(n8576), .C2(n8427), .A(n8426), .B(n8425), .ZN(n8437)
         );
  NOR2_X1 U9845 ( .A1(n8441), .A2(n8429), .ZN(n8431) );
  XNOR2_X1 U9846 ( .A(n8431), .B(n8430), .ZN(n8432) );
  OAI222_X1 U9847 ( .A1(n8491), .A2(n8435), .B1(n8434), .B2(n8433), .C1(n8432), 
        .C2(n8486), .ZN(n8575) );
  NAND2_X1 U9848 ( .A1(n8575), .A2(n9993), .ZN(n8436) );
  OAI211_X1 U9849 ( .C1(n8579), .C2(n8501), .A(n8437), .B(n8436), .ZN(P2_U3279) );
  INV_X1 U9850 ( .A(n8438), .ZN(n8439) );
  AOI21_X1 U9851 ( .B1(n8580), .B2(n8460), .A(n8439), .ZN(n8581) );
  INV_X1 U9852 ( .A(n8581), .ZN(n8458) );
  OAI21_X1 U9853 ( .B1(n4584), .B2(n8443), .A(n8440), .ZN(n8584) );
  INV_X1 U9854 ( .A(n8584), .ZN(n8448) );
  AOI21_X1 U9855 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8444) );
  NOR2_X1 U9856 ( .A1(n8444), .A2(n8486), .ZN(n8447) );
  OAI22_X1 U9857 ( .A1(n8490), .A2(n8491), .B1(n8445), .B2(n8434), .ZN(n8446)
         );
  AOI211_X1 U9858 ( .C1(n8448), .C2(n10061), .A(n8447), .B(n8446), .ZN(n8583)
         );
  OAI21_X1 U9859 ( .B1(n8449), .B2(n8584), .A(n8583), .ZN(n8450) );
  NAND2_X1 U9860 ( .A1(n8450), .A2(n9993), .ZN(n8457) );
  INV_X1 U9861 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8453) );
  OAI22_X1 U9862 ( .A1(n9993), .A2(n8453), .B1(n8452), .B2(n8451), .ZN(n8454)
         );
  AOI21_X1 U9863 ( .B1(n8580), .B2(n8455), .A(n8454), .ZN(n8456) );
  OAI211_X1 U9864 ( .C1(n8458), .C2(n9989), .A(n8457), .B(n8456), .ZN(P2_U3280) );
  XNOR2_X1 U9865 ( .A(n8459), .B(n8467), .ZN(n8589) );
  INV_X1 U9866 ( .A(n8460), .ZN(n8461) );
  AOI21_X1 U9867 ( .B1(n8585), .B2(n8462), .A(n8461), .ZN(n8586) );
  INV_X1 U9868 ( .A(n8463), .ZN(n8464) );
  AOI22_X1 U9869 ( .A1(n8496), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8464), .B2(
        n9991), .ZN(n8465) );
  OAI21_X1 U9870 ( .B1(n8466), .B2(n9988), .A(n8465), .ZN(n8475) );
  XNOR2_X1 U9871 ( .A(n8468), .B(n8467), .ZN(n8473) );
  AOI222_X1 U9872 ( .A1(n10004), .A2(n8473), .B1(n8472), .B2(n8471), .C1(n8470), .C2(n8469), .ZN(n8588) );
  NOR2_X1 U9873 ( .A1(n8588), .A2(n8496), .ZN(n8474) );
  AOI211_X1 U9874 ( .C1(n8586), .C2(n8499), .A(n8475), .B(n8474), .ZN(n8476)
         );
  OAI21_X1 U9875 ( .B1(n8589), .B2(n8501), .A(n8476), .ZN(P2_U3281) );
  INV_X1 U9876 ( .A(n8477), .ZN(n8478) );
  AOI21_X1 U9877 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n8594) );
  XNOR2_X1 U9878 ( .A(n8481), .B(n8590), .ZN(n8591) );
  INV_X1 U9879 ( .A(n8482), .ZN(n8483) );
  AOI22_X1 U9880 ( .A1(n8496), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8483), .B2(
        n9991), .ZN(n8484) );
  OAI21_X1 U9881 ( .B1(n8485), .B2(n9988), .A(n8484), .ZN(n8498) );
  NOR2_X1 U9882 ( .A1(n8487), .A2(n8486), .ZN(n8495) );
  OAI21_X1 U9883 ( .B1(n4572), .B2(n8489), .A(n8488), .ZN(n8494) );
  OAI22_X1 U9884 ( .A1(n8492), .A2(n8491), .B1(n8490), .B2(n8434), .ZN(n8493)
         );
  AOI21_X1 U9885 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(n8593) );
  NOR2_X1 U9886 ( .A1(n8593), .A2(n8496), .ZN(n8497) );
  AOI211_X1 U9887 ( .C1(n8591), .C2(n8499), .A(n8498), .B(n8497), .ZN(n8500)
         );
  OAI21_X1 U9888 ( .B1(n8594), .B2(n8501), .A(n8500), .ZN(P2_U3282) );
  NAND2_X1 U9889 ( .A1(n8502), .A2(n10073), .ZN(n8503) );
  OAI211_X1 U9890 ( .C1(n8504), .C2(n10065), .A(n8503), .B(n8507), .ZN(n8595)
         );
  MUX2_X1 U9891 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8595), .S(n10097), .Z(
        P2_U3551) );
  NAND3_X1 U9892 ( .A1(n8506), .A2(n10074), .A3(n8505), .ZN(n8508) );
  OAI211_X1 U9893 ( .C1(n8509), .C2(n10063), .A(n8508), .B(n8507), .ZN(n8596)
         );
  MUX2_X1 U9894 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8596), .S(n10097), .Z(
        P2_U3550) );
  NAND2_X1 U9895 ( .A1(n8510), .A2(n10069), .ZN(n8516) );
  OAI22_X1 U9896 ( .A1(n8512), .A2(n10065), .B1(n8511), .B2(n10063), .ZN(n8513) );
  NOR2_X1 U9897 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  NAND2_X1 U9898 ( .A1(n8516), .A2(n8515), .ZN(n8597) );
  MUX2_X1 U9899 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8597), .S(n10097), .Z(
        P2_U3549) );
  AOI22_X1 U9900 ( .A1(n8518), .A2(n10074), .B1(n10073), .B2(n8517), .ZN(n8519) );
  OAI21_X1 U9901 ( .B1(n8522), .B2(n10078), .A(n8521), .ZN(n8598) );
  MUX2_X1 U9902 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8598), .S(n10097), .Z(
        P2_U3548) );
  AOI22_X1 U9903 ( .A1(n8524), .A2(n10074), .B1(n10073), .B2(n8523), .ZN(n8525) );
  OAI211_X1 U9904 ( .C1(n8527), .C2(n10078), .A(n8526), .B(n8525), .ZN(n8599)
         );
  MUX2_X1 U9905 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8599), .S(n10097), .Z(
        P2_U3547) );
  AOI21_X1 U9906 ( .B1(n10073), .B2(n8529), .A(n8528), .ZN(n8530) );
  OAI211_X1 U9907 ( .C1(n8532), .C2(n10078), .A(n8531), .B(n8530), .ZN(n8600)
         );
  MUX2_X1 U9908 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8600), .S(n10097), .Z(
        P2_U3546) );
  AOI211_X1 U9909 ( .C1(n10073), .C2(n8535), .A(n8534), .B(n8533), .ZN(n8536)
         );
  OAI21_X1 U9910 ( .B1(n10078), .B2(n8537), .A(n8536), .ZN(n8601) );
  MUX2_X1 U9911 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8601), .S(n10097), .Z(
        P2_U3545) );
  AOI211_X1 U9912 ( .C1(n10073), .C2(n8540), .A(n8539), .B(n8538), .ZN(n8541)
         );
  OAI21_X1 U9913 ( .B1(n8542), .B2(n10078), .A(n8541), .ZN(n8602) );
  MUX2_X1 U9914 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8602), .S(n10097), .Z(
        P2_U3544) );
  AOI22_X1 U9915 ( .A1(n8544), .A2(n10074), .B1(n10073), .B2(n8543), .ZN(n8547) );
  NAND3_X1 U9916 ( .A1(n8545), .A2(n8328), .A3(n10069), .ZN(n8546) );
  NAND3_X1 U9917 ( .A1(n8548), .A2(n8547), .A3(n8546), .ZN(n8603) );
  MUX2_X1 U9918 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8603), .S(n10097), .Z(
        P2_U3543) );
  AOI22_X1 U9919 ( .A1(n8550), .A2(n10074), .B1(n10073), .B2(n8549), .ZN(n8551) );
  OAI211_X1 U9920 ( .C1(n8553), .C2(n10078), .A(n8552), .B(n8551), .ZN(n8604)
         );
  MUX2_X1 U9921 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8604), .S(n10097), .Z(
        P2_U3542) );
  INV_X1 U9922 ( .A(n8554), .ZN(n8558) );
  AOI22_X1 U9923 ( .A1(n8556), .A2(n10074), .B1(n10073), .B2(n8555), .ZN(n8557) );
  OAI211_X1 U9924 ( .C1(n10078), .C2(n8559), .A(n8558), .B(n8557), .ZN(n8605)
         );
  MUX2_X1 U9925 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8605), .S(n10097), .Z(
        P2_U3541) );
  AOI22_X1 U9926 ( .A1(n8561), .A2(n10074), .B1(n10073), .B2(n8560), .ZN(n8562) );
  OAI211_X1 U9927 ( .C1(n10078), .C2(n8564), .A(n8563), .B(n8562), .ZN(n8606)
         );
  MUX2_X1 U9928 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8606), .S(n10097), .Z(
        P2_U3540) );
  AOI211_X1 U9929 ( .C1(n10073), .C2(n8567), .A(n8566), .B(n8565), .ZN(n8568)
         );
  OAI21_X1 U9930 ( .B1(n10078), .B2(n8569), .A(n8568), .ZN(n8607) );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8607), .S(n10097), .Z(
        P2_U3539) );
  AOI22_X1 U9932 ( .A1(n8571), .A2(n10074), .B1(n10073), .B2(n8570), .ZN(n8572) );
  OAI211_X1 U9933 ( .C1(n10078), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8608)
         );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8608), .S(n10097), .Z(
        P2_U3538) );
  AOI211_X1 U9935 ( .C1(n10073), .C2(n8577), .A(n8576), .B(n8575), .ZN(n8578)
         );
  OAI21_X1 U9936 ( .B1(n8579), .B2(n10078), .A(n8578), .ZN(n8609) );
  MUX2_X1 U9937 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8609), .S(n10097), .Z(
        P2_U3537) );
  AOI22_X1 U9938 ( .A1(n8581), .A2(n10074), .B1(n10073), .B2(n8580), .ZN(n8582) );
  OAI211_X1 U9939 ( .C1(n10056), .C2(n8584), .A(n8583), .B(n8582), .ZN(n8610)
         );
  MUX2_X1 U9940 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8610), .S(n10097), .Z(
        P2_U3536) );
  AOI22_X1 U9941 ( .A1(n8586), .A2(n10074), .B1(n10073), .B2(n8585), .ZN(n8587) );
  OAI211_X1 U9942 ( .C1(n8589), .C2(n10078), .A(n8588), .B(n8587), .ZN(n8611)
         );
  MUX2_X1 U9943 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8611), .S(n10097), .Z(
        P2_U3535) );
  AOI22_X1 U9944 ( .A1(n8591), .A2(n10074), .B1(n10073), .B2(n8590), .ZN(n8592) );
  OAI211_X1 U9945 ( .C1(n8594), .C2(n10078), .A(n8593), .B(n8592), .ZN(n8612)
         );
  MUX2_X1 U9946 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8612), .S(n10097), .Z(
        P2_U3534) );
  MUX2_X1 U9947 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8595), .S(n10083), .Z(
        P2_U3519) );
  MUX2_X1 U9948 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8596), .S(n10083), .Z(
        P2_U3518) );
  MUX2_X1 U9949 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8597), .S(n10083), .Z(
        P2_U3517) );
  MUX2_X1 U9950 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8598), .S(n10083), .Z(
        P2_U3516) );
  MUX2_X1 U9951 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8599), .S(n10083), .Z(
        P2_U3515) );
  MUX2_X1 U9952 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8600), .S(n10083), .Z(
        P2_U3514) );
  MUX2_X1 U9953 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8601), .S(n10083), .Z(
        P2_U3513) );
  MUX2_X1 U9954 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8602), .S(n10083), .Z(
        P2_U3512) );
  MUX2_X1 U9955 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8603), .S(n10083), .Z(
        P2_U3511) );
  MUX2_X1 U9956 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8604), .S(n10083), .Z(
        P2_U3510) );
  MUX2_X1 U9957 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8605), .S(n10083), .Z(
        P2_U3509) );
  MUX2_X1 U9958 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8606), .S(n10083), .Z(
        P2_U3508) );
  MUX2_X1 U9959 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8607), .S(n10083), .Z(
        P2_U3507) );
  MUX2_X1 U9960 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8608), .S(n10083), .Z(
        P2_U3505) );
  MUX2_X1 U9961 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8609), .S(n10083), .Z(
        P2_U3502) );
  MUX2_X1 U9962 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8610), .S(n10083), .Z(
        P2_U3499) );
  MUX2_X1 U9963 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8611), .S(n10083), .Z(
        P2_U3496) );
  MUX2_X1 U9964 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8612), .S(n10083), .Z(
        P2_U3493) );
  INV_X1 U9965 ( .A(n8613), .ZN(n9592) );
  NOR4_X1 U9966 ( .A1(n6014), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6195), .A4(
        P2_U3152), .ZN(n8614) );
  AOI21_X1 U9967 ( .B1(n8623), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8614), .ZN(
        n8615) );
  OAI21_X1 U9968 ( .B1(n9592), .B2(n6488), .A(n8615), .ZN(P2_U3327) );
  INV_X1 U9969 ( .A(n8837), .ZN(n9594) );
  AOI22_X1 U9970 ( .A1(n8616), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8618), .ZN(n8617) );
  OAI21_X1 U9971 ( .B1(n9594), .B2(n6488), .A(n8617), .ZN(P2_U3328) );
  AOI22_X1 U9972 ( .A1(n8619), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8618), .ZN(n8620) );
  OAI21_X1 U9973 ( .B1(n8621), .B2(n6488), .A(n8620), .ZN(P2_U3329) );
  INV_X1 U9974 ( .A(n7719), .ZN(n9600) );
  AOI21_X1 U9975 ( .B1(n8623), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8622), .ZN(
        n8624) );
  OAI21_X1 U9976 ( .B1(n9600), .B2(n6488), .A(n8624), .ZN(P2_U3330) );
  MUX2_X1 U9977 ( .A(n8625), .B(n9960), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358)
         );
  XNOR2_X1 U9978 ( .A(n8628), .B(n8627), .ZN(n8629) );
  XNOR2_X1 U9979 ( .A(n8626), .B(n8629), .ZN(n8635) );
  INV_X1 U9980 ( .A(n9461), .ZN(n8811) );
  NAND2_X1 U9981 ( .A1(n8764), .A2(n9430), .ZN(n8632) );
  NOR2_X1 U9982 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8630), .ZN(n9758) );
  AOI21_X1 U9983 ( .B1(n8757), .B2(n9427), .A(n9758), .ZN(n8631) );
  OAI211_X1 U9984 ( .C1(n8811), .C2(n8755), .A(n8632), .B(n8631), .ZN(n8633)
         );
  AOI21_X1 U9985 ( .B1(n9150), .B2(n8770), .A(n8633), .ZN(n8634) );
  OAI21_X1 U9986 ( .B1(n8635), .B2(n8772), .A(n8634), .ZN(P1_U3213) );
  NAND2_X1 U9987 ( .A1(n8636), .A2(n8637), .ZN(n8638) );
  XOR2_X1 U9988 ( .A(n8639), .B(n8638), .Z(n8644) );
  NAND2_X1 U9989 ( .A1(n9266), .A2(n8757), .ZN(n8641) );
  INV_X1 U9990 ( .A(n9325), .ZN(n9162) );
  AOI22_X1 U9991 ( .A1(n9162), .A2(n8765), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8640) );
  OAI211_X1 U9992 ( .C1(n8733), .C2(n9297), .A(n8641), .B(n8640), .ZN(n8642)
         );
  AOI21_X1 U9993 ( .B1(n9522), .B2(n8770), .A(n8642), .ZN(n8643) );
  OAI21_X1 U9994 ( .B1(n8644), .B2(n8772), .A(n8643), .ZN(P1_U3214) );
  INV_X1 U9995 ( .A(n9542), .ZN(n9352) );
  INV_X1 U9996 ( .A(n8645), .ZN(n8649) );
  NOR3_X1 U9997 ( .A1(n8646), .A2(n8740), .A3(n8647), .ZN(n8648) );
  OAI21_X1 U9998 ( .B1(n8649), .B2(n8648), .A(n8751), .ZN(n8654) );
  INV_X1 U9999 ( .A(n9389), .ZN(n8782) );
  NOR2_X1 U10000 ( .A1(n8650), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9126) );
  AOI21_X1 U10001 ( .B1(n8757), .B2(n9358), .A(n9126), .ZN(n8651) );
  OAI21_X1 U10002 ( .B1(n8782), .B2(n8755), .A(n8651), .ZN(n8652) );
  AOI21_X1 U10003 ( .B1(n9350), .B2(n8764), .A(n8652), .ZN(n8653) );
  OAI211_X1 U10004 ( .C1(n9352), .C2(n8760), .A(n8654), .B(n8653), .ZN(
        P1_U3217) );
  AOI21_X1 U10005 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8663) );
  OAI22_X1 U10006 ( .A1(n9325), .A2(n8768), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8658), .ZN(n8659) );
  AOI21_X1 U10007 ( .B1(n8765), .B2(n9358), .A(n8659), .ZN(n8660) );
  OAI21_X1 U10008 ( .B1(n8733), .B2(n9321), .A(n8660), .ZN(n8661) );
  AOI21_X1 U10009 ( .B1(n9532), .B2(n8770), .A(n8661), .ZN(n8662) );
  OAI21_X1 U10010 ( .B1(n8663), .B2(n8772), .A(n8662), .ZN(P1_U3221) );
  INV_X1 U10011 ( .A(n9471), .ZN(n9663) );
  OAI21_X1 U10012 ( .B1(n8665), .B2(n4585), .A(n8664), .ZN(n8666) );
  NAND2_X1 U10013 ( .A1(n8666), .A2(n8751), .ZN(n8671) );
  NAND2_X1 U10014 ( .A1(n8757), .A2(n9461), .ZN(n8668) );
  OAI211_X1 U10015 ( .C1(n9143), .C2(n8755), .A(n8668), .B(n8667), .ZN(n8669)
         );
  AOI21_X1 U10016 ( .B1(n9467), .B2(n8764), .A(n8669), .ZN(n8670) );
  OAI211_X1 U10017 ( .C1(n9663), .C2(n8760), .A(n8671), .B(n8670), .ZN(
        P1_U3222) );
  OAI21_X1 U10018 ( .B1(n8674), .B2(n8672), .A(n8673), .ZN(n8675) );
  NAND2_X1 U10019 ( .A1(n8675), .A2(n8751), .ZN(n8680) );
  OAI22_X1 U10020 ( .A1(n9294), .A2(n8755), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8676), .ZN(n8678) );
  NOR2_X1 U10021 ( .A1(n9167), .A2(n8768), .ZN(n8677) );
  AOI211_X1 U10022 ( .C1(n9270), .C2(n8764), .A(n8678), .B(n8677), .ZN(n8679)
         );
  OAI211_X1 U10023 ( .C1(n9261), .C2(n8760), .A(n8680), .B(n8679), .ZN(
        P1_U3223) );
  INV_X1 U10024 ( .A(n9561), .ZN(n9399) );
  INV_X1 U10025 ( .A(n8681), .ZN(n8686) );
  AOI21_X1 U10026 ( .B1(n8684), .B2(n8682), .A(n8683), .ZN(n8685) );
  OAI21_X1 U10027 ( .B1(n8686), .B2(n8685), .A(n8751), .ZN(n8690) );
  INV_X1 U10028 ( .A(n9427), .ZN(n8821) );
  AOI22_X1 U10029 ( .A1(n8757), .A2(n9403), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8687) );
  OAI21_X1 U10030 ( .B1(n8821), .B2(n8755), .A(n8687), .ZN(n8688) );
  AOI21_X1 U10031 ( .B1(n9397), .B2(n8764), .A(n8688), .ZN(n8689) );
  OAI211_X1 U10032 ( .C1(n9399), .C2(n8760), .A(n8690), .B(n8689), .ZN(
        P1_U3224) );
  INV_X1 U10033 ( .A(n9555), .ZN(n9385) );
  OAI21_X1 U10034 ( .B1(n8693), .B2(n8691), .A(n8692), .ZN(n8694) );
  NAND2_X1 U10035 ( .A1(n8694), .A2(n8751), .ZN(n8698) );
  INV_X1 U10036 ( .A(n9419), .ZN(n8820) );
  NAND2_X1 U10037 ( .A1(n8757), .A2(n9389), .ZN(n8695) );
  NAND2_X1 U10038 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9800) );
  OAI211_X1 U10039 ( .C1(n8820), .C2(n8755), .A(n8695), .B(n9800), .ZN(n8696)
         );
  AOI21_X1 U10040 ( .B1(n9383), .B2(n8764), .A(n8696), .ZN(n8697) );
  OAI211_X1 U10041 ( .C1(n9385), .C2(n8760), .A(n8698), .B(n8697), .ZN(
        P1_U3226) );
  INV_X1 U10042 ( .A(n8699), .ZN(n8703) );
  AOI21_X1 U10043 ( .B1(n8636), .B2(n8701), .A(n8700), .ZN(n8702) );
  OAI21_X1 U10044 ( .B1(n8703), .B2(n8702), .A(n8751), .ZN(n8707) );
  AOI22_X1 U10045 ( .A1(n9313), .A2(n8765), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8704) );
  OAI21_X1 U10046 ( .B1(n8733), .B2(n9283), .A(n8704), .ZN(n8705) );
  AOI21_X1 U10047 ( .B1(n9254), .B2(n8757), .A(n8705), .ZN(n8706) );
  OAI211_X1 U10048 ( .C1(n9287), .C2(n8760), .A(n8707), .B(n8706), .ZN(
        P1_U3227) );
  INV_X1 U10049 ( .A(n9537), .ZN(n9339) );
  AND3_X1 U10050 ( .A1(n8645), .A2(n8710), .A3(n8709), .ZN(n8711) );
  OAI21_X1 U10051 ( .B1(n8708), .B2(n8711), .A(n8751), .ZN(n8716) );
  OAI22_X1 U10052 ( .A1(n9160), .A2(n8768), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8712), .ZN(n8714) );
  NOR2_X1 U10053 ( .A1(n8733), .A2(n9336), .ZN(n8713) );
  AOI211_X1 U10054 ( .C1(n8765), .C2(n9369), .A(n8714), .B(n8713), .ZN(n8715)
         );
  OAI211_X1 U10055 ( .C1(n9339), .C2(n8760), .A(n8716), .B(n8715), .ZN(
        P1_U3231) );
  XNOR2_X1 U10056 ( .A(n8719), .B(n8718), .ZN(n8720) );
  XNOR2_X1 U10057 ( .A(n8717), .B(n8720), .ZN(n8725) );
  NAND2_X1 U10058 ( .A1(n8764), .A2(n9451), .ZN(n8722) );
  AND2_X1 U10059 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9745) );
  AOI21_X1 U10060 ( .B1(n8757), .B2(n9418), .A(n9745), .ZN(n8721) );
  OAI211_X1 U10061 ( .C1(n9448), .C2(n8755), .A(n8722), .B(n8721), .ZN(n8723)
         );
  AOI21_X1 U10062 ( .B1(n9452), .B2(n8770), .A(n8723), .ZN(n8724) );
  OAI21_X1 U10063 ( .B1(n8725), .B2(n8772), .A(n8724), .ZN(P1_U3232) );
  NAND2_X1 U10064 ( .A1(n5108), .A2(n8726), .ZN(n8728) );
  XNOR2_X1 U10065 ( .A(n8728), .B(n8727), .ZN(n8736) );
  OAI22_X1 U10066 ( .A1(n9160), .A2(n8755), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8729), .ZN(n8730) );
  AOI21_X1 U10067 ( .B1(n8757), .B2(n9313), .A(n8730), .ZN(n8731) );
  OAI21_X1 U10068 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8734) );
  AOI21_X1 U10069 ( .B1(n9525), .B2(n8770), .A(n8734), .ZN(n8735) );
  OAI21_X1 U10070 ( .B1(n8736), .B2(n8772), .A(n8735), .ZN(P1_U3233) );
  INV_X1 U10071 ( .A(n8646), .ZN(n8741) );
  OAI21_X1 U10072 ( .B1(n8738), .B2(n8740), .A(n8737), .ZN(n8739) );
  OAI21_X1 U10073 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8742) );
  NAND2_X1 U10074 ( .A1(n8742), .A2(n8751), .ZN(n8746) );
  INV_X1 U10075 ( .A(n9403), .ZN(n8788) );
  NAND2_X1 U10076 ( .A1(n8757), .A2(n9369), .ZN(n8743) );
  NAND2_X1 U10077 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9815) );
  OAI211_X1 U10078 ( .C1(n8788), .C2(n8755), .A(n8743), .B(n9815), .ZN(n8744)
         );
  AOI21_X1 U10079 ( .B1(n9373), .B2(n8764), .A(n8744), .ZN(n8745) );
  OAI211_X1 U10080 ( .C1(n4707), .C2(n8760), .A(n8746), .B(n8745), .ZN(
        P1_U3236) );
  NOR2_X1 U10081 ( .A1(n8749), .A2(n4728), .ZN(n8750) );
  XNOR2_X1 U10082 ( .A(n8747), .B(n8750), .ZN(n8752) );
  NAND2_X1 U10083 ( .A1(n8752), .A2(n8751), .ZN(n8759) );
  INV_X1 U10084 ( .A(n9168), .ZN(n9255) );
  INV_X1 U10085 ( .A(n8753), .ZN(n9249) );
  AOI22_X1 U10086 ( .A1(n9249), .A2(n8764), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8754) );
  OAI21_X1 U10087 ( .B1(n9279), .B2(n8755), .A(n8754), .ZN(n8756) );
  AOI21_X1 U10088 ( .B1(n9255), .B2(n8757), .A(n8756), .ZN(n8758) );
  OAI211_X1 U10089 ( .C1(n9251), .C2(n8760), .A(n8759), .B(n8758), .ZN(
        P1_U3238) );
  NAND2_X1 U10090 ( .A1(n8682), .A2(n8761), .ZN(n8762) );
  XOR2_X1 U10091 ( .A(n8763), .B(n8762), .Z(n8773) );
  NAND2_X1 U10092 ( .A1(n8764), .A2(n9411), .ZN(n8767) );
  AND2_X1 U10093 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9774) );
  AOI21_X1 U10094 ( .B1(n8765), .B2(n9418), .A(n9774), .ZN(n8766) );
  OAI211_X1 U10095 ( .C1(n8820), .C2(n8768), .A(n8767), .B(n8766), .ZN(n8769)
         );
  AOI21_X1 U10096 ( .B1(n9565), .B2(n8770), .A(n8769), .ZN(n8771) );
  OAI21_X1 U10097 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(P1_U3239) );
  NAND2_X1 U10098 ( .A1(n8774), .A2(n8848), .ZN(n8776) );
  NAND2_X1 U10099 ( .A1(n8838), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8775) );
  INV_X1 U10100 ( .A(n9227), .ZN(n8973) );
  OR2_X1 U10101 ( .A1(n9492), .A2(n8973), .ZN(n8777) );
  NAND2_X1 U10102 ( .A1(n8777), .A2(n8961), .ZN(n9047) );
  NAND2_X1 U10103 ( .A1(n9522), .A2(n9280), .ZN(n8943) );
  INV_X1 U10104 ( .A(n8943), .ZN(n8778) );
  NAND2_X1 U10105 ( .A1(n9511), .A2(n9279), .ZN(n8983) );
  NAND2_X1 U10106 ( .A1(n9525), .A2(n9325), .ZN(n8985) );
  INV_X1 U10107 ( .A(n9358), .ZN(n9324) );
  NAND2_X1 U10108 ( .A1(n9537), .A2(n9324), .ZN(n8988) );
  INV_X1 U10109 ( .A(n8988), .ZN(n8779) );
  NAND2_X1 U10110 ( .A1(n8987), .A2(n8779), .ZN(n8780) );
  NAND2_X1 U10111 ( .A1(n9532), .A2(n9160), .ZN(n8986) );
  AND2_X1 U10112 ( .A1(n8780), .A2(n8986), .ZN(n8781) );
  AND2_X1 U10113 ( .A1(n8985), .A2(n8781), .ZN(n8935) );
  INV_X1 U10114 ( .A(n8935), .ZN(n8784) );
  INV_X1 U10115 ( .A(n9369), .ZN(n9157) );
  NAND2_X1 U10116 ( .A1(n9542), .A2(n9157), .ZN(n9188) );
  INV_X1 U10117 ( .A(n9188), .ZN(n9340) );
  OR2_X1 U10118 ( .A1(n8784), .A2(n9340), .ZN(n9038) );
  OR2_X1 U10119 ( .A1(n9555), .A2(n8788), .ZN(n9183) );
  NAND2_X1 U10120 ( .A1(n9187), .A2(n9183), .ZN(n8860) );
  NAND2_X1 U10121 ( .A1(n9548), .A2(n8782), .ZN(n8990) );
  NAND2_X1 U10122 ( .A1(n8860), .A2(n8990), .ZN(n8787) );
  OR2_X1 U10123 ( .A1(n9542), .A2(n9157), .ZN(n8989) );
  AND2_X1 U10124 ( .A1(n9189), .A2(n8989), .ZN(n8929) );
  AND2_X1 U10125 ( .A1(n8987), .A2(n8929), .ZN(n8783) );
  NAND2_X1 U10126 ( .A1(n9301), .A2(n9313), .ZN(n9194) );
  OAI211_X1 U10127 ( .C1(n8784), .C2(n8783), .A(n9194), .B(n9191), .ZN(n8785)
         );
  INV_X1 U10128 ( .A(n8785), .ZN(n8786) );
  OAI211_X1 U10129 ( .C1(n9038), .C2(n8787), .A(n8942), .B(n8786), .ZN(n9040)
         );
  NAND2_X1 U10130 ( .A1(n9555), .A2(n8788), .ZN(n8921) );
  NAND2_X1 U10131 ( .A1(n8990), .A2(n8921), .ZN(n8861) );
  NAND2_X1 U10132 ( .A1(n9561), .A2(n8820), .ZN(n9386) );
  INV_X1 U10133 ( .A(n9386), .ZN(n9182) );
  INV_X1 U10134 ( .A(n9418), .ZN(n9449) );
  NAND2_X1 U10135 ( .A1(n9150), .A2(n9449), .ZN(n8908) );
  NAND2_X1 U10136 ( .A1(n9452), .A2(n8811), .ZN(n9179) );
  AND2_X1 U10137 ( .A1(n8908), .A2(n9179), .ZN(n8914) );
  INV_X1 U10138 ( .A(n8914), .ZN(n8792) );
  NAND2_X1 U10139 ( .A1(n9471), .A2(n9448), .ZN(n8992) );
  INV_X1 U10140 ( .A(n8992), .ZN(n8791) );
  NAND2_X1 U10141 ( .A1(n9171), .A2(n8896), .ZN(n8892) );
  NAND2_X1 U10142 ( .A1(n8892), .A2(n9172), .ZN(n8789) );
  NAND2_X1 U10143 ( .A1(n9643), .A2(n9143), .ZN(n8905) );
  NAND2_X1 U10144 ( .A1(n8789), .A2(n8905), .ZN(n8790) );
  OR3_X1 U10145 ( .A1(n8792), .A2(n8791), .A3(n8790), .ZN(n8817) );
  INV_X1 U10146 ( .A(n8817), .ZN(n8793) );
  NAND2_X1 U10147 ( .A1(n9565), .A2(n8821), .ZN(n9181) );
  NAND4_X1 U10148 ( .A1(n8793), .A2(n9181), .A3(n8895), .A4(n8877), .ZN(n8794)
         );
  OR3_X1 U10149 ( .A1(n8861), .A2(n9182), .A3(n8794), .ZN(n9035) );
  INV_X1 U10150 ( .A(n8795), .ZN(n8797) );
  NAND2_X1 U10151 ( .A1(n4480), .A2(n6801), .ZN(n8796) );
  NAND3_X1 U10152 ( .A1(n8797), .A2(n8979), .A3(n8796), .ZN(n8798) );
  NAND2_X1 U10153 ( .A1(n8799), .A2(n8798), .ZN(n8801) );
  OAI21_X1 U10154 ( .B1(n8802), .B2(n8801), .A(n8800), .ZN(n8803) );
  NAND2_X1 U10155 ( .A1(n8803), .A2(n9026), .ZN(n8805) );
  NAND3_X1 U10156 ( .A1(n8805), .A2(n8804), .A3(n9028), .ZN(n8808) );
  INV_X1 U10157 ( .A(n9025), .ZN(n8874) );
  NOR2_X1 U10158 ( .A1(n9030), .A2(n8874), .ZN(n8807) );
  NAND2_X1 U10159 ( .A1(n8806), .A2(n8864), .ZN(n9031) );
  AOI21_X1 U10160 ( .B1(n8808), .B2(n8807), .A(n9031), .ZN(n8824) );
  INV_X1 U10161 ( .A(n8809), .ZN(n8810) );
  NOR2_X1 U10162 ( .A1(n8894), .A2(n8810), .ZN(n8893) );
  INV_X1 U10163 ( .A(n9150), .ZN(n9650) );
  AND2_X1 U10164 ( .A1(n9650), .A2(n9418), .ZN(n9415) );
  INV_X1 U10165 ( .A(n9415), .ZN(n8816) );
  OR2_X1 U10166 ( .A1(n9452), .A2(n8811), .ZN(n8991) );
  NAND2_X1 U10167 ( .A1(n9443), .A2(n9174), .ZN(n8812) );
  NAND2_X1 U10168 ( .A1(n8812), .A2(n8992), .ZN(n8813) );
  AND2_X1 U10169 ( .A1(n8991), .A2(n8813), .ZN(n8912) );
  INV_X1 U10170 ( .A(n8912), .ZN(n8814) );
  NAND2_X1 U10171 ( .A1(n8914), .A2(n8814), .ZN(n8815) );
  OAI211_X1 U10172 ( .C1(n8817), .C2(n8893), .A(n8816), .B(n8815), .ZN(n8819)
         );
  NOR2_X1 U10173 ( .A1(n8817), .A2(n9172), .ZN(n8818) );
  OAI21_X1 U10174 ( .B1(n8819), .B2(n8818), .A(n9181), .ZN(n8822) );
  OR2_X1 U10175 ( .A1(n9561), .A2(n8820), .ZN(n8922) );
  OR2_X1 U10176 ( .A1(n9565), .A2(n8821), .ZN(n8918) );
  AND3_X1 U10177 ( .A1(n8822), .A2(n8922), .A3(n8918), .ZN(n8823) );
  OR3_X1 U10178 ( .A1(n8861), .A2(n9182), .A3(n8823), .ZN(n9033) );
  OAI21_X1 U10179 ( .B1(n9035), .B2(n8824), .A(n9033), .ZN(n8825) );
  INV_X1 U10180 ( .A(n8825), .ZN(n8826) );
  NOR2_X1 U10181 ( .A1(n9038), .A2(n8826), .ZN(n8827) );
  NOR2_X1 U10182 ( .A1(n9040), .A2(n8827), .ZN(n8828) );
  NOR2_X1 U10183 ( .A1(n9042), .A2(n8828), .ZN(n8830) );
  AND2_X1 U10184 ( .A1(n9196), .A2(n8984), .ZN(n9041) );
  INV_X1 U10185 ( .A(n9041), .ZN(n8829) );
  OR3_X1 U10186 ( .A1(n9238), .A2(n8830), .A3(n8829), .ZN(n8831) );
  NOR2_X1 U10187 ( .A1(n9047), .A2(n8831), .ZN(n8846) );
  NAND2_X1 U10188 ( .A1(n9495), .A2(n9203), .ZN(n9198) );
  OAI21_X1 U10189 ( .B1(n9251), .B2(n9265), .A(n8958), .ZN(n8832) );
  NAND2_X1 U10190 ( .A1(n8832), .A2(n9221), .ZN(n8833) );
  AND2_X1 U10191 ( .A1(n9198), .A2(n8833), .ZN(n8834) );
  OR2_X1 U10192 ( .A1(n9047), .A2(n8834), .ZN(n8836) );
  NAND2_X1 U10193 ( .A1(n9492), .A2(n8973), .ZN(n8835) );
  AND2_X1 U10194 ( .A1(n8836), .A2(n8835), .ZN(n9044) );
  INV_X1 U10195 ( .A(n9044), .ZN(n8845) );
  NAND2_X1 U10196 ( .A1(n8837), .A2(n8848), .ZN(n8840) );
  NAND2_X1 U10197 ( .A1(n8838), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U10198 ( .A1(n5278), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U10199 ( .A1(n8851), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U10200 ( .A1(n8841), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8842) );
  AND3_X1 U10201 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n9201) );
  OR2_X1 U10202 ( .A1(n9486), .A2(n9201), .ZN(n9019) );
  OAI21_X1 U10203 ( .B1(n8846), .B2(n8845), .A(n9019), .ZN(n8847) );
  NAND2_X1 U10204 ( .A1(n9486), .A2(n9201), .ZN(n9018) );
  NAND2_X1 U10205 ( .A1(n8847), .A2(n9018), .ZN(n8855) );
  NAND2_X1 U10206 ( .A1(n8613), .A2(n8848), .ZN(n8850) );
  NAND2_X1 U10207 ( .A1(n8838), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U10208 ( .A1(n5278), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U10209 ( .A1(n8851), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U10210 ( .A1(n4482), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8852) );
  NAND3_X1 U10211 ( .A1(n8854), .A2(n8853), .A3(n8852), .ZN(n9069) );
  INV_X1 U10212 ( .A(n9069), .ZN(n9133) );
  NAND2_X1 U10213 ( .A1(n9482), .A2(n9133), .ZN(n9021) );
  NAND2_X1 U10214 ( .A1(n8855), .A2(n9021), .ZN(n8856) );
  OR2_X1 U10215 ( .A1(n9482), .A2(n9133), .ZN(n9022) );
  NAND2_X1 U10216 ( .A1(n8856), .A2(n9022), .ZN(n8857) );
  XNOR2_X1 U10217 ( .A(n8857), .B(n9327), .ZN(n9059) );
  NAND2_X1 U10218 ( .A1(n9019), .A2(n9069), .ZN(n8858) );
  NAND2_X1 U10219 ( .A1(n8858), .A2(n9482), .ZN(n9049) );
  INV_X1 U10220 ( .A(n9201), .ZN(n9070) );
  NAND2_X1 U10221 ( .A1(n9070), .A2(n9069), .ZN(n8859) );
  NAND2_X1 U10222 ( .A1(n9486), .A2(n8859), .ZN(n9045) );
  MUX2_X1 U10223 ( .A(n8861), .B(n8860), .S(n8969), .Z(n8862) );
  INV_X1 U10224 ( .A(n8862), .ZN(n8926) );
  AND4_X1 U10225 ( .A1(n8864), .A2(n8873), .A3(n8863), .A4(n8969), .ZN(n8865)
         );
  OAI21_X1 U10226 ( .B1(n9864), .B2(n8866), .A(n8865), .ZN(n8888) );
  NAND2_X1 U10227 ( .A1(n9868), .A2(n8969), .ZN(n8867) );
  INV_X1 U10228 ( .A(n8969), .ZN(n8971) );
  OAI22_X1 U10229 ( .A1(n8867), .A2(n9913), .B1(n8971), .B2(n9073), .ZN(n8871)
         );
  OAI21_X1 U10230 ( .B1(n8867), .B2(n9073), .A(n8882), .ZN(n8870) );
  NAND2_X1 U10231 ( .A1(n9074), .A2(n8971), .ZN(n8883) );
  OAI21_X1 U10232 ( .B1(n8883), .B2(n8868), .A(n9913), .ZN(n8869) );
  AOI22_X1 U10233 ( .A1(n8872), .A2(n8871), .B1(n8870), .B2(n8869), .ZN(n8887)
         );
  OAI211_X1 U10234 ( .C1(n8875), .C2(n8874), .A(n9028), .B(n8873), .ZN(n8880)
         );
  AND2_X1 U10235 ( .A1(n8876), .A2(n8971), .ZN(n8879) );
  NAND4_X1 U10236 ( .A1(n8880), .A2(n8879), .A3(n8878), .A4(n8877), .ZN(n8886)
         );
  NAND2_X1 U10237 ( .A1(n9073), .A2(n8971), .ZN(n8881) );
  OAI21_X1 U10238 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8884) );
  NAND2_X1 U10239 ( .A1(n8884), .A2(n9920), .ZN(n8885) );
  NAND4_X1 U10240 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n8891)
         );
  INV_X1 U10241 ( .A(n8896), .ZN(n8889) );
  NOR2_X1 U10242 ( .A1(n8889), .A2(n8894), .ZN(n9836) );
  AND2_X1 U10243 ( .A1(n4494), .A2(n8890), .ZN(n9002) );
  NAND3_X1 U10244 ( .A1(n8891), .A2(n9836), .A3(n9002), .ZN(n8904) );
  OAI211_X1 U10245 ( .C1(n8893), .C2(n8892), .A(n9443), .B(n9172), .ZN(n8901)
         );
  INV_X1 U10246 ( .A(n8894), .ZN(n8898) );
  NAND2_X1 U10247 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  NAND3_X1 U10248 ( .A1(n8898), .A2(n9172), .A3(n8897), .ZN(n8899) );
  NAND2_X1 U10249 ( .A1(n8899), .A2(n9171), .ZN(n8900) );
  MUX2_X1 U10250 ( .A(n8901), .B(n8900), .S(n8969), .Z(n8902) );
  INV_X1 U10251 ( .A(n8902), .ZN(n8903) );
  NAND4_X1 U10252 ( .A1(n8904), .A2(n9630), .A3(n8992), .A4(n8903), .ZN(n8913)
         );
  NAND2_X1 U10253 ( .A1(n8992), .A2(n8905), .ZN(n8906) );
  NAND2_X1 U10254 ( .A1(n8906), .A2(n9443), .ZN(n8907) );
  NAND3_X1 U10255 ( .A1(n8913), .A2(n8914), .A3(n8907), .ZN(n8911) );
  INV_X1 U10256 ( .A(n8991), .ZN(n8909) );
  OAI21_X1 U10257 ( .B1(n9415), .B2(n8909), .A(n8908), .ZN(n8910) );
  NAND2_X1 U10258 ( .A1(n8911), .A2(n8910), .ZN(n8917) );
  NAND2_X1 U10259 ( .A1(n8913), .A2(n8912), .ZN(n8915) );
  AOI21_X1 U10260 ( .B1(n8915), .B2(n8914), .A(n9415), .ZN(n8916) );
  MUX2_X1 U10261 ( .A(n8917), .B(n8916), .S(n8969), .Z(n8920) );
  NAND2_X1 U10262 ( .A1(n8918), .A2(n9181), .ZN(n9414) );
  NAND2_X1 U10263 ( .A1(n8922), .A2(n9386), .ZN(n9395) );
  INV_X1 U10264 ( .A(n9395), .ZN(n9402) );
  MUX2_X1 U10265 ( .A(n8918), .B(n9181), .S(n8971), .Z(n8919) );
  OAI211_X1 U10266 ( .C1(n8920), .C2(n9414), .A(n9402), .B(n8919), .ZN(n8924)
         );
  NAND2_X1 U10267 ( .A1(n9183), .A2(n8921), .ZN(n9380) );
  INV_X1 U10268 ( .A(n9380), .ZN(n9387) );
  MUX2_X1 U10269 ( .A(n8922), .B(n9386), .S(n8969), .Z(n8923) );
  NAND3_X1 U10270 ( .A1(n8924), .A2(n9387), .A3(n8923), .ZN(n8925) );
  NAND2_X1 U10271 ( .A1(n8926), .A2(n8925), .ZN(n8928) );
  NAND3_X1 U10272 ( .A1(n8928), .A2(n9187), .A3(n8989), .ZN(n8927) );
  NAND3_X1 U10273 ( .A1(n8927), .A2(n9188), .A3(n8988), .ZN(n8932) );
  NAND3_X1 U10274 ( .A1(n8928), .A2(n8990), .A3(n9188), .ZN(n8930) );
  NAND2_X1 U10275 ( .A1(n8930), .A2(n8929), .ZN(n8931) );
  MUX2_X1 U10276 ( .A(n8932), .B(n8931), .S(n8969), .Z(n8937) );
  INV_X1 U10277 ( .A(n8986), .ZN(n9310) );
  AOI21_X1 U10278 ( .B1(n8937), .B2(n9189), .A(n9310), .ZN(n8934) );
  NAND2_X1 U10279 ( .A1(n9191), .A2(n8987), .ZN(n8933) );
  OAI21_X1 U10280 ( .B1(n8934), .B2(n8933), .A(n8985), .ZN(n8940) );
  INV_X1 U10281 ( .A(n8987), .ZN(n8936) );
  OAI21_X1 U10282 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8938) );
  NAND2_X1 U10283 ( .A1(n8938), .A2(n9191), .ZN(n8939) );
  MUX2_X1 U10284 ( .A(n8940), .B(n8939), .S(n8969), .Z(n8945) );
  NAND2_X1 U10285 ( .A1(n9194), .A2(n8943), .ZN(n9291) );
  NOR2_X1 U10286 ( .A1(n9277), .A2(n9291), .ZN(n8944) );
  NAND2_X1 U10287 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NAND2_X1 U10288 ( .A1(n4545), .A2(n8946), .ZN(n8955) );
  OAI22_X1 U10289 ( .A1(n8955), .A2(n9505), .B1(n8971), .B2(n8983), .ZN(n8947)
         );
  NAND2_X1 U10290 ( .A1(n8947), .A2(n9167), .ZN(n8950) );
  AOI21_X1 U10291 ( .B1(n9251), .B2(n9195), .A(n9265), .ZN(n8948) );
  MUX2_X1 U10292 ( .A(n9251), .B(n8948), .S(n8971), .Z(n8949) );
  NAND2_X1 U10293 ( .A1(n8950), .A2(n8949), .ZN(n8957) );
  OAI21_X1 U10294 ( .B1(n9195), .B2(n9251), .A(n8958), .ZN(n8953) );
  NAND2_X1 U10295 ( .A1(n8983), .A2(n9265), .ZN(n8951) );
  NAND2_X1 U10296 ( .A1(n9221), .A2(n8951), .ZN(n8952) );
  MUX2_X1 U10297 ( .A(n8953), .B(n8952), .S(n8969), .Z(n8954) );
  OAI21_X1 U10298 ( .B1(n8955), .B2(n9238), .A(n8954), .ZN(n8956) );
  NAND2_X1 U10299 ( .A1(n8957), .A2(n8956), .ZN(n8960) );
  INV_X1 U10300 ( .A(n9222), .ZN(n9197) );
  MUX2_X1 U10301 ( .A(n8958), .B(n9221), .S(n8971), .Z(n8959) );
  NAND3_X1 U10302 ( .A1(n8960), .A2(n9197), .A3(n8959), .ZN(n8963) );
  MUX2_X1 U10303 ( .A(n9198), .B(n8961), .S(n8969), .Z(n8962) );
  AND2_X1 U10304 ( .A1(n8963), .A2(n8962), .ZN(n8972) );
  NAND3_X1 U10305 ( .A1(n9045), .A2(n8972), .A3(n9227), .ZN(n8964) );
  AND2_X1 U10306 ( .A1(n9049), .A2(n8964), .ZN(n8968) );
  NAND3_X1 U10307 ( .A1(n9049), .A2(n8972), .A3(n9492), .ZN(n8965) );
  NAND2_X1 U10308 ( .A1(n8965), .A2(n9045), .ZN(n8966) );
  NAND2_X1 U10309 ( .A1(n8966), .A2(n9021), .ZN(n8967) );
  MUX2_X1 U10310 ( .A(n8968), .B(n8967), .S(n8969), .Z(n8978) );
  AND2_X1 U10311 ( .A1(n9227), .A2(n8969), .ZN(n8970) );
  AOI21_X1 U10312 ( .B1(n9492), .B2(n8971), .A(n8970), .ZN(n8976) );
  INV_X1 U10313 ( .A(n8972), .ZN(n8974) );
  NAND3_X1 U10314 ( .A1(n8974), .A2(n9209), .A3(n8973), .ZN(n8975) );
  NAND4_X1 U10315 ( .A1(n9049), .A2(n8976), .A3(n8975), .A4(n9045), .ZN(n8977)
         );
  NAND2_X1 U10316 ( .A1(n8978), .A2(n8977), .ZN(n9058) );
  AND2_X1 U10317 ( .A1(n9022), .A2(n8979), .ZN(n9051) );
  INV_X1 U10318 ( .A(n9051), .ZN(n8981) );
  OR2_X1 U10319 ( .A1(n8981), .A2(n8980), .ZN(n9057) );
  NAND3_X1 U10320 ( .A1(n9058), .A2(n9051), .A3(n8982), .ZN(n9056) );
  INV_X1 U10321 ( .A(n9263), .ZN(n9013) );
  INV_X1 U10322 ( .A(n9277), .ZN(n9012) );
  NAND2_X1 U10323 ( .A1(n9191), .A2(n8985), .ZN(n9311) );
  NAND2_X1 U10324 ( .A1(n8987), .A2(n8986), .ZN(n9328) );
  INV_X1 U10325 ( .A(n9328), .ZN(n9009) );
  NAND2_X1 U10326 ( .A1(n8989), .A2(n9188), .ZN(n9354) );
  XNOR2_X1 U10327 ( .A(n9150), .B(n9449), .ZN(n9436) );
  NAND2_X1 U10328 ( .A1(n8991), .A2(n9179), .ZN(n9177) );
  INV_X1 U10329 ( .A(n9177), .ZN(n9442) );
  NOR2_X1 U10330 ( .A1(n8994), .A2(n8993), .ZN(n8998) );
  NAND4_X1 U10331 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n9001)
         );
  NOR4_X1 U10332 ( .A1(n9001), .A2(n9030), .A3(n9000), .A4(n8999), .ZN(n9003)
         );
  AND4_X1 U10333 ( .A1(n9003), .A2(n9836), .A3(n9002), .A4(n9630), .ZN(n9004)
         );
  NAND3_X1 U10334 ( .A1(n9442), .A2(n9475), .A3(n9004), .ZN(n9005) );
  NOR3_X1 U10335 ( .A1(n9414), .A2(n9436), .A3(n9005), .ZN(n9006) );
  NAND4_X1 U10336 ( .A1(n9366), .A2(n9402), .A3(n9387), .A4(n9006), .ZN(n9007)
         );
  NOR2_X1 U10337 ( .A1(n9354), .A2(n9007), .ZN(n9008) );
  NAND3_X1 U10338 ( .A1(n9009), .A2(n9342), .A3(n9008), .ZN(n9010) );
  NOR3_X1 U10339 ( .A1(n9291), .A2(n9311), .A3(n9010), .ZN(n9011) );
  NAND3_X1 U10340 ( .A1(n9013), .A2(n9012), .A3(n9011), .ZN(n9014) );
  OR3_X1 U10341 ( .A1(n9238), .A2(n9014), .A3(n9253), .ZN(n9015) );
  NOR2_X1 U10342 ( .A1(n9222), .A2(n9015), .ZN(n9016) );
  AND2_X1 U10343 ( .A1(n9199), .A2(n9016), .ZN(n9017) );
  AND2_X1 U10344 ( .A1(n9018), .A2(n9017), .ZN(n9020) );
  NAND4_X1 U10345 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n9024)
         );
  NAND2_X1 U10346 ( .A1(n9024), .A2(n9023), .ZN(n9054) );
  NAND3_X1 U10347 ( .A1(n9027), .A2(n9026), .A3(n9025), .ZN(n9029) );
  NAND2_X1 U10348 ( .A1(n9029), .A2(n9028), .ZN(n9032) );
  AOI21_X1 U10349 ( .B1(n9032), .B2(n7103), .A(n9031), .ZN(n9034) );
  OAI21_X1 U10350 ( .B1(n9035), .B2(n9034), .A(n9033), .ZN(n9036) );
  INV_X1 U10351 ( .A(n9036), .ZN(n9037) );
  NOR2_X1 U10352 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NOR2_X1 U10353 ( .A1(n9040), .A2(n9039), .ZN(n9043) );
  OAI211_X1 U10354 ( .C1(n9043), .C2(n9042), .A(n9221), .B(n9041), .ZN(n9046)
         );
  OAI211_X1 U10355 ( .C1(n9047), .C2(n9046), .A(n9045), .B(n9044), .ZN(n9048)
         );
  NAND2_X1 U10356 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  NAND2_X1 U10357 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NAND2_X1 U10358 ( .A1(n9052), .A2(n9054), .ZN(n9053) );
  MUX2_X1 U10359 ( .A(n9054), .B(n9053), .S(n9327), .Z(n9055) );
  INV_X1 U10360 ( .A(n9688), .ZN(n9131) );
  NAND2_X1 U10361 ( .A1(n9060), .A2(n9131), .ZN(n9066) );
  INV_X1 U10362 ( .A(n9061), .ZN(n9062) );
  OAI21_X1 U10363 ( .B1(n9063), .B2(n9062), .A(P1_B_REG_SCAN_IN), .ZN(n9064)
         );
  INV_X1 U10364 ( .A(n9064), .ZN(n9065) );
  OAI21_X1 U10365 ( .B1(n9067), .B2(n9066), .A(n9065), .ZN(n9068) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9069), .S(n9692), .Z(
        P1_U3586) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9070), .S(n9692), .Z(
        P1_U3585) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9227), .S(n9692), .Z(
        P1_U3584) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9169), .S(n9692), .Z(
        P1_U3583) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9255), .S(n9692), .Z(
        P1_U3582) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9265), .S(n9692), .Z(
        P1_U3581) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9254), .S(n9692), .Z(
        P1_U3580) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9266), .S(n9692), .Z(
        P1_U3579) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9162), .S(n9692), .Z(
        P1_U3577) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9343), .S(n9692), .Z(
        P1_U3576) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9358), .S(n9692), .Z(
        P1_U3575) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9369), .S(n9692), .Z(
        P1_U3574) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9389), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9403), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9419), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9427), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9418), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9461), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9634), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9462), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9633), .S(n9692), .Z(
        P1_U3565) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9071), .S(n9692), .Z(
        P1_U3564) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9072), .S(n9692), .Z(
        P1_U3563) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9074), .S(n9692), .Z(
        P1_U3561) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9075), .S(n9692), .Z(
        P1_U3560) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9076), .S(n9692), .Z(
        P1_U3559) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9077), .S(n9692), .Z(
        P1_U3558) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6850), .S(n9692), .Z(
        P1_U3557) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n4480), .S(n9692), .Z(
        P1_U3556) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6803), .S(n9692), .Z(
        P1_U3555) );
  OAI21_X1 U10397 ( .B1(n9080), .B2(n9079), .A(n9078), .ZN(n9081) );
  NAND2_X1 U10398 ( .A1(n9081), .A2(n9811), .ZN(n9092) );
  NOR2_X1 U10399 ( .A1(n9817), .A2(n9082), .ZN(n9083) );
  AOI211_X1 U10400 ( .C1(n9696), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9084), .B(
        n9083), .ZN(n9091) );
  AND3_X1 U10401 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(n9088) );
  OAI21_X1 U10402 ( .B1(n9089), .B2(n9088), .A(n9806), .ZN(n9090) );
  NAND3_X1 U10403 ( .A1(n9092), .A2(n9091), .A3(n9090), .ZN(P1_U3252) );
  AOI21_X1 U10404 ( .B1(n9094), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9093), .ZN(
        n9743) );
  NAND2_X1 U10405 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9746), .ZN(n9095) );
  OAI21_X1 U10406 ( .B1(n9746), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9095), .ZN(
        n9742) );
  NOR2_X1 U10407 ( .A1(n9743), .A2(n9742), .ZN(n9741) );
  AOI21_X1 U10408 ( .B1(n9746), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9741), .ZN(
        n9096) );
  NOR2_X1 U10409 ( .A1(n9096), .A2(n9761), .ZN(n9097) );
  INV_X1 U10410 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U10411 ( .A(n9761), .B(n9096), .ZN(n9756) );
  NOR2_X1 U10412 ( .A1(n9755), .A2(n9756), .ZN(n9754) );
  NOR2_X1 U10413 ( .A1(n9097), .A2(n9754), .ZN(n9098) );
  NOR2_X1 U10414 ( .A1(n9098), .A2(n9111), .ZN(n9099) );
  INV_X1 U10415 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U10416 ( .A(n9098), .B(n9111), .ZN(n9772) );
  NOR2_X1 U10417 ( .A1(n9771), .A2(n9772), .ZN(n9770) );
  NOR2_X1 U10418 ( .A1(n9099), .A2(n9770), .ZN(n9786) );
  XNOR2_X1 U10419 ( .A(n9789), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U10420 ( .A1(n9789), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U10421 ( .A1(n9782), .A2(n9100), .ZN(n9799) );
  INV_X1 U10422 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9101) );
  XNOR2_X1 U10423 ( .A(n9114), .B(n9101), .ZN(n9798) );
  NAND2_X1 U10424 ( .A1(n9799), .A2(n9798), .ZN(n9797) );
  NAND2_X1 U10425 ( .A1(n9114), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U10426 ( .A1(n9797), .A2(n9102), .ZN(n9814) );
  INV_X1 U10427 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9103) );
  MUX2_X1 U10428 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9103), .S(n9104), .Z(n9813) );
  NAND2_X1 U10429 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  NAND2_X1 U10430 ( .A1(n9104), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U10431 ( .A1(n9812), .A2(n9105), .ZN(n9106) );
  XNOR2_X1 U10432 ( .A(n9106), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9123) );
  INV_X1 U10433 ( .A(n9123), .ZN(n9120) );
  INV_X1 U10434 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9653) );
  INV_X1 U10435 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9659) );
  AOI21_X1 U10436 ( .B1(n9108), .B2(n9667), .A(n9107), .ZN(n9748) );
  MUX2_X1 U10437 ( .A(n9659), .B(P1_REG1_REG_13__SCAN_IN), .S(n9746), .Z(n9749) );
  NOR2_X1 U10438 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  AOI21_X1 U10439 ( .B1(n9109), .B2(n9659), .A(n9747), .ZN(n9765) );
  MUX2_X1 U10440 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9653), .S(n9761), .Z(n9764) );
  NOR2_X1 U10441 ( .A1(n9765), .A2(n9764), .ZN(n9763) );
  AOI21_X1 U10442 ( .B1(n9761), .B2(n9653), .A(n9763), .ZN(n9110) );
  NAND2_X1 U10443 ( .A1(n9775), .A2(n9110), .ZN(n9112) );
  XNOR2_X1 U10444 ( .A(n9111), .B(n9110), .ZN(n9777) );
  NAND2_X1 U10445 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U10446 ( .A1(n9112), .A2(n9776), .ZN(n9791) );
  INV_X1 U10447 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9113) );
  XNOR2_X1 U10448 ( .A(n9789), .B(n9113), .ZN(n9792) );
  AOI22_X1 U10449 ( .A1(n9791), .A2(n9792), .B1(n9789), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n9804) );
  XNOR2_X1 U10450 ( .A(n9114), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9805) );
  INV_X1 U10451 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9115) );
  OAI22_X1 U10452 ( .A1(n9804), .A2(n9805), .B1(n9802), .B2(n9115), .ZN(n9822)
         );
  INV_X1 U10453 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10454 ( .A1(n9818), .A2(n9116), .ZN(n9117) );
  OAI21_X1 U10455 ( .B1(n9818), .B2(n9116), .A(n9117), .ZN(n9821) );
  NOR2_X1 U10456 ( .A1(n9822), .A2(n9821), .ZN(n9820) );
  INV_X1 U10457 ( .A(n9117), .ZN(n9118) );
  NOR2_X1 U10458 ( .A1(n9820), .A2(n9118), .ZN(n9119) );
  XOR2_X1 U10459 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9119), .Z(n9121) );
  AOI22_X1 U10460 ( .A1(n9120), .A2(n9811), .B1(n9121), .B2(n9806), .ZN(n9125)
         );
  OAI21_X1 U10461 ( .B1(n9121), .B2(n9823), .A(n9817), .ZN(n9122) );
  AOI21_X1 U10462 ( .B1(n9123), .B2(n9723), .A(n9122), .ZN(n9124) );
  MUX2_X1 U10463 ( .A(n9125), .B(n9124), .S(n9863), .Z(n9128) );
  INV_X1 U10464 ( .A(n9126), .ZN(n9127) );
  OAI211_X1 U10465 ( .C1(n9129), .C2(n9828), .A(n9128), .B(n9127), .ZN(
        P1_U3260) );
  INV_X1 U10466 ( .A(n9452), .ZN(n9654) );
  NAND2_X1 U10467 ( .A1(n9465), .A2(n9654), .ZN(n9450) );
  OR2_X2 U10468 ( .A1(n9428), .A2(n9565), .ZN(n9409) );
  NAND2_X1 U10469 ( .A1(n9334), .A2(n9161), .ZN(n9318) );
  OR2_X2 U10470 ( .A1(n9318), .A2(n9525), .ZN(n9305) );
  AND2_X2 U10471 ( .A1(n9219), .A2(n9241), .ZN(n9215) );
  NAND2_X1 U10472 ( .A1(n9209), .A2(n9215), .ZN(n9206) );
  NOR2_X1 U10473 ( .A1(n9486), .A2(n9206), .ZN(n9130) );
  XOR2_X1 U10474 ( .A(n9482), .B(n9130), .Z(n9484) );
  NAND2_X1 U10475 ( .A1(n9131), .A2(P1_B_REG_SCAN_IN), .ZN(n9132) );
  NAND2_X1 U10476 ( .A1(n9635), .A2(n9132), .ZN(n9202) );
  NOR2_X1 U10477 ( .A1(n9133), .A2(n9202), .ZN(n9485) );
  INV_X1 U10478 ( .A(n9485), .ZN(n9134) );
  NOR2_X1 U10479 ( .A1(n9134), .A2(n9640), .ZN(n9137) );
  AOI21_X1 U10480 ( .B1(n9640), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9137), .ZN(
        n9136) );
  NAND2_X1 U10481 ( .A1(n9482), .A2(n9644), .ZN(n9135) );
  OAI211_X1 U10482 ( .C1(n9484), .C2(n9455), .A(n9136), .B(n9135), .ZN(
        P1_U3261) );
  XNOR2_X1 U10483 ( .A(n9486), .B(n9206), .ZN(n9488) );
  AOI21_X1 U10484 ( .B1(n9640), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9137), .ZN(
        n9139) );
  NAND2_X1 U10485 ( .A1(n9486), .A2(n9644), .ZN(n9138) );
  OAI211_X1 U10486 ( .C1(n9488), .C2(n9455), .A(n9139), .B(n9138), .ZN(
        P1_U3262) );
  OR2_X1 U10487 ( .A1(n9140), .A2(n9633), .ZN(n9141) );
  NAND2_X1 U10488 ( .A1(n9624), .A2(n9668), .ZN(n9144) );
  NAND2_X1 U10489 ( .A1(n9471), .A2(n9634), .ZN(n9146) );
  OR2_X1 U10490 ( .A1(n9452), .A2(n9461), .ZN(n9147) );
  NAND2_X1 U10491 ( .A1(n9452), .A2(n9461), .ZN(n9148) );
  AND2_X1 U10492 ( .A1(n9150), .A2(n9418), .ZN(n9151) );
  NAND2_X1 U10493 ( .A1(n9565), .A2(n9427), .ZN(n9152) );
  NAND2_X1 U10494 ( .A1(n9153), .A2(n9152), .ZN(n9394) );
  NAND2_X1 U10495 ( .A1(n9561), .A2(n9419), .ZN(n9154) );
  OR2_X1 U10496 ( .A1(n9555), .A2(n9403), .ZN(n9155) );
  NAND2_X1 U10497 ( .A1(n9156), .A2(n9155), .ZN(n9363) );
  NOR2_X1 U10498 ( .A1(n9542), .A2(n9369), .ZN(n9158) );
  NAND2_X1 U10499 ( .A1(n9309), .A2(n9325), .ZN(n9164) );
  NOR2_X1 U10500 ( .A1(n9522), .A2(n9313), .ZN(n9165) );
  NOR2_X1 U10501 ( .A1(n9287), .A2(n9294), .ZN(n9166) );
  XNOR2_X1 U10502 ( .A(n9170), .B(n9199), .ZN(n9489) );
  INV_X1 U10503 ( .A(n9489), .ZN(n9213) );
  NAND2_X1 U10504 ( .A1(n9631), .A2(n9630), .ZN(n9175) );
  NAND2_X1 U10505 ( .A1(n9175), .A2(n9174), .ZN(n9459) );
  NAND2_X1 U10506 ( .A1(n9459), .A2(n9475), .ZN(n9444) );
  INV_X1 U10507 ( .A(n9443), .ZN(n9176) );
  NOR2_X1 U10508 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  NOR2_X1 U10509 ( .A1(n9414), .A2(n9415), .ZN(n9180) );
  NAND2_X1 U10510 ( .A1(n9416), .A2(n9181), .ZN(n9401) );
  NAND2_X1 U10511 ( .A1(n9401), .A2(n9402), .ZN(n9400) );
  NOR2_X1 U10512 ( .A1(n9380), .A2(n9182), .ZN(n9185) );
  INV_X1 U10513 ( .A(n9183), .ZN(n9184) );
  INV_X1 U10514 ( .A(n9366), .ZN(n9186) );
  INV_X1 U10515 ( .A(n9187), .ZN(n9355) );
  NAND2_X1 U10516 ( .A1(n9342), .A2(n9188), .ZN(n9190) );
  INV_X1 U10517 ( .A(n9191), .ZN(n9192) );
  OAI21_X1 U10518 ( .B1(n9292), .B2(n9291), .A(n9194), .ZN(n9276) );
  NAND2_X1 U10519 ( .A1(n9239), .A2(n9235), .ZN(n9220) );
  NAND3_X1 U10520 ( .A1(n9220), .A2(n9197), .A3(n9221), .ZN(n9226) );
  NAND2_X1 U10521 ( .A1(n9226), .A2(n9198), .ZN(n9200) );
  INV_X1 U10522 ( .A(n9204), .ZN(n9205) );
  OAI21_X1 U10523 ( .B1(n9209), .B2(n9215), .A(n9206), .ZN(n9490) );
  NOR2_X1 U10524 ( .A1(n9490), .A2(n9455), .ZN(n9211) );
  AOI22_X1 U10525 ( .A1(n9207), .A2(n9861), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9640), .ZN(n9208) );
  OAI21_X1 U10526 ( .B1(n9209), .B2(n9845), .A(n9208), .ZN(n9210) );
  AOI211_X1 U10527 ( .C1(n9491), .C2(n9874), .A(n9211), .B(n9210), .ZN(n9212)
         );
  OAI21_X1 U10528 ( .B1(n9213), .B2(n9477), .A(n9212), .ZN(P1_U3355) );
  INV_X1 U10529 ( .A(n9241), .ZN(n9216) );
  AOI21_X1 U10530 ( .B1(n9495), .B2(n9216), .A(n9215), .ZN(n9496) );
  AOI22_X1 U10531 ( .A1(n9217), .A2(n9861), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9640), .ZN(n9218) );
  OAI21_X1 U10532 ( .B1(n9219), .B2(n9845), .A(n9218), .ZN(n9233) );
  INV_X1 U10533 ( .A(n9220), .ZN(n9224) );
  INV_X1 U10534 ( .A(n9221), .ZN(n9223) );
  OAI21_X1 U10535 ( .B1(n9224), .B2(n9223), .A(n9222), .ZN(n9225) );
  NAND2_X1 U10536 ( .A1(n9226), .A2(n9225), .ZN(n9231) );
  NAND2_X1 U10537 ( .A1(n9255), .A2(n9632), .ZN(n9229) );
  NAND2_X1 U10538 ( .A1(n9227), .A2(n9635), .ZN(n9228) );
  AOI211_X1 U10539 ( .C1(n9496), .C2(n9833), .A(n9233), .B(n9232), .ZN(n9234)
         );
  OAI21_X1 U10540 ( .B1(n9477), .B2(n9499), .A(n9234), .ZN(P1_U3263) );
  XNOR2_X1 U10541 ( .A(n9236), .B(n9235), .ZN(n9504) );
  NOR2_X1 U10542 ( .A1(n9237), .A2(n9845), .ZN(n9245) );
  XNOR2_X1 U10543 ( .A(n9239), .B(n9238), .ZN(n9240) );
  AOI222_X1 U10544 ( .A1(n9840), .A2(n9240), .B1(n9169), .B2(n9635), .C1(n9265), .C2(n9632), .ZN(n9503) );
  AOI211_X1 U10545 ( .C1(n9501), .C2(n9248), .A(n9934), .B(n9241), .ZN(n9500)
         );
  AOI22_X1 U10546 ( .A1(n9500), .A2(n9327), .B1(n9861), .B2(n9242), .ZN(n9243)
         );
  AOI21_X1 U10547 ( .B1(n9503), .B2(n9243), .A(n9640), .ZN(n9244) );
  AOI211_X1 U10548 ( .C1(n9640), .C2(P1_REG2_REG_27__SCAN_IN), .A(n9245), .B(
        n9244), .ZN(n9246) );
  OAI21_X1 U10549 ( .B1(n9504), .B2(n9477), .A(n9246), .ZN(P1_U3264) );
  XNOR2_X1 U10550 ( .A(n9247), .B(n9253), .ZN(n9509) );
  AOI21_X1 U10551 ( .B1(n9505), .B2(n9268), .A(n4705), .ZN(n9506) );
  AOI22_X1 U10552 ( .A1(n9249), .A2(n9861), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9640), .ZN(n9250) );
  OAI21_X1 U10553 ( .B1(n9251), .B2(n9845), .A(n9250), .ZN(n9258) );
  XOR2_X1 U10554 ( .A(n9253), .B(n9252), .Z(n9256) );
  AOI222_X1 U10555 ( .A1(n9840), .A2(n9256), .B1(n9255), .B2(n9635), .C1(n9254), .C2(n9632), .ZN(n9508) );
  NOR2_X1 U10556 ( .A1(n9508), .A2(n9640), .ZN(n9257) );
  AOI211_X1 U10557 ( .C1(n9506), .C2(n9833), .A(n9258), .B(n9257), .ZN(n9259)
         );
  OAI21_X1 U10558 ( .B1(n9477), .B2(n9509), .A(n9259), .ZN(P1_U3265) );
  XOR2_X1 U10559 ( .A(n9263), .B(n9260), .Z(n9514) );
  NOR2_X1 U10560 ( .A1(n9261), .A2(n9845), .ZN(n9273) );
  NOR2_X1 U10561 ( .A1(n4489), .A2(n9262), .ZN(n9264) );
  XNOR2_X1 U10562 ( .A(n9264), .B(n9263), .ZN(n9267) );
  AOI222_X1 U10563 ( .A1(n9840), .A2(n9267), .B1(n9266), .B2(n9632), .C1(n9265), .C2(n9635), .ZN(n9513) );
  INV_X1 U10564 ( .A(n9281), .ZN(n9269) );
  AOI211_X1 U10565 ( .C1(n9511), .C2(n9269), .A(n9934), .B(n4701), .ZN(n9510)
         );
  AOI22_X1 U10566 ( .A1(n9510), .A2(n9327), .B1(n9861), .B2(n9270), .ZN(n9271)
         );
  AOI21_X1 U10567 ( .B1(n9513), .B2(n9271), .A(n9640), .ZN(n9272) );
  AOI211_X1 U10568 ( .C1(n9640), .C2(P1_REG2_REG_25__SCAN_IN), .A(n9273), .B(
        n9272), .ZN(n9274) );
  OAI21_X1 U10569 ( .B1(n9514), .B2(n9477), .A(n9274), .ZN(P1_U3266) );
  XNOR2_X1 U10570 ( .A(n9275), .B(n9277), .ZN(n9519) );
  AOI21_X1 U10571 ( .B1(n9277), .B2(n9276), .A(n4489), .ZN(n9278) );
  OAI222_X1 U10572 ( .A1(n9871), .A2(n9280), .B1(n9869), .B2(n9279), .C1(n9866), .C2(n9278), .ZN(n9515) );
  INV_X1 U10573 ( .A(n9295), .ZN(n9282) );
  AOI211_X1 U10574 ( .C1(n9517), .C2(n9282), .A(n9934), .B(n9281), .ZN(n9516)
         );
  INV_X1 U10575 ( .A(n9376), .ZN(n9296) );
  NAND2_X1 U10576 ( .A1(n9516), .A2(n9296), .ZN(n9286) );
  INV_X1 U10577 ( .A(n9283), .ZN(n9284) );
  AOI22_X1 U10578 ( .A1(n9284), .A2(n9861), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9640), .ZN(n9285) );
  OAI211_X1 U10579 ( .C1(n9287), .C2(n9845), .A(n9286), .B(n9285), .ZN(n9288)
         );
  AOI21_X1 U10580 ( .B1(n9515), .B2(n9874), .A(n9288), .ZN(n9289) );
  OAI21_X1 U10581 ( .B1(n9519), .B2(n9477), .A(n9289), .ZN(P1_U3267) );
  XOR2_X1 U10582 ( .A(n9290), .B(n9291), .Z(n9524) );
  XNOR2_X1 U10583 ( .A(n9292), .B(n9291), .ZN(n9293) );
  OAI222_X1 U10584 ( .A1(n9871), .A2(n9325), .B1(n9869), .B2(n9294), .C1(n9866), .C2(n9293), .ZN(n9520) );
  AOI211_X1 U10585 ( .C1(n9522), .C2(n9305), .A(n9934), .B(n9295), .ZN(n9521)
         );
  NAND2_X1 U10586 ( .A1(n9521), .A2(n9296), .ZN(n9300) );
  INV_X1 U10587 ( .A(n9297), .ZN(n9298) );
  AOI22_X1 U10588 ( .A1(n9298), .A2(n9861), .B1(n9640), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9299) );
  OAI211_X1 U10589 ( .C1(n9301), .C2(n9845), .A(n9300), .B(n9299), .ZN(n9302)
         );
  AOI21_X1 U10590 ( .B1(n9520), .B2(n9874), .A(n9302), .ZN(n9303) );
  OAI21_X1 U10591 ( .B1(n9524), .B2(n9477), .A(n9303), .ZN(P1_U3268) );
  XNOR2_X1 U10592 ( .A(n9304), .B(n9311), .ZN(n9529) );
  INV_X1 U10593 ( .A(n9305), .ZN(n9306) );
  AOI21_X1 U10594 ( .B1(n9525), .B2(n9318), .A(n9306), .ZN(n9526) );
  AOI22_X1 U10595 ( .A1(n9640), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9307), .B2(
        n9861), .ZN(n9308) );
  OAI21_X1 U10596 ( .B1(n9309), .B2(n9845), .A(n9308), .ZN(n9316) );
  NOR2_X1 U10597 ( .A1(n4518), .A2(n9310), .ZN(n9312) );
  XNOR2_X1 U10598 ( .A(n9312), .B(n9311), .ZN(n9314) );
  AOI222_X1 U10599 ( .A1(n9840), .A2(n9314), .B1(n9343), .B2(n9632), .C1(n9313), .C2(n9635), .ZN(n9528) );
  NOR2_X1 U10600 ( .A1(n9528), .A2(n9640), .ZN(n9315) );
  AOI211_X1 U10601 ( .C1(n9526), .C2(n9833), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI21_X1 U10602 ( .B1(n9477), .B2(n9529), .A(n9317), .ZN(P1_U3269) );
  INV_X1 U10603 ( .A(n9334), .ZN(n9320) );
  INV_X1 U10604 ( .A(n9318), .ZN(n9319) );
  AOI211_X1 U10605 ( .C1(n9532), .C2(n9320), .A(n9934), .B(n9319), .ZN(n9531)
         );
  NOR2_X1 U10606 ( .A1(n9321), .A2(n9847), .ZN(n9326) );
  AOI21_X1 U10607 ( .B1(n9328), .B2(n9322), .A(n4518), .ZN(n9323) );
  OAI222_X1 U10608 ( .A1(n9869), .A2(n9325), .B1(n9871), .B2(n9324), .C1(n9866), .C2(n9323), .ZN(n9530) );
  AOI211_X1 U10609 ( .C1(n9531), .C2(n9327), .A(n9326), .B(n9530), .ZN(n9332)
         );
  AOI22_X1 U10610 ( .A1(n9532), .A2(n9644), .B1(n9640), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9331) );
  OR2_X1 U10611 ( .A1(n9329), .A2(n9328), .ZN(n9534) );
  INV_X1 U10612 ( .A(n9477), .ZN(n9437) );
  NAND3_X1 U10613 ( .A1(n9534), .A2(n9533), .A3(n9437), .ZN(n9330) );
  OAI211_X1 U10614 ( .C1(n9332), .C2(n9640), .A(n9331), .B(n9330), .ZN(
        P1_U3270) );
  XOR2_X1 U10615 ( .A(n9342), .B(n9333), .Z(n9541) );
  INV_X1 U10616 ( .A(n9349), .ZN(n9335) );
  AOI21_X1 U10617 ( .B1(n9537), .B2(n9335), .A(n9334), .ZN(n9538) );
  INV_X1 U10618 ( .A(n9336), .ZN(n9337) );
  AOI22_X1 U10619 ( .A1(n9640), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9337), .B2(
        n9861), .ZN(n9338) );
  OAI21_X1 U10620 ( .B1(n9339), .B2(n9845), .A(n9338), .ZN(n9346) );
  NOR2_X1 U10621 ( .A1(n9353), .A2(n9340), .ZN(n9341) );
  XOR2_X1 U10622 ( .A(n9342), .B(n9341), .Z(n9344) );
  AOI222_X1 U10623 ( .A1(n9840), .A2(n9344), .B1(n9369), .B2(n9632), .C1(n9343), .C2(n9635), .ZN(n9540) );
  NOR2_X1 U10624 ( .A1(n9540), .A2(n9640), .ZN(n9345) );
  AOI211_X1 U10625 ( .C1(n9538), .C2(n9833), .A(n9346), .B(n9345), .ZN(n9347)
         );
  OAI21_X1 U10626 ( .B1(n9477), .B2(n9541), .A(n9347), .ZN(P1_U3271) );
  XOR2_X1 U10627 ( .A(n9348), .B(n9354), .Z(n9546) );
  AOI21_X1 U10628 ( .B1(n9542), .B2(n4570), .A(n9349), .ZN(n9543) );
  AOI22_X1 U10629 ( .A1(n9640), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9350), .B2(
        n9861), .ZN(n9351) );
  OAI21_X1 U10630 ( .B1(n9352), .B2(n9845), .A(n9351), .ZN(n9361) );
  OAI21_X1 U10631 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(n9357) );
  NAND2_X1 U10632 ( .A1(n4929), .A2(n9357), .ZN(n9359) );
  AOI222_X1 U10633 ( .A1(n9840), .A2(n9359), .B1(n9389), .B2(n9632), .C1(n9358), .C2(n9635), .ZN(n9545) );
  NOR2_X1 U10634 ( .A1(n9545), .A2(n9640), .ZN(n9360) );
  AOI211_X1 U10635 ( .C1(n9543), .C2(n9833), .A(n9361), .B(n9360), .ZN(n9362)
         );
  OAI21_X1 U10636 ( .B1(n9477), .B2(n9546), .A(n9362), .ZN(P1_U3272) );
  AND2_X1 U10637 ( .A1(n9363), .A2(n9366), .ZN(n9364) );
  OR2_X1 U10638 ( .A1(n9365), .A2(n9364), .ZN(n9547) );
  XNOR2_X1 U10639 ( .A(n9367), .B(n9366), .ZN(n9368) );
  NAND2_X1 U10640 ( .A1(n9368), .A2(n9840), .ZN(n9371) );
  AOI22_X1 U10641 ( .A1(n9635), .A2(n9369), .B1(n9403), .B2(n9632), .ZN(n9370)
         );
  NAND2_X1 U10642 ( .A1(n9371), .A2(n9370), .ZN(n9552) );
  AOI21_X1 U10643 ( .B1(n9381), .B2(n9548), .A(n9934), .ZN(n9372) );
  NAND2_X1 U10644 ( .A1(n9372), .A2(n4570), .ZN(n9550) );
  AOI22_X1 U10645 ( .A1(n9640), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9373), .B2(
        n9861), .ZN(n9375) );
  NAND2_X1 U10646 ( .A1(n9548), .A2(n9644), .ZN(n9374) );
  OAI211_X1 U10647 ( .C1(n9550), .C2(n9376), .A(n9375), .B(n9374), .ZN(n9377)
         );
  AOI21_X1 U10648 ( .B1(n9552), .B2(n9874), .A(n9377), .ZN(n9378) );
  OAI21_X1 U10649 ( .B1(n9547), .B2(n9477), .A(n9378), .ZN(P1_U3273) );
  XNOR2_X1 U10650 ( .A(n9379), .B(n9380), .ZN(n9559) );
  INV_X1 U10651 ( .A(n9396), .ZN(n9382) );
  AOI21_X1 U10652 ( .B1(n9555), .B2(n9382), .A(n4709), .ZN(n9556) );
  AOI22_X1 U10653 ( .A1(n9640), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9383), .B2(
        n9861), .ZN(n9384) );
  OAI21_X1 U10654 ( .B1(n9385), .B2(n9845), .A(n9384), .ZN(n9392) );
  NAND2_X1 U10655 ( .A1(n9400), .A2(n9386), .ZN(n9388) );
  XNOR2_X1 U10656 ( .A(n9388), .B(n9387), .ZN(n9390) );
  AOI222_X1 U10657 ( .A1(n9840), .A2(n9390), .B1(n9389), .B2(n9635), .C1(n9419), .C2(n9632), .ZN(n9558) );
  NOR2_X1 U10658 ( .A1(n9558), .A2(n9640), .ZN(n9391) );
  AOI211_X1 U10659 ( .C1(n9556), .C2(n9833), .A(n9392), .B(n9391), .ZN(n9393)
         );
  OAI21_X1 U10660 ( .B1(n9477), .B2(n9559), .A(n9393), .ZN(P1_U3274) );
  XNOR2_X1 U10661 ( .A(n9394), .B(n9395), .ZN(n9564) );
  AOI211_X1 U10662 ( .C1(n9561), .C2(n9409), .A(n9934), .B(n9396), .ZN(n9560)
         );
  AOI22_X1 U10663 ( .A1(n9640), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9397), .B2(
        n9861), .ZN(n9398) );
  OAI21_X1 U10664 ( .B1(n9399), .B2(n9845), .A(n9398), .ZN(n9406) );
  OAI21_X1 U10665 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9404) );
  AOI222_X1 U10666 ( .A1(n9840), .A2(n9404), .B1(n9403), .B2(n9635), .C1(n9427), .C2(n9632), .ZN(n9563) );
  NOR2_X1 U10667 ( .A1(n9563), .A2(n9640), .ZN(n9405) );
  AOI211_X1 U10668 ( .C1(n9560), .C2(n9433), .A(n9406), .B(n9405), .ZN(n9407)
         );
  OAI21_X1 U10669 ( .B1(n9477), .B2(n9564), .A(n9407), .ZN(P1_U3275) );
  XOR2_X1 U10670 ( .A(n9408), .B(n9414), .Z(n9569) );
  INV_X1 U10671 ( .A(n9409), .ZN(n9410) );
  AOI21_X1 U10672 ( .B1(n9565), .B2(n9428), .A(n9410), .ZN(n9566) );
  INV_X1 U10673 ( .A(n9565), .ZN(n9413) );
  AOI22_X1 U10674 ( .A1(n9640), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9411), .B2(
        n9861), .ZN(n9412) );
  OAI21_X1 U10675 ( .B1(n9413), .B2(n9845), .A(n9412), .ZN(n9422) );
  OAI21_X1 U10676 ( .B1(n4567), .B2(n9415), .A(n9414), .ZN(n9417) );
  NAND2_X1 U10677 ( .A1(n9417), .A2(n9416), .ZN(n9420) );
  AOI222_X1 U10678 ( .A1(n9840), .A2(n9420), .B1(n9419), .B2(n9635), .C1(n9418), .C2(n9632), .ZN(n9568) );
  NOR2_X1 U10679 ( .A1(n9568), .A2(n9640), .ZN(n9421) );
  AOI211_X1 U10680 ( .C1(n9566), .C2(n9833), .A(n9422), .B(n9421), .ZN(n9423)
         );
  OAI21_X1 U10681 ( .B1(n9569), .B2(n9477), .A(n9423), .ZN(P1_U3276) );
  AND2_X1 U10682 ( .A1(n9461), .A2(n9632), .ZN(n9426) );
  AOI211_X1 U10683 ( .C1(n9436), .C2(n9424), .A(n9866), .B(n4567), .ZN(n9425)
         );
  AOI211_X1 U10684 ( .C1(n9635), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9649)
         );
  INV_X1 U10685 ( .A(n9450), .ZN(n9429) );
  OAI211_X1 U10686 ( .C1(n9429), .C2(n9650), .A(n9856), .B(n9428), .ZN(n9648)
         );
  INV_X1 U10687 ( .A(n9648), .ZN(n9434) );
  AOI22_X1 U10688 ( .A1(n9640), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9430), .B2(
        n9861), .ZN(n9431) );
  OAI21_X1 U10689 ( .B1(n9650), .B2(n9845), .A(n9431), .ZN(n9432) );
  AOI21_X1 U10690 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9439) );
  XOR2_X1 U10691 ( .A(n9435), .B(n9436), .Z(n9652) );
  NAND2_X1 U10692 ( .A1(n9652), .A2(n9437), .ZN(n9438) );
  OAI211_X1 U10693 ( .C1(n9649), .C2(n9640), .A(n9439), .B(n9438), .ZN(
        P1_U3277) );
  XNOR2_X1 U10694 ( .A(n9440), .B(n9442), .ZN(n9658) );
  INV_X1 U10695 ( .A(n9658), .ZN(n9458) );
  INV_X1 U10696 ( .A(n9441), .ZN(n9446) );
  AOI21_X1 U10697 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(n9445) );
  NOR2_X1 U10698 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  OAI222_X1 U10699 ( .A1(n9869), .A2(n9449), .B1(n9871), .B2(n9448), .C1(n9866), .C2(n9447), .ZN(n9656) );
  OAI21_X1 U10700 ( .B1(n9465), .B2(n9654), .A(n9450), .ZN(n9655) );
  AOI22_X1 U10701 ( .A1(n9640), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9451), .B2(
        n9861), .ZN(n9454) );
  NAND2_X1 U10702 ( .A1(n9452), .A2(n9644), .ZN(n9453) );
  OAI211_X1 U10703 ( .C1(n9655), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9456)
         );
  AOI21_X1 U10704 ( .B1(n9656), .B2(n9874), .A(n9456), .ZN(n9457) );
  OAI21_X1 U10705 ( .B1(n9477), .B2(n9458), .A(n9457), .ZN(P1_U3278) );
  XNOR2_X1 U10706 ( .A(n9459), .B(n5064), .ZN(n9460) );
  NAND2_X1 U10707 ( .A1(n9460), .A2(n9840), .ZN(n9464) );
  AOI22_X1 U10708 ( .A1(n9632), .A2(n9462), .B1(n9461), .B2(n9635), .ZN(n9463)
         );
  NAND2_X1 U10709 ( .A1(n9464), .A2(n9463), .ZN(n9665) );
  OAI21_X1 U10710 ( .B1(n4587), .B2(n9663), .A(n9856), .ZN(n9466) );
  OR2_X1 U10711 ( .A1(n9466), .A2(n9465), .ZN(n9662) );
  INV_X1 U10712 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9469) );
  INV_X1 U10713 ( .A(n9467), .ZN(n9468) );
  OAI22_X1 U10714 ( .A1(n9874), .A2(n9469), .B1(n9468), .B2(n9847), .ZN(n9470)
         );
  AOI21_X1 U10715 ( .B1(n9471), .B2(n9644), .A(n9470), .ZN(n9472) );
  OAI21_X1 U10716 ( .B1(n9662), .B2(n9473), .A(n9472), .ZN(n9480) );
  INV_X1 U10717 ( .A(n9474), .ZN(n9478) );
  AND2_X1 U10718 ( .A1(n9476), .A2(n9475), .ZN(n9661) );
  NOR3_X1 U10719 ( .A1(n9478), .A2(n9661), .A3(n9477), .ZN(n9479) );
  AOI211_X1 U10720 ( .C1(n9874), .C2(n9665), .A(n9480), .B(n9479), .ZN(n9481)
         );
  INV_X1 U10721 ( .A(n9481), .ZN(P1_U3279) );
  AOI21_X1 U10722 ( .B1(n9482), .B2(n9647), .A(n9485), .ZN(n9483) );
  OAI21_X1 U10723 ( .B1(n9484), .B2(n9934), .A(n9483), .ZN(n9570) );
  MUX2_X1 U10724 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9570), .S(n9948), .Z(
        P1_U3554) );
  AOI21_X1 U10725 ( .B1(n9486), .B2(n9647), .A(n9485), .ZN(n9487) );
  OAI21_X1 U10726 ( .B1(n9488), .B2(n9934), .A(n9487), .ZN(n9571) );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9571), .S(n9948), .Z(
        P1_U3553) );
  NAND2_X1 U10728 ( .A1(n9489), .A2(n9924), .ZN(n9494) );
  NAND2_X1 U10729 ( .A1(n9494), .A2(n9493), .ZN(n9572) );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9572), .S(n9948), .Z(
        P1_U3552) );
  AOI22_X1 U10731 ( .A1(n9496), .A2(n9856), .B1(n9647), .B2(n9495), .ZN(n9497)
         );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9573), .S(n9948), .Z(
        P1_U3551) );
  AOI21_X1 U10733 ( .B1(n9647), .B2(n9501), .A(n9500), .ZN(n9502) );
  OAI211_X1 U10734 ( .C1(n9504), .C2(n9660), .A(n9503), .B(n9502), .ZN(n9574)
         );
  MUX2_X1 U10735 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9574), .S(n9948), .Z(
        P1_U3550) );
  AOI22_X1 U10736 ( .A1(n9506), .A2(n9856), .B1(n9647), .B2(n9505), .ZN(n9507)
         );
  OAI211_X1 U10737 ( .C1(n9509), .C2(n9660), .A(n9508), .B(n9507), .ZN(n9575)
         );
  MUX2_X1 U10738 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9575), .S(n9948), .Z(
        P1_U3549) );
  AOI21_X1 U10739 ( .B1(n9647), .B2(n9511), .A(n9510), .ZN(n9512) );
  OAI211_X1 U10740 ( .C1(n9514), .C2(n9660), .A(n9513), .B(n9512), .ZN(n9576)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9576), .S(n9948), .Z(
        P1_U3548) );
  AOI211_X1 U10742 ( .C1(n9647), .C2(n9517), .A(n9516), .B(n9515), .ZN(n9518)
         );
  OAI21_X1 U10743 ( .B1(n9660), .B2(n9519), .A(n9518), .ZN(n9577) );
  MUX2_X1 U10744 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9577), .S(n9948), .Z(
        P1_U3547) );
  AOI211_X1 U10745 ( .C1(n9647), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9523)
         );
  OAI21_X1 U10746 ( .B1(n9524), .B2(n9660), .A(n9523), .ZN(n9578) );
  MUX2_X1 U10747 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9578), .S(n9948), .Z(
        P1_U3546) );
  AOI22_X1 U10748 ( .A1(n9526), .A2(n9856), .B1(n9647), .B2(n9525), .ZN(n9527)
         );
  OAI211_X1 U10749 ( .C1(n9529), .C2(n9660), .A(n9528), .B(n9527), .ZN(n9579)
         );
  MUX2_X1 U10750 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9579), .S(n9948), .Z(
        P1_U3545) );
  AOI211_X1 U10751 ( .C1(n9647), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9536)
         );
  NAND3_X1 U10752 ( .A1(n9534), .A2(n9533), .A3(n9924), .ZN(n9535) );
  NAND2_X1 U10753 ( .A1(n9536), .A2(n9535), .ZN(n9580) );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9580), .S(n9948), .Z(
        P1_U3544) );
  AOI22_X1 U10755 ( .A1(n9538), .A2(n9856), .B1(n9647), .B2(n9537), .ZN(n9539)
         );
  OAI211_X1 U10756 ( .C1(n9541), .C2(n9660), .A(n9540), .B(n9539), .ZN(n9581)
         );
  MUX2_X1 U10757 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9581), .S(n9948), .Z(
        P1_U3543) );
  AOI22_X1 U10758 ( .A1(n9543), .A2(n9856), .B1(n9647), .B2(n9542), .ZN(n9544)
         );
  OAI211_X1 U10759 ( .C1(n9546), .C2(n9660), .A(n9545), .B(n9544), .ZN(n9582)
         );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9582), .S(n9948), .Z(
        P1_U3542) );
  OR2_X1 U10761 ( .A1(n9547), .A2(n9660), .ZN(n9554) );
  NAND2_X1 U10762 ( .A1(n9548), .A2(n9647), .ZN(n9549) );
  NAND2_X1 U10763 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  NOR2_X1 U10764 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  NAND2_X1 U10765 ( .A1(n9554), .A2(n9553), .ZN(n9583) );
  MUX2_X1 U10766 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9583), .S(n9948), .Z(
        P1_U3541) );
  AOI22_X1 U10767 ( .A1(n9556), .A2(n9856), .B1(n9647), .B2(n9555), .ZN(n9557)
         );
  OAI211_X1 U10768 ( .C1(n9559), .C2(n9660), .A(n9558), .B(n9557), .ZN(n9584)
         );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9584), .S(n9948), .Z(
        P1_U3540) );
  AOI21_X1 U10770 ( .B1(n9647), .B2(n9561), .A(n9560), .ZN(n9562) );
  OAI211_X1 U10771 ( .C1(n9564), .C2(n9660), .A(n9563), .B(n9562), .ZN(n9585)
         );
  MUX2_X1 U10772 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9585), .S(n9948), .Z(
        P1_U3539) );
  AOI22_X1 U10773 ( .A1(n9566), .A2(n9856), .B1(n9647), .B2(n9565), .ZN(n9567)
         );
  OAI211_X1 U10774 ( .C1(n9569), .C2(n9660), .A(n9568), .B(n9567), .ZN(n9586)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9586), .S(n9948), .Z(
        P1_U3538) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9570), .S(n9906), .Z(
        P1_U3522) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9571), .S(n9906), .Z(
        P1_U3521) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9572), .S(n9906), .Z(
        P1_U3520) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9574), .S(n9906), .Z(
        P1_U3518) );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9575), .S(n9906), .Z(
        P1_U3517) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9576), .S(n9906), .Z(
        P1_U3516) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9577), .S(n9906), .Z(
        P1_U3515) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9578), .S(n9906), .Z(
        P1_U3514) );
  MUX2_X1 U10784 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9579), .S(n9906), .Z(
        P1_U3513) );
  MUX2_X1 U10785 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9580), .S(n9906), .Z(
        P1_U3512) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9581), .S(n9906), .Z(
        P1_U3511) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9582), .S(n9906), .Z(
        P1_U3510) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9583), .S(n9906), .Z(
        P1_U3508) );
  MUX2_X1 U10789 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9584), .S(n9906), .Z(
        P1_U3505) );
  MUX2_X1 U10790 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9585), .S(n9906), .Z(
        P1_U3502) );
  MUX2_X1 U10791 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9586), .S(n9906), .Z(
        P1_U3499) );
  NOR2_X1 U10792 ( .A1(n9587), .A2(n9881), .ZN(n9878) );
  MUX2_X1 U10793 ( .A(P1_D_REG_0__SCAN_IN), .B(n9588), .S(n9878), .Z(P1_U3440)
         );
  INV_X1 U10794 ( .A(n5127), .ZN(n9589) );
  NOR4_X1 U10795 ( .A1(n9589), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5453), .ZN(n9590) );
  AOI21_X1 U10796 ( .B1(n9597), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9590), .ZN(
        n9591) );
  OAI21_X1 U10797 ( .B1(n9592), .B2(n9599), .A(n9591), .ZN(P1_U3322) );
  INV_X1 U10798 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10427) );
  OAI222_X1 U10799 ( .A1(n9595), .A2(n10427), .B1(n9599), .B2(n9594), .C1(
        P1_U3084), .C2(n9593), .ZN(P1_U3323) );
  AOI21_X1 U10800 ( .B1(n9597), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9596), .ZN(
        n9598) );
  OAI21_X1 U10801 ( .B1(n9600), .B2(n9599), .A(n9598), .ZN(P1_U3325) );
  MUX2_X1 U10802 ( .A(n9601), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10803 ( .A1(n9966), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9614) );
  AOI211_X1 U10804 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(n9606)
         );
  AOI21_X1 U10805 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9613) );
  OAI211_X1 U10806 ( .C1(n9611), .C2(n9610), .A(n9964), .B(n9609), .ZN(n9612)
         );
  NAND3_X1 U10807 ( .A1(n9614), .A2(n9613), .A3(n9612), .ZN(P2_U3247) );
  NOR2_X1 U10808 ( .A1(n9615), .A2(n10078), .ZN(n9620) );
  OAI22_X1 U10809 ( .A1(n9617), .A2(n10065), .B1(n9616), .B2(n10063), .ZN(
        n9618) );
  AOI211_X1 U10810 ( .C1(n9620), .C2(n8194), .A(n9619), .B(n9618), .ZN(n9622)
         );
  AOI22_X1 U10811 ( .A1(n10097), .A2(n9622), .B1(n6257), .B2(n10095), .ZN(
        P2_U3533) );
  INV_X1 U10812 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9621) );
  AOI22_X1 U10813 ( .A1(n10083), .A2(n9622), .B1(n9621), .B2(n10081), .ZN(
        P2_U3490) );
  INV_X1 U10814 ( .A(n9630), .ZN(n9623) );
  XNOR2_X1 U10815 ( .A(n9624), .B(n9623), .ZN(n9671) );
  AND2_X1 U10816 ( .A1(n9625), .A2(n9643), .ZN(n9626) );
  OR2_X1 U10817 ( .A1(n9626), .A2(n4587), .ZN(n9669) );
  INV_X1 U10818 ( .A(n9669), .ZN(n9627) );
  AOI22_X1 U10819 ( .A1(n9671), .A2(n9834), .B1(n9833), .B2(n9627), .ZN(n9646)
         );
  INV_X1 U10820 ( .A(n9628), .ZN(n9629) );
  OAI22_X1 U10821 ( .A1(n9874), .A2(n6736), .B1(n9629), .B2(n9847), .ZN(n9642)
         );
  XNOR2_X1 U10822 ( .A(n9631), .B(n9630), .ZN(n9637) );
  AOI22_X1 U10823 ( .A1(n9635), .A2(n9634), .B1(n9633), .B2(n9632), .ZN(n9636)
         );
  OAI21_X1 U10824 ( .B1(n9637), .B2(n9866), .A(n9636), .ZN(n9638) );
  AOI21_X1 U10825 ( .B1(n9671), .B2(n9639), .A(n9638), .ZN(n9673) );
  NOR2_X1 U10826 ( .A1(n9673), .A2(n9640), .ZN(n9641) );
  AOI211_X1 U10827 ( .C1(n9644), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9645)
         );
  NAND2_X1 U10828 ( .A1(n9646), .A2(n9645), .ZN(P1_U3280) );
  INV_X1 U10829 ( .A(n9647), .ZN(n9932) );
  OAI211_X1 U10830 ( .C1(n9650), .C2(n9932), .A(n9649), .B(n9648), .ZN(n9651)
         );
  AOI21_X1 U10831 ( .B1(n9924), .B2(n9652), .A(n9651), .ZN(n9676) );
  AOI22_X1 U10832 ( .A1(n9948), .A2(n9676), .B1(n9653), .B2(n9957), .ZN(
        P1_U3537) );
  OAI22_X1 U10833 ( .A1(n9655), .A2(n9934), .B1(n9654), .B2(n9932), .ZN(n9657)
         );
  AOI211_X1 U10834 ( .C1(n9658), .C2(n9924), .A(n9657), .B(n9656), .ZN(n9678)
         );
  AOI22_X1 U10835 ( .A1(n9948), .A2(n9678), .B1(n9659), .B2(n9957), .ZN(
        P1_U3536) );
  NOR2_X1 U10836 ( .A1(n9661), .A2(n9660), .ZN(n9666) );
  OAI21_X1 U10837 ( .B1(n9663), .B2(n9932), .A(n9662), .ZN(n9664) );
  AOI211_X1 U10838 ( .C1(n9666), .C2(n9474), .A(n9665), .B(n9664), .ZN(n9680)
         );
  AOI22_X1 U10839 ( .A1(n9948), .A2(n9680), .B1(n9667), .B2(n9957), .ZN(
        P1_U3535) );
  OAI22_X1 U10840 ( .A1(n9669), .A2(n9934), .B1(n9668), .B2(n9932), .ZN(n9670)
         );
  AOI21_X1 U10841 ( .B1(n9671), .B2(n9939), .A(n9670), .ZN(n9672) );
  AND2_X1 U10842 ( .A1(n9673), .A2(n9672), .ZN(n9682) );
  AOI22_X1 U10843 ( .A1(n9948), .A2(n9682), .B1(n9674), .B2(n9957), .ZN(
        P1_U3534) );
  INV_X1 U10844 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U10845 ( .A1(n9906), .A2(n9676), .B1(n9675), .B2(n9940), .ZN(
        P1_U3496) );
  INV_X1 U10846 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10847 ( .A1(n9906), .A2(n9678), .B1(n9677), .B2(n9940), .ZN(
        P1_U3493) );
  INV_X1 U10848 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U10849 ( .A1(n9906), .A2(n9680), .B1(n9679), .B2(n9940), .ZN(
        P1_U3490) );
  INV_X1 U10850 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U10851 ( .A1(n9906), .A2(n9682), .B1(n9681), .B2(n9940), .ZN(
        P1_U3487) );
  XNOR2_X1 U10852 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10853 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10854 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9702) );
  OAI211_X1 U10855 ( .C1(n9685), .C2(n9684), .A(n9811), .B(n9683), .ZN(n9686)
         );
  OAI21_X1 U10856 ( .B1(n9817), .B2(n9687), .A(n9686), .ZN(n9695) );
  MUX2_X1 U10857 ( .A(n9690), .B(n9689), .S(n9688), .Z(n9693) );
  OAI211_X1 U10858 ( .C1(n9693), .C2(n5923), .A(n9692), .B(n9691), .ZN(n9717)
         );
  INV_X1 U10859 ( .A(n9717), .ZN(n9694) );
  AOI211_X1 U10860 ( .C1(n9696), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9695), .B(
        n9694), .ZN(n9701) );
  XOR2_X1 U10861 ( .A(n9698), .B(n9697), .Z(n9699) );
  NAND2_X1 U10862 ( .A1(n9806), .A2(n9699), .ZN(n9700) );
  OAI211_X1 U10863 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9702), .A(n9701), .B(
        n9700), .ZN(P1_U3243) );
  INV_X1 U10864 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U10865 ( .A1(n9790), .A2(n9703), .ZN(n9709) );
  OAI21_X1 U10866 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  NAND2_X1 U10867 ( .A1(n9811), .A2(n9707), .ZN(n9708) );
  OAI211_X1 U10868 ( .C1(n9828), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9711)
         );
  INV_X1 U10869 ( .A(n9711), .ZN(n9719) );
  OAI21_X1 U10870 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9715) );
  NAND2_X1 U10871 ( .A1(n9806), .A2(n9715), .ZN(n9716) );
  NAND4_X1 U10872 ( .A1(n9719), .A2(n9718), .A3(n9717), .A4(n9716), .ZN(
        P1_U3245) );
  INV_X1 U10873 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9740) );
  INV_X1 U10874 ( .A(n9727), .ZN(n9722) );
  NAND2_X1 U10875 ( .A1(n9790), .A2(n9722), .ZN(n9738) );
  INV_X1 U10876 ( .A(n9720), .ZN(n9721) );
  NAND3_X1 U10877 ( .A1(n9723), .A2(n9722), .A3(n9721), .ZN(n9726) );
  INV_X1 U10878 ( .A(n9724), .ZN(n9725) );
  AND2_X1 U10879 ( .A1(n9726), .A2(n9725), .ZN(n9737) );
  NAND3_X1 U10880 ( .A1(n9728), .A2(n6606), .A3(n9727), .ZN(n9729) );
  NAND3_X1 U10881 ( .A1(n9811), .A2(n9730), .A3(n9729), .ZN(n9736) );
  NAND2_X1 U10882 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  NAND3_X1 U10883 ( .A1(n9806), .A2(n9734), .A3(n9733), .ZN(n9735) );
  AND4_X1 U10884 ( .A1(n9738), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(n9739)
         );
  OAI21_X1 U10885 ( .B1(n9828), .B2(n9740), .A(n9739), .ZN(P1_U3249) );
  INV_X1 U10886 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9753) );
  AOI211_X1 U10887 ( .C1(n9743), .C2(n9742), .A(n9741), .B(n9784), .ZN(n9744)
         );
  AOI211_X1 U10888 ( .C1(n9790), .C2(n9746), .A(n9745), .B(n9744), .ZN(n9752)
         );
  AOI21_X1 U10889 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9750) );
  OR2_X1 U10890 ( .A1(n9823), .A2(n9750), .ZN(n9751) );
  OAI211_X1 U10891 ( .C1(n9753), .C2(n9828), .A(n9752), .B(n9751), .ZN(
        P1_U3254) );
  INV_X1 U10892 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9769) );
  AOI21_X1 U10893 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  NAND2_X1 U10894 ( .A1(n9811), .A2(n9757), .ZN(n9760) );
  INV_X1 U10895 ( .A(n9758), .ZN(n9759) );
  OAI211_X1 U10896 ( .C1(n9817), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9762)
         );
  INV_X1 U10897 ( .A(n9762), .ZN(n9768) );
  AOI21_X1 U10898 ( .B1(n9765), .B2(n9764), .A(n9763), .ZN(n9766) );
  OR2_X1 U10899 ( .A1(n9823), .A2(n9766), .ZN(n9767) );
  OAI211_X1 U10900 ( .C1(n9769), .C2(n9828), .A(n9768), .B(n9767), .ZN(
        P1_U3255) );
  INV_X1 U10901 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9780) );
  AOI211_X1 U10902 ( .C1(n9772), .C2(n9771), .A(n9770), .B(n9784), .ZN(n9773)
         );
  AOI211_X1 U10903 ( .C1(n9790), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9779)
         );
  OAI211_X1 U10904 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9777), .A(n9806), .B(
        n9776), .ZN(n9778) );
  OAI211_X1 U10905 ( .C1(n9828), .C2(n9780), .A(n9779), .B(n9778), .ZN(
        P1_U3256) );
  INV_X1 U10906 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9796) );
  NOR2_X1 U10907 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9781), .ZN(n9788) );
  INV_X1 U10908 ( .A(n9782), .ZN(n9783) );
  AOI211_X1 U10909 ( .C1(n9786), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9787)
         );
  AOI211_X1 U10910 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9795)
         );
  XOR2_X1 U10911 ( .A(n9792), .B(n9791), .Z(n9793) );
  NAND2_X1 U10912 ( .A1(n9793), .A2(n9806), .ZN(n9794) );
  OAI211_X1 U10913 ( .C1(n9828), .C2(n9796), .A(n9795), .B(n9794), .ZN(
        P1_U3257) );
  INV_X1 U10914 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9810) );
  OAI211_X1 U10915 ( .C1(n9799), .C2(n9798), .A(n9797), .B(n9811), .ZN(n9801)
         );
  OAI211_X1 U10916 ( .C1(n9802), .C2(n9817), .A(n9801), .B(n9800), .ZN(n9803)
         );
  INV_X1 U10917 ( .A(n9803), .ZN(n9809) );
  XOR2_X1 U10918 ( .A(n9805), .B(n9804), .Z(n9807) );
  NAND2_X1 U10919 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  OAI211_X1 U10920 ( .C1(n9828), .C2(n9810), .A(n9809), .B(n9808), .ZN(
        P1_U3258) );
  INV_X1 U10921 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9827) );
  OAI211_X1 U10922 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9816)
         );
  OAI211_X1 U10923 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9819)
         );
  INV_X1 U10924 ( .A(n9819), .ZN(n9826) );
  AOI21_X1 U10925 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9824) );
  OR2_X1 U10926 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  OAI211_X1 U10927 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(
        P1_U3259) );
  XOR2_X1 U10928 ( .A(n9829), .B(n9836), .Z(n9844) );
  INV_X1 U10929 ( .A(n9844), .ZN(n9938) );
  OAI21_X1 U10930 ( .B1(n9831), .B2(n9933), .A(n9830), .ZN(n9935) );
  INV_X1 U10931 ( .A(n9935), .ZN(n9832) );
  AOI22_X1 U10932 ( .A1(n9938), .A2(n9834), .B1(n9833), .B2(n9832), .ZN(n9853)
         );
  XOR2_X1 U10933 ( .A(n9836), .B(n9835), .Z(n9841) );
  OAI22_X1 U10934 ( .A1(n9838), .A2(n9871), .B1(n9837), .B2(n9869), .ZN(n9839)
         );
  AOI21_X1 U10935 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9842) );
  OAI21_X1 U10936 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9936) );
  NOR2_X1 U10937 ( .A1(n9845), .A2(n9933), .ZN(n9851) );
  INV_X1 U10938 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9849) );
  INV_X1 U10939 ( .A(n9846), .ZN(n9848) );
  OAI22_X1 U10940 ( .A1(n9874), .A2(n9849), .B1(n9848), .B2(n9847), .ZN(n9850)
         );
  AOI211_X1 U10941 ( .C1(n9936), .C2(n9874), .A(n9851), .B(n9850), .ZN(n9852)
         );
  NAND2_X1 U10942 ( .A1(n9853), .A2(n9852), .ZN(P1_U3282) );
  XOR2_X1 U10943 ( .A(n9854), .B(n9865), .Z(n9911) );
  OAI211_X1 U10944 ( .C1(n9857), .C2(n9908), .A(n9856), .B(n9855), .ZN(n9907)
         );
  AOI22_X1 U10945 ( .A1(n9861), .A2(n9860), .B1(n9859), .B2(n9858), .ZN(n9862)
         );
  OAI21_X1 U10946 ( .B1(n9907), .B2(n9863), .A(n9862), .ZN(n9872) );
  XOR2_X1 U10947 ( .A(n9865), .B(n9864), .Z(n9867) );
  OAI222_X1 U10948 ( .A1(n9871), .A2(n9870), .B1(n9869), .B2(n9868), .C1(n9867), .C2(n9866), .ZN(n9909) );
  AOI211_X1 U10949 ( .C1(n9873), .C2(n9911), .A(n9872), .B(n9909), .ZN(n9875)
         );
  AOI22_X1 U10950 ( .A1(n9640), .A2(n9876), .B1(n9875), .B2(n9874), .ZN(
        P1_U3286) );
  AND2_X1 U10951 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9877), .ZN(P1_U3292) );
  AND2_X1 U10952 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9877), .ZN(P1_U3293) );
  AND2_X1 U10953 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9877), .ZN(P1_U3294) );
  AND2_X1 U10954 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9877), .ZN(P1_U3295) );
  AND2_X1 U10955 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9877), .ZN(P1_U3296) );
  AND2_X1 U10956 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9877), .ZN(P1_U3297) );
  AND2_X1 U10957 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9877), .ZN(P1_U3298) );
  AND2_X1 U10958 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9877), .ZN(P1_U3299) );
  AND2_X1 U10959 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9877), .ZN(P1_U3300) );
  AND2_X1 U10960 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9877), .ZN(P1_U3301) );
  AND2_X1 U10961 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9877), .ZN(P1_U3302) );
  AND2_X1 U10962 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9877), .ZN(P1_U3303) );
  AND2_X1 U10963 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9877), .ZN(P1_U3304) );
  AND2_X1 U10964 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9877), .ZN(P1_U3305) );
  AND2_X1 U10965 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9877), .ZN(P1_U3306) );
  AND2_X1 U10966 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9877), .ZN(P1_U3307) );
  AND2_X1 U10967 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9877), .ZN(P1_U3308) );
  AND2_X1 U10968 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9877), .ZN(P1_U3309) );
  AND2_X1 U10969 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9877), .ZN(P1_U3310) );
  AND2_X1 U10970 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9877), .ZN(P1_U3311) );
  AND2_X1 U10971 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9877), .ZN(P1_U3312) );
  AND2_X1 U10972 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9877), .ZN(P1_U3313) );
  AND2_X1 U10973 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9877), .ZN(P1_U3314) );
  AND2_X1 U10974 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9877), .ZN(P1_U3315) );
  AND2_X1 U10975 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9877), .ZN(P1_U3316) );
  AND2_X1 U10976 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9877), .ZN(P1_U3317) );
  AND2_X1 U10977 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9877), .ZN(P1_U3318) );
  INV_X1 U10978 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10472) );
  NOR2_X1 U10979 ( .A1(n9878), .A2(n10472), .ZN(P1_U3319) );
  INV_X1 U10980 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U10981 ( .A1(n9878), .A2(n10338), .ZN(P1_U3320) );
  INV_X1 U10982 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10496) );
  NOR2_X1 U10983 ( .A1(n9878), .A2(n10496), .ZN(P1_U3321) );
  INV_X1 U10984 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9880) );
  AOI21_X1 U10985 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(P1_U3441) );
  INV_X1 U10986 ( .A(n9882), .ZN(n9886) );
  OAI21_X1 U10987 ( .B1(n6801), .B2(n9932), .A(n9883), .ZN(n9885) );
  AOI211_X1 U10988 ( .C1(n9939), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9942)
         );
  INV_X1 U10989 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9887) );
  AOI22_X1 U10990 ( .A1(n9906), .A2(n9942), .B1(n9887), .B2(n9940), .ZN(
        P1_U3457) );
  OAI22_X1 U10991 ( .A1(n9889), .A2(n9934), .B1(n9888), .B2(n9932), .ZN(n9891)
         );
  AOI211_X1 U10992 ( .C1(n9939), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9944)
         );
  INV_X1 U10993 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U10994 ( .A1(n9906), .A2(n9944), .B1(n9893), .B2(n9940), .ZN(
        P1_U3460) );
  OAI22_X1 U10995 ( .A1(n9895), .A2(n9934), .B1(n9894), .B2(n9932), .ZN(n9897)
         );
  AOI211_X1 U10996 ( .C1(n9939), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9945)
         );
  INV_X1 U10997 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10998 ( .A1(n9906), .A2(n9945), .B1(n9899), .B2(n9940), .ZN(
        P1_U3463) );
  OAI22_X1 U10999 ( .A1(n9901), .A2(n9934), .B1(n9900), .B2(n9932), .ZN(n9903)
         );
  AOI211_X1 U11000 ( .C1(n9939), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9947)
         );
  INV_X1 U11001 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U11002 ( .A1(n9906), .A2(n9947), .B1(n9905), .B2(n9940), .ZN(
        P1_U3466) );
  OAI21_X1 U11003 ( .B1(n9908), .B2(n9932), .A(n9907), .ZN(n9910) );
  AOI211_X1 U11004 ( .C1(n9924), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9950)
         );
  INV_X1 U11005 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U11006 ( .A1(n9906), .A2(n9950), .B1(n9912), .B2(n9940), .ZN(
        P1_U3469) );
  OAI22_X1 U11007 ( .A1(n9914), .A2(n9934), .B1(n9913), .B2(n9932), .ZN(n9916)
         );
  AOI211_X1 U11008 ( .C1(n9939), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9952)
         );
  INV_X1 U11009 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U11010 ( .A1(n9906), .A2(n9952), .B1(n9918), .B2(n9940), .ZN(
        P1_U3472) );
  OAI21_X1 U11011 ( .B1(n9920), .B2(n9932), .A(n9919), .ZN(n9922) );
  AOI211_X1 U11012 ( .C1(n9924), .C2(n9923), .A(n9922), .B(n9921), .ZN(n9954)
         );
  INV_X1 U11013 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U11014 ( .A1(n9906), .A2(n9954), .B1(n9925), .B2(n9940), .ZN(
        P1_U3475) );
  OAI21_X1 U11015 ( .B1(n9927), .B2(n9932), .A(n9926), .ZN(n9929) );
  AOI211_X1 U11016 ( .C1(n9939), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9956)
         );
  INV_X1 U11017 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U11018 ( .A1(n9906), .A2(n9956), .B1(n9931), .B2(n9940), .ZN(
        P1_U3478) );
  OAI22_X1 U11019 ( .A1(n9935), .A2(n9934), .B1(n9933), .B2(n9932), .ZN(n9937)
         );
  AOI211_X1 U11020 ( .C1(n9939), .C2(n9938), .A(n9937), .B(n9936), .ZN(n9959)
         );
  INV_X1 U11021 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U11022 ( .A1(n9906), .A2(n9959), .B1(n9941), .B2(n9940), .ZN(
        P1_U3481) );
  AOI22_X1 U11023 ( .A1(n9948), .A2(n9942), .B1(n6501), .B2(n9957), .ZN(
        P1_U3524) );
  AOI22_X1 U11024 ( .A1(n9948), .A2(n9944), .B1(n9943), .B2(n9957), .ZN(
        P1_U3525) );
  AOI22_X1 U11025 ( .A1(n9948), .A2(n9945), .B1(n6500), .B2(n9957), .ZN(
        P1_U3526) );
  AOI22_X1 U11026 ( .A1(n9948), .A2(n9947), .B1(n9946), .B2(n9957), .ZN(
        P1_U3527) );
  AOI22_X1 U11027 ( .A1(n9948), .A2(n9950), .B1(n9949), .B2(n9957), .ZN(
        P1_U3528) );
  AOI22_X1 U11028 ( .A1(n9948), .A2(n9952), .B1(n9951), .B2(n9957), .ZN(
        P1_U3529) );
  AOI22_X1 U11029 ( .A1(n9948), .A2(n9954), .B1(n9953), .B2(n9957), .ZN(
        P1_U3530) );
  AOI22_X1 U11030 ( .A1(n9948), .A2(n9956), .B1(n9955), .B2(n9957), .ZN(
        P1_U3531) );
  AOI22_X1 U11031 ( .A1(n9948), .A2(n9959), .B1(n9958), .B2(n9957), .ZN(
        P1_U3532) );
  OAI211_X1 U11032 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9962), .A(n9961), .B(
        n9960), .ZN(n9963) );
  AOI21_X1 U11033 ( .B1(n9965), .B2(n6049), .A(n9963), .ZN(n9970) );
  AOI22_X1 U11034 ( .A1(n9965), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9964), .ZN(n9969) );
  AOI22_X1 U11035 ( .A1(n9966), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9967) );
  OAI221_X1 U11036 ( .B1(n9970), .B2(n9969), .C1(n9970), .C2(n9968), .A(n9967), 
        .ZN(P2_U3245) );
  INV_X1 U11037 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9984) );
  INV_X1 U11038 ( .A(n9971), .ZN(n9979) );
  INV_X1 U11039 ( .A(n9972), .ZN(n9978) );
  INV_X1 U11040 ( .A(n9973), .ZN(n9976) );
  AOI22_X1 U11041 ( .A1(n9991), .A2(n9976), .B1(n9975), .B2(n9974), .ZN(n9977)
         );
  OAI211_X1 U11042 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(n9981)
         );
  AOI21_X1 U11043 ( .B1(n9986), .B2(n9982), .A(n9981), .ZN(n9983) );
  AOI22_X1 U11044 ( .A1(n8496), .A2(n9984), .B1(n9983), .B2(n9993), .ZN(
        P2_U3291) );
  NAND2_X1 U11045 ( .A1(n6761), .A2(n9985), .ZN(n10010) );
  OAI21_X1 U11046 ( .B1(n9986), .B2(n10004), .A(n10010), .ZN(n9987) );
  AND2_X1 U11047 ( .A1(n9987), .A2(n10005), .ZN(n9994) );
  AOI21_X1 U11048 ( .B1(n9989), .B2(n9988), .A(n10007), .ZN(n9990) );
  AOI21_X1 U11049 ( .B1(n9991), .B2(P2_REG3_REG_0__SCAN_IN), .A(n9990), .ZN(
        n9992) );
  OAI221_X1 U11050 ( .B1(n8289), .B2(n9994), .C1(n9993), .C2(n6049), .A(n9992), 
        .ZN(P2_U3296) );
  INV_X1 U11051 ( .A(n9995), .ZN(n9997) );
  NAND2_X1 U11052 ( .A1(n9997), .A2(n9996), .ZN(n10000) );
  AND2_X1 U11053 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10000), .ZN(P2_U3297) );
  AND2_X1 U11054 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10000), .ZN(P2_U3298) );
  AND2_X1 U11055 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10000), .ZN(P2_U3299) );
  AND2_X1 U11056 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10000), .ZN(P2_U3300) );
  AND2_X1 U11057 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10000), .ZN(P2_U3301) );
  AND2_X1 U11058 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10000), .ZN(P2_U3302) );
  AND2_X1 U11059 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10000), .ZN(P2_U3303) );
  AND2_X1 U11060 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10000), .ZN(P2_U3304) );
  AND2_X1 U11061 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10000), .ZN(P2_U3305) );
  AND2_X1 U11062 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10000), .ZN(P2_U3306) );
  AND2_X1 U11063 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10000), .ZN(P2_U3307) );
  AND2_X1 U11064 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10000), .ZN(P2_U3308) );
  AND2_X1 U11065 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10000), .ZN(P2_U3309) );
  AND2_X1 U11066 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10000), .ZN(P2_U3310) );
  AND2_X1 U11067 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10000), .ZN(P2_U3311) );
  AND2_X1 U11068 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10000), .ZN(P2_U3312) );
  AND2_X1 U11069 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10000), .ZN(P2_U3313) );
  AND2_X1 U11070 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10000), .ZN(P2_U3314) );
  AND2_X1 U11071 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10000), .ZN(P2_U3315) );
  AND2_X1 U11072 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10000), .ZN(P2_U3316) );
  AND2_X1 U11073 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10000), .ZN(P2_U3317) );
  AND2_X1 U11074 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10000), .ZN(P2_U3318) );
  AND2_X1 U11075 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10000), .ZN(P2_U3319) );
  AND2_X1 U11076 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10000), .ZN(P2_U3320) );
  AND2_X1 U11077 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10000), .ZN(P2_U3321) );
  AND2_X1 U11078 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10000), .ZN(P2_U3322) );
  AND2_X1 U11079 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10000), .ZN(P2_U3323) );
  AND2_X1 U11080 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10000), .ZN(P2_U3324) );
  AND2_X1 U11081 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10000), .ZN(P2_U3325) );
  AND2_X1 U11082 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10000), .ZN(P2_U3326) );
  AOI22_X1 U11083 ( .A1(n9999), .A2(n10000), .B1(n10003), .B2(n9998), .ZN(
        P2_U3437) );
  AOI22_X1 U11084 ( .A1(n10003), .A2(n10002), .B1(n10001), .B2(n10000), .ZN(
        P2_U3438) );
  NAND2_X1 U11085 ( .A1(n10010), .A2(n10004), .ZN(n10006) );
  OAI211_X1 U11086 ( .C1(n10008), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10009) );
  AOI21_X1 U11087 ( .B1(n10069), .B2(n10010), .A(n10009), .ZN(n10085) );
  AOI22_X1 U11088 ( .A1(n10083), .A2(n10085), .B1(n6050), .B2(n10081), .ZN(
        P2_U3451) );
  OAI22_X1 U11089 ( .A1(n10012), .A2(n10065), .B1(n10011), .B2(n10063), .ZN(
        n10014) );
  AOI211_X1 U11090 ( .C1(n10069), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10086) );
  AOI22_X1 U11091 ( .A1(n10083), .A2(n10086), .B1(n6062), .B2(n10081), .ZN(
        P2_U3457) );
  INV_X1 U11092 ( .A(n10056), .ZN(n10039) );
  NAND2_X1 U11093 ( .A1(n10021), .A2(n10039), .ZN(n10017) );
  OAI211_X1 U11094 ( .C1(n10018), .C2(n10063), .A(n10017), .B(n10016), .ZN(
        n10019) );
  AOI211_X1 U11095 ( .C1(n10061), .C2(n10021), .A(n10020), .B(n10019), .ZN(
        n10087) );
  AOI22_X1 U11096 ( .A1(n10083), .A2(n10087), .B1(n6073), .B2(n10081), .ZN(
        P2_U3460) );
  OAI21_X1 U11097 ( .B1(n10023), .B2(n10063), .A(n10022), .ZN(n10025) );
  AOI211_X1 U11098 ( .C1(n10069), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10088) );
  INV_X1 U11099 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11100 ( .A1(n10083), .A2(n10088), .B1(n10027), .B2(n10081), .ZN(
        P2_U3463) );
  OAI211_X1 U11101 ( .C1(n10030), .C2(n10063), .A(n10029), .B(n10028), .ZN(
        n10031) );
  AOI21_X1 U11102 ( .B1(n10069), .B2(n10032), .A(n10031), .ZN(n10089) );
  AOI22_X1 U11103 ( .A1(n10083), .A2(n10089), .B1(n6116), .B2(n10081), .ZN(
        P2_U3469) );
  NAND2_X1 U11104 ( .A1(n10033), .A2(n10073), .ZN(n10034) );
  OAI211_X1 U11105 ( .C1(n10065), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10037) );
  AOI21_X1 U11106 ( .B1(n10038), .B2(n10069), .A(n10037), .ZN(n10090) );
  AOI22_X1 U11107 ( .A1(n10083), .A2(n10090), .B1(n6135), .B2(n10081), .ZN(
        P2_U3472) );
  AND2_X1 U11108 ( .A1(n10040), .A2(n10039), .ZN(n10044) );
  OAI22_X1 U11109 ( .A1(n10042), .A2(n10065), .B1(n10041), .B2(n10063), .ZN(
        n10043) );
  NOR3_X1 U11110 ( .A1(n10045), .A2(n10044), .A3(n10043), .ZN(n10091) );
  AOI22_X1 U11111 ( .A1(n10083), .A2(n10091), .B1(n6155), .B2(n10081), .ZN(
        P2_U3475) );
  INV_X1 U11112 ( .A(n10052), .ZN(n10050) );
  AOI21_X1 U11113 ( .B1(n10073), .B2(n10047), .A(n10046), .ZN(n10048) );
  OAI211_X1 U11114 ( .C1(n10050), .C2(n10056), .A(n10049), .B(n10048), .ZN(
        n10051) );
  AOI21_X1 U11115 ( .B1(n10061), .B2(n10052), .A(n10051), .ZN(n10092) );
  AOI22_X1 U11116 ( .A1(n10083), .A2(n10092), .B1(n6176), .B2(n10081), .ZN(
        P2_U3478) );
  OAI211_X1 U11117 ( .C1(n10055), .C2(n10063), .A(n10054), .B(n10053), .ZN(
        n10059) );
  INV_X1 U11118 ( .A(n10060), .ZN(n10057) );
  NOR2_X1 U11119 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  AOI211_X1 U11120 ( .C1(n10061), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10093) );
  AOI22_X1 U11121 ( .A1(n10083), .A2(n10093), .B1(n6204), .B2(n10081), .ZN(
        P2_U3481) );
  INV_X1 U11122 ( .A(n10062), .ZN(n10070) );
  OAI22_X1 U11123 ( .A1(n10066), .A2(n10065), .B1(n10064), .B2(n10063), .ZN(
        n10067) );
  AOI211_X1 U11124 ( .C1(n10070), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10094) );
  INV_X1 U11125 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U11126 ( .A1(n10083), .A2(n10094), .B1(n10071), .B2(n10081), .ZN(
        P2_U3484) );
  AOI22_X1 U11127 ( .A1(n10075), .A2(n10074), .B1(n10073), .B2(n10072), .ZN(
        n10076) );
  OAI211_X1 U11128 ( .C1(n10079), .C2(n10078), .A(n10077), .B(n10076), .ZN(
        n10080) );
  INV_X1 U11129 ( .A(n10080), .ZN(n10096) );
  INV_X1 U11130 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11131 ( .A1(n10083), .A2(n10096), .B1(n10082), .B2(n10081), .ZN(
        P2_U3487) );
  AOI22_X1 U11132 ( .A1(n10097), .A2(n10085), .B1(n10084), .B2(n10095), .ZN(
        P2_U3520) );
  AOI22_X1 U11133 ( .A1(n10097), .A2(n10086), .B1(n7134), .B2(n10095), .ZN(
        P2_U3522) );
  AOI22_X1 U11134 ( .A1(n10097), .A2(n10087), .B1(n7129), .B2(n10095), .ZN(
        P2_U3523) );
  AOI22_X1 U11135 ( .A1(n10097), .A2(n10088), .B1(n7128), .B2(n10095), .ZN(
        P2_U3524) );
  AOI22_X1 U11136 ( .A1(n10097), .A2(n10089), .B1(n7172), .B2(n10095), .ZN(
        P2_U3526) );
  AOI22_X1 U11137 ( .A1(n10097), .A2(n10090), .B1(n7170), .B2(n10095), .ZN(
        P2_U3527) );
  AOI22_X1 U11138 ( .A1(n10097), .A2(n10091), .B1(n7169), .B2(n10095), .ZN(
        P2_U3528) );
  AOI22_X1 U11139 ( .A1(n10097), .A2(n10092), .B1(n7168), .B2(n10095), .ZN(
        P2_U3529) );
  AOI22_X1 U11140 ( .A1(n10097), .A2(n10093), .B1(n7179), .B2(n10095), .ZN(
        P2_U3530) );
  AOI22_X1 U11141 ( .A1(n10097), .A2(n10094), .B1(n7271), .B2(n10095), .ZN(
        P2_U3531) );
  AOI22_X1 U11142 ( .A1(n10097), .A2(n10096), .B1(n7275), .B2(n10095), .ZN(
        P2_U3532) );
  NAND3_X1 U11143 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10100) );
  AND2_X1 U11144 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10098) );
  NOR2_X1 U11145 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10098), .ZN(n10099) );
  INV_X1 U11146 ( .A(n10099), .ZN(n10116) );
  NAND2_X1 U11147 ( .A1(n10101), .A2(n10100), .ZN(n10115) );
  OAI222_X1 U11148 ( .A1(n10101), .A2(n10100), .B1(n10101), .B2(n10116), .C1(
        n10099), .C2(n10115), .ZN(ADD_1071_U5) );
  XOR2_X1 U11149 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NOR2_X1 U11150 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n10102) );
  AOI21_X1 U11151 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10102), .ZN(n10121) );
  NOR2_X1 U11152 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n10103) );
  AOI21_X1 U11153 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10103), .ZN(n10124) );
  NOR2_X1 U11154 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n10104) );
  AOI21_X1 U11155 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10104), .ZN(n10127) );
  NOR2_X1 U11156 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10105) );
  AOI21_X1 U11157 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10105), .ZN(n10130) );
  NOR2_X1 U11158 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10106) );
  AOI21_X1 U11159 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10106), .ZN(n10133) );
  NOR2_X1 U11160 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10107) );
  AOI21_X1 U11161 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10107), .ZN(n10136) );
  NOR2_X1 U11162 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10108) );
  AOI21_X1 U11163 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10108), .ZN(n10139) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10109) );
  AOI21_X1 U11165 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10109), .ZN(n10142) );
  NOR2_X1 U11166 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n10110) );
  AOI21_X1 U11167 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10110), .ZN(n10526) );
  NOR2_X1 U11168 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n10111) );
  AOI21_X1 U11169 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10111), .ZN(n10541) );
  NOR2_X1 U11170 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10112) );
  AOI21_X1 U11171 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10112), .ZN(n10529) );
  NOR2_X1 U11172 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10113) );
  AOI21_X1 U11173 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10113), .ZN(n10544) );
  NOR2_X1 U11174 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10114) );
  AOI21_X1 U11175 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10114), .ZN(n10535) );
  NAND2_X1 U11176 ( .A1(n10116), .A2(n10115), .ZN(n10532) );
  NAND2_X1 U11177 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10117) );
  OAI21_X1 U11178 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10117), .ZN(n10531) );
  NOR2_X1 U11179 ( .A1(n10532), .A2(n10531), .ZN(n10530) );
  AOI21_X1 U11180 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10530), .ZN(n10547) );
  NAND2_X1 U11181 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10118) );
  OAI21_X1 U11182 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10118), .ZN(n10546) );
  NOR2_X1 U11183 ( .A1(n10547), .A2(n10546), .ZN(n10545) );
  AOI21_X1 U11184 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10545), .ZN(n10550) );
  NOR2_X1 U11185 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10119) );
  AOI21_X1 U11186 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10119), .ZN(n10549) );
  NAND2_X1 U11187 ( .A1(n10550), .A2(n10549), .ZN(n10548) );
  OAI21_X1 U11188 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10548), .ZN(n10534) );
  NAND2_X1 U11189 ( .A1(n10535), .A2(n10534), .ZN(n10533) );
  OAI21_X1 U11190 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10533), .ZN(n10543) );
  NAND2_X1 U11191 ( .A1(n10544), .A2(n10543), .ZN(n10542) );
  OAI21_X1 U11192 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10542), .ZN(n10528) );
  NAND2_X1 U11193 ( .A1(n10529), .A2(n10528), .ZN(n10527) );
  OAI21_X1 U11194 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10527), .ZN(n10540) );
  NAND2_X1 U11195 ( .A1(n10541), .A2(n10540), .ZN(n10539) );
  OAI21_X1 U11196 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10539), .ZN(n10525) );
  NAND2_X1 U11197 ( .A1(n10526), .A2(n10525), .ZN(n10524) );
  OAI21_X1 U11198 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10524), .ZN(n10141) );
  NAND2_X1 U11199 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U11200 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10140), .ZN(n10138) );
  NAND2_X1 U11201 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  OAI21_X1 U11202 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10137), .ZN(n10135) );
  NAND2_X1 U11203 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U11204 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10134), .ZN(n10132) );
  NAND2_X1 U11205 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  OAI21_X1 U11206 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10131), .ZN(n10129) );
  NAND2_X1 U11207 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  OAI21_X1 U11208 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10128), .ZN(n10126) );
  NAND2_X1 U11209 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  OAI21_X1 U11210 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10125), .ZN(n10123) );
  NAND2_X1 U11211 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  OAI21_X1 U11212 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10122), .ZN(n10120) );
  NAND2_X1 U11213 ( .A1(n10121), .A2(n10120), .ZN(n10144) );
  OAI21_X1 U11214 ( .B1(n10121), .B2(n10120), .A(n10144), .ZN(ADD_1071_U56) );
  OAI21_X1 U11215 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(ADD_1071_U57) );
  OAI21_X1 U11216 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1071_U58) );
  OAI21_X1 U11217 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(ADD_1071_U59) );
  OAI21_X1 U11218 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(ADD_1071_U60) );
  OAI21_X1 U11219 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(ADD_1071_U61) );
  OAI21_X1 U11220 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(ADD_1071_U62) );
  OAI21_X1 U11221 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1071_U63) );
  NOR2_X1 U11222 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .ZN(n10143) );
  AOI21_X1 U11223 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10143), .ZN(n10538) );
  OAI21_X1 U11224 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10144), .ZN(n10537) );
  NAND2_X1 U11225 ( .A1(n10538), .A2(n10537), .ZN(n10536) );
  OAI21_X1 U11226 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10536), .ZN(n10523) );
  OAI22_X1 U11227 ( .A1(SI_16_), .A2(keyinput_g16), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n10145) );
  AOI221_X1 U11228 ( .B1(SI_16_), .B2(keyinput_g16), .C1(keyinput_g29), .C2(
        SI_3_), .A(n10145), .ZN(n10152) );
  OAI22_X1 U11229 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g94), .B1(
        keyinput_g14), .B2(SI_18_), .ZN(n10146) );
  AOI221_X1 U11230 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .C1(SI_18_), 
        .C2(keyinput_g14), .A(n10146), .ZN(n10151) );
  OAI22_X1 U11231 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_g122), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n10147) );
  AOI221_X1 U11232 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g79), .C2(P2_DATAO_REG_17__SCAN_IN), .A(n10147), .ZN(n10150)
         );
  OAI22_X1 U11233 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n10148) );
  AOI221_X1 U11234 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g61), .C2(P2_REG3_REG_6__SCAN_IN), .A(n10148), .ZN(n10149) );
  NAND4_X1 U11235 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10180) );
  OAI22_X1 U11236 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10153) );
  AOI221_X1 U11237 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        keyinput_g60), .C2(P2_REG3_REG_18__SCAN_IN), .A(n10153), .ZN(n10160)
         );
  OAI22_X1 U11238 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n10154) );
  AOI221_X1 U11239 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10154), .ZN(n10159)
         );
  OAI22_X1 U11240 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g126), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput_g121), .ZN(n10155) );
  AOI221_X1 U11241 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g121), .C2(P1_IR_REG_30__SCAN_IN), .A(n10155), .ZN(n10158) );
  OAI22_X1 U11242 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10156) );
  AOI221_X1 U11243 ( .B1(SI_23_), .B2(keyinput_g9), .C1(keyinput_g56), .C2(
        P2_REG3_REG_13__SCAN_IN), .A(n10156), .ZN(n10157) );
  NAND4_X1 U11244 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10179) );
  OAI22_X1 U11245 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_g92), .B1(
        keyinput_g33), .B2(P2_RD_REG_SCAN_IN), .ZN(n10161) );
  AOI221_X1 U11246 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_g92), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n10161), .ZN(n10168) );
  OAI22_X1 U11247 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g106), .B1(
        keyinput_g75), .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n10162) );
  AOI221_X1 U11248 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g106), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n10162), .ZN(n10167)
         );
  OAI22_X1 U11249 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        keyinput_g46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n10163) );
  AOI221_X1 U11250 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n10163), .ZN(n10166)
         );
  OAI22_X1 U11251 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g93), .B1(
        keyinput_g74), .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10164) );
  AOI221_X1 U11252 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n10164), .ZN(n10165)
         );
  NAND4_X1 U11253 ( .A1(n10168), .A2(n10167), .A3(n10166), .A4(n10165), .ZN(
        n10178) );
  OAI22_X1 U11254 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g58), .B2(P2_REG3_REG_11__SCAN_IN), .ZN(n10169) );
  AOI221_X1 U11255 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10169), .ZN(n10176)
         );
  OAI22_X1 U11256 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g104), .B1(SI_20_), .B2(keyinput_g12), .ZN(n10170) );
  AOI221_X1 U11257 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g12), .C2(SI_20_), .A(n10170), .ZN(n10175) );
  OAI22_X1 U11258 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_g71), .B1(
        keyinput_g55), .B2(P2_REG3_REG_20__SCAN_IN), .ZN(n10171) );
  AOI221_X1 U11259 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n10171), .ZN(n10174)
         );
  OAI22_X1 U11260 ( .A1(SI_12_), .A2(keyinput_g20), .B1(keyinput_g0), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10172) );
  AOI221_X1 U11261 ( .B1(SI_12_), .B2(keyinput_g20), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_g0), .A(n10172), .ZN(n10173) );
  NAND4_X1 U11262 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NOR4_X1 U11263 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10519) );
  OAI22_X1 U11264 ( .A1(SI_17_), .A2(keyinput_g15), .B1(keyinput_g53), .B2(
        P2_REG3_REG_9__SCAN_IN), .ZN(n10181) );
  AOI221_X1 U11265 ( .B1(SI_17_), .B2(keyinput_g15), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n10181), .ZN(n10188) );
  OAI22_X1 U11266 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g111), .B1(
        keyinput_g70), .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10182) );
  AOI221_X1 U11267 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g111), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_g70), .A(n10182), .ZN(n10187)
         );
  OAI22_X1 U11268 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_g117), .B1(
        keyinput_g13), .B2(SI_19_), .ZN(n10183) );
  AOI221_X1 U11269 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_g117), .C1(
        SI_19_), .C2(keyinput_g13), .A(n10183), .ZN(n10186) );
  OAI22_X1 U11270 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g124), .B1(SI_0_), 
        .B2(keyinput_g32), .ZN(n10184) );
  AOI221_X1 U11271 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g32), .C2(SI_0_), .A(n10184), .ZN(n10185) );
  NAND4_X1 U11272 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10311) );
  OAI22_X1 U11273 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g114), .B1(
        keyinput_g44), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10189) );
  AOI221_X1 U11274 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n10189), .ZN(n10214) );
  OAI22_X1 U11275 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g103), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n10190) );
  AOI221_X1 U11276 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g40), .C2(P2_REG3_REG_3__SCAN_IN), .A(n10190), .ZN(n10193) );
  OAI22_X1 U11277 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g113), .B1(
        keyinput_g63), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n10191) );
  AOI221_X1 U11278 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g113), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n10191), .ZN(n10192)
         );
  OAI211_X1 U11279 ( .C1(n10472), .C2(keyinput_g127), .A(n10193), .B(n10192), 
        .ZN(n10194) );
  AOI21_X1 U11280 ( .B1(n10472), .B2(keyinput_g127), .A(n10194), .ZN(n10213)
         );
  AOI22_X1 U11281 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .ZN(n10195) );
  OAI221_X1 U11282 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n10195), .ZN(n10202)
         );
  AOI22_X1 U11283 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P1_D_REG_0__SCAN_IN), 
        .B2(keyinput_g123), .ZN(n10196) );
  OAI221_X1 U11284 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P1_D_REG_0__SCAN_IN), 
        .C2(keyinput_g123), .A(n10196), .ZN(n10201) );
  AOI22_X1 U11285 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_g100), .ZN(n10197) );
  OAI221_X1 U11286 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_g100), .A(n10197), .ZN(n10200) );
  AOI22_X1 U11287 ( .A1(SI_7_), .A2(keyinput_g25), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .ZN(n10198) );
  OAI221_X1 U11288 ( .B1(SI_7_), .B2(keyinput_g25), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_g81), .A(n10198), .ZN(n10199)
         );
  NOR4_X1 U11289 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10212) );
  AOI22_X1 U11290 ( .A1(SI_21_), .A2(keyinput_g11), .B1(P1_IR_REG_25__SCAN_IN), 
        .B2(keyinput_g116), .ZN(n10203) );
  OAI221_X1 U11291 ( .B1(SI_21_), .B2(keyinput_g11), .C1(P1_IR_REG_25__SCAN_IN), .C2(keyinput_g116), .A(n10203), .ZN(n10210) );
  AOI22_X1 U11292 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P1_IR_REG_27__SCAN_IN), 
        .B2(keyinput_g118), .ZN(n10204) );
  OAI221_X1 U11293 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P1_IR_REG_27__SCAN_IN), 
        .C2(keyinput_g118), .A(n10204), .ZN(n10209) );
  AOI22_X1 U11294 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P1_IR_REG_0__SCAN_IN), 
        .B2(keyinput_g91), .ZN(n10205) );
  OAI221_X1 U11295 ( .B1(SI_30_), .B2(keyinput_g2), .C1(P1_IR_REG_0__SCAN_IN), 
        .C2(keyinput_g91), .A(n10205), .ZN(n10208) );
  AOI22_X1 U11296 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g99), .ZN(n10206) );
  OAI221_X1 U11297 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g99), .A(n10206), .ZN(n10207) );
  NOR4_X1 U11298 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10211) );
  NAND4_X1 U11299 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10310) );
  AOI22_X1 U11300 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P1_IR_REG_10__SCAN_IN), 
        .B2(keyinput_g101), .ZN(n10215) );
  OAI221_X1 U11301 ( .B1(SI_10_), .B2(keyinput_g22), .C1(P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n10215), .ZN(n10223) );
  AOI22_X1 U11302 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(SI_2_), .B2(keyinput_g30), .ZN(n10216) );
  OAI221_X1 U11303 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        SI_2_), .C2(keyinput_g30), .A(n10216), .ZN(n10222) );
  AOI22_X1 U11304 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_g96), .ZN(n10217) );
  OAI221_X1 U11305 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_g96), .A(n10217), .ZN(n10221) );
  INV_X1 U11306 ( .A(SI_11_), .ZN(n10219) );
  AOI22_X1 U11307 ( .A1(n10219), .A2(keyinput_g21), .B1(keyinput_g47), .B2(
        n10473), .ZN(n10218) );
  OAI221_X1 U11308 ( .B1(n10219), .B2(keyinput_g21), .C1(n10473), .C2(
        keyinput_g47), .A(n10218), .ZN(n10220) );
  NOR4_X1 U11309 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10259) );
  AOI22_X1 U11310 ( .A1(n5766), .A2(keyinput_g73), .B1(keyinput_g52), .B2(
        n10356), .ZN(n10224) );
  OAI221_X1 U11311 ( .B1(n5766), .B2(keyinput_g73), .C1(n10356), .C2(
        keyinput_g52), .A(n10224), .ZN(n10232) );
  AOI22_X1 U11312 ( .A1(n10470), .A2(keyinput_g39), .B1(n10455), .B2(
        keyinput_g45), .ZN(n10225) );
  OAI221_X1 U11313 ( .B1(n10470), .B2(keyinput_g39), .C1(n10455), .C2(
        keyinput_g45), .A(n10225), .ZN(n10231) );
  XNOR2_X1 U11314 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_g69), .ZN(n10229) );
  XNOR2_X1 U11315 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g109), .ZN(n10228)
         );
  XNOR2_X1 U11316 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g110), .ZN(n10227)
         );
  XNOR2_X1 U11317 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_g108), .ZN(n10226)
         );
  NAND4_X1 U11318 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10230) );
  NOR3_X1 U11319 ( .A1(n10232), .A2(n10231), .A3(n10230), .ZN(n10258) );
  AOI22_X1 U11320 ( .A1(n10380), .A2(keyinput_g51), .B1(keyinput_g54), .B2(
        n10234), .ZN(n10233) );
  OAI221_X1 U11321 ( .B1(n10380), .B2(keyinput_g51), .C1(n10234), .C2(
        keyinput_g54), .A(n10233), .ZN(n10243) );
  AOI22_X1 U11322 ( .A1(n10236), .A2(keyinput_g83), .B1(n10324), .B2(
        keyinput_g6), .ZN(n10235) );
  OAI221_X1 U11323 ( .B1(n10236), .B2(keyinput_g83), .C1(n10324), .C2(
        keyinput_g6), .A(n10235), .ZN(n10242) );
  INV_X1 U11324 ( .A(SI_24_), .ZN(n10327) );
  AOI22_X1 U11325 ( .A1(n10327), .A2(keyinput_g8), .B1(keyinput_g66), .B2(
        n10427), .ZN(n10237) );
  OAI221_X1 U11326 ( .B1(n10327), .B2(keyinput_g8), .C1(n10427), .C2(
        keyinput_g66), .A(n10237), .ZN(n10241) );
  AOI22_X1 U11327 ( .A1(n10330), .A2(keyinput_g77), .B1(keyinput_g87), .B2(
        n10239), .ZN(n10238) );
  OAI221_X1 U11328 ( .B1(n10330), .B2(keyinput_g77), .C1(n10239), .C2(
        keyinput_g87), .A(n10238), .ZN(n10240) );
  NOR4_X1 U11329 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10257) );
  AOI22_X1 U11330 ( .A1(n10323), .A2(keyinput_g90), .B1(n10245), .B2(
        keyinput_g82), .ZN(n10244) );
  OAI221_X1 U11331 ( .B1(n10323), .B2(keyinput_g90), .C1(n10245), .C2(
        keyinput_g82), .A(n10244), .ZN(n10255) );
  AOI22_X1 U11332 ( .A1(n10248), .A2(keyinput_g18), .B1(n10247), .B2(
        keyinput_g105), .ZN(n10246) );
  OAI221_X1 U11333 ( .B1(n10248), .B2(keyinput_g18), .C1(n10247), .C2(
        keyinput_g105), .A(n10246), .ZN(n10254) );
  XNOR2_X1 U11334 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10252) );
  XNOR2_X1 U11335 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_g80), .ZN(n10251) );
  XNOR2_X1 U11336 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g120), .ZN(n10250)
         );
  XNOR2_X1 U11337 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n10249) );
  NAND4_X1 U11338 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10253) );
  NOR3_X1 U11339 ( .A1(n10255), .A2(n10254), .A3(n10253), .ZN(n10256) );
  NAND4_X1 U11340 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10309) );
  AOI22_X1 U11341 ( .A1(n10326), .A2(keyinput_g78), .B1(keyinput_g41), .B2(
        n10426), .ZN(n10260) );
  OAI221_X1 U11342 ( .B1(n10326), .B2(keyinput_g78), .C1(n10426), .C2(
        keyinput_g41), .A(n10260), .ZN(n10264) );
  XNOR2_X1 U11343 ( .A(n10261), .B(keyinput_g97), .ZN(n10263) );
  XNOR2_X1 U11344 ( .A(n10460), .B(keyinput_g62), .ZN(n10262) );
  NOR3_X1 U11345 ( .A1(n10264), .A2(n10263), .A3(n10262), .ZN(n10268) );
  XNOR2_X1 U11346 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g102), .ZN(n10267)
         );
  XNOR2_X1 U11347 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g107), .ZN(n10266)
         );
  XNOR2_X1 U11348 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_g84), .ZN(n10265) );
  NAND4_X1 U11349 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10270) );
  XNOR2_X1 U11350 ( .A(n10496), .B(keyinput_g125), .ZN(n10269) );
  NOR2_X1 U11351 ( .A1(n10270), .A2(n10269), .ZN(n10307) );
  INV_X1 U11352 ( .A(SI_31_), .ZN(n10272) );
  AOI22_X1 U11353 ( .A1(n10273), .A2(keyinput_g89), .B1(keyinput_g1), .B2(
        n10272), .ZN(n10271) );
  OAI221_X1 U11354 ( .B1(n10273), .B2(keyinput_g89), .C1(n10272), .C2(
        keyinput_g1), .A(n10271), .ZN(n10282) );
  AOI22_X1 U11355 ( .A1(n6137), .A2(keyinput_g35), .B1(n10442), .B2(
        keyinput_g24), .ZN(n10274) );
  OAI221_X1 U11356 ( .B1(n6137), .B2(keyinput_g35), .C1(n10442), .C2(
        keyinput_g24), .A(n10274), .ZN(n10281) );
  AOI22_X1 U11357 ( .A1(n10352), .A2(keyinput_g5), .B1(keyinput_g17), .B2(
        n10276), .ZN(n10275) );
  OAI221_X1 U11358 ( .B1(n10352), .B2(keyinput_g5), .C1(n10276), .C2(
        keyinput_g17), .A(n10275), .ZN(n10280) );
  XNOR2_X1 U11359 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g95), .ZN(n10278) );
  XNOR2_X1 U11360 ( .A(SI_25_), .B(keyinput_g7), .ZN(n10277) );
  NAND2_X1 U11361 ( .A1(n10278), .A2(n10277), .ZN(n10279) );
  NOR4_X1 U11362 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10306) );
  AOI22_X1 U11363 ( .A1(P2_U3152), .A2(keyinput_g34), .B1(n7588), .B2(
        keyinput_g4), .ZN(n10283) );
  OAI221_X1 U11364 ( .B1(P2_U3152), .B2(keyinput_g34), .C1(n7588), .C2(
        keyinput_g4), .A(n10283), .ZN(n10292) );
  AOI22_X1 U11365 ( .A1(n10285), .A2(keyinput_g59), .B1(n10469), .B2(
        keyinput_g23), .ZN(n10284) );
  OAI221_X1 U11366 ( .B1(n10285), .B2(keyinput_g59), .C1(n10469), .C2(
        keyinput_g23), .A(n10284), .ZN(n10291) );
  XNOR2_X1 U11367 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .ZN(n10289)
         );
  XNOR2_X1 U11368 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .ZN(n10288)
         );
  XNOR2_X1 U11369 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g115), .ZN(n10287)
         );
  XNOR2_X1 U11370 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_g68), .ZN(n10286) );
  NAND4_X1 U11371 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10290) );
  NOR3_X1 U11372 ( .A1(n10292), .A2(n10291), .A3(n10290), .ZN(n10305) );
  INV_X1 U11373 ( .A(SI_6_), .ZN(n10342) );
  AOI22_X1 U11374 ( .A1(n10294), .A2(keyinput_g72), .B1(keyinput_g26), .B2(
        n10342), .ZN(n10293) );
  OAI221_X1 U11375 ( .B1(n10294), .B2(keyinput_g72), .C1(n10342), .C2(
        keyinput_g26), .A(n10293), .ZN(n10303) );
  AOI22_X1 U11376 ( .A1(n10476), .A2(keyinput_g88), .B1(n10296), .B2(
        keyinput_g19), .ZN(n10295) );
  OAI221_X1 U11377 ( .B1(n10476), .B2(keyinput_g88), .C1(n10296), .C2(
        keyinput_g19), .A(n10295), .ZN(n10302) );
  XNOR2_X1 U11378 ( .A(SI_5_), .B(keyinput_g27), .ZN(n10300) );
  XNOR2_X1 U11379 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n10299) );
  XNOR2_X1 U11380 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g112), .ZN(n10298)
         );
  XNOR2_X1 U11381 ( .A(SI_22_), .B(keyinput_g10), .ZN(n10297) );
  NAND4_X1 U11382 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10301) );
  NOR3_X1 U11383 ( .A1(n10303), .A2(n10302), .A3(n10301), .ZN(n10304) );
  NAND4_X1 U11384 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  NOR4_X1 U11385 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10518) );
  XNOR2_X1 U11386 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f98), .ZN(n10315) );
  XNOR2_X1 U11387 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10314) );
  XNOR2_X1 U11388 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_f102), .ZN(n10313)
         );
  XNOR2_X1 U11389 ( .A(SI_15_), .B(keyinput_f17), .ZN(n10312) );
  NAND4_X1 U11390 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10321) );
  XNOR2_X1 U11391 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f116), .ZN(n10319)
         );
  XNOR2_X1 U11392 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f101), .ZN(n10318)
         );
  XNOR2_X1 U11393 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f95), .ZN(n10317) );
  XNOR2_X1 U11394 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_f71), .ZN(n10316) );
  NAND4_X1 U11395 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  NOR2_X1 U11396 ( .A1(n10321), .A2(n10320), .ZN(n10512) );
  AOI22_X1 U11397 ( .A1(n10324), .A2(keyinput_f6), .B1(keyinput_f90), .B2(
        n10323), .ZN(n10322) );
  OAI221_X1 U11398 ( .B1(n10324), .B2(keyinput_f6), .C1(n10323), .C2(
        keyinput_f90), .A(n10322), .ZN(n10336) );
  AOI22_X1 U11399 ( .A1(n10327), .A2(keyinput_f8), .B1(keyinput_f78), .B2(
        n10326), .ZN(n10325) );
  OAI221_X1 U11400 ( .B1(n10327), .B2(keyinput_f8), .C1(n10326), .C2(
        keyinput_f78), .A(n10325), .ZN(n10335) );
  INV_X1 U11401 ( .A(SI_17_), .ZN(n10329) );
  AOI22_X1 U11402 ( .A1(n10330), .A2(keyinput_f77), .B1(keyinput_f15), .B2(
        n10329), .ZN(n10328) );
  OAI221_X1 U11403 ( .B1(n10330), .B2(keyinput_f77), .C1(n10329), .C2(
        keyinput_f15), .A(n10328), .ZN(n10334) );
  XOR2_X1 U11404 ( .A(n6371), .B(keyinput_f60), .Z(n10332) );
  XNOR2_X1 U11405 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_f118), .ZN(n10331)
         );
  NAND2_X1 U11406 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  NOR4_X1 U11407 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10511) );
  OAI22_X1 U11408 ( .A1(n10339), .A2(keyinput_f100), .B1(n10338), .B2(
        keyinput_f126), .ZN(n10337) );
  AOI221_X1 U11409 ( .B1(n10339), .B2(keyinput_f100), .C1(keyinput_f126), .C2(
        n10338), .A(n10337), .ZN(n10350) );
  OAI22_X1 U11410 ( .A1(n10342), .A2(keyinput_f26), .B1(n10341), .B2(
        keyinput_f61), .ZN(n10340) );
  AOI221_X1 U11411 ( .B1(n10342), .B2(keyinput_f26), .C1(keyinput_f61), .C2(
        n10341), .A(n10340), .ZN(n10349) );
  INV_X1 U11412 ( .A(SI_30_), .ZN(n10344) );
  OAI22_X1 U11413 ( .A1(n10345), .A2(keyinput_f9), .B1(n10344), .B2(
        keyinput_f2), .ZN(n10343) );
  AOI221_X1 U11414 ( .B1(n10345), .B2(keyinput_f9), .C1(keyinput_f2), .C2(
        n10344), .A(n10343), .ZN(n10348) );
  OAI22_X1 U11415 ( .A1(n6219), .A2(keyinput_f58), .B1(n6137), .B2(
        keyinput_f35), .ZN(n10346) );
  AOI221_X1 U11416 ( .B1(n6219), .B2(keyinput_f58), .C1(keyinput_f35), .C2(
        n6137), .A(n10346), .ZN(n10347) );
  NAND4_X1 U11417 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10365) );
  INV_X1 U11418 ( .A(SI_0_), .ZN(n10353) );
  AOI22_X1 U11419 ( .A1(n10353), .A2(keyinput_f32), .B1(n10352), .B2(
        keyinput_f5), .ZN(n10351) );
  OAI221_X1 U11420 ( .B1(n10353), .B2(keyinput_f32), .C1(n10352), .C2(
        keyinput_f5), .A(n10351), .ZN(n10364) );
  AOI22_X1 U11421 ( .A1(n10356), .A2(keyinput_f52), .B1(n10355), .B2(
        keyinput_f13), .ZN(n10354) );
  OAI221_X1 U11422 ( .B1(n10356), .B2(keyinput_f52), .C1(n10355), .C2(
        keyinput_f13), .A(n10354), .ZN(n10363) );
  XOR2_X1 U11423 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .Z(n10361) );
  XOR2_X1 U11424 ( .A(SI_11_), .B(keyinput_f21), .Z(n10360) );
  XOR2_X1 U11425 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f121), .Z(n10359) );
  XNOR2_X1 U11426 ( .A(n10357), .B(keyinput_f27), .ZN(n10358) );
  OR4_X1 U11427 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NOR4_X1 U11428 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10510) );
  OAI22_X1 U11429 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_f74), .B1(
        keyinput_f25), .B2(SI_7_), .ZN(n10366) );
  AOI221_X1 U11430 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .C1(
        SI_7_), .C2(keyinput_f25), .A(n10366), .ZN(n10373) );
  OAI22_X1 U11431 ( .A1(SI_28_), .A2(keyinput_f4), .B1(keyinput_f44), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10367) );
  AOI221_X1 U11432 ( .B1(SI_28_), .B2(keyinput_f4), .C1(P2_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n10367), .ZN(n10372) );
  OAI22_X1 U11433 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f104), .B1(
        keyinput_f50), .B2(P2_REG3_REG_17__SCAN_IN), .ZN(n10368) );
  AOI221_X1 U11434 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n10368), .ZN(n10371)
         );
  OAI22_X1 U11435 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f119), .B1(
        keyinput_f1), .B2(SI_31_), .ZN(n10369) );
  AOI221_X1 U11436 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f119), .C1(
        SI_31_), .C2(keyinput_f1), .A(n10369), .ZN(n10370) );
  NAND4_X1 U11437 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10508) );
  OAI22_X1 U11438 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_f106), .B1(
        keyinput_f89), .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n10374) );
  AOI221_X1 U11439 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_f106), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n10374), .ZN(n10400)
         );
  OAI22_X1 U11440 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f124), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n10375) );
  AOI221_X1 U11441 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .C1(
        keyinput_f67), .C2(P2_DATAO_REG_29__SCAN_IN), .A(n10375), .ZN(n10378)
         );
  OAI22_X1 U11442 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_f70), .B1(
        keyinput_f79), .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n10376) );
  AOI221_X1 U11443 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_f79), .A(n10376), .ZN(n10377)
         );
  OAI211_X1 U11444 ( .C1(n10380), .C2(keyinput_f51), .A(n10378), .B(n10377), 
        .ZN(n10379) );
  AOI21_X1 U11445 ( .B1(n10380), .B2(keyinput_f51), .A(n10379), .ZN(n10399) );
  AOI22_X1 U11446 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        SI_14_), .B2(keyinput_f18), .ZN(n10381) );
  OAI221_X1 U11447 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        SI_14_), .C2(keyinput_f18), .A(n10381), .ZN(n10388) );
  AOI22_X1 U11448 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_f85), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_f94), .ZN(n10382) );
  OAI221_X1 U11449 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_f94), .A(n10382), .ZN(n10387) );
  AOI22_X1 U11450 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P1_IR_REG_22__SCAN_IN), 
        .B2(keyinput_f113), .ZN(n10383) );
  OAI221_X1 U11451 ( .B1(SI_3_), .B2(keyinput_f29), .C1(P1_IR_REG_22__SCAN_IN), 
        .C2(keyinput_f113), .A(n10383), .ZN(n10386) );
  AOI22_X1 U11452 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_f123), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .ZN(n10384) );
  OAI221_X1 U11453 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f96), .A(n10384), .ZN(n10385) );
  NOR4_X1 U11454 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10398) );
  AOI22_X1 U11455 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .ZN(n10389) );
  OAI221_X1 U11456 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_f82), .A(n10389), .ZN(n10396)
         );
  AOI22_X1 U11457 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n10390) );
  OAI221_X1 U11458 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n10390), .ZN(n10395)
         );
  AOI22_X1 U11459 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_f84), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_f112), .ZN(n10391) );
  OAI221_X1 U11460 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_f112), .A(n10391), .ZN(n10394) );
  AOI22_X1 U11461 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n10392) );
  OAI221_X1 U11462 ( .B1(SI_29_), .B2(keyinput_f3), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10392), .ZN(n10393) );
  NOR4_X1 U11463 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  NAND4_X1 U11464 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10507) );
  AOI22_X1 U11465 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_f93), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .ZN(n10401) );
  OAI221_X1 U11466 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_f93), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f108), .A(n10401), .ZN(n10408) );
  AOI22_X1 U11467 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10402) );
  OAI221_X1 U11468 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10402), .ZN(n10407)
         );
  AOI22_X1 U11469 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_f115), .ZN(n10403) );
  OAI221_X1 U11470 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_f115), .A(n10403), .ZN(n10406) );
  AOI22_X1 U11471 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_f73), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10404) );
  OAI221_X1 U11472 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_f69), .A(n10404), .ZN(n10405)
         );
  NOR4_X1 U11473 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10440) );
  AOI22_X1 U11474 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_f105), .ZN(n10409) );
  OAI221_X1 U11475 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_f105), .A(n10409), .ZN(n10416) );
  AOI22_X1 U11476 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .ZN(n10410) );
  OAI221_X1 U11477 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n10410), .ZN(n10415)
         );
  AOI22_X1 U11478 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n10411) );
  OAI221_X1 U11479 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n10411), .ZN(n10414)
         );
  AOI22_X1 U11480 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_13_), .B2(
        keyinput_f19), .ZN(n10412) );
  OAI221_X1 U11481 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_13_), .C2(
        keyinput_f19), .A(n10412), .ZN(n10413) );
  NOR4_X1 U11482 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10439) );
  AOI22_X1 U11483 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_f91), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .ZN(n10417) );
  OAI221_X1 U11484 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_f91), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_f109), .A(n10417), .ZN(n10424) );
  AOI22_X1 U11485 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_f64), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10418) );
  OAI221_X1 U11486 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_f64), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10418), .ZN(n10423)
         );
  AOI22_X1 U11487 ( .A1(SI_2_), .A2(keyinput_f30), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10419) );
  OAI221_X1 U11488 ( .B1(SI_2_), .B2(keyinput_f30), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10419), .ZN(n10422)
         );
  AOI22_X1 U11489 ( .A1(SI_20_), .A2(keyinput_f12), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_f110), .ZN(n10420) );
  OAI221_X1 U11490 ( .B1(SI_20_), .B2(keyinput_f12), .C1(P1_IR_REG_19__SCAN_IN), .C2(keyinput_f110), .A(n10420), .ZN(n10421) );
  NOR4_X1 U11491 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10438) );
  AOI22_X1 U11492 ( .A1(n10427), .A2(keyinput_f66), .B1(n10426), .B2(
        keyinput_f41), .ZN(n10425) );
  OAI221_X1 U11493 ( .B1(n10427), .B2(keyinput_f66), .C1(n10426), .C2(
        keyinput_f41), .A(n10425), .ZN(n10436) );
  AOI22_X1 U11494 ( .A1(SI_22_), .A2(keyinput_f10), .B1(P1_IR_REG_26__SCAN_IN), 
        .B2(keyinput_f117), .ZN(n10428) );
  OAI221_X1 U11495 ( .B1(SI_22_), .B2(keyinput_f10), .C1(P1_IR_REG_26__SCAN_IN), .C2(keyinput_f117), .A(n10428), .ZN(n10435) );
  XNOR2_X1 U11496 ( .A(n10429), .B(keyinput_f7), .ZN(n10433) );
  XNOR2_X1 U11497 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f107), .ZN(n10432)
         );
  XNOR2_X1 U11498 ( .A(SI_10_), .B(keyinput_f22), .ZN(n10431) );
  XNOR2_X1 U11499 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_f114), .ZN(n10430)
         );
  NAND4_X1 U11500 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  NOR3_X1 U11501 ( .A1(n10436), .A2(n10435), .A3(n10434), .ZN(n10437) );
  NAND4_X1 U11502 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10506) );
  AOI22_X1 U11503 ( .A1(n10442), .A2(keyinput_f24), .B1(keyinput_f56), .B2(
        n7286), .ZN(n10441) );
  OAI221_X1 U11504 ( .B1(n10442), .B2(keyinput_f24), .C1(n7286), .C2(
        keyinput_f56), .A(n10441), .ZN(n10452) );
  AOI22_X1 U11505 ( .A1(n10445), .A2(keyinput_f80), .B1(n10444), .B2(
        keyinput_f16), .ZN(n10443) );
  OAI221_X1 U11506 ( .B1(n10445), .B2(keyinput_f80), .C1(n10444), .C2(
        keyinput_f16), .A(n10443), .ZN(n10451) );
  XOR2_X1 U11507 ( .A(n6178), .B(keyinput_f53), .Z(n10449) );
  XNOR2_X1 U11508 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f97), .ZN(n10448) );
  XNOR2_X1 U11509 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n10447)
         );
  XNOR2_X1 U11510 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f111), .ZN(n10446)
         );
  NAND4_X1 U11511 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10450) );
  NOR3_X1 U11512 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n10504) );
  AOI22_X1 U11513 ( .A1(n10455), .A2(keyinput_f45), .B1(n10454), .B2(
        keyinput_f99), .ZN(n10453) );
  OAI221_X1 U11514 ( .B1(n10455), .B2(keyinput_f45), .C1(n10454), .C2(
        keyinput_f99), .A(n10453), .ZN(n10467) );
  AOI22_X1 U11515 ( .A1(n10458), .A2(keyinput_f65), .B1(n10457), .B2(
        keyinput_f40), .ZN(n10456) );
  OAI221_X1 U11516 ( .B1(n10458), .B2(keyinput_f65), .C1(n10457), .C2(
        keyinput_f40), .A(n10456), .ZN(n10466) );
  AOI22_X1 U11517 ( .A1(n10461), .A2(keyinput_f38), .B1(n10460), .B2(
        keyinput_f62), .ZN(n10459) );
  OAI221_X1 U11518 ( .B1(n10461), .B2(keyinput_f38), .C1(n10460), .C2(
        keyinput_f62), .A(n10459), .ZN(n10465) );
  XNOR2_X1 U11519 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_f83), .ZN(n10463) );
  XNOR2_X1 U11520 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10462) );
  NAND2_X1 U11521 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  NOR4_X1 U11522 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10503) );
  AOI22_X1 U11523 ( .A1(n10470), .A2(keyinput_f39), .B1(n10469), .B2(
        keyinput_f23), .ZN(n10468) );
  OAI221_X1 U11524 ( .B1(n10470), .B2(keyinput_f39), .C1(n10469), .C2(
        keyinput_f23), .A(n10468), .ZN(n10483) );
  AOI22_X1 U11525 ( .A1(n10473), .A2(keyinput_f47), .B1(n10472), .B2(
        keyinput_f127), .ZN(n10471) );
  OAI221_X1 U11526 ( .B1(n10473), .B2(keyinput_f47), .C1(n10472), .C2(
        keyinput_f127), .A(n10471), .ZN(n10482) );
  INV_X1 U11527 ( .A(SI_18_), .ZN(n10475) );
  AOI22_X1 U11528 ( .A1(n10476), .A2(keyinput_f88), .B1(n10475), .B2(
        keyinput_f14), .ZN(n10474) );
  OAI221_X1 U11529 ( .B1(n10476), .B2(keyinput_f88), .C1(n10475), .C2(
        keyinput_f14), .A(n10474), .ZN(n10481) );
  AOI22_X1 U11530 ( .A1(n10479), .A2(keyinput_f103), .B1(keyinput_f37), .B2(
        n10478), .ZN(n10477) );
  OAI221_X1 U11531 ( .B1(n10479), .B2(keyinput_f103), .C1(n10478), .C2(
        keyinput_f37), .A(n10477), .ZN(n10480) );
  NOR4_X1 U11532 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10502) );
  AOI22_X1 U11533 ( .A1(n10486), .A2(keyinput_f11), .B1(keyinput_f46), .B2(
        n10485), .ZN(n10484) );
  OAI221_X1 U11534 ( .B1(n10486), .B2(keyinput_f11), .C1(n10485), .C2(
        keyinput_f46), .A(n10484), .ZN(n10487) );
  INV_X1 U11535 ( .A(n10487), .ZN(n10500) );
  AOI22_X1 U11536 ( .A1(n10490), .A2(keyinput_f75), .B1(keyinput_f57), .B2(
        n10489), .ZN(n10488) );
  OAI221_X1 U11537 ( .B1(n10490), .B2(keyinput_f75), .C1(n10489), .C2(
        keyinput_f57), .A(n10488), .ZN(n10491) );
  INV_X1 U11538 ( .A(n10491), .ZN(n10499) );
  XNOR2_X1 U11539 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f122), .ZN(n10494)
         );
  XNOR2_X1 U11540 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f92), .ZN(n10493) );
  XNOR2_X1 U11541 ( .A(keyinput_f49), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n10492)
         );
  AND3_X1 U11542 ( .A1(n10494), .A2(n10493), .A3(n10492), .ZN(n10498) );
  INV_X1 U11543 ( .A(keyinput_f125), .ZN(n10495) );
  XNOR2_X1 U11544 ( .A(n10496), .B(n10495), .ZN(n10497) );
  AND4_X1 U11545 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10501) );
  NAND4_X1 U11546 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10505) );
  NOR4_X1 U11547 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  NAND4_X1 U11548 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10514) );
  AOI21_X1 U11549 ( .B1(keyinput_f42), .B2(n10514), .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10516) );
  INV_X1 U11550 ( .A(keyinput_f42), .ZN(n10513) );
  AOI21_X1 U11551 ( .B1(n10514), .B2(n10513), .A(keyinput_g42), .ZN(n10515) );
  AOI22_X1 U11552 ( .A1(keyinput_g42), .A2(n10516), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(n10515), .ZN(n10517) );
  AOI21_X1 U11553 ( .B1(n10519), .B2(n10518), .A(n10517), .ZN(n10521) );
  XNOR2_X1 U11554 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10520) );
  XNOR2_X1 U11555 ( .A(n10521), .B(n10520), .ZN(n10522) );
  XNOR2_X1 U11556 ( .A(n10523), .B(n10522), .ZN(ADD_1071_U4) );
  OAI21_X1 U11557 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(ADD_1071_U47) );
  OAI21_X1 U11558 ( .B1(n10529), .B2(n10528), .A(n10527), .ZN(ADD_1071_U49) );
  AOI21_X1 U11559 ( .B1(n10532), .B2(n10531), .A(n10530), .ZN(ADD_1071_U54) );
  OAI21_X1 U11560 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(ADD_1071_U51) );
  OAI21_X1 U11561 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(ADD_1071_U55) );
  OAI21_X1 U11562 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(ADD_1071_U48) );
  OAI21_X1 U11563 ( .B1(n10544), .B2(n10543), .A(n10542), .ZN(ADD_1071_U50) );
  AOI21_X1 U11564 ( .B1(n10547), .B2(n10546), .A(n10545), .ZN(ADD_1071_U53) );
  OAI21_X1 U11565 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(ADD_1071_U52) );
  INV_X1 U5001 ( .A(n6811), .ZN(n5172) );
  AND2_X1 U5102 ( .A1(n5031), .A2(n4533), .ZN(n4484) );
  NAND2_X1 U5930 ( .A1(n7760), .A2(n7759), .ZN(n7812) );
  AOI211_X1 U6176 ( .C1(n6358), .C2(n6357), .A(n7810), .B(n6356), .ZN(n6382)
         );
  NAND2_X2 U7842 ( .A1(n6367), .A2(n6355), .ZN(n7810) );
endmodule

