

module b17_C_gen_AntiSAT_k_128_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12541, n12542, n12543, n12544, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270;

  MUX2_X1 U11075 ( .A(n19097), .B(n19096), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19099) );
  INV_X1 U11076 ( .A(n20319), .ZN(n20361) );
  INV_X1 U11077 ( .A(n18255), .ZN(n18226) );
  NAND2_X1 U11078 ( .A1(n14614), .A2(n14604), .ZN(n14603) );
  OR2_X1 U11079 ( .A1(n15293), .A2(n15287), .ZN(n15285) );
  NOR3_X1 U11080 ( .A1(n17737), .A2(n17712), .A3(n17625), .ZN(n17714) );
  AND2_X1 U11081 ( .A1(n13718), .A2(n13929), .ZN(n16083) );
  NAND2_X1 U11082 ( .A1(n10642), .A2(n9827), .ZN(n20452) );
  INV_X1 U11083 ( .A(n14510), .ZN(n12760) );
  NOR2_X2 U11084 ( .A1(n18610), .A2(n18642), .ZN(n11702) );
  INV_X1 U11085 ( .A(n12648), .ZN(n14516) );
  NAND2_X1 U11086 ( .A1(n10550), .A2(n10549), .ZN(n10784) );
  INV_X2 U11087 ( .A(n12298), .ZN(n16070) );
  CLKBUF_X2 U11088 ( .A(n11971), .Z(n14506) );
  CLKBUF_X2 U11089 ( .A(n12755), .Z(n9648) );
  AND2_X2 U11090 ( .A1(n11824), .A2(n12026), .ZN(n12072) );
  AND2_X2 U11092 ( .A1(n12018), .A2(n12026), .ZN(n12150) );
  INV_X1 U11093 ( .A(n11550), .ZN(n17770) );
  INV_X1 U11094 ( .A(n17333), .ZN(n17575) );
  INV_X1 U11095 ( .A(n17522), .ZN(n16196) );
  CLKBUF_X2 U11096 ( .A(n11551), .Z(n17574) );
  INV_X2 U11097 ( .A(n16179), .ZN(n11513) );
  AND2_X1 U11098 ( .A1(n10282), .A2(n10281), .ZN(n10215) );
  NOR2_X1 U11099 ( .A1(n9970), .A2(n10343), .ZN(n9969) );
  BUF_X2 U11100 ( .A(n10283), .Z(n9672) );
  AND2_X2 U11101 ( .A1(n15992), .A2(n16709), .ZN(n11899) );
  AND3_X1 U11102 ( .A1(n14224), .A2(n10226), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10227) );
  OAI22_X1 U11103 ( .A1(n16828), .A2(n13436), .B1(n13426), .B2(n13437), .ZN(
        n20840) );
  NAND2_X2 U11104 ( .A1(n16364), .A2(n13386), .ZN(n13437) );
  NAND2_X2 U11105 ( .A1(n16364), .A2(n13623), .ZN(n13436) );
  INV_X1 U11107 ( .A(n21270), .ZN(n9632) );
  INV_X1 U11108 ( .A(n10350), .ZN(n11297) );
  NOR2_X2 U11109 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10233) );
  AND3_X1 U11110 ( .A1(n10409), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10241) );
  INV_X1 U11111 ( .A(n11422), .ZN(n11284) );
  INV_X1 U11112 ( .A(n11406), .ZN(n10518) );
  NAND2_X1 U11113 ( .A1(n10033), .A2(n11910), .ZN(n13163) );
  AND2_X1 U11114 ( .A1(n13243), .A2(n10231), .ZN(n10363) );
  NOR2_X1 U11115 ( .A1(n10789), .A2(n10757), .ZN(n10791) );
  NAND2_X1 U11116 ( .A1(n13638), .A2(n13213), .ZN(n16260) );
  NOR2_X1 U11117 ( .A1(n14992), .A2(n14990), .ZN(n16330) );
  AND2_X1 U11118 ( .A1(n9946), .A2(n9737), .ZN(n14950) );
  INV_X2 U11119 ( .A(n14158), .ZN(n9817) );
  AND2_X1 U11120 ( .A1(n12862), .A2(n10396), .ZN(n10405) );
  CLKBUF_X2 U11121 ( .A(n11970), .Z(n14510) );
  NOR2_X1 U11122 ( .A1(n13720), .A2(n19612), .ZN(n13716) );
  OR2_X1 U11123 ( .A1(n11460), .A2(n9869), .ZN(n10220) );
  INV_X1 U11124 ( .A(n14164), .ZN(n14204) );
  NAND2_X1 U11125 ( .A1(n9801), .A2(n10843), .ZN(n13532) );
  XNOR2_X1 U11127 ( .A(n9948), .B(n12681), .ZN(n13693) );
  NAND2_X1 U11128 ( .A1(n13444), .A2(n12035), .ZN(n13484) );
  NAND2_X1 U11129 ( .A1(n12489), .A2(n19650), .ZN(n12619) );
  NAND2_X1 U11130 ( .A1(n11999), .A2(n12007), .ZN(n11998) );
  XNOR2_X1 U11131 ( .A(n9843), .B(n9927), .ZN(n14472) );
  NAND4_X2 U11132 ( .A1(n12594), .A2(n12593), .A3(n12592), .A4(n12591), .ZN(
        n14497) );
  BUF_X1 U11133 ( .A(n11919), .Z(n19659) );
  AND2_X1 U11134 ( .A1(n9881), .A2(n9879), .ZN(n18036) );
  NOR2_X1 U11135 ( .A1(n13213), .A2(n13635), .ZN(n16253) );
  CLKBUF_X3 U11136 ( .A(n13693), .Z(n9676) );
  CLKBUF_X3 U11137 ( .A(n19433), .Z(n9647) );
  NOR2_X1 U11138 ( .A1(n15479), .A2(n15478), .ZN(n15480) );
  NOR2_X2 U11139 ( .A1(n13484), .A2(n10048), .ZN(n15307) );
  NAND2_X1 U11140 ( .A1(n15307), .A2(n12162), .ZN(n16592) );
  INV_X1 U11142 ( .A(n17271), .ZN(n9731) );
  NAND2_X2 U11143 ( .A1(n19229), .A2(n19235), .ZN(n17302) );
  OR2_X1 U11144 ( .A1(n17789), .A2(n17660), .ZN(n17661) );
  NOR2_X2 U11145 ( .A1(n17746), .A2(n11542), .ZN(n18142) );
  INV_X1 U11146 ( .A(n16946), .ZN(n18610) );
  INV_X1 U11147 ( .A(n20327), .ZN(n14732) );
  XNOR2_X1 U11148 ( .A(n14167), .B(n14166), .ZN(n15017) );
  OR2_X1 U11149 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n14332), .ZN(n9633) );
  NAND2_X1 U11150 ( .A1(n10232), .A2(n13458), .ZN(n11422) );
  INV_X2 U11151 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U11152 ( .A1(n11879), .A2(n11878), .ZN(n11911) );
  AND3_X1 U11153 ( .A1(n9679), .A2(n9729), .A3(n9972), .ZN(n9634) );
  INV_X2 U11154 ( .A(n11418), .ZN(n11338) );
  OR2_X2 U11155 ( .A1(n17765), .A2(n11550), .ZN(n11549) );
  AND3_X2 U11156 ( .A1(n9732), .A2(n11520), .A3(n10001), .ZN(n11550) );
  NAND3_X2 U11157 ( .A1(n11498), .A2(n11497), .A3(n11496), .ZN(n11736) );
  INV_X1 U11159 ( .A(n10810), .ZN(n10421) );
  NAND2_X1 U11160 ( .A1(n10397), .A2(n10810), .ZN(n13299) );
  NOR2_X2 U11161 ( .A1(n13995), .A2(n13994), .ZN(n10093) );
  NAND2_X1 U11162 ( .A1(n10241), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10337) );
  AND2_X2 U11165 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15992) );
  AND2_X4 U11166 ( .A1(n15978), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9635) );
  NOR4_X2 U11167 ( .A1(n14543), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21201), 
        .A4(n21182), .ZN(n14185) );
  INV_X1 U11168 ( .A(n11911), .ZN(n9636) );
  BUF_X4 U11169 ( .A(n12025), .Z(n9637) );
  BUF_X4 U11170 ( .A(n12025), .Z(n9638) );
  NAND2_X2 U11172 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n9868), .ZN(
        n11458) );
  XNOR2_X2 U11173 ( .A(n10592), .B(n13314), .ZN(n13310) );
  NAND2_X2 U11174 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  AND2_X1 U11175 ( .A1(n15992), .A2(n16709), .ZN(n9641) );
  INV_X1 U11176 ( .A(n11406), .ZN(n9673) );
  AND3_X2 U11177 ( .A1(n11808), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9642) );
  AND3_X2 U11178 ( .A1(n12397), .A2(n16709), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9643) );
  NOR2_X4 U11180 ( .A1(n16745), .A2(n16918), .ZN(n18248) );
  AND2_X1 U11181 ( .A1(n15977), .A2(n12397), .ZN(n9645) );
  AND2_X1 U11182 ( .A1(n15977), .A2(n12397), .ZN(n9646) );
  AND2_X1 U11183 ( .A1(n15977), .A2(n12397), .ZN(n9660) );
  AND2_X4 U11184 ( .A1(n15977), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12020) );
  AND2_X4 U11185 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15977) );
  CLKBUF_X1 U11186 ( .A(n14575), .Z(n14576) );
  AOI211_X1 U11187 ( .C1(n15655), .C2(n19595), .A(n15413), .B(n15412), .ZN(
        n15414) );
  CLKBUF_X1 U11188 ( .A(n14590), .Z(n14601) );
  NAND2_X1 U11189 ( .A1(n10208), .A2(n14307), .ZN(n14427) );
  AND2_X1 U11190 ( .A1(n14635), .A2(n14182), .ZN(n14584) );
  NOR2_X1 U11191 ( .A1(n14991), .A2(n10733), .ZN(n9983) );
  OR2_X1 U11192 ( .A1(n15144), .A2(n10738), .ZN(n14992) );
  XNOR2_X1 U11193 ( .A(n16352), .B(n15021), .ZN(n15003) );
  INV_X4 U11194 ( .A(n10723), .ZN(n16352) );
  AND2_X1 U11195 ( .A1(n13715), .A2(n13929), .ZN(n19628) );
  NAND2_X1 U11196 ( .A1(n18036), .A2(n18383), .ZN(n18035) );
  OAI22_X1 U11197 ( .A1(n18259), .A2(n18462), .B1(n18084), .B2(n18460), .ZN(
        n18127) );
  OAI22_X1 U11198 ( .A1(n15939), .A2(n15938), .B1(n14233), .B2(n12619), .ZN(
        n15926) );
  AND2_X1 U11199 ( .A1(n13689), .A2(n12007), .ZN(n14053) );
  NAND2_X1 U11200 ( .A1(n12451), .A2(n11857), .ZN(n13164) );
  INV_X2 U11201 ( .A(n10406), .ZN(n13634) );
  BUF_X1 U11202 ( .A(n11927), .Z(n9670) );
  INV_X2 U11203 ( .A(n11914), .ZN(n11906) );
  INV_X1 U11204 ( .A(n16039), .ZN(n11927) );
  AND2_X1 U11205 ( .A1(n11843), .A2(n11842), .ZN(n13155) );
  AND4_X1 U11206 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10316) );
  CLKBUF_X3 U11207 ( .A(n11554), .Z(n9653) );
  INV_X4 U11208 ( .A(n10220), .ZN(n17572) );
  INV_X1 U11210 ( .A(n9654), .ZN(n11425) );
  INV_X1 U11211 ( .A(n10380), .ZN(n9649) );
  INV_X1 U11212 ( .A(n11487), .ZN(n17257) );
  AND2_X2 U11213 ( .A1(n9638), .A2(n12026), .ZN(n12073) );
  NOR2_X1 U11214 ( .A1(n10238), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10252) );
  INV_X2 U11215 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14224) );
  INV_X2 U11216 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19229) );
  INV_X2 U11217 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16709) );
  NOR2_X4 U11218 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15994) );
  AND2_X1 U11219 ( .A1(n14534), .A2(n14533), .ZN(n14879) );
  AND2_X1 U11220 ( .A1(n9910), .A2(n9909), .ZN(n14898) );
  OAI21_X1 U11221 ( .B1(n14562), .B2(n14547), .A(n14546), .ZN(n14891) );
  NOR2_X1 U11222 ( .A1(n14892), .A2(n9885), .ZN(n14888) );
  OAI21_X1 U11223 ( .B1(n14576), .B2(n14577), .A(n14561), .ZN(n14906) );
  AND2_X1 U11224 ( .A1(n9956), .A2(n9952), .ZN(n9951) );
  AOI21_X1 U11225 ( .B1(n9887), .B2(n15074), .A(n14886), .ZN(n9886) );
  AOI21_X1 U11226 ( .B1(n9887), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14885), .ZN(n14892) );
  AND2_X1 U11227 ( .A1(n14575), .A2(n9911), .ZN(n14562) );
  OR2_X1 U11228 ( .A1(n14192), .A2(n15066), .ZN(n10747) );
  NOR2_X1 U11229 ( .A1(n15420), .A2(n15647), .ZN(n9889) );
  NAND2_X1 U11230 ( .A1(n14909), .A2(n9754), .ZN(n10146) );
  AND2_X1 U11231 ( .A1(n14909), .A2(n9693), .ZN(n9935) );
  NOR2_X1 U11232 ( .A1(n15783), .A2(n9807), .ZN(n15799) );
  NAND2_X1 U11233 ( .A1(n14921), .A2(n10743), .ZN(n14883) );
  AND2_X1 U11234 ( .A1(n15905), .A2(n9700), .ZN(n15419) );
  OAI21_X1 U11235 ( .B1(n15542), .B2(n15541), .A(n15493), .ZN(n15533) );
  AND2_X1 U11236 ( .A1(n15905), .A2(n15872), .ZN(n15622) );
  NAND2_X1 U11237 ( .A1(n9798), .A2(n9832), .ZN(n14907) );
  AND2_X1 U11238 ( .A1(n9736), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U11239 ( .A1(n12328), .A2(n12327), .ZN(n15253) );
  AOI21_X1 U11240 ( .B1(n16800), .B2(n18150), .A(n16759), .ZN(n16760) );
  XNOR2_X1 U11241 ( .A(n14511), .B(n10124), .ZN(n16587) );
  NAND2_X1 U11242 ( .A1(n9946), .A2(n9947), .ZN(n14976) );
  OR2_X1 U11243 ( .A1(n12302), .A2(n12301), .ZN(n10217) );
  NAND2_X1 U11244 ( .A1(n15266), .A2(n15265), .ZN(n15264) );
  AND2_X1 U11245 ( .A1(n14318), .A2(n9740), .ZN(n9844) );
  OR2_X1 U11246 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  XNOR2_X1 U11247 ( .A(n14316), .B(n15940), .ZN(n15937) );
  AND2_X1 U11248 ( .A1(n9878), .A2(n9877), .ZN(n17891) );
  NAND2_X1 U11249 ( .A1(n14312), .A2(n19411), .ZN(n14316) );
  AOI21_X1 U11250 ( .B1(n12225), .B2(n10046), .A(n12249), .ZN(n10044) );
  AND2_X1 U11251 ( .A1(n9714), .A2(n12248), .ZN(n12225) );
  AND2_X1 U11252 ( .A1(n10040), .A2(n10037), .ZN(n9714) );
  AND2_X1 U11253 ( .A1(n14681), .A2(n14181), .ZN(n14635) );
  NAND2_X1 U11254 ( .A1(n9884), .A2(n9727), .ZN(n14991) );
  NOR2_X1 U11255 ( .A1(n9943), .A2(n10727), .ZN(n9942) );
  AND3_X1 U11256 ( .A1(n9905), .A2(n13656), .A3(n9760), .ZN(n9903) );
  NAND2_X1 U11257 ( .A1(n15003), .A2(n10732), .ZN(n15145) );
  AND2_X1 U11258 ( .A1(n10851), .A2(n10850), .ZN(n13541) );
  NAND2_X1 U11259 ( .A1(n17950), .A2(n18310), .ZN(n17949) );
  AOI21_X1 U11260 ( .B1(n10842), .B2(n11010), .A(n10841), .ZN(n13533) );
  OAI211_X1 U11261 ( .C1(n10856), .C2(n11031), .A(n10855), .B(n10854), .ZN(
        n13656) );
  NOR2_X1 U11262 ( .A1(n15323), .A2(n15322), .ZN(n12653) );
  NAND2_X1 U11263 ( .A1(n13305), .A2(n12017), .ZN(n13444) );
  OR2_X1 U11264 ( .A1(n14656), .A2(n14174), .ZN(n14620) );
  AOI21_X1 U11265 ( .B1(n10863), .B2(n11010), .A(n10862), .ZN(n13810) );
  AND2_X1 U11266 ( .A1(n17997), .A2(n17983), .ZN(n18025) );
  NAND2_X1 U11267 ( .A1(n13307), .A2(n13306), .ZN(n13305) );
  AND2_X1 U11268 ( .A1(n11989), .A2(n13885), .ZN(n13307) );
  XNOR2_X1 U11269 ( .A(n10722), .B(n10710), .ZN(n10863) );
  OR2_X1 U11270 ( .A1(n12016), .A2(n11988), .ZN(n11989) );
  NAND2_X1 U11271 ( .A1(n13715), .A2(n16001), .ZN(n13746) );
  NAND2_X1 U11272 ( .A1(n13723), .A2(n13722), .ZN(n20055) );
  AND2_X1 U11273 ( .A1(n13716), .A2(n16001), .ZN(n14287) );
  NAND2_X1 U11274 ( .A1(n10662), .A2(n9820), .ZN(n10722) );
  AND2_X1 U11275 ( .A1(n13710), .A2(n14031), .ZN(n13715) );
  NAND2_X1 U11276 ( .A1(n11986), .A2(n11985), .ZN(n12016) );
  INV_X1 U11277 ( .A(n13720), .ZN(n13723) );
  OR2_X1 U11278 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  OR2_X1 U11279 ( .A1(n20447), .A2(n20441), .ZN(n15154) );
  XNOR2_X1 U11280 ( .A(n13227), .B(n10588), .ZN(n13234) );
  AND2_X1 U11281 ( .A1(n11581), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U11282 ( .A1(n13226), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13227) );
  NAND2_X2 U11283 ( .A1(n14865), .A2(n13300), .ZN(n14869) );
  AND2_X1 U11284 ( .A1(n12855), .A2(n20300), .ZN(n12931) );
  NAND2_X1 U11285 ( .A1(n10581), .A2(n10580), .ZN(n13226) );
  NAND3_X1 U11286 ( .A1(n9823), .A2(n9825), .A3(n9822), .ZN(n20663) );
  AND2_X1 U11287 ( .A1(n12821), .A2(n9761), .ZN(n15236) );
  AND2_X1 U11288 ( .A1(n13815), .A2(n13814), .ZN(n13912) );
  XNOR2_X1 U11289 ( .A(n10537), .B(n10535), .ZN(n10804) );
  NAND2_X1 U11290 ( .A1(n18170), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18169) );
  OR2_X1 U11291 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  NAND2_X2 U11292 ( .A1(n10800), .A2(n10799), .ZN(n16254) );
  NOR2_X2 U11293 ( .A1(n14351), .A2(n14347), .ZN(n14373) );
  INV_X1 U11294 ( .A(n18499), .ZN(n18312) );
  NOR2_X2 U11295 ( .A1(n16037), .A2(n19782), .ZN(n16038) );
  CLKBUF_X1 U11296 ( .A(n10812), .Z(n14221) );
  AND2_X1 U11297 ( .A1(n10465), .A2(n10463), .ZN(n10528) );
  AND2_X1 U11298 ( .A1(n15959), .A2(n12566), .ZN(n15939) );
  AND2_X1 U11299 ( .A1(n12679), .A2(n11981), .ZN(n12681) );
  OR2_X1 U11300 ( .A1(n11980), .A2(n11979), .ZN(n12679) );
  NAND2_X1 U11301 ( .A1(n13338), .A2(n13337), .ZN(n13545) );
  AOI21_X2 U11302 ( .B1(n14514), .B2(n16735), .A(n10021), .ZN(n19433) );
  INV_X1 U11303 ( .A(n14097), .ZN(n19062) );
  INV_X1 U11304 ( .A(n19390), .ZN(n19459) );
  AOI21_X2 U11305 ( .B1(n19053), .B2(n19046), .A(n19052), .ZN(n19047) );
  NAND2_X1 U11306 ( .A1(n10415), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10430) );
  XNOR2_X1 U11307 ( .A(n9711), .B(n12792), .ZN(n14514) );
  NAND2_X1 U11308 ( .A1(n10408), .A2(n10135), .ZN(n9900) );
  INV_X2 U11309 ( .A(n17618), .ZN(n17596) );
  NOR2_X1 U11310 ( .A1(n13317), .A2(n13316), .ZN(n13338) );
  NAND2_X1 U11311 ( .A1(n19046), .A2(n14096), .ZN(n18593) );
  NAND2_X1 U11312 ( .A1(n18215), .A2(n18216), .ZN(n18214) );
  AOI211_X2 U11313 ( .C1(n19256), .C2(n11718), .A(n16945), .B(n17838), .ZN(
        n19046) );
  AND3_X1 U11314 ( .A1(n11952), .A2(n11951), .A3(n10222), .ZN(n11954) );
  NAND2_X1 U11315 ( .A1(n14326), .A2(n12704), .ZN(n14332) );
  NOR2_X2 U11316 ( .A1(n16917), .A2(n11717), .ZN(n16945) );
  NAND2_X1 U11317 ( .A1(n15996), .A2(n9810), .ZN(n13150) );
  NAND2_X1 U11318 ( .A1(n18547), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18546) );
  XNOR2_X1 U11319 ( .A(n11570), .B(n11569), .ZN(n18547) );
  NOR2_X1 U11320 ( .A1(n15172), .A2(n12791), .ZN(n15185) );
  NOR2_X1 U11321 ( .A1(n19272), .A2(n14087), .ZN(n19051) );
  NAND2_X1 U11322 ( .A1(n9811), .A2(n11929), .ZN(n11933) );
  OR2_X1 U11323 ( .A1(n14163), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12889) );
  AOI21_X1 U11324 ( .B1(n14218), .B2(n13405), .A(n10405), .ZN(n10401) );
  NAND2_X1 U11325 ( .A1(n11957), .A2(n13151), .ZN(n15996) );
  AND2_X1 U11326 ( .A1(n10403), .A2(n13638), .ZN(n10138) );
  NAND2_X1 U11327 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  NOR2_X1 U11328 ( .A1(n15184), .A2(n19322), .ZN(n15183) );
  NOR4_X1 U11329 ( .A1(n18619), .A2(n18623), .A3(n11713), .A4(n11703), .ZN(
        n11723) );
  OR2_X1 U11330 ( .A1(n12676), .A2(n12446), .ZN(n11950) );
  NAND2_X1 U11331 ( .A1(n9932), .A2(n11866), .ZN(n13154) );
  INV_X1 U11332 ( .A(n14218), .ZN(n13260) );
  OAI21_X1 U11333 ( .B1(n12619), .B2(n13105), .A(n12488), .ZN(n13057) );
  NAND2_X1 U11334 ( .A1(n12492), .A2(n10053), .ZN(n13056) );
  INV_X1 U11335 ( .A(n10404), .ZN(n9650) );
  AND2_X1 U11336 ( .A1(n12860), .A2(n10225), .ZN(n12861) );
  NAND2_X4 U11337 ( .A1(n13213), .A2(n13635), .ZN(n14158) );
  NAND2_X2 U11338 ( .A1(n13170), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12696) );
  AND2_X1 U11339 ( .A1(n13030), .A2(n13151), .ZN(n12472) );
  INV_X2 U11340 ( .A(n17729), .ZN(n18642) );
  INV_X1 U11341 ( .A(n13635), .ZN(n13638) );
  AND2_X1 U11342 ( .A1(n11937), .A2(n12471), .ZN(n13170) );
  AND2_X1 U11343 ( .A1(n12449), .A2(n19659), .ZN(n11857) );
  NOR2_X1 U11344 ( .A1(n11907), .A2(n11916), .ZN(n11924) );
  NAND2_X2 U11345 ( .A1(n12666), .A2(n12489), .ZN(n12648) );
  AND4_X2 U11346 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10810) );
  NAND4_X1 U11347 ( .A1(n9634), .A2(n9969), .A3(n10352), .A4(n9971), .ZN(
        n10406) );
  NOR2_X2 U11348 ( .A1(n10369), .A2(n10368), .ZN(n10225) );
  NAND2_X1 U11349 ( .A1(n11936), .A2(n11906), .ZN(n11866) );
  NAND3_X1 U11350 ( .A1(n11617), .A2(n11616), .A3(n11615), .ZN(n18632) );
  NAND2_X1 U11351 ( .A1(n11927), .A2(n9636), .ZN(n12435) );
  INV_X1 U11352 ( .A(n13081), .ZN(n13178) );
  NAND2_X1 U11353 ( .A1(n11844), .A2(n12485), .ZN(n11908) );
  INV_X1 U11354 ( .A(n11928), .ZN(n12666) );
  CLKBUF_X3 U11355 ( .A(n12485), .Z(n19650) );
  NOR2_X2 U11356 ( .A1(n11597), .A2(n11596), .ZN(n19256) );
  INV_X2 U11357 ( .A(U212), .ZN(n16864) );
  OR2_X2 U11358 ( .A1(n16865), .A2(n16807), .ZN(n16867) );
  AND4_X1 U11359 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10250) );
  INV_X2 U11360 ( .A(n13881), .ZN(n11844) );
  INV_X1 U11361 ( .A(n13155), .ZN(n19646) );
  OR2_X1 U11362 ( .A1(n12504), .A2(n12503), .ZN(n13117) );
  NAND2_X1 U11363 ( .A1(n11856), .A2(n11855), .ZN(n11919) );
  AND2_X1 U11364 ( .A1(n9977), .A2(n10344), .ZN(n9971) );
  AND4_X1 U11365 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10224) );
  NOR2_X1 U11366 ( .A1(n10285), .A2(n10284), .ZN(n10294) );
  AND4_X1 U11367 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10273) );
  NOR2_X1 U11368 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  AND2_X1 U11369 ( .A1(n9838), .A2(n9837), .ZN(n11830) );
  AND2_X1 U11370 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n9970) );
  CLKBUF_X1 U11371 ( .A(n19195), .Z(n19189) );
  NAND2_X1 U11372 ( .A1(n10351), .A2(n10345), .ZN(n9973) );
  NAND2_X2 U11373 ( .A1(n21031), .A2(n20979), .ZN(n21025) );
  NAND2_X2 U11374 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21031), .ZN(n21028) );
  OAI21_X1 U11375 ( .B1(n11872), .B2(n11871), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11879) );
  NAND3_X1 U11376 ( .A1(n11896), .A2(n11895), .A3(n11894), .ZN(n11905) );
  NAND2_X2 U11377 ( .A1(n20229), .A2(n20183), .ZN(n20232) );
  INV_X1 U11378 ( .A(n10337), .ZN(n9665) );
  NAND2_X2 U11379 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20229), .ZN(n20228) );
  INV_X1 U11380 ( .A(n11359), .ZN(n10379) );
  CLKBUF_X1 U11381 ( .A(n13460), .Z(n9656) );
  BUF_X2 U11382 ( .A(n11551), .Z(n16191) );
  INV_X1 U11383 ( .A(n11464), .ZN(n17333) );
  NAND2_X2 U11384 ( .A1(n19265), .A2(n19132), .ZN(n19180) );
  AND2_X1 U11385 ( .A1(n11898), .A2(n11897), .ZN(n11903) );
  AND3_X1 U11386 ( .A1(n11893), .A2(n12026), .A3(n11892), .ZN(n11896) );
  AND2_X2 U11387 ( .A1(n13243), .A2(n10243), .ZN(n10447) );
  AND2_X1 U11388 ( .A1(n10252), .A2(n13243), .ZN(n11086) );
  INV_X2 U11389 ( .A(n21073), .ZN(n21031) );
  NAND2_X1 U11390 ( .A1(n13262), .A2(n13461), .ZN(n13460) );
  AND2_X2 U11391 ( .A1(n12018), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12098) );
  AND2_X2 U11392 ( .A1(n9658), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12579) );
  BUF_X4 U11393 ( .A(n11486), .Z(n9651) );
  AND2_X2 U11394 ( .A1(n9659), .A2(n12026), .ZN(n12569) );
  NAND2_X1 U11395 ( .A1(n10227), .A2(n13461), .ZN(n10359) );
  INV_X2 U11396 ( .A(n16906), .ZN(n16908) );
  NAND2_X1 U11397 ( .A1(n10252), .A2(n13243), .ZN(n11418) );
  BUF_X2 U11398 ( .A(n11640), .Z(n17455) );
  BUF_X2 U11399 ( .A(n11638), .Z(n9652) );
  NAND2_X1 U11400 ( .A1(n13262), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10551) );
  INV_X1 U11401 ( .A(n10495), .ZN(n9654) );
  NOR2_X1 U11402 ( .A1(n13264), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10243) );
  AND2_X1 U11403 ( .A1(n9695), .A2(n9819), .ZN(n10350) );
  AND2_X1 U11404 ( .A1(n14224), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10232) );
  AND2_X1 U11405 ( .A1(n10238), .A2(n13258), .ZN(n10242) );
  NAND2_X1 U11406 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11463) );
  INV_X2 U11407 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19235) );
  AND2_X2 U11408 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13263) );
  NAND2_X2 U11409 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19065) );
  NOR2_X1 U11410 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10239) );
  INV_X4 U11411 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12397) );
  NAND2_X1 U11412 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12781) );
  AND2_X1 U11413 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U11414 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13258) );
  NOR2_X2 U11415 ( .A1(n15317), .A2(n15318), .ZN(n10132) );
  AOI22_X2 U11416 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19953), .B1(
        n14241), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13706) );
  AND2_X2 U11417 ( .A1(n10407), .A2(n11775), .ZN(n10412) );
  NOR2_X4 U11418 ( .A1(n11461), .A2(n11465), .ZN(n11509) );
  NAND2_X1 U11419 ( .A1(n11879), .A2(n11878), .ZN(n9655) );
  INV_X2 U11420 ( .A(n11911), .ZN(n12298) );
  BUF_X4 U11421 ( .A(n13460), .Z(n9657) );
  AND2_X2 U11422 ( .A1(n15978), .A2(n12397), .ZN(n9658) );
  AND2_X2 U11423 ( .A1(n15978), .A2(n12397), .ZN(n9659) );
  AND2_X2 U11424 ( .A1(n15978), .A2(n12397), .ZN(n12231) );
  XNOR2_X2 U11425 ( .A(n14195), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15045) );
  NOR2_X2 U11426 ( .A1(n14194), .A2(n14193), .ZN(n14195) );
  AND2_X1 U11427 ( .A1(n15977), .A2(n12397), .ZN(n9661) );
  INV_X1 U11428 ( .A(n9661), .ZN(n9662) );
  AND2_X1 U11430 ( .A1(n15977), .A2(n12397), .ZN(n12019) );
  CLKBUF_X1 U11431 ( .A(n11422), .Z(n9664) );
  AND2_X2 U11432 ( .A1(n13716), .A2(n13929), .ZN(n14292) );
  INV_X1 U11433 ( .A(n9675), .ZN(n13785) );
  NAND2_X1 U11434 ( .A1(n11933), .A2(n12298), .ZN(n9810) );
  NAND2_X1 U11435 ( .A1(n10401), .A2(n10400), .ZN(n10420) );
  NAND2_X2 U11436 ( .A1(n13718), .A2(n16001), .ZN(n14296) );
  NOR2_X2 U11437 ( .A1(n17302), .A2(n11458), .ZN(n9666) );
  AND2_X2 U11438 ( .A1(n12856), .A2(n10397), .ZN(n10399) );
  NAND3_X4 U11439 ( .A1(n9783), .A2(n10250), .A3(n9782), .ZN(n10397) );
  NAND3_X4 U11440 ( .A1(n10215), .A2(n10294), .A3(n10293), .ZN(n13412) );
  XNOR2_X1 U11441 ( .A(n11991), .B(n11990), .ZN(n9667) );
  XNOR2_X1 U11442 ( .A(n11991), .B(n11990), .ZN(n9668) );
  OAI21_X2 U11444 ( .B1(n15952), .B2(n15951), .A(n14277), .ZN(n15936) );
  AOI211_X2 U11445 ( .C1(n19597), .C2(n19342), .A(n15548), .B(n15547), .ZN(
        n15549) );
  OAI21_X2 U11446 ( .B1(n10604), .B2(n13314), .A(n10603), .ZN(n13369) );
  NAND2_X1 U11447 ( .A1(n13548), .A2(n10531), .ZN(n13238) );
  OAI21_X1 U11448 ( .B1(n13307), .B2(n13306), .A(n13305), .ZN(n20248) );
  BUF_X2 U11449 ( .A(n13693), .Z(n9675) );
  XNOR2_X2 U11450 ( .A(n14266), .B(n14265), .ZN(n14418) );
  OAI211_X2 U11451 ( .C1(n15533), .C2(n15495), .A(n15519), .B(n15517), .ZN(
        n15509) );
  NAND2_X1 U11452 ( .A1(n10239), .A2(n13263), .ZN(n10495) );
  NAND2_X1 U11453 ( .A1(n16592), .A2(n10043), .ZN(n10035) );
  OAI211_X1 U11454 ( .C1(n16592), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n15296) );
  AND2_X1 U11455 ( .A1(n11926), .A2(n11938), .ZN(n12755) );
  NAND2_X1 U11456 ( .A1(n10227), .A2(n13461), .ZN(n9671) );
  INV_X4 U11457 ( .A(n10389), .ZN(n10644) );
  INV_X2 U11458 ( .A(n10359), .ZN(n10389) );
  NAND2_X1 U11459 ( .A1(n10252), .A2(n13263), .ZN(n10283) );
  AND3_X1 U11460 ( .A1(n13155), .A2(n11915), .A3(n11914), .ZN(n11920) );
  NAND2_X1 U11461 ( .A1(n11906), .A2(n11915), .ZN(n13156) );
  INV_X1 U11462 ( .A(n11359), .ZN(n9674) );
  NAND2_X1 U11463 ( .A1(n10045), .A2(n10044), .ZN(n10047) );
  AND2_X2 U11464 ( .A1(n13243), .A2(n10239), .ZN(n10452) );
  NOR2_X4 U11465 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13243) );
  NOR2_X1 U11466 ( .A1(n14224), .A2(n10136), .ZN(n10135) );
  NOR2_X1 U11467 ( .A1(n10426), .A2(n12861), .ZN(n9796) );
  NAND2_X1 U11468 ( .A1(n14281), .A2(n14280), .ZN(n14308) );
  INV_X1 U11469 ( .A(n10707), .ZN(n9967) );
  NOR2_X1 U11470 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U11471 ( .A1(n12453), .A2(n9723), .ZN(n11936) );
  AOI21_X1 U11472 ( .B1(n11955), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11964), .ZN(n11967) );
  NOR2_X1 U11473 ( .A1(n9655), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12489) );
  AOI21_X1 U11474 ( .B1(n19076), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11674), .ZN(n11680) );
  AND2_X1 U11475 ( .A1(n11688), .A2(n11681), .ZN(n11674) );
  OAI22_X1 U11476 ( .A1(n9868), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19081), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U11477 ( .A1(n9799), .A2(n9757), .ZN(n14612) );
  INV_X1 U11478 ( .A(n14660), .ZN(n9799) );
  INV_X1 U11479 ( .A(n10154), .ZN(n10153) );
  INV_X1 U11480 ( .A(n13810), .ZN(n9902) );
  NAND2_X1 U11481 ( .A1(n10810), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11031) );
  AND2_X1 U11482 ( .A1(n9964), .A2(n10728), .ZN(n9790) );
  AND2_X2 U11483 ( .A1(n15008), .A2(n10730), .ZN(n9984) );
  AOI21_X1 U11484 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20254), .A(
        n12401), .ZN(n12403) );
  NOR2_X1 U11485 ( .A1(n12426), .A2(n12400), .ZN(n12401) );
  OR2_X1 U11486 ( .A1(n16537), .A2(n14402), .ZN(n14411) );
  INV_X1 U11487 ( .A(n9914), .ZN(n9913) );
  OAI21_X1 U11488 ( .B1(n9918), .B2(n15698), .A(n9915), .ZN(n9914) );
  INV_X1 U11489 ( .A(n15457), .ZN(n9915) );
  NOR2_X1 U11490 ( .A1(n15464), .A2(n9921), .ZN(n9920) );
  INV_X1 U11491 ( .A(n9923), .ZN(n9921) );
  NOR2_X1 U11492 ( .A1(n10202), .A2(n15586), .ZN(n10196) );
  AND4_X1 U11493 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12592) );
  AND4_X1 U11494 ( .A1(n12590), .A2(n12589), .A3(n12588), .A4(n12587), .ZN(
        n12591) );
  AOI22_X1 U11495 ( .A1(n9648), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11973) );
  AND2_X1 U11496 ( .A1(n13057), .A2(n13056), .ZN(n12509) );
  AND2_X1 U11497 ( .A1(n17950), .A2(n10007), .ZN(n9856) );
  NOR2_X1 U11498 ( .A1(n18289), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10007) );
  XNOR2_X1 U11499 ( .A(n17765), .B(n11550), .ZN(n11566) );
  NAND2_X1 U11500 ( .A1(n9831), .A2(n16352), .ZN(n14936) );
  NAND2_X1 U11501 ( .A1(n14950), .A2(n15133), .ZN(n9831) );
  AND2_X1 U11502 ( .A1(n16330), .A2(n9684), .ZN(n9947) );
  NAND2_X1 U11503 ( .A1(n10147), .A2(n10145), .ZN(n9794) );
  INV_X1 U11504 ( .A(n14871), .ZN(n10145) );
  NAND2_X1 U11505 ( .A1(n10144), .A2(n10147), .ZN(n10748) );
  INV_X1 U11506 ( .A(n10146), .ZN(n10144) );
  OR3_X1 U11507 ( .A1(n13254), .A2(n13253), .A3(n13252), .ZN(n16230) );
  NAND2_X1 U11508 ( .A1(n9710), .A2(n14406), .ZN(n14502) );
  NAND2_X2 U11509 ( .A1(n11911), .A2(n16039), .ZN(n13081) );
  AND2_X1 U11510 ( .A1(n19537), .A2(n12656), .ZN(n13058) );
  NAND2_X1 U11511 ( .A1(n12653), .A2(n12652), .ZN(n14518) );
  INV_X1 U11512 ( .A(n14497), .ZN(n14233) );
  AOI21_X1 U11513 ( .B1(n10189), .B2(n10192), .A(n10187), .ZN(n15405) );
  AND2_X1 U11514 ( .A1(n10191), .A2(n10190), .ZN(n10189) );
  NOR2_X1 U11515 ( .A1(n10188), .A2(n14489), .ZN(n10187) );
  AND2_X1 U11516 ( .A1(n10193), .A2(n15416), .ZN(n10190) );
  NAND2_X1 U11517 ( .A1(n14484), .A2(n14489), .ZN(n9843) );
  INV_X1 U11518 ( .A(n13901), .ZN(n10057) );
  INV_X1 U11519 ( .A(n13765), .ZN(n10059) );
  NAND2_X1 U11520 ( .A1(n13145), .A2(n13144), .ZN(n13181) );
  AOI21_X1 U11521 ( .B1(n19612), .B2(n13086), .A(n12004), .ZN(n13096) );
  INV_X1 U11522 ( .A(n19286), .ZN(n13144) );
  INV_X1 U11523 ( .A(n20098), .ZN(n19782) );
  OR2_X1 U11524 ( .A1(n17271), .A2(n16976), .ZN(n10086) );
  OR2_X1 U11525 ( .A1(n16986), .A2(n10087), .ZN(n10085) );
  OR2_X1 U11526 ( .A1(n16976), .A2(n17902), .ZN(n10087) );
  NAND2_X1 U11527 ( .A1(n16775), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16762) );
  NAND2_X1 U11528 ( .A1(n9999), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9998) );
  AOI21_X1 U11529 ( .B1(n18155), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n9991), .ZN(n9990) );
  INV_X1 U11530 ( .A(n16795), .ZN(n9991) );
  AOI21_X1 U11531 ( .B1(n9864), .B2(n18195), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U11532 ( .A1(n18214), .A2(n9862), .ZN(n9866) );
  NOR2_X1 U11533 ( .A1(n18195), .A2(n9864), .ZN(n9862) );
  NAND2_X1 U11534 ( .A1(n18546), .A2(n11571), .ZN(n18215) );
  INV_X1 U11535 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16735) );
  INV_X1 U11536 ( .A(n14512), .ZN(n10124) );
  AND2_X1 U11537 ( .A1(n19537), .A2(n12666), .ZN(n19495) );
  INV_X1 U11538 ( .A(n9957), .ZN(n9956) );
  OAI21_X1 U11539 ( .B1(n15704), .B2(n16665), .A(n9958), .ZN(n9957) );
  AOI21_X1 U11540 ( .B1(n16565), .B2(n19597), .A(n15463), .ZN(n9958) );
  NAND2_X1 U11541 ( .A1(n15799), .A2(n9806), .ZN(n9805) );
  NAND2_X1 U11542 ( .A1(n19617), .A2(n15800), .ZN(n9806) );
  INV_X1 U11543 ( .A(n16756), .ZN(n17746) );
  AND2_X1 U11544 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U11545 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n9818) );
  INV_X1 U11546 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11382) );
  AOI21_X1 U11547 ( .B1(n11926), .B2(n9687), .A(n9758), .ZN(n9950) );
  AND2_X1 U11548 ( .A1(n10761), .A2(n10762), .ZN(n10759) );
  OAI211_X1 U11549 ( .C1(n12856), .C2(n16260), .A(n9797), .B(n13240), .ZN(
        n10426) );
  INV_X1 U11550 ( .A(n10370), .ZN(n9797) );
  INV_X1 U11551 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11329) );
  INV_X1 U11552 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11132) );
  INV_X1 U11553 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11326) );
  INV_X1 U11554 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11327) );
  AND2_X1 U11555 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10231) );
  INV_X1 U11556 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11256) );
  INV_X1 U11557 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10508) );
  OR2_X1 U11558 ( .A1(n11418), .A2(n10253), .ZN(n10257) );
  NOR2_X1 U11559 ( .A1(n14267), .A2(n10175), .ZN(n10171) );
  INV_X1 U11560 ( .A(n14309), .ZN(n10175) );
  AND2_X1 U11561 ( .A1(n13753), .A2(n13940), .ZN(n9933) );
  AND4_X1 U11562 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12593) );
  AND2_X1 U11563 ( .A1(n12395), .A2(n12394), .ZN(n12428) );
  OR2_X1 U11564 ( .A1(n13065), .A2(n12429), .ZN(n12395) );
  NOR2_X1 U11565 ( .A1(n17752), .A2(n11545), .ZN(n11543) );
  INV_X1 U11566 ( .A(n17749), .ZN(n11544) );
  NOR2_X1 U11567 ( .A1(n17760), .A2(n11549), .ZN(n11546) );
  INV_X1 U11568 ( .A(n17756), .ZN(n11547) );
  INV_X1 U11569 ( .A(n14626), .ZN(n10106) );
  NAND2_X1 U11570 ( .A1(n13260), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11438) );
  OR2_X1 U11571 ( .A1(n9762), .A2(n14761), .ZN(n9908) );
  INV_X1 U11572 ( .A(n14752), .ZN(n10152) );
  NAND2_X1 U11573 ( .A1(n14909), .A2(n10742), .ZN(n14192) );
  OR2_X1 U11574 ( .A1(n10099), .A2(n14593), .ZN(n10097) );
  INV_X1 U11575 ( .A(n14564), .ZN(n10099) );
  NOR2_X1 U11576 ( .A1(n14638), .A2(n10108), .ZN(n10107) );
  INV_X1 U11577 ( .A(n14650), .ZN(n10108) );
  INV_X1 U11578 ( .A(n9965), .ZN(n9964) );
  INV_X1 U11579 ( .A(n14154), .ZN(n14113) );
  NAND2_X1 U11580 ( .A1(n14204), .A2(n9817), .ZN(n14154) );
  NOR2_X1 U11581 ( .A1(n10505), .A2(n10532), .ZN(n10504) );
  NAND2_X1 U11582 ( .A1(n10408), .A2(n10134), .ZN(n10133) );
  NAND2_X1 U11583 ( .A1(n10531), .A2(n10441), .ZN(n9781) );
  NOR2_X1 U11584 ( .A1(n13475), .A2(n10440), .ZN(n9824) );
  NAND2_X1 U11585 ( .A1(n10399), .A2(n14164), .ZN(n13240) );
  AND2_X1 U11586 ( .A1(n10399), .A2(n13634), .ZN(n10403) );
  INV_X1 U11587 ( .A(n10420), .ZN(n12872) );
  NAND2_X1 U11588 ( .A1(n20663), .A2(n10532), .ZN(n10566) );
  NAND2_X1 U11589 ( .A1(n10381), .A2(n9934), .ZN(n10388) );
  NAND2_X1 U11590 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n9934) );
  OAI22_X1 U11591 ( .A1(n9672), .A2(n11327), .B1(n10495), .B2(n11326), .ZN(
        n10285) );
  NAND2_X1 U11592 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U11593 ( .A1(n9786), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9785) );
  AOI22_X1 U11594 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9788), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n9787) );
  AND2_X1 U11595 ( .A1(n10545), .A2(n20894), .ZN(n20664) );
  NOR2_X1 U11596 ( .A1(n14415), .A2(n10184), .ZN(n10183) );
  AND2_X1 U11597 ( .A1(n14320), .A2(n13493), .ZN(n14326) );
  NAND2_X1 U11598 ( .A1(n10171), .A2(n14313), .ZN(n10173) );
  NAND2_X1 U11599 ( .A1(n13897), .A2(n13898), .ZN(n14268) );
  AND2_X1 U11600 ( .A1(n12824), .A2(n14009), .ZN(n10075) );
  NOR2_X1 U11601 ( .A1(n15275), .A2(n10128), .ZN(n10127) );
  INV_X1 U11602 ( .A(n15267), .ZN(n10128) );
  NAND2_X1 U11603 ( .A1(n10122), .A2(n13872), .ZN(n10121) );
  INV_X1 U11604 ( .A(n13516), .ZN(n10122) );
  NAND2_X1 U11605 ( .A1(n10072), .A2(n15357), .ZN(n10071) );
  INV_X1 U11606 ( .A(n15371), .ZN(n10072) );
  INV_X1 U11607 ( .A(n15363), .ZN(n10073) );
  AND2_X1 U11608 ( .A1(n12621), .A2(n12620), .ZN(n15234) );
  INV_X1 U11609 ( .A(n16637), .ZN(n9961) );
  NAND2_X1 U11610 ( .A1(n14336), .A2(n10204), .ZN(n10203) );
  NOR2_X1 U11611 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  INV_X1 U11612 ( .A(n13489), .ZN(n10120) );
  INV_X1 U11613 ( .A(n13526), .ZN(n10118) );
  NAND2_X1 U11614 ( .A1(n14428), .A2(n14497), .ZN(n14434) );
  INV_X1 U11615 ( .A(n14427), .ZN(n14428) );
  INV_X1 U11616 ( .A(n11967), .ZN(n11965) );
  NAND2_X1 U11617 ( .A1(n11994), .A2(n11993), .ZN(n11996) );
  NOR2_X1 U11618 ( .A1(n12511), .A2(n12510), .ZN(n12527) );
  OR2_X1 U11619 ( .A1(n9676), .A2(n13700), .ZN(n14237) );
  NOR2_X1 U11620 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19235), .ZN(
        n11681) );
  OR2_X1 U11621 ( .A1(n17302), .A2(n9867), .ZN(n11462) );
  NAND2_X1 U11622 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  NOR4_X1 U11623 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n19235), .ZN(n11640) );
  INV_X1 U11624 ( .A(n11510), .ZN(n17522) );
  NOR3_X1 U11625 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n11465), .ZN(n11486) );
  NAND2_X1 U11626 ( .A1(n11519), .A2(n10003), .ZN(n10002) );
  NAND2_X1 U11627 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10003) );
  NAND2_X1 U11628 ( .A1(n11709), .A2(n17622), .ZN(n11714) );
  NOR2_X1 U11629 ( .A1(n9852), .A2(n17939), .ZN(n11587) );
  NAND2_X1 U11630 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  NAND2_X1 U11631 ( .A1(n18142), .A2(n18272), .ZN(n9853) );
  AND2_X1 U11632 ( .A1(n17729), .A2(n18619), .ZN(n11724) );
  NAND2_X1 U11633 ( .A1(n18169), .A2(n11577), .ZN(n11580) );
  NAND2_X1 U11634 ( .A1(n11546), .A2(n11547), .ZN(n11545) );
  AOI21_X1 U11635 ( .B1(n11680), .B2(n11679), .A(n11678), .ZN(n11690) );
  INV_X1 U11636 ( .A(n10397), .ZN(n10295) );
  AND2_X1 U11637 ( .A1(n10159), .A2(n14698), .ZN(n10158) );
  AOI21_X1 U11638 ( .B1(n14064), .B2(n11170), .A(n10904), .ZN(n13991) );
  NAND2_X1 U11639 ( .A1(n13328), .A2(n10826), .ZN(n13325) );
  NAND2_X1 U11640 ( .A1(n10166), .A2(n10162), .ZN(n14189) );
  NOR2_X1 U11641 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  INV_X1 U11642 ( .A(n14190), .ZN(n10163) );
  NAND2_X1 U11643 ( .A1(n14562), .A2(n14547), .ZN(n14546) );
  AND2_X1 U11644 ( .A1(n14962), .A2(n10741), .ZN(n14975) );
  NAND2_X1 U11645 ( .A1(n10839), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10846) );
  INV_X1 U11646 ( .A(n14192), .ZN(n10745) );
  NOR2_X1 U11647 ( .A1(n14872), .A2(n15066), .ZN(n9937) );
  AND2_X1 U11648 ( .A1(n14550), .A2(n14535), .ZN(n14537) );
  NOR2_X2 U11649 ( .A1(n14603), .A2(n10096), .ZN(n14550) );
  OR3_X1 U11650 ( .A1(n14579), .A2(n10097), .A3(n10098), .ZN(n10096) );
  INV_X1 U11651 ( .A(n14548), .ZN(n10098) );
  NAND2_X1 U11652 ( .A1(n14909), .A2(n14883), .ZN(n9887) );
  NOR3_X1 U11653 ( .A1(n14603), .A2(n14579), .A3(n10097), .ZN(n14566) );
  AND2_X1 U11654 ( .A1(n9983), .A2(n9742), .ZN(n9834) );
  NAND2_X1 U11655 ( .A1(n14757), .A2(n10101), .ZN(n10100) );
  NOR2_X1 U11656 ( .A1(n14683), .A2(n10102), .ZN(n10101) );
  NAND2_X1 U11657 ( .A1(n10093), .A2(n10092), .ZN(n14781) );
  INV_X1 U11658 ( .A(n14071), .ZN(n10092) );
  INV_X1 U11659 ( .A(n10719), .ZN(n9943) );
  NAND2_X1 U11660 ( .A1(n9835), .A2(n10671), .ZN(n13663) );
  NAND2_X1 U11661 ( .A1(n10607), .A2(n10606), .ZN(n13531) );
  OR2_X1 U11662 ( .A1(n20453), .A2(n10567), .ZN(n20609) );
  NOR2_X1 U11663 ( .A1(n10306), .A2(n10305), .ZN(n10317) );
  NOR2_X1 U11664 ( .A1(n20807), .A2(n20582), .ZN(n20725) );
  NOR2_X1 U11665 ( .A1(n20719), .A2(n20582), .ZN(n20869) );
  NAND2_X1 U11666 ( .A1(n10532), .A2(n13387), .ZN(n20582) );
  INV_X1 U11667 ( .A(n13554), .ZN(n20902) );
  NOR2_X1 U11668 ( .A1(n21061), .A2(n13209), .ZN(n16271) );
  AOI221_X1 U11669 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12403), 
        .C1(n12444), .C2(n12403), .A(n12402), .ZN(n13070) );
  OR2_X1 U11670 ( .A1(n14502), .A2(n14401), .ZN(n16537) );
  INV_X1 U11671 ( .A(n10025), .ZN(n15181) );
  OR2_X1 U11672 ( .A1(n10213), .A2(n15722), .ZN(n15724) );
  AND2_X1 U11673 ( .A1(n15308), .A2(n15306), .ZN(n12162) );
  AND2_X1 U11674 ( .A1(n15926), .A2(n10064), .ZN(n15864) );
  AND2_X1 U11675 ( .A1(n10065), .A2(n12609), .ZN(n10064) );
  AND2_X1 U11676 ( .A1(n15895), .A2(n15865), .ZN(n12609) );
  INV_X1 U11677 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U11678 ( .A1(n15285), .A2(n10125), .ZN(n15269) );
  INV_X1 U11679 ( .A(n10127), .ZN(n10125) );
  NAND2_X1 U11680 ( .A1(n15905), .A2(n9894), .ZN(n14471) );
  NOR2_X1 U11681 ( .A1(n15285), .A2(n15275), .ZN(n15276) );
  NAND2_X1 U11682 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  OR2_X1 U11683 ( .A1(n9682), .A2(n9913), .ZN(n9850) );
  NAND2_X1 U11684 ( .A1(n9682), .A2(n9919), .ZN(n9849) );
  NAND2_X1 U11685 ( .A1(n9744), .A2(n9924), .ZN(n9923) );
  INV_X1 U11686 ( .A(n15476), .ZN(n9924) );
  NAND2_X1 U11687 ( .A1(n15781), .A2(n9701), .ZN(n15522) );
  NAND2_X1 U11688 ( .A1(n15633), .A2(n9844), .ZN(n10197) );
  NOR2_X1 U11689 ( .A1(n14345), .A2(n10199), .ZN(n10198) );
  NOR2_X1 U11690 ( .A1(n15617), .A2(n10205), .ZN(n10204) );
  NAND2_X1 U11691 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  INV_X1 U11692 ( .A(n15917), .ZN(n10206) );
  AND2_X1 U11693 ( .A1(n15633), .A2(n9845), .ZN(n15615) );
  AND2_X1 U11694 ( .A1(n14318), .A2(n9846), .ZN(n9845) );
  AND2_X1 U11695 ( .A1(n10057), .A2(n15960), .ZN(n10056) );
  NAND2_X1 U11696 ( .A1(n10054), .A2(n10058), .ZN(n13900) );
  NAND2_X1 U11697 ( .A1(n11998), .A2(n12001), .ZN(n19612) );
  AND2_X1 U11698 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11983), .ZN(
        n19839) );
  NOR2_X1 U11699 ( .A1(n20258), .A2(n20267), .ZN(n19667) );
  NAND2_X1 U11700 ( .A1(n20258), .A2(n20265), .ZN(n19781) );
  NAND2_X1 U11701 ( .A1(n11884), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11891) );
  NAND2_X1 U11702 ( .A1(n11889), .A2(n12026), .ZN(n11890) );
  AND2_X1 U11703 ( .A1(n20258), .A2(n20267), .ZN(n20045) );
  INV_X1 U11704 ( .A(n20045), .ZN(n20241) );
  OR2_X1 U11705 ( .A1(n16732), .A2(n16027), .ZN(n16028) );
  AND2_X1 U11706 ( .A1(n16747), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16775) );
  NOR2_X1 U11707 ( .A1(n11637), .A2(n11636), .ZN(n16946) );
  BUF_X1 U11708 ( .A(n11640), .Z(n17576) );
  NOR4_X2 U11709 ( .A1(n16946), .A2(n11715), .A3(n18627), .A4(n11714), .ZN(
        n17838) );
  NOR2_X1 U11710 ( .A1(n16781), .A2(n16777), .ZN(n16747) );
  OR2_X1 U11711 ( .A1(n17900), .A2(n17892), .ZN(n16781) );
  AND2_X1 U11712 ( .A1(n17919), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17894) );
  INV_X1 U11713 ( .A(n16748), .ZN(n17919) );
  NOR2_X1 U11714 ( .A1(n10081), .A2(n10079), .ZN(n10078) );
  NAND2_X1 U11715 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11716 ( .A1(n11585), .A2(n9855), .ZN(n17923) );
  NOR2_X1 U11717 ( .A1(n10004), .A2(n9856), .ZN(n9855) );
  NAND2_X1 U11718 ( .A1(n10005), .A2(n9756), .ZN(n10004) );
  NAND2_X1 U11719 ( .A1(n11580), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18460) );
  NAND2_X1 U11720 ( .A1(n18460), .A2(n18142), .ZN(n9988) );
  NAND2_X1 U11721 ( .A1(n9987), .A2(n18460), .ZN(n18164) );
  NOR2_X1 U11722 ( .A1(n9860), .A2(n9858), .ZN(n9857) );
  AND2_X1 U11723 ( .A1(n18214), .A2(n9863), .ZN(n9860) );
  NAND2_X1 U11724 ( .A1(n18237), .A2(n11567), .ZN(n11570) );
  XNOR2_X1 U11725 ( .A(n11566), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18239) );
  NAND2_X1 U11726 ( .A1(n18238), .A2(n18239), .ZN(n18237) );
  INV_X1 U11727 ( .A(n18627), .ZN(n11712) );
  INV_X1 U11728 ( .A(n20345), .ZN(n20377) );
  NAND2_X2 U11729 ( .A1(n13284), .A2(n13283), .ZN(n14770) );
  OR2_X1 U11730 ( .A1(n13282), .A2(n14158), .ZN(n13283) );
  OR2_X1 U11731 ( .A1(n13281), .A2(n20294), .ZN(n13284) );
  OAI21_X1 U11732 ( .B1(n14531), .B2(n14190), .A(n14189), .ZN(n14217) );
  NAND2_X1 U11733 ( .A1(n14561), .A2(n14563), .ZN(n9910) );
  INV_X1 U11734 ( .A(n14562), .ZN(n9909) );
  XNOR2_X1 U11735 ( .A(n10139), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15044) );
  NAND2_X1 U11736 ( .A1(n10750), .A2(n10749), .ZN(n10139) );
  AND2_X1 U11737 ( .A1(n12881), .A2(n12880), .ZN(n16445) );
  AND2_X1 U11738 ( .A1(n12931), .A2(n12930), .ZN(n20438) );
  INV_X1 U11739 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20690) );
  INV_X1 U11740 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20862) );
  INV_X1 U11741 ( .A(n20959), .ZN(n20945) );
  XNOR2_X1 U11742 ( .A(n12392), .B(n12391), .ZN(n12678) );
  OR2_X1 U11743 ( .A1(n16506), .A2(n19538), .ZN(n12673) );
  NAND2_X1 U11744 ( .A1(n15325), .A2(n15324), .ZN(n16516) );
  OR2_X1 U11745 ( .A1(n13016), .A2(n13160), .ZN(n12473) );
  AND2_X1 U11746 ( .A1(n19537), .A2(n12486), .ZN(n16619) );
  NOR2_X1 U11747 ( .A1(n15441), .A2(n16664), .ZN(n9954) );
  OR2_X1 U11748 ( .A1(n19288), .A2(n9636), .ZN(n16665) );
  INV_X1 U11749 ( .A(n16664), .ZN(n19595) );
  XNOR2_X1 U11750 ( .A(n14518), .B(n14517), .ZN(n16500) );
  XNOR2_X1 U11751 ( .A(n9889), .B(n14509), .ZN(n14527) );
  OR2_X1 U11752 ( .A1(n14526), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U11753 ( .A1(n14523), .A2(n14524), .ZN(n10062) );
  XOR2_X1 U11754 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14503), .Z(
        n14504) );
  NAND2_X1 U11755 ( .A1(n10185), .A2(n14489), .ZN(n15417) );
  NAND2_X1 U11756 ( .A1(n10192), .A2(n10186), .ZN(n10185) );
  XNOR2_X1 U11757 ( .A(n9841), .B(n14416), .ZN(n14470) );
  OAI21_X1 U11758 ( .B1(n14472), .B2(n14486), .A(n9842), .ZN(n9841) );
  NAND2_X1 U11759 ( .A1(n9843), .A2(n9927), .ZN(n9842) );
  NAND2_X1 U11760 ( .A1(n9851), .A2(n9918), .ZN(n15459) );
  OR2_X1 U11761 ( .A1(n14387), .A2(n9919), .ZN(n9851) );
  NAND2_X1 U11762 ( .A1(n9809), .A2(n9808), .ZN(n9807) );
  NAND2_X1 U11763 ( .A1(n15785), .A2(n15784), .ZN(n9808) );
  OR2_X1 U11764 ( .A1(n13181), .A2(n13147), .ZN(n16677) );
  AND2_X1 U11765 ( .A1(n13173), .A2(n20289), .ZN(n19611) );
  INV_X1 U11766 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20254) );
  NAND2_X1 U11767 ( .A1(n12010), .A2(n12009), .ZN(n14054) );
  NAND2_X1 U11768 ( .A1(n14053), .A2(n13086), .ZN(n12010) );
  AND2_X1 U11769 ( .A1(n10086), .A2(n17271), .ZN(n10084) );
  INV_X1 U11770 ( .A(n17286), .ZN(n17305) );
  INV_X1 U11771 ( .A(n17314), .ZN(n17280) );
  INV_X1 U11772 ( .A(n17315), .ZN(n17285) );
  AND2_X1 U11773 ( .A1(n9997), .A2(n9995), .ZN(n16800) );
  NAND2_X1 U11774 ( .A1(n18575), .A2(n18406), .ZN(n18509) );
  OR2_X1 U11775 ( .A1(n10771), .A2(n10770), .ZN(n10774) );
  NAND2_X1 U11776 ( .A1(n14236), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14239) );
  INV_X1 U11777 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11207) );
  INV_X1 U11778 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11243) );
  INV_X1 U11779 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11246) );
  INV_X1 U11780 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U11781 ( .A1(n11866), .A2(n11906), .ZN(n10031) );
  INV_X1 U11782 ( .A(n11866), .ZN(n10032) );
  AND4_X1 U11783 ( .A1(n14291), .A2(n14290), .A3(n14289), .A4(n14288), .ZN(
        n14302) );
  NOR2_X1 U11784 ( .A1(n14249), .A2(n14248), .ZN(n14260) );
  AOI22_X1 U11785 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13704), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13705) );
  OR2_X1 U11786 ( .A1(n11679), .A2(n11680), .ZN(n11675) );
  INV_X1 U11787 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11352) );
  NOR2_X1 U11788 ( .A1(n13991), .A2(n10151), .ZN(n10150) );
  INV_X1 U11789 ( .A(n14067), .ZN(n10151) );
  INV_X1 U11790 ( .A(n9672), .ZN(n11392) );
  INV_X1 U11791 ( .A(n9657), .ZN(n11412) );
  INV_X1 U11792 ( .A(n11420), .ZN(n11393) );
  NAND2_X1 U11793 ( .A1(n10662), .A2(n10661), .ZN(n10148) );
  NAND2_X1 U11794 ( .A1(n9817), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U11795 ( .A1(n10420), .A2(n13634), .ZN(n9795) );
  NOR2_X1 U11796 ( .A1(n10409), .A2(n10136), .ZN(n10134) );
  NAND2_X1 U11797 ( .A1(n10408), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U11798 ( .A1(n9828), .A2(n10567), .ZN(n10642) );
  NAND2_X1 U11799 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n9977) );
  INV_X1 U11800 ( .A(n9656), .ZN(n9786) );
  INV_X1 U11801 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11419) );
  INV_X1 U11802 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11407) );
  INV_X1 U11803 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11421) );
  NAND2_X1 U11804 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n9882) );
  INV_X1 U11805 ( .A(n12696), .ZN(n11971) );
  OR2_X1 U11806 ( .A1(n12565), .A2(n12564), .ZN(n12810) );
  INV_X1 U11807 ( .A(n13942), .ZN(n14281) );
  OR2_X1 U11808 ( .A1(n12414), .A2(n12413), .ZN(n14278) );
  AOI22_X1 U11809 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n14295), .B1(
        n16083), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13719) );
  AND2_X1 U11810 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  AND2_X1 U11811 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10169) );
  AOI21_X1 U11812 ( .B1(n12581), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n10170), .ZN(n12497) );
  OR2_X1 U11813 ( .A1(n12424), .A2(n12423), .ZN(n12531) );
  INV_X1 U11814 ( .A(n13156), .ZN(n13151) );
  NAND2_X1 U11815 ( .A1(n11908), .A2(n11914), .ZN(n11934) );
  XNOR2_X1 U11816 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12425) );
  NAND2_X1 U11817 ( .A1(n12399), .A2(n12398), .ZN(n12426) );
  AOI21_X1 U11818 ( .B1(n9646), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12026), .ZN(n11813) );
  NOR2_X1 U11819 ( .A1(n11463), .A2(n11465), .ZN(n11510) );
  NOR2_X1 U11820 ( .A1(n11463), .A2(n17302), .ZN(n11464) );
  NAND2_X1 U11821 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n9869), .ZN(
        n11461) );
  AOI221_X1 U11822 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10758), 
        .C1(n16486), .C2(n10758), .A(n10756), .ZN(n11781) );
  NAND2_X1 U11823 ( .A1(n10167), .A2(n10165), .ZN(n10164) );
  INV_X1 U11824 ( .A(n14563), .ZN(n10165) );
  NOR2_X1 U11825 ( .A1(n14532), .A2(n10168), .ZN(n10167) );
  INV_X1 U11826 ( .A(n14547), .ZN(n10168) );
  NAND2_X1 U11827 ( .A1(n14647), .A2(n10157), .ZN(n10156) );
  INV_X1 U11828 ( .A(n14661), .ZN(n10157) );
  OR2_X1 U11829 ( .A1(n10723), .A2(n10734), .ZN(n9684) );
  NOR2_X1 U11830 ( .A1(n10993), .A2(n10160), .ZN(n10159) );
  INV_X1 U11831 ( .A(n14721), .ZN(n10160) );
  AOI21_X1 U11832 ( .B1(n10723), .B2(n15023), .A(n14937), .ZN(n9832) );
  NAND2_X1 U11833 ( .A1(n14948), .A2(n10723), .ZN(n9798) );
  NAND2_X1 U11834 ( .A1(n10103), .A2(n14753), .ZN(n10102) );
  INV_X1 U11835 ( .A(n14699), .ZN(n10103) );
  INV_X1 U11836 ( .A(n15145), .ZN(n9884) );
  NOR2_X1 U11837 ( .A1(n9821), .A2(n10693), .ZN(n9820) );
  INV_X1 U11838 ( .A(n10661), .ZN(n9821) );
  AND3_X1 U11839 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10535) );
  NAND2_X1 U11840 ( .A1(n9830), .A2(n9829), .ZN(n10537) );
  NAND2_X1 U11841 ( .A1(n9735), .A2(n10575), .ZN(n9829) );
  INV_X1 U11842 ( .A(n10598), .ZN(n10143) );
  INV_X1 U11843 ( .A(n10550), .ZN(n10142) );
  INV_X1 U11844 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U11845 ( .A1(n10300), .A2(n9833), .ZN(n10306) );
  OR2_X1 U11846 ( .A1(n10334), .A2(n10333), .ZN(n10223) );
  OR2_X1 U11847 ( .A1(n11422), .A2(n11257), .ZN(n10320) );
  NOR2_X1 U11848 ( .A1(n10259), .A2(n10258), .ZN(n10274) );
  OAI21_X1 U11849 ( .B1(n21068), .B2(n13383), .A(n13382), .ZN(n13387) );
  OR2_X1 U11850 ( .A1(n12521), .A2(n12520), .ZN(n12806) );
  NAND2_X1 U11851 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  NOR2_X1 U11852 ( .A1(n10179), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10177) );
  INV_X1 U11853 ( .A(n14392), .ZN(n10178) );
  NAND2_X1 U11854 ( .A1(n15288), .A2(n15278), .ZN(n10179) );
  OR2_X1 U11855 ( .A1(n14369), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14390) );
  AND2_X1 U11856 ( .A1(n9681), .A2(n9759), .ZN(n10180) );
  NOR2_X1 U11857 ( .A1(n14000), .A2(n10182), .ZN(n10181) );
  NAND2_X1 U11858 ( .A1(n14335), .A2(n14342), .ZN(n14344) );
  NOR2_X1 U11859 ( .A1(n14268), .A2(n10174), .ZN(n14315) );
  NOR2_X1 U11860 ( .A1(n14268), .A2(n14267), .ZN(n14310) );
  NAND2_X1 U11861 ( .A1(n13126), .A2(n13127), .ZN(n13756) );
  AOI211_X1 U11862 ( .C1(n12330), .C2(n12326), .A(n13443), .B(n12369), .ZN(
        n12327) );
  NAND2_X1 U11863 ( .A1(n15294), .A2(n10046), .ZN(n10045) );
  INV_X1 U11864 ( .A(n15281), .ZN(n10046) );
  INV_X1 U11865 ( .A(n16588), .ZN(n10039) );
  NOR2_X1 U11866 ( .A1(n16591), .A2(n10042), .ZN(n10041) );
  INV_X1 U11867 ( .A(n15301), .ZN(n10042) );
  AND2_X1 U11868 ( .A1(n10066), .A2(n15908), .ZN(n10065) );
  NOR2_X1 U11869 ( .A1(n13869), .A2(n10067), .ZN(n10066) );
  INV_X1 U11870 ( .A(n15925), .ZN(n10067) );
  INV_X1 U11871 ( .A(n11936), .ZN(n12471) );
  NAND2_X1 U11872 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n10015), .ZN(
        n10014) );
  NOR2_X1 U11873 ( .A1(n15431), .A2(n10016), .ZN(n10015) );
  NOR2_X1 U11874 ( .A1(n15467), .A2(n10020), .ZN(n10019) );
  NOR2_X1 U11875 ( .A1(n15176), .A2(n19335), .ZN(n10025) );
  NOR2_X1 U11876 ( .A1(n15624), .A2(n10024), .ZN(n10023) );
  INV_X1 U11877 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10024) );
  INV_X1 U11878 ( .A(n15416), .ZN(n10188) );
  NAND2_X1 U11879 ( .A1(n14487), .A2(n15662), .ZN(n10193) );
  NAND2_X1 U11880 ( .A1(n10194), .A2(n10195), .ZN(n10191) );
  AND2_X1 U11881 ( .A1(n9699), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9894) );
  NAND2_X1 U11882 ( .A1(n9913), .A2(n9916), .ZN(n9848) );
  NAND2_X1 U11883 ( .A1(n9917), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9916) );
  INV_X1 U11884 ( .A(n9919), .ZN(n9917) );
  OR2_X1 U11885 ( .A1(n19336), .A2(n14384), .ZN(n15493) );
  INV_X1 U11886 ( .A(n13986), .ZN(n10109) );
  OR3_X1 U11887 ( .A1(n15245), .A2(n14233), .A3(n15800), .ZN(n15490) );
  NOR2_X1 U11888 ( .A1(n12818), .A2(n10111), .ZN(n10110) );
  INV_X1 U11889 ( .A(n15603), .ZN(n10111) );
  INV_X1 U11890 ( .A(n10204), .ZN(n10199) );
  INV_X1 U11891 ( .A(n16645), .ZN(n9846) );
  NOR2_X1 U11892 ( .A1(n12551), .A2(n12550), .ZN(n14262) );
  INV_X1 U11893 ( .A(n12619), .ZN(n12553) );
  OAI21_X1 U11894 ( .B1(n9813), .B2(n13937), .A(n13939), .ZN(n13946) );
  NAND2_X1 U11895 ( .A1(n12794), .A2(n12448), .ZN(n12465) );
  NAND2_X1 U11896 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  NOR2_X1 U11897 ( .A1(n13019), .A2(n12459), .ZN(n15991) );
  NAND2_X1 U11898 ( .A1(n13164), .A2(n11914), .ZN(n9932) );
  AOI22_X1 U11899 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11892) );
  AOI21_X1 U11900 ( .B1(n12020), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12026), .ZN(n11898) );
  NAND3_X1 U11901 ( .A1(n20243), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20098), 
        .ZN(n16041) );
  NAND2_X1 U11902 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20281), .ZN(
        n12429) );
  INV_X1 U11903 ( .A(n12445), .ZN(n13132) );
  NAND2_X1 U11904 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19235), .ZN(
        n11465) );
  NAND2_X1 U11905 ( .A1(n18616), .A2(n11724), .ZN(n11715) );
  NOR2_X1 U11906 ( .A1(n17134), .A2(n10091), .ZN(n10090) );
  NAND2_X1 U11907 ( .A1(n18025), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10005) );
  AND2_X1 U11908 ( .A1(n10009), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10006) );
  NAND2_X1 U11909 ( .A1(n10012), .A2(n10010), .ZN(n10009) );
  AND2_X1 U11910 ( .A1(n10011), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10010) );
  INV_X1 U11911 ( .A(n18325), .ZN(n10012) );
  NOR2_X1 U11912 ( .A1(n18018), .A2(n17964), .ZN(n10011) );
  INV_X1 U11913 ( .A(n18460), .ZN(n18066) );
  NAND2_X1 U11914 ( .A1(n18182), .A2(n11574), .ZN(n11575) );
  NOR2_X1 U11915 ( .A1(n11746), .A2(n18198), .ZN(n11748) );
  INV_X1 U11916 ( .A(n14096), .ZN(n19048) );
  NOR2_X1 U11917 ( .A1(n11627), .A2(n11626), .ZN(n11709) );
  NAND2_X1 U11918 ( .A1(n10882), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10921) );
  INV_X1 U11919 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20322) );
  NOR2_X1 U11920 ( .A1(n13790), .A2(n13792), .ZN(n20366) );
  INV_X1 U11921 ( .A(n13651), .ZN(n13791) );
  AND2_X1 U11922 ( .A1(n13650), .A2(n13649), .ZN(n13683) );
  INV_X1 U11923 ( .A(n14121), .ZN(n14165) );
  AND2_X1 U11924 ( .A1(n14664), .A2(n9755), .ZN(n14614) );
  INV_X1 U11925 ( .A(n14615), .ZN(n10105) );
  NAND2_X1 U11926 ( .A1(n14664), .A2(n9747), .ZN(n14628) );
  AND2_X1 U11927 ( .A1(n14677), .A2(n14662), .ZN(n14664) );
  NAND2_X1 U11928 ( .A1(n9817), .A2(n13817), .ZN(n12908) );
  NAND2_X1 U11929 ( .A1(n11784), .A2(n11783), .ZN(n13253) );
  AND2_X1 U11930 ( .A1(n20769), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11443) );
  NAND2_X1 U11931 ( .A1(n11374), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11440) );
  NOR2_X1 U11932 ( .A1(n14563), .A2(n9912), .ZN(n9911) );
  INV_X1 U11933 ( .A(n14577), .ZN(n9912) );
  OR2_X1 U11934 ( .A1(n11320), .A2(n14915), .ZN(n11321) );
  NAND2_X1 U11935 ( .A1(n11267), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11320) );
  AND2_X1 U11936 ( .A1(n11194), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11195) );
  INV_X1 U11937 ( .A(n11193), .ZN(n11194) );
  NAND2_X1 U11938 ( .A1(n14637), .A2(n10155), .ZN(n10154) );
  INV_X1 U11939 ( .A(n10156), .ZN(n10155) );
  AOI21_X1 U11940 ( .B1(n11200), .B2(n11199), .A(n11198), .ZN(n14625) );
  NAND2_X1 U11941 ( .A1(n9907), .A2(n11100), .ZN(n9906) );
  INV_X1 U11942 ( .A(n9908), .ZN(n9907) );
  CLKBUF_X1 U11943 ( .A(n14612), .Z(n14624) );
  NAND2_X1 U11944 ( .A1(n11144), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11193) );
  AND2_X1 U11945 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n11075), .ZN(
        n11076) );
  NAND2_X1 U11946 ( .A1(n11076), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11143) );
  INV_X1 U11947 ( .A(n11071), .ZN(n11075) );
  NOR2_X1 U11948 ( .A1(n11034), .A2(n11033), .ZN(n11035) );
  NAND2_X1 U11949 ( .A1(n11013), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11034) );
  NOR2_X1 U11950 ( .A1(n10994), .A2(n14713), .ZN(n11013) );
  OR2_X1 U11951 ( .A1(n10973), .A2(n14724), .ZN(n10994) );
  INV_X1 U11952 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14724) );
  AND2_X1 U11953 ( .A1(n10925), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10926) );
  NAND2_X1 U11954 ( .A1(n10926), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10973) );
  NOR2_X1 U11955 ( .A1(n10921), .A2(n20322), .ZN(n10925) );
  INV_X1 U11956 ( .A(n13991), .ZN(n10149) );
  AND2_X1 U11957 ( .A1(n10852), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10858) );
  NOR2_X1 U11958 ( .A1(n10846), .A2(n16376), .ZN(n10852) );
  INV_X1 U11959 ( .A(n13533), .ZN(n10843) );
  INV_X1 U11960 ( .A(n13323), .ZN(n9801) );
  AND2_X1 U11961 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10827), .ZN(
        n10839) );
  NAND2_X1 U11962 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10828) );
  INV_X1 U11963 ( .A(n13231), .ZN(n10825) );
  NAND2_X1 U11964 ( .A1(n10745), .A2(n10744), .ZN(n14903) );
  NOR3_X1 U11965 ( .A1(n14603), .A2(n14579), .A3(n14593), .ZN(n14578) );
  NAND2_X1 U11966 ( .A1(n14664), .A2(n10107), .ZN(n14640) );
  NAND2_X1 U11967 ( .A1(n14664), .A2(n14650), .ZN(n14652) );
  AND2_X1 U11968 ( .A1(n16330), .A2(n9691), .ZN(n9945) );
  NOR2_X2 U11969 ( .A1(n9705), .A2(n14675), .ZN(n14677) );
  NOR2_X1 U11970 ( .A1(n10723), .A2(n10739), .ZN(n14990) );
  NOR3_X1 U11971 ( .A1(n14708), .A2(n10104), .A3(n14699), .ZN(n14760) );
  NOR2_X1 U11972 ( .A1(n14708), .A2(n14699), .ZN(n14758) );
  NAND2_X1 U11973 ( .A1(n9817), .A2(n14114), .ZN(n14115) );
  OR2_X1 U11974 ( .A1(n14710), .A2(n14711), .ZN(n14708) );
  NAND2_X1 U11975 ( .A1(n14780), .A2(n12926), .ZN(n14710) );
  INV_X1 U11976 ( .A(n9940), .ZN(n9939) );
  NAND2_X1 U11977 ( .A1(n9966), .A2(n9790), .ZN(n9789) );
  OAI21_X1 U11978 ( .B1(n9942), .B2(n9941), .A(n10729), .ZN(n9940) );
  NAND2_X1 U11979 ( .A1(n9817), .A2(n20323), .ZN(n12914) );
  NAND2_X1 U11980 ( .A1(n13912), .A2(n13911), .ZN(n13995) );
  AND2_X1 U11981 ( .A1(n12907), .A2(n12906), .ZN(n13658) );
  NOR2_X1 U11982 ( .A1(n13659), .A2(n13658), .ZN(n13815) );
  AND2_X1 U11983 ( .A1(n12899), .A2(n12898), .ZN(n13544) );
  NAND2_X1 U11984 ( .A1(n9817), .A2(n12900), .ZN(n12901) );
  NAND2_X1 U11985 ( .A1(n10095), .A2(n10094), .ZN(n13659) );
  NOR2_X1 U11986 ( .A1(n13543), .A2(n13544), .ZN(n10094) );
  INV_X1 U11987 ( .A(n13545), .ZN(n10095) );
  NAND2_X1 U11988 ( .A1(n9962), .A2(n10640), .ZN(n9793) );
  XNOR2_X1 U11989 ( .A(n10605), .B(n10572), .ZN(n13370) );
  INV_X1 U11990 ( .A(n20442), .ZN(n15151) );
  NAND2_X1 U11991 ( .A1(n13286), .A2(n9817), .ZN(n13285) );
  NOR2_X1 U11992 ( .A1(n12876), .A2(n12875), .ZN(n20441) );
  AND2_X1 U11993 ( .A1(n14204), .A2(n14150), .ZN(n14121) );
  NAND2_X1 U11994 ( .A1(n10812), .A2(n10532), .ZN(n10574) );
  NAND2_X1 U11995 ( .A1(n10541), .A2(n10540), .ZN(n10596) );
  INV_X1 U11996 ( .A(n20452), .ZN(n13498) );
  NAND2_X1 U11997 ( .A1(n13475), .A2(n10440), .ZN(n9825) );
  AND2_X2 U11998 ( .A1(n13263), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13262) );
  INV_X1 U11999 ( .A(n20294), .ZN(n20300) );
  NOR2_X1 U12000 ( .A1(n10378), .A2(n10377), .ZN(n10394) );
  NOR2_X1 U12001 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  NOR2_X1 U12002 ( .A1(n10230), .A2(n10249), .ZN(n9782) );
  OR2_X1 U12003 ( .A1(n13553), .A2(n13552), .ZN(n20454) );
  OR2_X1 U12004 ( .A1(n13474), .A2(n13473), .ZN(n16244) );
  OR2_X1 U12005 ( .A1(n14493), .A2(n14492), .ZN(n14498) );
  INV_X1 U12006 ( .A(n14493), .ZN(n14490) );
  NOR3_X1 U12007 ( .A1(n14393), .A2(n14392), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n14408) );
  NAND2_X1 U12008 ( .A1(n14373), .A2(n15208), .ZN(n14369) );
  NAND2_X1 U12009 ( .A1(n13865), .A2(n19650), .ZN(n14406) );
  NAND2_X1 U12010 ( .A1(n14335), .A2(n9681), .ZN(n14362) );
  NOR2_X1 U12011 ( .A1(n14268), .A2(n10173), .ZN(n13865) );
  NOR2_X2 U12012 ( .A1(n14268), .A2(n9719), .ZN(n14320) );
  INV_X1 U12013 ( .A(n13864), .ZN(n10172) );
  NAND2_X1 U12014 ( .A1(n11969), .A2(n10211), .ZN(n10210) );
  INV_X1 U12015 ( .A(n11990), .ZN(n10211) );
  XNOR2_X1 U12016 ( .A(n10047), .B(n12275), .ZN(n15274) );
  NOR3_X1 U12017 ( .A1(n15724), .A2(n10073), .A3(n15371), .ZN(n15365) );
  NOR2_X1 U12018 ( .A1(n15724), .A2(n15371), .ZN(n15372) );
  INV_X1 U12019 ( .A(n15234), .ZN(n10074) );
  NAND2_X1 U12020 ( .A1(n12821), .A2(n9746), .ZN(n15810) );
  AND2_X1 U12021 ( .A1(n12821), .A2(n10075), .ZN(n15812) );
  AND2_X1 U12022 ( .A1(n15926), .A2(n10065), .ZN(n15906) );
  INV_X1 U12023 ( .A(n11919), .ZN(n12453) );
  NAND2_X1 U12024 ( .A1(n14516), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10053) );
  INV_X1 U12025 ( .A(n12968), .ZN(n16042) );
  NOR2_X1 U12026 ( .A1(n15191), .A2(n10014), .ZN(n15423) );
  NAND2_X1 U12027 ( .A1(n10129), .A2(n10127), .ZN(n10126) );
  NOR2_X1 U12028 ( .A1(n14442), .A2(n10130), .ZN(n10129) );
  INV_X1 U12029 ( .A(n14473), .ZN(n10130) );
  NOR2_X1 U12030 ( .A1(n15191), .A2(n15431), .ZN(n15190) );
  OR2_X1 U12031 ( .A1(n15187), .A2(n15169), .ZN(n15191) );
  NAND2_X1 U12032 ( .A1(n15185), .A2(n10018), .ZN(n15187) );
  AND2_X1 U12033 ( .A1(n9697), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10018) );
  NAND2_X1 U12034 ( .A1(n15185), .A2(n9697), .ZN(n15189) );
  NAND2_X1 U12035 ( .A1(n15185), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15186) );
  NAND2_X1 U12036 ( .A1(n10025), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15184) );
  AND2_X1 U12037 ( .A1(n15173), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15177) );
  NOR2_X1 U12038 ( .A1(n14005), .A2(n14004), .ZN(n15173) );
  NAND2_X1 U12039 ( .A1(n12788), .A2(n10022), .ZN(n14005) );
  AND2_X1 U12040 ( .A1(n9680), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U12041 ( .A1(n12788), .A2(n9680), .ZN(n12790) );
  INV_X1 U12042 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U12043 ( .A1(n12788), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12787) );
  NOR2_X1 U12044 ( .A1(n12785), .A2(n19389), .ZN(n12788) );
  NOR2_X1 U12045 ( .A1(n13526), .A2(n10121), .ZN(n13873) );
  NOR2_X1 U12046 ( .A1(n12784), .A2(n12692), .ZN(n12786) );
  NAND2_X1 U12047 ( .A1(n12786), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12785) );
  NOR2_X1 U12048 ( .A1(n13526), .A2(n13516), .ZN(n13871) );
  OAI211_X1 U12049 ( .C1(n15958), .C2(n14417), .A(n9815), .B(n14424), .ZN(
        n15946) );
  OR2_X1 U12050 ( .A1(n15954), .A2(n14307), .ZN(n14424) );
  NAND2_X1 U12051 ( .A1(n15946), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15945) );
  NOR2_X1 U12052 ( .A1(n12781), .A2(n14040), .ZN(n12783) );
  AND2_X1 U12053 ( .A1(n10191), .A2(n10193), .ZN(n10186) );
  NAND2_X1 U12054 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  NOR2_X1 U12055 ( .A1(n10073), .A2(n15347), .ZN(n10069) );
  INV_X1 U12056 ( .A(n10071), .ZN(n10070) );
  AND2_X1 U12057 ( .A1(n14403), .A2(n14411), .ZN(n15440) );
  OR2_X1 U12058 ( .A1(n14409), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15446) );
  NOR2_X1 U12059 ( .A1(n14410), .A2(n15690), .ZN(n15447) );
  AOI21_X1 U12060 ( .B1(n9920), .B2(n9926), .A(n9689), .ZN(n9918) );
  INV_X1 U12061 ( .A(n9920), .ZN(n9919) );
  OR2_X1 U12062 ( .A1(n15205), .A2(n15302), .ZN(n15479) );
  OR2_X1 U12063 ( .A1(n15747), .A2(n15712), .ZN(n15741) );
  NOR2_X1 U12064 ( .A1(n15311), .A2(n15310), .ZN(n15309) );
  NAND2_X1 U12065 ( .A1(n10132), .A2(n10131), .ZN(n15311) );
  INV_X1 U12066 ( .A(n15225), .ZN(n10131) );
  INV_X1 U12067 ( .A(n15815), .ZN(n9809) );
  NAND2_X1 U12068 ( .A1(n9960), .A2(n15788), .ZN(n9959) );
  INV_X1 U12069 ( .A(n14436), .ZN(n9960) );
  NAND2_X1 U12070 ( .A1(n15604), .A2(n10110), .ZN(n13987) );
  NAND2_X1 U12071 ( .A1(n15604), .A2(n15603), .ZN(n15606) );
  NOR2_X1 U12072 ( .A1(n15889), .A2(n10117), .ZN(n10116) );
  INV_X1 U12073 ( .A(n10119), .ZN(n10117) );
  NAND2_X1 U12074 ( .A1(n10118), .A2(n10119), .ZN(n15890) );
  AND2_X1 U12075 ( .A1(n14338), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15917) );
  NAND2_X1 U12076 ( .A1(n15926), .A2(n15925), .ZN(n15924) );
  NAND2_X1 U12077 ( .A1(n15633), .A2(n14318), .ZN(n16642) );
  AND2_X1 U12078 ( .A1(n12568), .A2(n12567), .ZN(n15938) );
  NAND2_X1 U12079 ( .A1(n14418), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15954) );
  AOI211_X1 U12080 ( .C1(n15782), .C2(n13769), .A(n13768), .B(n15786), .ZN(
        n15941) );
  CLKBUF_X1 U12081 ( .A(n12465), .Z(n12466) );
  NAND2_X1 U12082 ( .A1(n11982), .A2(n20153), .ZN(n12008) );
  NAND2_X1 U12083 ( .A1(n13279), .A2(n12015), .ZN(n13306) );
  INV_X1 U12084 ( .A(n12435), .ZN(n13030) );
  NAND2_X1 U12085 ( .A1(n20248), .A2(n20276), .ZN(n19697) );
  OR2_X1 U12086 ( .A1(n20248), .A2(n20276), .ZN(n16105) );
  INV_X1 U12087 ( .A(n19667), .ZN(n19671) );
  OR2_X1 U12088 ( .A1(n20248), .A2(n19456), .ZN(n16104) );
  INV_X1 U12089 ( .A(n19781), .ZN(n16106) );
  INV_X1 U12090 ( .A(n16105), .ZN(n19946) );
  NAND2_X1 U12091 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20098), .ZN(n19637) );
  INV_X1 U12092 ( .A(n16104), .ZN(n20046) );
  NOR2_X2 U12093 ( .A1(n16040), .A2(n16041), .ZN(n19657) );
  INV_X1 U12094 ( .A(n14295), .ZN(n20096) );
  INV_X1 U12095 ( .A(n19637), .ZN(n19658) );
  OR2_X1 U12096 ( .A1(n13070), .A2(n12464), .ZN(n16698) );
  AND2_X1 U12097 ( .A1(n12463), .A2(n12462), .ZN(n12464) );
  NOR2_X1 U12098 ( .A1(n11928), .A2(n13881), .ZN(n11921) );
  AOI21_X1 U12099 ( .B1(n11686), .B2(n11690), .A(n11689), .ZN(n19039) );
  OAI22_X1 U12100 ( .A1(n17056), .A2(n9731), .B1(n10077), .B2(n9731), .ZN(
        n17036) );
  INV_X1 U12101 ( .A(n17972), .ZN(n10077) );
  NOR2_X1 U12102 ( .A1(n17036), .A2(n17957), .ZN(n17035) );
  NOR2_X1 U12103 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17251), .ZN(n17236) );
  INV_X1 U12104 ( .A(n17308), .ZN(n17294) );
  NOR2_X1 U12105 ( .A1(n19249), .A2(n16946), .ZN(n16949) );
  NOR2_X1 U12106 ( .A1(n11465), .A2(n11458), .ZN(n11551) );
  INV_X1 U12107 ( .A(n18632), .ZN(n17622) );
  NOR3_X1 U12108 ( .A1(n16299), .A2(n18610), .A3(n16745), .ZN(n16302) );
  NOR2_X1 U12109 ( .A1(n11518), .A2(n10002), .ZN(n10001) );
  NOR2_X1 U12110 ( .A1(n14100), .A2(n19254), .ZN(n17776) );
  INV_X1 U12111 ( .A(n16747), .ZN(n16749) );
  NAND2_X1 U12112 ( .A1(n17894), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17900) );
  AND2_X1 U12113 ( .A1(n16941), .A2(n9692), .ZN(n17930) );
  NOR2_X1 U12114 ( .A1(n18031), .A2(n18032), .ZN(n16941) );
  AND2_X1 U12115 ( .A1(n10090), .A2(n18095), .ZN(n10089) );
  AND3_X1 U12116 ( .A1(n10089), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18190), .ZN(n18041) );
  INV_X1 U12117 ( .A(n18009), .ZN(n18105) );
  AND2_X1 U12118 ( .A1(n18190), .A2(n10090), .ZN(n18120) );
  NOR2_X1 U12119 ( .A1(n18202), .A2(n18201), .ZN(n18190) );
  INV_X1 U12120 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17274) );
  AND2_X1 U12121 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18213) );
  INV_X1 U12122 ( .A(n19256), .ZN(n16745) );
  INV_X1 U12123 ( .A(n16289), .ZN(n9994) );
  NOR2_X1 U12124 ( .A1(n18142), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9993) );
  NAND2_X1 U12125 ( .A1(n17907), .A2(n18142), .ZN(n16285) );
  NAND2_X1 U12126 ( .A1(n11673), .A2(n18142), .ZN(n9878) );
  INV_X1 U12127 ( .A(n17906), .ZN(n9877) );
  AND2_X1 U12128 ( .A1(n10008), .A2(n17949), .ZN(n11586) );
  NOR2_X1 U12129 ( .A1(n18025), .A2(n10009), .ZN(n10008) );
  INV_X1 U12130 ( .A(n18410), .ZN(n17937) );
  INV_X1 U12131 ( .A(n11584), .ZN(n17950) );
  NAND2_X1 U12132 ( .A1(n18372), .A2(n18066), .ZN(n18324) );
  NAND2_X1 U12133 ( .A1(n11582), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9881) );
  NAND2_X1 U12134 ( .A1(n18142), .A2(n18398), .ZN(n9880) );
  INV_X1 U12135 ( .A(n18048), .ZN(n18372) );
  NOR2_X1 U12136 ( .A1(n11758), .A2(n18162), .ZN(n18462) );
  NOR2_X1 U12137 ( .A1(n18163), .A2(n18502), .ZN(n18162) );
  XNOR2_X1 U12138 ( .A(n11575), .B(n9986), .ZN(n18170) );
  INV_X1 U12139 ( .A(n11576), .ZN(n9986) );
  NOR2_X1 U12140 ( .A1(n18188), .A2(n18522), .ZN(n18187) );
  NOR2_X1 U12141 ( .A1(n18200), .A2(n18199), .ZN(n18198) );
  INV_X1 U12142 ( .A(n19039), .ZN(n16915) );
  NAND2_X1 U12143 ( .A1(n18246), .A2(n18253), .ZN(n18245) );
  OR2_X1 U12144 ( .A1(n11707), .A2(n11701), .ZN(n19041) );
  INV_X1 U12145 ( .A(n16304), .ZN(n18254) );
  AND2_X1 U12146 ( .A1(n16304), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18253) );
  INV_X1 U12147 ( .A(n19051), .ZN(n19068) );
  INV_X1 U12148 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19076) );
  NAND2_X1 U12149 ( .A1(n11670), .A2(n11669), .ZN(n18627) );
  AOI211_X1 U12150 ( .C1(n17455), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n11668), .B(n11667), .ZN(n11669) );
  INV_X1 U12151 ( .A(n18636), .ZN(n18981) );
  AND2_X1 U12152 ( .A1(n13651), .A2(n13643), .ZN(n20319) );
  AND2_X1 U12153 ( .A1(n13651), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20365) );
  INV_X1 U12154 ( .A(n13683), .ZN(n13790) );
  AND2_X1 U12155 ( .A1(n13650), .A2(n13636), .ZN(n20345) );
  INV_X1 U12156 ( .A(n14765), .ZN(n14784) );
  INV_X1 U12157 ( .A(n14824), .ZN(n14848) );
  INV_X1 U12158 ( .A(n14865), .ZN(n14847) );
  OR2_X1 U12159 ( .A1(n14847), .A2(n13300), .ZN(n14868) );
  AND2_X1 U12160 ( .A1(n13212), .A2(n13211), .ZN(n20381) );
  INV_X1 U12161 ( .A(n13820), .ZN(n20421) );
  OAI21_X1 U12162 ( .B1(n14948), .B2(n15023), .A(n10723), .ZN(n14935) );
  INV_X1 U12163 ( .A(n16370), .ZN(n16361) );
  INV_X1 U12164 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16376) );
  INV_X1 U12165 ( .A(n16375), .ZN(n16351) );
  NAND2_X1 U12166 ( .A1(n10745), .A2(n9937), .ZN(n9936) );
  OR2_X1 U12167 ( .A1(n14537), .A2(n14536), .ZN(n15059) );
  NAND2_X1 U12168 ( .A1(n9982), .A2(n10748), .ZN(n14874) );
  OAI21_X1 U12169 ( .B1(n14902), .B2(n10747), .A(n16352), .ZN(n9982) );
  OR2_X1 U12170 ( .A1(n14550), .A2(n14549), .ZN(n15070) );
  INV_X1 U12171 ( .A(n9886), .ZN(n9885) );
  OR2_X1 U12172 ( .A1(n15116), .A2(n15036), .ZN(n15093) );
  NAND2_X1 U12173 ( .A1(n9938), .A2(n10728), .ZN(n14061) );
  NAND2_X1 U12174 ( .A1(n9944), .A2(n9942), .ZN(n9938) );
  NAND2_X1 U12175 ( .A1(n9968), .A2(n10707), .ZN(n13965) );
  NAND2_X1 U12176 ( .A1(n13663), .A2(n13662), .ZN(n9968) );
  NAND2_X1 U12177 ( .A1(n13285), .A2(n9816), .ZN(n13686) );
  OR2_X1 U12178 ( .A1(n13286), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U12179 ( .A1(n12931), .A2(n16249), .ZN(n20442) );
  INV_X1 U12180 ( .A(n20431), .ZN(n20439) );
  INV_X1 U12181 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20722) );
  INV_X1 U12182 ( .A(n21045), .ZN(n21043) );
  NOR2_X1 U12183 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21040) );
  OAI21_X1 U12184 ( .B1(n20599), .B2(n20583), .A(n20869), .ZN(n20601) );
  NOR2_X2 U12185 ( .A1(n20609), .A2(n20697), .ZN(n20655) );
  INV_X1 U12186 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13394) );
  INV_X1 U12187 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13398) );
  INV_X1 U12188 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13440) );
  INV_X1 U12189 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13404) );
  AOI21_X1 U12190 ( .B1(n13385), .B2(n13388), .A(n13384), .ZN(n13441) );
  OAI211_X1 U12191 ( .C1(n20685), .C2(n20811), .A(n20669), .B(n20725), .ZN(
        n20687) );
  OAI21_X1 U12192 ( .B1(n20730), .B2(n20729), .A(n20728), .ZN(n20760) );
  INV_X1 U12193 ( .A(n20802), .ZN(n20759) );
  OR2_X1 U12194 ( .A1(n20778), .A2(n20777), .ZN(n20846) );
  NOR2_X1 U12195 ( .A1(n13554), .A2(n20454), .ZN(n20853) );
  OAI21_X1 U12196 ( .B1(n20816), .B2(n20815), .A(n20814), .ZN(n20855) );
  AOI22_X1 U12197 ( .A1(n20808), .A2(n20815), .B1(n20807), .B2(n20806), .ZN(
        n20859) );
  INV_X1 U12198 ( .A(n20723), .ZN(n20899) );
  NOR2_X1 U12199 ( .A1(n20582), .A2(n13826), .ZN(n20898) );
  INV_X1 U12200 ( .A(n20820), .ZN(n20913) );
  NOR2_X1 U12201 ( .A1(n20582), .A2(n14841), .ZN(n20912) );
  INV_X1 U12202 ( .A(n20827), .ZN(n20919) );
  INV_X1 U12203 ( .A(n20739), .ZN(n20925) );
  NOR2_X1 U12204 ( .A1(n20582), .A2(n13822), .ZN(n20924) );
  INV_X1 U12205 ( .A(n20743), .ZN(n20931) );
  NOR2_X1 U12206 ( .A1(n20582), .A2(n14825), .ZN(n20930) );
  INV_X1 U12207 ( .A(n20747), .ZN(n20937) );
  INV_X1 U12208 ( .A(n20845), .ZN(n20943) );
  NOR2_X1 U12209 ( .A1(n20582), .A2(n13657), .ZN(n20942) );
  INV_X1 U12210 ( .A(n20948), .ZN(n20955) );
  INV_X1 U12211 ( .A(n20756), .ZN(n20953) );
  NAND2_X1 U12212 ( .A1(n20902), .A2(n20455), .ZN(n20959) );
  OR2_X1 U12213 ( .A1(n20961), .A2(n10532), .ZN(n20294) );
  INV_X1 U12214 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16490) );
  NAND2_X1 U12215 ( .A1(n19315), .A2(n19316), .ZN(n19314) );
  AND2_X1 U12216 ( .A1(n19282), .A2(n12815), .ZN(n19448) );
  NAND2_X1 U12217 ( .A1(n19433), .A2(n10218), .ZN(n15220) );
  INV_X1 U12218 ( .A(n19425), .ZN(n19444) );
  NAND2_X1 U12219 ( .A1(n12797), .A2(n12796), .ZN(n19443) );
  AND2_X1 U12220 ( .A1(n14509), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12221 ( .A1(n9696), .A2(n10049), .ZN(n10048) );
  INV_X1 U12222 ( .A(n19472), .ZN(n10049) );
  NOR2_X1 U12223 ( .A1(n9753), .A2(n13485), .ZN(n10052) );
  NAND2_X1 U12224 ( .A1(n10051), .A2(n9696), .ZN(n19471) );
  AND2_X1 U12225 ( .A1(n19490), .A2(n19659), .ZN(n19487) );
  AND2_X1 U12226 ( .A1(n12677), .A2(n13144), .ZN(n19490) );
  INV_X1 U12227 ( .A(n19487), .ZN(n19481) );
  NOR2_X1 U12228 ( .A1(n15282), .A2(n15281), .ZN(n15280) );
  NOR2_X1 U12229 ( .A1(n15294), .A2(n12225), .ZN(n15282) );
  AND2_X1 U12230 ( .A1(n13058), .A2(n12968), .ZN(n19497) );
  AND2_X1 U12231 ( .A1(n19551), .A2(n19538), .ZN(n19529) );
  INV_X1 U12232 ( .A(n19538), .ZN(n19547) );
  NAND2_X1 U12233 ( .A1(n15390), .A2(n13059), .ZN(n19522) );
  NOR2_X1 U12234 ( .A1(n19558), .A2(n19572), .ZN(n19557) );
  BUF_X1 U12236 ( .A(n19557), .Z(n19588) );
  OR2_X1 U12237 ( .A1(n15269), .A2(n15268), .ZN(n16540) );
  NAND2_X1 U12238 ( .A1(n14433), .A2(n14432), .ZN(n16638) );
  INV_X1 U12239 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U12240 ( .A1(n19288), .A2(n13080), .ZN(n16670) );
  CLKBUF_X1 U12241 ( .A(n16662), .Z(n19592) );
  AND2_X1 U12242 ( .A1(n16670), .A2(n20264), .ZN(n19597) );
  INV_X1 U12243 ( .A(n16661), .ZN(n19603) );
  INV_X1 U12244 ( .A(n19612), .ZN(n14031) );
  INV_X1 U12245 ( .A(n16670), .ZN(n19593) );
  AND2_X1 U12246 ( .A1(n16670), .A2(n13108), .ZN(n16661) );
  INV_X1 U12247 ( .A(n19597), .ZN(n15640) );
  INV_X1 U12248 ( .A(n16665), .ZN(n19598) );
  NAND2_X1 U12249 ( .A1(n9922), .A2(n9923), .ZN(n15465) );
  NAND2_X1 U12250 ( .A1(n14387), .A2(n9925), .ZN(n9922) );
  NAND2_X1 U12251 ( .A1(n10197), .A2(n10201), .ZN(n15588) );
  NAND2_X1 U12252 ( .A1(n10200), .A2(n10204), .ZN(n15599) );
  OR2_X1 U12253 ( .A1(n15615), .A2(n14336), .ZN(n10200) );
  NOR2_X1 U12254 ( .A1(n12529), .A2(n10055), .ZN(n15961) );
  NAND2_X1 U12255 ( .A1(n10058), .A2(n10057), .ZN(n10055) );
  XNOR2_X1 U12256 ( .A(n9813), .B(n9812), .ZN(n13787) );
  INV_X1 U12257 ( .A(n13937), .ZN(n9812) );
  INV_X1 U12258 ( .A(n19456), .ZN(n20276) );
  INV_X1 U12259 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20272) );
  INV_X1 U12260 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20262) );
  NAND2_X1 U12261 ( .A1(n11997), .A2(n12015), .ZN(n13277) );
  NOR2_X1 U12262 ( .A1(n12529), .A2(n12528), .ZN(n13766) );
  AOI221_X1 U12263 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16740), .C1(n16297), .C2(
        n16740), .A(n20098), .ZN(n20279) );
  CLKBUF_X1 U12264 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n15984) );
  AND2_X1 U12265 ( .A1(n13099), .A2(n13098), .ZN(n20265) );
  NOR2_X1 U12266 ( .A1(n19671), .A2(n19697), .ZN(n19693) );
  OR2_X1 U12267 ( .A1(n19709), .A2(n19782), .ZN(n19727) );
  OAI21_X1 U12268 ( .B1(n19738), .B2(n19737), .A(n19736), .ZN(n19756) );
  AND2_X1 U12269 ( .A1(n19666), .A2(n19961), .ZN(n19760) );
  AND2_X1 U12270 ( .A1(n19666), .A2(n16106), .ZN(n19817) );
  NOR2_X1 U12271 ( .A1(n19697), .A2(n20241), .ZN(n19868) );
  INV_X1 U12272 ( .A(n19868), .ZN(n19880) );
  OAI21_X1 U12273 ( .B1(n19839), .B2(n20153), .A(n19838), .ZN(n19877) );
  AOI22_X1 U12274 ( .A1(n16066), .A2(n16065), .B1(n16064), .B2(n19955), .ZN(
        n19897) );
  NOR2_X1 U12275 ( .A1(n16104), .A2(n20244), .ZN(n19975) );
  INV_X1 U12276 ( .A(n19975), .ZN(n19983) );
  INV_X1 U12277 ( .A(n20109), .ZN(n20023) );
  INV_X1 U12278 ( .A(n20127), .ZN(n20031) );
  OAI21_X1 U12279 ( .B1(n20059), .B2(n20058), .A(n20057), .ZN(n20086) );
  INV_X1 U12280 ( .A(n20070), .ZN(n20112) );
  INV_X1 U12281 ( .A(n20073), .ZN(n20118) );
  AND2_X1 U12282 ( .A1(n19646), .A2(n19658), .ZN(n20122) );
  AND2_X1 U12283 ( .A1(n19650), .A2(n19658), .ZN(n20128) );
  INV_X1 U12284 ( .A(n20134), .ZN(n20147) );
  INV_X1 U12285 ( .A(n20044), .ZN(n20146) );
  OR2_X1 U12286 ( .A1(n20162), .A2(n19955), .ZN(n19286) );
  AND2_X1 U12287 ( .A1(n16702), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16732) );
  INV_X1 U12288 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n20154) );
  INV_X1 U12289 ( .A(n19258), .ZN(n19272) );
  AND2_X1 U12290 ( .A1(n10088), .A2(n17271), .ZN(n16975) );
  INV_X1 U12291 ( .A(n10088), .ZN(n16985) );
  NAND2_X1 U12292 ( .A1(n16948), .A2(n16949), .ZN(n17308) );
  NOR2_X1 U12293 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17060), .ZN(n17049) );
  NOR2_X1 U12294 ( .A1(n17051), .A2(n17972), .ZN(n17050) );
  NOR2_X1 U12295 ( .A1(n17056), .A2(n9731), .ZN(n17051) );
  NOR2_X1 U12296 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17102), .ZN(n17093) );
  NOR2_X1 U12297 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17176), .ZN(n17160) );
  NOR2_X1 U12298 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17198), .ZN(n17180) );
  NOR2_X2 U12299 ( .A1(n19206), .A2(n17255), .ZN(n17286) );
  NAND4_X1 U12300 ( .A1(n18491), .A2(n19249), .A3(n19109), .A4(n19098), .ZN(
        n17318) );
  NOR2_X1 U12301 ( .A1(n17424), .A2(n17448), .ZN(n17437) );
  AOI211_X1 U12302 ( .C1(n11487), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n11646), .B(n11645), .ZN(n11647) );
  INV_X1 U12303 ( .A(n17641), .ZN(n17636) );
  NOR3_X1 U12304 ( .A1(n17800), .A2(n17802), .A3(n17696), .ZN(n17685) );
  INV_X1 U12305 ( .A(n17691), .ZN(n17696) );
  NOR2_X1 U12306 ( .A1(n17763), .A2(n17622), .ZN(n17701) );
  AND2_X1 U12307 ( .A1(n17729), .A2(n16303), .ZN(n17715) );
  NOR2_X1 U12308 ( .A1(n11540), .A2(n11539), .ZN(n17749) );
  NOR2_X1 U12309 ( .A1(n11530), .A2(n11529), .ZN(n17756) );
  INV_X1 U12310 ( .A(n11736), .ZN(n17760) );
  NOR2_X1 U12311 ( .A1(n11508), .A2(n11507), .ZN(n17765) );
  INV_X1 U12312 ( .A(n17771), .ZN(n17766) );
  INV_X1 U12313 ( .A(n17715), .ZN(n17763) );
  INV_X1 U12314 ( .A(n17764), .ZN(n17775) );
  NOR2_X1 U12315 ( .A1(n19071), .A2(n17763), .ZN(n17772) );
  CLKBUF_X1 U12316 ( .A(n17884), .Z(n17877) );
  INV_X1 U12317 ( .A(n17887), .ZN(n17878) );
  NOR2_X1 U12318 ( .A1(n16758), .A2(n18084), .ZN(n16759) );
  NAND2_X1 U12319 ( .A1(n17891), .A2(n17890), .ZN(n9876) );
  NOR2_X1 U12320 ( .A1(n18017), .A2(n17905), .ZN(n9873) );
  NAND2_X1 U12321 ( .A1(n17904), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U12322 ( .A1(n18115), .A2(n17902), .ZN(n9872) );
  INV_X1 U12323 ( .A(n17894), .ZN(n17893) );
  NAND2_X1 U12324 ( .A1(n16941), .A2(n10078), .ZN(n17960) );
  NAND2_X1 U12325 ( .A1(n16941), .A2(n9683), .ZN(n17993) );
  NAND3_X1 U12326 ( .A1(n18041), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18031) );
  NAND2_X1 U12327 ( .A1(n10089), .A2(n18190), .ZN(n18073) );
  NOR2_X1 U12328 ( .A1(n18226), .A2(n18156), .ZN(n18189) );
  AND2_X1 U12329 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18157) );
  NAND2_X1 U12330 ( .A1(n18190), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18171) );
  INV_X1 U12331 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18201) );
  NOR2_X1 U12332 ( .A1(n16918), .A2(n19256), .ZN(n18228) );
  INV_X1 U12333 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18236) );
  INV_X1 U12334 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19216) );
  OAI21_X1 U12335 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19250), .A(n16918), 
        .ZN(n18255) );
  INV_X1 U12336 ( .A(n9854), .ZN(n17922) );
  OR4_X1 U12337 ( .A1(n18025), .A2(n18325), .A3(n18262), .A4(n18018), .ZN(
        n17954) );
  NAND2_X1 U12338 ( .A1(n18079), .A2(n18372), .ZN(n18410) );
  NOR2_X1 U12339 ( .A1(n18062), .A2(n9988), .ZN(n18154) );
  AND2_X1 U12340 ( .A1(n9866), .A2(n9861), .ZN(n18184) );
  NAND2_X1 U12341 ( .A1(n18196), .A2(n18195), .ZN(n18194) );
  NAND2_X1 U12342 ( .A1(n18214), .A2(n11572), .ZN(n18196) );
  INV_X1 U12343 ( .A(n11568), .ZN(n11569) );
  CLKBUF_X1 U12344 ( .A(n18491), .Z(n18591) );
  INV_X1 U12345 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19085) );
  AOI211_X1 U12346 ( .C1(n19251), .C2(n19069), .A(n18609), .B(n14105), .ZN(
        n19236) );
  CLKBUF_X1 U12347 ( .A(n16896), .Z(n16902) );
  AOI211_X1 U12348 ( .C1(n20346), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14212), .B(
        n14211), .ZN(n14216) );
  NOR2_X1 U12349 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  NOR2_X1 U12350 ( .A1(n14770), .A2(n14736), .ZN(n9898) );
  NOR2_X1 U12351 ( .A1(n15078), .A2(n14765), .ZN(n9899) );
  OAI21_X1 U12352 ( .B1(n15044), .B2(n16349), .A(n9734), .ZN(P1_U2968) );
  AND2_X1 U12353 ( .A1(n15043), .A2(n15042), .ZN(n9791) );
  AND2_X1 U12354 ( .A1(n12673), .A2(n12672), .ZN(n12674) );
  OAI211_X1 U12355 ( .C1(n14530), .C2(n16665), .A(n9890), .B(n9888), .ZN(
        P2_U2983) );
  NAND2_X1 U12356 ( .A1(n14527), .A2(n19595), .ZN(n9888) );
  INV_X1 U12357 ( .A(n14515), .ZN(n9891) );
  NAND2_X1 U12358 ( .A1(n9954), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9952) );
  AND2_X1 U12359 ( .A1(n10063), .A2(n10060), .ZN(n14529) );
  OR2_X1 U12360 ( .A1(n16500), .A2(n16677), .ZN(n10063) );
  NAND2_X1 U12361 ( .A1(n15669), .A2(n15668), .ZN(n15670) );
  OAI21_X1 U12362 ( .B1(n14470), .B2(n15974), .A(n14469), .ZN(P2_U3018) );
  NAND2_X1 U12363 ( .A1(n9955), .A2(n15462), .ZN(n15707) );
  OR2_X1 U12364 ( .A1(n15798), .A2(n15974), .ZN(n9803) );
  INV_X1 U12365 ( .A(n15797), .ZN(n9802) );
  NAND2_X1 U12366 ( .A1(n9805), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9804) );
  OR2_X1 U12367 ( .A1(n16972), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10076) );
  AOI211_X1 U12368 ( .C1(n16968), .C2(n17278), .A(n16967), .B(n16966), .ZN(
        n16971) );
  NAND2_X1 U12369 ( .A1(n9874), .A2(n9870), .ZN(P3_U2802) );
  OR2_X1 U12370 ( .A1(n9875), .A2(n17889), .ZN(n9874) );
  NOR3_X1 U12371 ( .A1(n9873), .A2(n17901), .A3(n9871), .ZN(n9870) );
  NAND2_X1 U12372 ( .A1(n9876), .A2(n18150), .ZN(n9875) );
  OR2_X1 U12373 ( .A1(n16804), .A2(n18435), .ZN(n9985) );
  INV_X4 U12374 ( .A(n11462), .ZN(n17537) );
  NOR2_X1 U12375 ( .A1(n14697), .A2(n14761), .ZN(n9677) );
  NAND2_X1 U12376 ( .A1(n9751), .A2(n9800), .ZN(n13655) );
  INV_X1 U12377 ( .A(n10337), .ZN(n9788) );
  AND4_X1 U12378 ( .A1(n10028), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12379 ( .A1(n13150), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11970) );
  NAND2_X1 U12380 ( .A1(n10542), .A2(n10443), .ZN(n13257) );
  AND2_X1 U12381 ( .A1(n13809), .A2(n9770), .ZN(n13992) );
  NAND2_X1 U12382 ( .A1(n9677), .A2(n14752), .ZN(n14685) );
  AND2_X1 U12383 ( .A1(n10346), .A2(n9818), .ZN(n9679) );
  AND2_X1 U12384 ( .A1(n10023), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9680) );
  AND2_X1 U12385 ( .A1(n10181), .A2(n14227), .ZN(n9681) );
  AND2_X1 U12386 ( .A1(n9918), .A2(n15698), .ZN(n9682) );
  AND2_X1 U12387 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9683) );
  INV_X1 U12388 ( .A(n11572), .ZN(n9864) );
  AND2_X1 U12389 ( .A1(n10110), .A2(n10109), .ZN(n9685) );
  AND2_X1 U12390 ( .A1(n14722), .A2(n14721), .ZN(n9686) );
  AND2_X1 U12391 ( .A1(n9904), .A2(n9751), .ZN(n13809) );
  AND2_X1 U12392 ( .A1(n11938), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9687) );
  AND2_X1 U12393 ( .A1(n15498), .A2(n9738), .ZN(n9688) );
  AND3_X1 U12394 ( .A1(n14396), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14497), .ZN(n9689) );
  AND2_X1 U12395 ( .A1(n10058), .A2(n10056), .ZN(n9690) );
  AND2_X1 U12396 ( .A1(n9684), .A2(n9768), .ZN(n9691) );
  AND2_X1 U12397 ( .A1(n10078), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9692) );
  AND2_X1 U12398 ( .A1(n10742), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9693) );
  AND2_X1 U12399 ( .A1(n9685), .A2(n14018), .ZN(n9694) );
  AND2_X1 U12400 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9695) );
  INV_X2 U12401 ( .A(n10517), .ZN(n11230) );
  INV_X1 U12402 ( .A(n11384), .ZN(n11337) );
  INV_X1 U12403 ( .A(n12877), .ZN(n9836) );
  NAND2_X1 U12404 ( .A1(n10040), .A2(n10041), .ZN(n15300) );
  AND2_X1 U12405 ( .A1(n10052), .A2(n10050), .ZN(n9696) );
  AND2_X1 U12406 ( .A1(n10019), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9697) );
  INV_X1 U12407 ( .A(n13532), .ZN(n9800) );
  INV_X1 U12408 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14040) );
  NOR2_X1 U12409 ( .A1(n18155), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9698) );
  AND2_X1 U12410 ( .A1(n14440), .A2(n9895), .ZN(n9699) );
  AND2_X1 U12411 ( .A1(n9894), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9700) );
  AND2_X1 U12412 ( .A1(n9771), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9701) );
  AND2_X1 U12413 ( .A1(n9701), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9702) );
  AND2_X1 U12414 ( .A1(n9702), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9703) );
  NOR2_X4 U12415 ( .A1(n19065), .A2(n11463), .ZN(n11487) );
  OR2_X1 U12416 ( .A1(n19659), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9704) );
  NOR2_X1 U12417 ( .A1(n11461), .A2(n17302), .ZN(n11554) );
  AND2_X2 U12418 ( .A1(n11899), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12036) );
  INV_X1 U12419 ( .A(n9984), .ZN(n12829) );
  INV_X1 U12420 ( .A(n9647), .ZN(n19416) );
  NOR2_X2 U12421 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11460), .ZN(
        n11553) );
  OR2_X1 U12422 ( .A1(n14708), .A2(n10100), .ZN(n9705) );
  OR2_X1 U12423 ( .A1(n15285), .A2(n10126), .ZN(n9706) );
  OR2_X1 U12424 ( .A1(n15724), .A2(n10068), .ZN(n9707) );
  NAND2_X1 U12425 ( .A1(n9964), .A2(n9966), .ZN(n9944) );
  NAND2_X1 U12426 ( .A1(n14779), .A2(n10954), .ZN(n14722) );
  OR2_X1 U12427 ( .A1(n15222), .A2(n15221), .ZN(n9708) );
  NOR2_X1 U12428 ( .A1(n13105), .A2(n16070), .ZN(n9709) );
  AND2_X2 U12429 ( .A1(n12383), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12142) );
  OR2_X1 U12430 ( .A1(n14393), .A2(n10176), .ZN(n9710) );
  NAND2_X1 U12431 ( .A1(n11919), .A2(n11830), .ZN(n11928) );
  OR3_X1 U12432 ( .A1(n15191), .A2(n10014), .A3(n10013), .ZN(n9711) );
  NOR2_X1 U12433 ( .A1(n14660), .A2(n10156), .ZN(n9712) );
  AND2_X1 U12434 ( .A1(n14335), .A2(n10181), .ZN(n9713) );
  NOR2_X1 U12435 ( .A1(n14612), .A2(n14613), .ZN(n14600) );
  NAND2_X1 U12436 ( .A1(n15269), .A2(n14473), .ZN(n14441) );
  NOR2_X1 U12437 ( .A1(n14697), .A2(n9908), .ZN(n9715) );
  AND2_X1 U12438 ( .A1(n15781), .A2(n9702), .ZN(n9716) );
  AND2_X1 U12439 ( .A1(n15905), .A2(n9699), .ZN(n9717) );
  OR2_X1 U12440 ( .A1(n14603), .A2(n14593), .ZN(n9718) );
  NAND2_X1 U12441 ( .A1(n9789), .A2(n9939), .ZN(n15008) );
  NAND2_X1 U12442 ( .A1(n9984), .A2(n9834), .ZN(n9946) );
  NAND2_X1 U12443 ( .A1(n9781), .A2(n10439), .ZN(n10542) );
  OR2_X1 U12444 ( .A1(n10173), .A2(n10172), .ZN(n9719) );
  INV_X1 U12445 ( .A(n18195), .ZN(n9865) );
  NAND2_X1 U12446 ( .A1(n14387), .A2(n9688), .ZN(n15475) );
  AND2_X1 U12447 ( .A1(n10575), .A2(n10532), .ZN(n9720) );
  AND2_X1 U12448 ( .A1(n13717), .A2(n16001), .ZN(n14295) );
  NOR2_X1 U12449 ( .A1(n14660), .A2(n10154), .ZN(n9721) );
  OAI21_X1 U12450 ( .B1(n10543), .B2(n13264), .A(n10438), .ZN(n10439) );
  OR3_X1 U12451 ( .A1(n15724), .A2(n10071), .A3(n10073), .ZN(n9722) );
  NAND2_X1 U12452 ( .A1(n15905), .A2(n14440), .ZN(n15462) );
  AND2_X1 U12453 ( .A1(n13163), .A2(n11912), .ZN(n11945) );
  AND3_X1 U12454 ( .A1(n13881), .A2(n11830), .A3(n13155), .ZN(n9723) );
  OR3_X1 U12455 ( .A1(n14393), .A2(n14392), .A3(n10179), .ZN(n9724) );
  NAND2_X1 U12456 ( .A1(n15936), .A2(n15937), .ZN(n15633) );
  INV_X1 U12457 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12458 ( .A1(n14306), .A2(n14305), .ZN(n14423) );
  INV_X1 U12459 ( .A(n14423), .ZN(n14307) );
  NAND2_X1 U12460 ( .A1(n14722), .A2(n10159), .ZN(n10161) );
  AND2_X1 U12461 ( .A1(n10311), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n9725) );
  AND3_X1 U12462 ( .A1(n11814), .A2(n11813), .A3(n11812), .ZN(n9726) );
  INV_X1 U12463 ( .A(n9926), .ZN(n9925) );
  NAND2_X1 U12464 ( .A1(n9688), .A2(n9744), .ZN(n9926) );
  NAND2_X1 U12465 ( .A1(n10723), .A2(n16417), .ZN(n9727) );
  NAND2_X1 U12466 ( .A1(n14722), .A2(n10158), .ZN(n14697) );
  INV_X1 U12467 ( .A(n10202), .ZN(n10201) );
  OAI21_X1 U12468 ( .B1(n14345), .B2(n10203), .A(n15598), .ZN(n10202) );
  AND2_X1 U12469 ( .A1(n9883), .A2(n9882), .ZN(n9728) );
  OR2_X1 U12470 ( .A1(n11422), .A2(n9975), .ZN(n9729) );
  AND2_X1 U12471 ( .A1(n9691), .A2(n15137), .ZN(n9730) );
  NAND2_X1 U12472 ( .A1(n12889), .A2(n12888), .ZN(n12891) );
  AND4_X1 U12474 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n9732) );
  AND2_X2 U12475 ( .A1(n11818), .A2(n11817), .ZN(n13881) );
  AND2_X1 U12476 ( .A1(n12467), .A2(n11935), .ZN(n9733) );
  INV_X1 U12477 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13429) );
  INV_X1 U12478 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13572) );
  INV_X1 U12479 ( .A(n10081), .ZN(n10080) );
  NAND2_X1 U12480 ( .A1(n9683), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10081) );
  INV_X1 U12481 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11206) );
  INV_X1 U12482 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13591) );
  AND2_X1 U12483 ( .A1(n11457), .A2(n11456), .ZN(n9734) );
  AND3_X1 U12484 ( .A1(n9733), .A2(n11934), .A3(n9893), .ZN(n11957) );
  NAND2_X1 U12485 ( .A1(n10573), .A2(n10720), .ZN(n9735) );
  OR2_X1 U12486 ( .A1(n16587), .A2(n15640), .ZN(n9736) );
  AND2_X1 U12487 ( .A1(n16330), .A2(n9730), .ZN(n9737) );
  AND2_X1 U12488 ( .A1(n14386), .A2(n15507), .ZN(n9738) );
  AND2_X1 U12489 ( .A1(n9946), .A2(n9945), .ZN(n9739) );
  AND2_X1 U12490 ( .A1(n10198), .A2(n9846), .ZN(n9740) );
  AND2_X1 U12491 ( .A1(n14417), .A2(n15954), .ZN(n9741) );
  INV_X1 U12492 ( .A(n10728), .ZN(n9941) );
  OR2_X1 U12493 ( .A1(n13956), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10728) );
  NAND2_X1 U12494 ( .A1(n10723), .A2(n10740), .ZN(n9742) );
  INV_X1 U12495 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11217) );
  INV_X1 U12496 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11212) );
  NOR2_X1 U12497 ( .A1(n14660), .A2(n14661), .ZN(n9743) );
  INV_X1 U12498 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10226) );
  INV_X1 U12499 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11245) );
  INV_X1 U12500 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U12501 ( .A1(n10138), .A2(n12872), .ZN(n11775) );
  NOR2_X1 U12502 ( .A1(n13484), .A2(n13485), .ZN(n13486) );
  OR3_X1 U12503 ( .A1(n16220), .A2(n14233), .A3(n15729), .ZN(n9744) );
  AND2_X1 U12504 ( .A1(n12821), .A2(n12824), .ZN(n12822) );
  AND2_X1 U12505 ( .A1(n15864), .A2(n15852), .ZN(n12821) );
  NAND2_X1 U12506 ( .A1(n15183), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15172) );
  NAND2_X1 U12507 ( .A1(n15309), .A2(n15206), .ZN(n15205) );
  AND2_X1 U12508 ( .A1(n15926), .A2(n10066), .ZN(n9745) );
  INV_X1 U12509 ( .A(n13475), .ZN(n9826) );
  AND2_X1 U12510 ( .A1(n10075), .A2(n15811), .ZN(n9746) );
  AND2_X1 U12511 ( .A1(n10107), .A2(n10106), .ZN(n9747) );
  AND2_X1 U12512 ( .A1(n12788), .A2(n10023), .ZN(n9748) );
  NOR2_X1 U12513 ( .A1(n13532), .A2(n13541), .ZN(n13540) );
  NAND2_X1 U12514 ( .A1(n13809), .A2(n10881), .ZN(n13906) );
  NOR2_X1 U12515 ( .A1(n16592), .A2(n16591), .ZN(n15299) );
  OR2_X1 U12516 ( .A1(n14872), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9749) );
  AND2_X1 U12517 ( .A1(n15604), .A2(n9685), .ZN(n9750) );
  INV_X1 U12518 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U12519 ( .A1(n9944), .A2(n10719), .ZN(n13955) );
  AND2_X1 U12520 ( .A1(n15604), .A2(n9694), .ZN(n14017) );
  AND2_X1 U12521 ( .A1(n9905), .A2(n13656), .ZN(n9751) );
  INV_X1 U12522 ( .A(n14485), .ZN(n9927) );
  OR3_X1 U12523 ( .A1(n14708), .A2(n10104), .A3(n10102), .ZN(n9752) );
  AND2_X1 U12524 ( .A1(n11831), .A2(n11916), .ZN(n12452) );
  NOR2_X1 U12525 ( .A1(n12057), .A2(n12056), .ZN(n9753) );
  AND2_X1 U12526 ( .A1(n10742), .A2(n10746), .ZN(n9754) );
  AND2_X1 U12527 ( .A1(n9747), .A2(n10105), .ZN(n9755) );
  NAND2_X1 U12528 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NOR2_X1 U12529 ( .A1(n9698), .A2(n10006), .ZN(n9756) );
  AND2_X1 U12530 ( .A1(n10153), .A2(n14625), .ZN(n9757) );
  INV_X1 U12531 ( .A(n10132), .ZN(n15316) );
  AND2_X1 U12532 ( .A1(n14123), .A2(n14122), .ZN(n14757) );
  INV_X1 U12533 ( .A(n10137), .ZN(n12846) );
  NAND2_X1 U12534 ( .A1(n12872), .A2(n10403), .ZN(n10137) );
  AND2_X1 U12535 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9758) );
  AND2_X1 U12536 ( .A1(n11172), .A2(n11171), .ZN(n14637) );
  OR2_X1 U12537 ( .A1(n19650), .A2(n19467), .ZN(n9759) );
  AND2_X1 U12538 ( .A1(n10881), .A2(n10150), .ZN(n9760) );
  AND2_X1 U12539 ( .A1(n9746), .A2(n10074), .ZN(n9761) );
  OR2_X1 U12540 ( .A1(n14686), .A2(n10152), .ZN(n9762) );
  AND2_X1 U12541 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n9763) );
  INV_X1 U12542 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12686) );
  OR2_X1 U12543 ( .A1(n18947), .A2(n18847), .ZN(n18636) );
  NOR2_X1 U12544 ( .A1(n12528), .A2(n10059), .ZN(n10058) );
  INV_X1 U12545 ( .A(n13484), .ZN(n10051) );
  INV_X1 U12546 ( .A(n18142), .ZN(n18155) );
  NOR2_X1 U12547 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11580), .ZN(
        n18062) );
  INV_X1 U12548 ( .A(n14342), .ZN(n10182) );
  INV_X1 U12549 ( .A(n12248), .ZN(n10043) );
  NOR3_X1 U12550 ( .A1(n15191), .A2(n10017), .A3(n15431), .ZN(n14445) );
  AND2_X1 U12551 ( .A1(n18142), .A2(n9994), .ZN(n9764) );
  INV_X1 U12553 ( .A(n10093), .ZN(n14072) );
  AND2_X1 U12554 ( .A1(n10051), .A2(n10052), .ZN(n9765) );
  AND2_X1 U12555 ( .A1(n19382), .A2(n14341), .ZN(n15881) );
  INV_X1 U12556 ( .A(n19617), .ZN(n15786) );
  OR2_X1 U12557 ( .A1(n13195), .A2(n15785), .ZN(n19617) );
  AND2_X1 U12558 ( .A1(n15185), .A2(n10019), .ZN(n9766) );
  INV_X1 U12559 ( .A(n10038), .ZN(n10037) );
  NAND2_X1 U12560 ( .A1(n10041), .A2(n10039), .ZN(n10038) );
  INV_X1 U12561 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10017) );
  INV_X1 U12562 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10083) );
  INV_X1 U12563 ( .A(n14198), .ZN(n9896) );
  INV_X1 U12564 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n9975) );
  AND2_X1 U12565 ( .A1(n16941), .A2(n10080), .ZN(n9767) );
  INV_X1 U12566 ( .A(n14231), .ZN(n10184) );
  AND2_X1 U12567 ( .A1(n16393), .A2(n16398), .ZN(n9768) );
  OR2_X1 U12568 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18142), .ZN(
        n9769) );
  AND2_X1 U12569 ( .A1(n10881), .A2(n10149), .ZN(n9770) );
  INV_X1 U12570 ( .A(n13618), .ZN(n10050) );
  INV_X1 U12571 ( .A(n14458), .ZN(n9895) );
  AND2_X1 U12572 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9771) );
  INV_X1 U12573 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10082) );
  INV_X1 U12574 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10016) );
  INV_X1 U12575 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10091) );
  INV_X1 U12576 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9979) );
  INV_X1 U12577 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10020) );
  OAI222_X1 U12578 ( .A1(n14769), .A2(n14217), .B1(n14770), .B2(n14208), .C1(
        n15046), .C2(n14765), .ZN(P1_U2842) );
  NAND2_X2 U12579 ( .A1(n14770), .A2(n14198), .ZN(n14769) );
  NOR2_X1 U12580 ( .A1(n20281), .A2(n19788), .ZN(n9772) );
  INV_X1 U12581 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20281) );
  AND2_X1 U12582 ( .A1(n16028), .A2(n16735), .ZN(n20098) );
  AOI21_X1 U12583 ( .B1(n16501), .B2(n19613), .A(n10061), .ZN(n10060) );
  NAND2_X1 U12584 ( .A1(n15645), .A2(n19613), .ZN(n15653) );
  NAND2_X1 U12585 ( .A1(n15667), .A2(n19613), .ZN(n15668) );
  NOR3_X2 U12586 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19103), .A3(
        n18822), .ZN(n18794) );
  INV_X1 U12587 ( .A(n20920), .ZN(n9773) );
  INV_X1 U12588 ( .A(n9773), .ZN(n9774) );
  INV_X1 U12589 ( .A(n20944), .ZN(n9775) );
  INV_X1 U12590 ( .A(n9775), .ZN(n9776) );
  INV_X1 U12591 ( .A(n20810), .ZN(n9777) );
  INV_X1 U12592 ( .A(n9777), .ZN(n9778) );
  OAI22_X2 U12593 ( .A1(n16824), .A2(n13436), .B1(n21218), .B2(n13437), .ZN(
        n20852) );
  AOI22_X2 U12594 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19656), .ZN(n20121) );
  NOR2_X2 U12595 ( .A1(n16042), .A2(n16041), .ZN(n19656) );
  NOR3_X2 U12596 ( .A1(n19103), .A2(n19076), .A3(n18731), .ZN(n18703) );
  CLKBUF_X1 U12597 ( .A(n12994), .Z(n9779) );
  NAND2_X1 U12598 ( .A1(n12799), .A2(n12795), .ZN(n12936) );
  NOR3_X1 U12599 ( .A1(n12936), .A2(n12298), .A3(n20175), .ZN(n12994) );
  OAI22_X2 U12600 ( .A1(n16830), .A2(n13436), .B1(n13414), .B2(n13437), .ZN(
        n20836) );
  CLKBUF_X1 U12601 ( .A(n20888), .Z(n9780) );
  OAI21_X1 U12602 ( .B1(n14797), .B2(n14769), .A(n9897), .ZN(P1_U2845) );
  OAI21_X2 U12603 ( .B1(n20452), .B2(n10757), .A(n10571), .ZN(n10605) );
  NAND2_X1 U12604 ( .A1(n9824), .A2(n9781), .ZN(n9823) );
  NOR2_X2 U12605 ( .A1(n9784), .A2(n9725), .ZN(n9783) );
  NAND3_X1 U12606 ( .A1(n10240), .A2(n9787), .A3(n9785), .ZN(n9784) );
  OR2_X2 U12607 ( .A1(n13663), .A2(n9967), .ZN(n9966) );
  OAI21_X1 U12608 ( .B1(n15044), .B2(n20431), .A(n9791), .ZN(P1_U3000) );
  NAND2_X1 U12609 ( .A1(n9793), .A2(n16369), .ZN(n9835) );
  XNOR2_X1 U12610 ( .A(n9793), .B(n9792), .ZN(n16478) );
  INV_X1 U12611 ( .A(n16369), .ZN(n9792) );
  NOR2_X2 U12612 ( .A1(n9794), .A2(n10146), .ZN(n14193) );
  AND2_X2 U12613 ( .A1(n10744), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10147) );
  NAND2_X2 U12614 ( .A1(n14883), .A2(n10723), .ZN(n10744) );
  OAI211_X1 U12615 ( .C1(n12848), .C2(n13260), .A(n9796), .B(n9795), .ZN(
        n10402) );
  NAND2_X2 U12616 ( .A1(n14907), .A2(n14936), .ZN(n14921) );
  NAND2_X2 U12617 ( .A1(n14976), .A2(n14975), .ZN(n14948) );
  OR2_X2 U12618 ( .A1(n14697), .A2(n9906), .ZN(n14660) );
  NAND3_X1 U12619 ( .A1(n9800), .A2(n9903), .A3(n9902), .ZN(n10932) );
  NOR2_X2 U12620 ( .A1(n14590), .A2(n14591), .ZN(n14575) );
  OAI21_X1 U12621 ( .B1(n20453), .B2(n11031), .A(n10822), .ZN(n10823) );
  NAND2_X2 U12622 ( .A1(n10596), .A2(n10595), .ZN(n20453) );
  INV_X1 U12623 ( .A(n10594), .ZN(n10541) );
  NAND3_X1 U12624 ( .A1(n9804), .A2(n9803), .A3(n9802), .ZN(P2_U3029) );
  INV_X1 U12625 ( .A(n12465), .ZN(n9811) );
  OAI21_X2 U12626 ( .B1(n9813), .B2(n14497), .A(n14043), .ZN(n13934) );
  XNOR2_X2 U12627 ( .A(n9840), .B(n9839), .ZN(n9813) );
  INV_X2 U12628 ( .A(n11830), .ZN(n12485) );
  AND2_X2 U12629 ( .A1(n15787), .A2(n15791), .ZN(n15781) );
  NAND2_X2 U12630 ( .A1(n9814), .A2(n9959), .ZN(n15787) );
  NAND4_X1 U12631 ( .A1(n14433), .A2(n14432), .A3(n9961), .A4(n15788), .ZN(
        n9814) );
  NAND2_X2 U12632 ( .A1(n14431), .A2(n16675), .ZN(n14432) );
  NAND2_X2 U12633 ( .A1(n14430), .A2(n15630), .ZN(n14433) );
  NAND2_X2 U12634 ( .A1(n15945), .A2(n14426), .ZN(n15632) );
  NAND2_X1 U12635 ( .A1(n9741), .A2(n15958), .ZN(n9815) );
  NAND2_X2 U12636 ( .A1(n14921), .A2(n16352), .ZN(n14909) );
  NAND2_X2 U12637 ( .A1(n14164), .A2(n9817), .ZN(n14163) );
  NAND2_X4 U12638 ( .A1(n10722), .A2(n10721), .ZN(n10723) );
  NAND3_X1 U12639 ( .A1(n13475), .A2(n10531), .A3(n10441), .ZN(n9822) );
  NAND2_X1 U12640 ( .A1(n10596), .A2(n13494), .ZN(n9827) );
  INV_X1 U12641 ( .A(n10567), .ZN(n13494) );
  INV_X1 U12642 ( .A(n10596), .ZN(n9828) );
  NAND2_X1 U12643 ( .A1(n10812), .A2(n9720), .ZN(n9830) );
  INV_X2 U12644 ( .A(n10350), .ZN(n11365) );
  NAND2_X1 U12645 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n9833) );
  NAND3_X1 U12646 ( .A1(n9650), .A2(n9836), .A3(n10405), .ZN(n11772) );
  NAND4_X1 U12647 ( .A1(n9650), .A2(n10405), .A3(n9836), .A4(n13213), .ZN(
        n12928) );
  NOR2_X1 U12648 ( .A1(n10404), .A2(n12877), .ZN(n10802) );
  NAND2_X1 U12649 ( .A1(n11823), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9838) );
  NAND2_X1 U12650 ( .A1(n11829), .A2(n12026), .ZN(n9837) );
  NAND2_X1 U12651 ( .A1(n13934), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13935) );
  NAND2_X1 U12652 ( .A1(n13754), .A2(n13753), .ZN(n9839) );
  NAND2_X1 U12653 ( .A1(n13941), .A2(n13940), .ZN(n9840) );
  AOI21_X2 U12654 ( .B1(n14387), .B2(n9850), .A(n9847), .ZN(n15450) );
  OR2_X2 U12655 ( .A1(n17923), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9854) );
  NAND2_X1 U12656 ( .A1(n9866), .A2(n9857), .ZN(n18182) );
  NAND2_X1 U12657 ( .A1(n18183), .A2(n9859), .ZN(n9858) );
  NAND2_X1 U12658 ( .A1(n9863), .A2(n9865), .ZN(n9859) );
  OAI21_X1 U12659 ( .B1(n18214), .B2(n9865), .A(n9863), .ZN(n9861) );
  NAND3_X1 U12660 ( .A1(n11562), .A2(n11564), .A3(n11563), .ZN(n16304) );
  INV_X2 U12661 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9868) );
  NOR2_X2 U12662 ( .A1(n17891), .A2(n17890), .ZN(n17889) );
  NAND2_X2 U12663 ( .A1(n18035), .A2(n18155), .ZN(n17997) );
  NAND2_X1 U12664 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9883) );
  AND4_X2 U12665 ( .A1(n10567), .A2(n10540), .A3(n10541), .A4(n10641), .ZN(
        n10662) );
  NAND2_X1 U12666 ( .A1(n9892), .A2(n11906), .ZN(n9893) );
  NAND3_X1 U12667 ( .A1(n11844), .A2(n9636), .A3(n14328), .ZN(n9892) );
  INV_X2 U12668 ( .A(n10337), .ZN(n10380) );
  AOI21_X2 U12669 ( .B1(n10421), .B2(n10295), .A(n9896), .ZN(n10424) );
  NAND2_X2 U12670 ( .A1(n9900), .A2(n10417), .ZN(n10465) );
  NAND3_X2 U12671 ( .A1(n9901), .A2(n10412), .A3(n10414), .ZN(n10408) );
  OR2_X2 U12672 ( .A1(n12928), .A2(n12837), .ZN(n10414) );
  INV_X1 U12673 ( .A(n10402), .ZN(n9901) );
  INV_X1 U12674 ( .A(n13541), .ZN(n9905) );
  NOR2_X1 U12675 ( .A1(n13810), .A2(n13532), .ZN(n9904) );
  NAND2_X1 U12676 ( .A1(n14575), .A2(n14577), .ZN(n14561) );
  NAND3_X1 U12677 ( .A1(n13717), .A2(n13929), .A3(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n9928) );
  NAND3_X1 U12678 ( .A1(n13718), .A2(n13929), .A3(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9929) );
  NAND3_X1 U12679 ( .A1(n13733), .A2(n13734), .A3(n9930), .ZN(n9931) );
  AND2_X1 U12680 ( .A1(n13717), .A2(n13929), .ZN(n19953) );
  NOR2_X1 U12681 ( .A1(n13739), .A2(n9931), .ZN(n13750) );
  AND2_X2 U12682 ( .A1(n10197), .A2(n10196), .ZN(n15560) );
  NAND3_X1 U12683 ( .A1(n13941), .A2(n13754), .A3(n9933), .ZN(n13942) );
  NAND4_X1 U12684 ( .A1(n13730), .A2(n13731), .A3(n13729), .A4(n13728), .ZN(
        n13941) );
  AND2_X4 U12685 ( .A1(n10241), .A2(n13461), .ZN(n11359) );
  INV_X2 U12686 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13461) );
  AND2_X2 U12687 ( .A1(n9935), .A2(n10744), .ZN(n14902) );
  NOR2_X1 U12688 ( .A1(n14902), .A2(n9936), .ZN(n14194) );
  OAI21_X2 U12689 ( .B1(n13238), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10533), 
        .ZN(n10803) );
  NAND2_X1 U12690 ( .A1(n9983), .A2(n9984), .ZN(n14980) );
  AOI21_X1 U12691 ( .B1(n9948), .B2(n12681), .A(n12680), .ZN(n13894) );
  NAND2_X2 U12692 ( .A1(n10210), .A2(n11974), .ZN(n9948) );
  NAND2_X1 U12693 ( .A1(n11926), .A2(n16039), .ZN(n12794) );
  NAND2_X1 U12694 ( .A1(n13150), .A2(n9763), .ZN(n9949) );
  NAND3_X1 U12695 ( .A1(n9950), .A2(n9949), .A3(n11939), .ZN(n11943) );
  OR2_X1 U12696 ( .A1(n15466), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9955) );
  NAND2_X1 U12697 ( .A1(n9953), .A2(n9951), .ZN(P2_U2990) );
  NAND2_X1 U12698 ( .A1(n15466), .A2(n9954), .ZN(n9953) );
  NAND3_X1 U12699 ( .A1(n14433), .A2(n14432), .A3(n9961), .ZN(n16640) );
  NAND2_X2 U12700 ( .A1(n16640), .A2(n14436), .ZN(n15905) );
  NAND2_X1 U12701 ( .A1(n15781), .A2(n9703), .ZN(n15487) );
  AND2_X1 U12702 ( .A1(n15781), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15545) );
  NAND2_X1 U12703 ( .A1(n13531), .A2(n13530), .ZN(n9962) );
  NAND2_X1 U12704 ( .A1(n10602), .A2(n10601), .ZN(n9963) );
  NAND2_X1 U12705 ( .A1(n13310), .A2(n9963), .ZN(n10603) );
  XNOR2_X1 U12706 ( .A(n13310), .B(n9963), .ZN(n13336) );
  OAI21_X1 U12707 ( .B1(n13662), .B2(n9967), .A(n13966), .ZN(n9965) );
  INV_X2 U12708 ( .A(n10551), .ZN(n9976) );
  NAND3_X1 U12709 ( .A1(n14204), .A2(n12887), .A3(n9978), .ZN(n12888) );
  NAND2_X1 U12710 ( .A1(n14902), .A2(n16352), .ZN(n9981) );
  NAND3_X1 U12711 ( .A1(n9981), .A2(n10748), .A3(n9980), .ZN(n10750) );
  AOI21_X1 U12712 ( .B1(n10747), .B2(n16352), .A(n9749), .ZN(n9980) );
  NAND3_X1 U12713 ( .A1(n16802), .A2(n16803), .A3(n9985), .ZN(P3_U2831) );
  NAND3_X1 U12714 ( .A1(n19229), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11460) );
  AND2_X2 U12715 ( .A1(n9987), .A2(n9988), .ZN(n18061) );
  INV_X1 U12716 ( .A(n18062), .ZN(n9987) );
  INV_X1 U12717 ( .A(n16284), .ZN(n9992) );
  NAND2_X1 U12718 ( .A1(n17907), .A2(n9764), .ZN(n16754) );
  NAND3_X1 U12719 ( .A1(n16754), .A2(n9990), .A3(n9989), .ZN(n9996) );
  NAND2_X1 U12720 ( .A1(n16284), .A2(n18155), .ZN(n9989) );
  NAND2_X1 U12721 ( .A1(n9992), .A2(n9993), .ZN(n16752) );
  NAND2_X1 U12722 ( .A1(n16752), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10000) );
  NAND2_X1 U12723 ( .A1(n9996), .A2(n16755), .ZN(n9995) );
  NAND3_X1 U12724 ( .A1(n10000), .A2(n9998), .A3(n9769), .ZN(n9997) );
  NAND2_X1 U12725 ( .A1(n16754), .A2(n19218), .ZN(n9999) );
  NAND2_X1 U12726 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10027) );
  NAND3_X1 U12727 ( .A1(n10028), .A2(n10026), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12784) );
  NOR2_X1 U12728 ( .A1(n12686), .A2(n10027), .ZN(n10026) );
  INV_X1 U12729 ( .A(n12781), .ZN(n10028) );
  NAND3_X1 U12730 ( .A1(n10028), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12782) );
  NAND3_X1 U12731 ( .A1(n13164), .A2(n13178), .A3(n10031), .ZN(n10030) );
  NAND4_X1 U12732 ( .A1(n10030), .A2(n10029), .A3(n13163), .A4(n11912), .ZN(
        n11913) );
  NAND3_X1 U12733 ( .A1(n10031), .A2(n13178), .A3(n10032), .ZN(n10029) );
  AND2_X2 U12734 ( .A1(n13029), .A2(n9670), .ZN(n10033) );
  INV_X1 U12735 ( .A(n16592), .ZN(n10040) );
  NAND2_X1 U12736 ( .A1(n10038), .A2(n10043), .ZN(n10034) );
  NAND2_X1 U12737 ( .A1(n10037), .A2(n12248), .ZN(n10036) );
  INV_X1 U12738 ( .A(n10047), .ZN(n12276) );
  NAND2_X1 U12739 ( .A1(n13881), .A2(n12485), .ZN(n11916) );
  NAND3_X1 U12740 ( .A1(n11997), .A2(n12015), .A3(n12014), .ZN(n13279) );
  INV_X1 U12741 ( .A(n12529), .ZN(n10054) );
  NAND2_X1 U12742 ( .A1(n10054), .A2(n9690), .ZN(n15959) );
  NAND3_X1 U12743 ( .A1(n16971), .A2(n16970), .A3(n10076), .ZN(P3_U2641) );
  XNOR2_X2 U12744 ( .A(n16762), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17271) );
  NAND2_X1 U12745 ( .A1(n10085), .A2(n10086), .ZN(n16974) );
  NAND2_X1 U12746 ( .A1(n10085), .A2(n10084), .ZN(n16963) );
  OR2_X1 U12747 ( .A1(n16986), .A2(n17902), .ZN(n10088) );
  OR2_X1 U12748 ( .A1(n11772), .A2(n14158), .ZN(n10407) );
  NOR2_X2 U12749 ( .A1(n14781), .A2(n14782), .ZN(n14780) );
  INV_X1 U12750 ( .A(n14757), .ZN(n10104) );
  NAND2_X1 U12751 ( .A1(n10114), .A2(n10112), .ZN(n11914) );
  NAND2_X1 U12752 ( .A1(n10113), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10112) );
  NAND4_X1 U12753 ( .A1(n11861), .A2(n11859), .A3(n11858), .A4(n11860), .ZN(
        n10113) );
  NAND2_X1 U12754 ( .A1(n10115), .A2(n12026), .ZN(n10114) );
  NAND4_X1 U12755 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11865), .ZN(
        n10115) );
  NAND2_X1 U12756 ( .A1(n10118), .A2(n10116), .ZN(n15892) );
  AND2_X2 U12757 ( .A1(n11944), .A2(n10123), .ZN(n11999) );
  NAND2_X1 U12758 ( .A1(n11998), .A2(n10123), .ZN(n11968) );
  NAND2_X1 U12759 ( .A1(n11941), .A2(n11940), .ZN(n10123) );
  NAND2_X1 U12760 ( .A1(n10133), .A2(n10411), .ZN(n10416) );
  INV_X1 U12761 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U12762 ( .A1(n10140), .A2(n10141), .ZN(n10462) );
  NAND3_X1 U12763 ( .A1(n10542), .A2(n10136), .A3(n10443), .ZN(n10140) );
  NAND2_X1 U12764 ( .A1(n10148), .A2(n10693), .ZN(n10694) );
  NAND2_X1 U12765 ( .A1(n10663), .A2(n10148), .ZN(n10844) );
  NAND2_X1 U12766 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  INV_X1 U12767 ( .A(n10161), .ZN(n14696) );
  NOR2_X1 U12768 ( .A1(n14561), .A2(n10164), .ZN(n14531) );
  INV_X1 U12769 ( .A(n14561), .ZN(n10166) );
  NOR2_X4 U12770 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15978) );
  AOI21_X1 U12771 ( .B1(n12150), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n10169), .ZN(n12479) );
  AND2_X1 U12772 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10170) );
  INV_X1 U12773 ( .A(n10171), .ZN(n10174) );
  NOR2_X1 U12774 ( .A1(n14393), .A2(n14392), .ZN(n14397) );
  NAND2_X1 U12775 ( .A1(n14335), .A2(n10180), .ZN(n14355) );
  NAND2_X1 U12776 ( .A1(n14502), .A2(n14231), .ZN(n14414) );
  NAND2_X1 U12777 ( .A1(n14502), .A2(n10183), .ZN(n14493) );
  NAND2_X1 U12778 ( .A1(n14484), .A2(n10194), .ZN(n10192) );
  INV_X1 U12779 ( .A(n14488), .ZN(n10194) );
  AND2_X1 U12780 ( .A1(n14485), .A2(n14486), .ZN(n10195) );
  INV_X1 U12781 ( .A(n15881), .ZN(n10207) );
  NAND3_X1 U12782 ( .A1(n14427), .A2(n14233), .A3(n10209), .ZN(n14312) );
  NAND2_X1 U12783 ( .A1(n14308), .A2(n14423), .ZN(n10209) );
  INV_X1 U12784 ( .A(n14308), .ZN(n10208) );
  AND2_X1 U12785 ( .A1(n14427), .A2(n10209), .ZN(n14417) );
  NAND2_X1 U12786 ( .A1(n11969), .A2(n11974), .ZN(n11991) );
  NAND3_X1 U12787 ( .A1(n13412), .A2(n13213), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10789) );
  NAND2_X1 U12788 ( .A1(n14546), .A2(n14532), .ZN(n14533) );
  XNOR2_X1 U12789 ( .A(n14207), .B(n14206), .ZN(n15046) );
  INV_X1 U12790 ( .A(n13551), .ZN(n13552) );
  NAND2_X1 U12791 ( .A1(n10825), .A2(n10824), .ZN(n13328) );
  OR2_X1 U12792 ( .A1(n20453), .A2(n13494), .ZN(n13554) );
  NAND2_X1 U12793 ( .A1(n13498), .A2(n20453), .ZN(n20778) );
  OR2_X1 U12794 ( .A1(n20453), .A2(n10757), .ZN(n10602) );
  NAND2_X1 U12795 ( .A1(n14193), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10749) );
  OR2_X1 U12796 ( .A1(n11406), .A2(n10260), .ZN(n10261) );
  NAND2_X1 U12797 ( .A1(n12856), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10550) );
  INV_X1 U12798 ( .A(n10495), .ZN(n10620) );
  OR2_X1 U12799 ( .A1(n20412), .A2(n13635), .ZN(n13820) );
  OAI21_X1 U12800 ( .B1(n10551), .B2(n11407), .A(n10296), .ZN(n10297) );
  NOR2_X1 U12801 ( .A1(n13156), .A2(n13081), .ZN(n11937) );
  NAND3_X1 U12802 ( .A1(n11936), .A2(n12298), .A3(n11908), .ZN(n13152) );
  NAND2_X1 U12803 ( .A1(n14017), .A2(n15232), .ZN(n15317) );
  INV_X1 U12804 ( .A(n13873), .ZN(n13874) );
  NAND2_X1 U12805 ( .A1(n15480), .A2(n15291), .ZN(n15293) );
  OR2_X1 U12806 ( .A1(n15615), .A2(n15614), .ZN(n15914) );
  NAND2_X1 U12807 ( .A1(n13524), .A2(n13525), .ZN(n13526) );
  AOI22_X1 U12808 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U12809 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11359), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10286) );
  OR2_X1 U12810 ( .A1(n13299), .A2(n13412), .ZN(n10319) );
  INV_X1 U12811 ( .A(n10297), .ZN(n10298) );
  XNOR2_X1 U12812 ( .A(n10462), .B(n10461), .ZN(n10594) );
  AND2_X4 U12813 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10242), .ZN(
        n10338) );
  NAND2_X1 U12814 ( .A1(n9676), .A2(n19454), .ZN(n13720) );
  NOR2_X1 U12815 ( .A1(n9676), .A2(n14053), .ZN(n13710) );
  AND2_X1 U12816 ( .A1(n9676), .A2(n13701), .ZN(n13718) );
  NOR2_X1 U12817 ( .A1(n20864), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10212) );
  OR2_X1 U12818 ( .A1(n15380), .A2(n15379), .ZN(n10213) );
  NAND2_X1 U12819 ( .A1(n13595), .A2(n13013), .ZN(n21059) );
  INV_X1 U12820 ( .A(n10818), .ZN(n13628) );
  INV_X1 U12821 ( .A(n13628), .ZN(n11170) );
  AND2_X1 U12822 ( .A1(n12666), .A2(n13881), .ZN(n10214) );
  AND2_X1 U12823 ( .A1(n11916), .A2(n11915), .ZN(n10216) );
  OR2_X1 U12824 ( .A1(n19339), .A2(n15543), .ZN(n10218) );
  INV_X1 U12825 ( .A(n18084), .ZN(n18165) );
  NOR2_X1 U12826 ( .A1(n14198), .A2(n20769), .ZN(n10857) );
  INV_X1 U12827 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12791) );
  INV_X1 U12828 ( .A(n14672), .ZN(n11100) );
  INV_X1 U12829 ( .A(n11031), .ZN(n11010) );
  OR2_X1 U12830 ( .A1(n15648), .A2(n15647), .ZN(n10219) );
  NAND2_X1 U12831 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10221) );
  NOR2_X1 U12832 ( .A1(n19065), .A2(n11461), .ZN(n11638) );
  AND2_X1 U12833 ( .A1(n11950), .A2(n11949), .ZN(n10222) );
  NAND2_X1 U12834 ( .A1(n13704), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14238) );
  AOI22_X1 U12835 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n10295), .B1(n13635), 
        .B2(n10784), .ZN(n10775) );
  INV_X1 U12836 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U12837 ( .A1(n14243), .A2(n14242), .ZN(n14244) );
  INV_X1 U12838 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11173) );
  INV_X1 U12839 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11330) );
  INV_X1 U12840 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11131) );
  INV_X1 U12841 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U12842 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11812) );
  OR2_X1 U12843 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20722), .ZN(
        n10753) );
  INV_X1 U12844 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11426) );
  INV_X1 U12845 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11353) );
  OR2_X1 U12846 ( .A1(n9657), .A2(n10354), .ZN(n10355) );
  AOI22_X1 U12847 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14234), .B1(
        n14235), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13734) );
  INV_X1 U12848 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13709) );
  NAND2_X1 U12849 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10265) );
  INV_X1 U12850 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11151) );
  INV_X1 U12851 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U12852 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9661), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U12853 ( .A1(n13634), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10549) );
  INV_X1 U12854 ( .A(n10767), .ZN(n10764) );
  INV_X1 U12855 ( .A(n13909), .ZN(n10881) );
  INV_X1 U12856 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11257) );
  INV_X1 U12857 ( .A(n11265), .ZN(n11266) );
  INV_X1 U12858 ( .A(n10504), .ZN(n10720) );
  NAND2_X1 U12859 ( .A1(n10530), .A2(n10529), .ZN(n13548) );
  INV_X1 U12860 ( .A(n12425), .ZN(n12400) );
  NOR2_X1 U12861 ( .A1(n13081), .A2(n16735), .ZN(n11938) );
  INV_X1 U12862 ( .A(n14279), .ZN(n14265) );
  AOI22_X1 U12863 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11881) );
  AOI21_X1 U12864 ( .B1(n20862), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10759), .ZN(n10758) );
  NAND2_X1 U12865 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10312) );
  INV_X1 U12866 ( .A(n14707), .ZN(n10993) );
  NOR2_X1 U12867 ( .A1(n11373), .A2(n14896), .ZN(n11374) );
  AND2_X1 U12868 ( .A1(n11266), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11267) );
  OR2_X1 U12869 ( .A1(n10932), .A2(n10931), .ZN(n10954) );
  NOR2_X1 U12870 ( .A1(n10460), .A2(n10459), .ZN(n10598) );
  AND2_X1 U12871 ( .A1(n16070), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U12872 ( .A1(n13702), .A2(n13086), .ZN(n11994) );
  INV_X1 U12873 ( .A(n12378), .ZN(n12384) );
  NAND2_X1 U12874 ( .A1(n15177), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15176) );
  INV_X1 U12875 ( .A(n12809), .ZN(n13755) );
  AND2_X1 U12876 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11734), .ZN(
        n11746) );
  INV_X1 U12877 ( .A(n11702), .ZN(n11713) );
  OR4_X1 U12878 ( .A1(n13792), .A2(n20984), .A3(n13373), .A4(n13791), .ZN(
        n20351) );
  AND2_X1 U12879 ( .A1(n14120), .A2(n14119), .ZN(n14699) );
  AND2_X1 U12880 ( .A1(n12910), .A2(n12909), .ZN(n13814) );
  INV_X1 U12881 ( .A(n10992), .ZN(n11192) );
  AND2_X1 U12882 ( .A1(n11441), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11451) );
  OR2_X1 U12883 ( .A1(n11321), .A2(n14580), .ZN(n11373) );
  NOR2_X1 U12884 ( .A1(n11143), .A2(n11142), .ZN(n11144) );
  INV_X1 U12885 ( .A(n11438), .ZN(n11402) );
  AND2_X1 U12886 ( .A1(n10858), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10882) );
  AND2_X1 U12887 ( .A1(n14131), .A2(n14130), .ZN(n14675) );
  AND2_X1 U12888 ( .A1(n12920), .A2(n12919), .ZN(n14071) );
  OR2_X1 U12889 ( .A1(n10856), .A2(n10757), .ZN(n10705) );
  NAND2_X1 U12890 ( .A1(n10548), .A2(n10547), .ZN(n13475) );
  AND3_X1 U12891 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n10532), .A3(n13387), 
        .ZN(n13432) );
  OR2_X1 U12892 ( .A1(n12534), .A2(n12533), .ZN(n13765) );
  OR2_X1 U12893 ( .A1(n12033), .A2(n12032), .ZN(n19479) );
  AND2_X1 U12894 ( .A1(n16735), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13086) );
  AND2_X1 U12895 ( .A1(n12248), .A2(n12247), .ZN(n12249) );
  NOR2_X1 U12896 ( .A1(n15659), .A2(n15663), .ZN(n15665) );
  AND2_X1 U12897 ( .A1(n14317), .A2(n15634), .ZN(n14318) );
  OAI21_X1 U12898 ( .B1(n13934), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13933), .ZN(n13936) );
  AND4_X1 U12899 ( .A1(n12573), .A2(n12572), .A3(n12571), .A4(n12570), .ZN(
        n12594) );
  OR2_X1 U12900 ( .A1(n13181), .A2(n16701), .ZN(n15782) );
  NAND2_X1 U12901 ( .A1(n16946), .A2(n16745), .ZN(n11717) );
  OR2_X1 U12902 ( .A1(n18366), .A2(n17905), .ZN(n11765) );
  INV_X1 U12903 ( .A(n19047), .ZN(n19070) );
  OR2_X1 U12904 ( .A1(n14572), .A2(n14184), .ZN(n14543) );
  INV_X1 U12905 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14713) );
  INV_X1 U12906 ( .A(n20365), .ZN(n20321) );
  INV_X1 U12907 ( .A(n21059), .ZN(n13644) );
  OR3_X1 U12908 ( .A1(n21059), .A2(n13631), .A3(n13630), .ZN(n13651) );
  NAND2_X1 U12909 ( .A1(n11195), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11265) );
  INV_X1 U12910 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11033) );
  INV_X1 U12911 ( .A(n10857), .ZN(n10992) );
  AND4_X1 U12912 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n13909) );
  INV_X1 U12913 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10751) );
  INV_X1 U12914 ( .A(n15154), .ZN(n16447) );
  NOR2_X1 U12915 ( .A1(n16447), .A2(n13292), .ZN(n15022) );
  NAND2_X1 U12916 ( .A1(n16254), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U12917 ( .A1(n20452), .A2(n20453), .ZN(n20555) );
  INV_X1 U12918 ( .A(n20631), .ZN(n20604) );
  OR2_X1 U12919 ( .A1(n20778), .A2(n20697), .ZN(n20757) );
  OR2_X1 U12920 ( .A1(n13553), .A2(n13551), .ZN(n20697) );
  AOI21_X1 U12921 ( .B1(n20690), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20582), 
        .ZN(n20906) );
  NAND2_X1 U12922 ( .A1(n13553), .A2(n13552), .ZN(n20777) );
  NAND2_X1 U12923 ( .A1(n13132), .A2(n12447), .ZN(n16702) );
  AND3_X1 U12924 ( .A1(n12539), .A2(n12538), .A3(n12537), .ZN(n13901) );
  NAND2_X1 U12925 ( .A1(n11996), .A2(n11995), .ZN(n12015) );
  NAND2_X1 U12926 ( .A1(n15272), .A2(n12277), .ZN(n12300) );
  OR2_X1 U12927 ( .A1(n13985), .A2(n13984), .ZN(n14021) );
  AND3_X1 U12928 ( .A1(n12599), .A2(n12598), .A3(n12597), .ZN(n13869) );
  INV_X1 U12929 ( .A(n19495), .ZN(n15390) );
  OAI21_X1 U12930 ( .B1(n12665), .B2(n12664), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12968) );
  NAND2_X1 U12931 ( .A1(n13894), .A2(n13893), .ZN(n13895) );
  NOR2_X1 U12932 ( .A1(n15651), .A2(n15650), .ZN(n15652) );
  NOR3_X1 U12933 ( .A1(n15666), .A2(n15665), .A3(n15664), .ZN(n15669) );
  OR2_X1 U12934 ( .A1(n16526), .A2(n14233), .ZN(n14485) );
  OR2_X1 U12935 ( .A1(n14376), .A2(n15748), .ZN(n15507) );
  OR2_X1 U12936 ( .A1(n14383), .A2(n14382), .ZN(n15584) );
  OR3_X1 U12937 ( .A1(n19362), .A2(n14233), .A3(n15858), .ZN(n15597) );
  NOR2_X1 U12938 ( .A1(n15914), .A2(n15915), .ZN(n15913) );
  AND2_X1 U12939 ( .A1(n13774), .A2(n13773), .ZN(n14456) );
  INV_X1 U12940 ( .A(n19613), .ZN(n15927) );
  OR2_X1 U12941 ( .A1(n14282), .A2(n16024), .ZN(n16036) );
  INV_X1 U12942 ( .A(n19839), .ZN(n19873) );
  INV_X1 U12943 ( .A(n20265), .ZN(n20267) );
  NOR2_X1 U12944 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17128), .ZN(n17113) );
  NOR2_X1 U12945 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17218), .ZN(n17210) );
  NOR2_X1 U12946 ( .A1(n16744), .A2(n14087), .ZN(n14102) );
  NOR2_X1 U12947 ( .A1(n17791), .A2(n17666), .ZN(n17665) );
  NAND2_X1 U12948 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18189), .ZN(n18044) );
  AND2_X1 U12949 ( .A1(n11765), .A2(n17897), .ZN(n11766) );
  NAND2_X1 U12950 ( .A1(n11543), .A2(n11544), .ZN(n11542) );
  INV_X1 U12951 ( .A(n18324), .ZN(n18402) );
  INV_X1 U12952 ( .A(n18462), .ZN(n18079) );
  NOR2_X1 U12953 ( .A1(n19051), .A2(n18593), .ZN(n18475) );
  OR2_X1 U12954 ( .A1(n19230), .A2(n19110), .ZN(n18608) );
  NAND2_X1 U12955 ( .A1(n19048), .A2(n19046), .ZN(n14097) );
  INV_X1 U12956 ( .A(n11711), .ZN(n18616) );
  NAND2_X1 U12957 ( .A1(n19256), .A2(n18312), .ZN(n18304) );
  NOR2_X1 U12958 ( .A1(n15046), .A2(n20377), .ZN(n14211) );
  OR2_X1 U12959 ( .A1(n14620), .A2(n14176), .ZN(n14588) );
  NOR2_X1 U12960 ( .A1(n14688), .A2(n21010), .ZN(n14681) );
  NOR2_X1 U12961 ( .A1(n16329), .A2(n14180), .ZN(n14715) );
  AND2_X1 U12962 ( .A1(n13651), .A2(n13632), .ZN(n20327) );
  INV_X1 U12963 ( .A(n20363), .ZN(n20346) );
  OR2_X1 U12964 ( .A1(n13683), .A2(n13791), .ZN(n20352) );
  INV_X1 U12965 ( .A(n14770), .ZN(n14783) );
  INV_X1 U12966 ( .A(n14840), .ZN(n14850) );
  NAND2_X1 U12967 ( .A1(n13253), .A2(n20300), .ZN(n11788) );
  INV_X1 U12968 ( .A(n13627), .ZN(n13846) );
  NAND2_X1 U12969 ( .A1(n11035), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11071) );
  AND2_X1 U12970 ( .A1(n16264), .A2(n20300), .ZN(n20302) );
  OR2_X1 U12971 ( .A1(n15098), .A2(n15039), .ZN(n15080) );
  OR2_X1 U12972 ( .A1(n15109), .A2(n15037), .ZN(n15098) );
  OAI21_X1 U12973 ( .B1(n15150), .B2(n20442), .A(n15105), .ZN(n16418) );
  INV_X1 U12974 ( .A(n20438), .ZN(n16466) );
  OR2_X1 U12975 ( .A1(n15154), .A2(n15151), .ZN(n16416) );
  AND2_X1 U12976 ( .A1(n12931), .A2(n16232), .ZN(n20447) );
  OAI22_X1 U12977 ( .A1(n20466), .A2(n20465), .B1(n20578), .B2(n20665), .ZN(
        n20489) );
  INV_X1 U12978 ( .A(n20555), .ZN(n20499) );
  AND2_X1 U12979 ( .A1(n20499), .A2(n20498), .ZN(n20542) );
  NOR2_X2 U12980 ( .A1(n20555), .A2(n20860), .ZN(n20571) );
  NOR2_X2 U12981 ( .A1(n20555), .A2(n20777), .ZN(n20600) );
  INV_X1 U12982 ( .A(n20609), .ZN(n20576) );
  OAI21_X1 U12983 ( .B1(n20639), .B2(n20638), .A(n20637), .ZN(n20657) );
  INV_X1 U12984 ( .A(n20454), .ZN(n20661) );
  INV_X1 U12985 ( .A(n20757), .ZN(n20752) );
  NAND2_X1 U12986 ( .A1(n13553), .A2(n13551), .ZN(n20860) );
  INV_X1 U12987 ( .A(n20846), .ZN(n20854) );
  INV_X1 U12988 ( .A(n20907), .ZN(n20901) );
  OAI211_X1 U12989 ( .C1(n20871), .C2(n20889), .A(n20870), .B(n20869), .ZN(
        n20891) );
  NOR2_X1 U12990 ( .A1(n20582), .A2(n14835), .ZN(n20918) );
  NOR2_X1 U12991 ( .A1(n20582), .A2(n14820), .ZN(n20936) );
  NOR2_X1 U12992 ( .A1(n20582), .A2(n13812), .ZN(n20951) );
  INV_X1 U12993 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20971) );
  NAND2_X1 U12994 ( .A1(n16520), .A2(n16521), .ZN(n16519) );
  NAND2_X1 U12995 ( .A1(n16532), .A2(n16533), .ZN(n16531) );
  NAND2_X1 U12996 ( .A1(n16555), .A2(n16556), .ZN(n16554) );
  NAND2_X1 U12997 ( .A1(n16581), .A2(n16582), .ZN(n16580) );
  NAND2_X1 U12998 ( .A1(n19330), .A2(n19331), .ZN(n19329) );
  NAND2_X1 U12999 ( .A1(n15220), .A2(n15536), .ZN(n15219) );
  OR3_X1 U13000 ( .A1(n19282), .A2(n19592), .A3(n12802), .ZN(n19425) );
  INV_X1 U13001 ( .A(n19453), .ZN(n19437) );
  NOR2_X1 U13002 ( .A1(n16698), .A2(n19286), .ZN(n12799) );
  OR2_X1 U13003 ( .A1(n12160), .A2(n12159), .ZN(n13973) );
  NOR2_X1 U13004 ( .A1(n14054), .A2(n13055), .ZN(n19456) );
  AND2_X1 U13005 ( .A1(n13058), .A2(n16042), .ZN(n19496) );
  INV_X1 U13006 ( .A(n19537), .ZN(n19546) );
  INV_X1 U13007 ( .A(n16495), .ZN(n13008) );
  NAND2_X1 U13008 ( .A1(n15653), .A2(n15652), .ZN(n15654) );
  AND2_X1 U13009 ( .A1(n14353), .A2(n15490), .ZN(n15550) );
  NOR2_X1 U13010 ( .A1(n16673), .A2(n16672), .ZN(n15922) );
  INV_X1 U13011 ( .A(n16677), .ZN(n19604) );
  AND2_X1 U13012 ( .A1(n13279), .A2(n13278), .ZN(n20258) );
  OAI21_X1 U13013 ( .B1(n19631), .B2(n19630), .A(n19629), .ZN(n19662) );
  INV_X1 U13014 ( .A(n19704), .ZN(n19726) );
  INV_X1 U13015 ( .A(n19961), .ZN(n20244) );
  NAND2_X1 U13016 ( .A1(n16036), .A2(n16033), .ZN(n19777) );
  INV_X1 U13017 ( .A(n19810), .ZN(n19800) );
  OR3_X1 U13018 ( .A1(n16051), .A2(n16053), .A3(n19782), .ZN(n19826) );
  AND2_X1 U13019 ( .A1(n20248), .A2(n19456), .ZN(n19666) );
  INV_X1 U13020 ( .A(n19871), .ZN(n19896) );
  INV_X1 U13021 ( .A(n19925), .ZN(n19914) );
  NOR2_X2 U13022 ( .A1(n19671), .A2(n16105), .ZN(n19942) );
  NOR2_X1 U13023 ( .A1(n20258), .A2(n20265), .ZN(n19961) );
  INV_X1 U13024 ( .A(n19990), .ZN(n20015) );
  NOR2_X1 U13025 ( .A1(n16104), .A2(n19781), .ZN(n20040) );
  INV_X1 U13026 ( .A(n20135), .ZN(n20079) );
  INV_X1 U13027 ( .A(n20062), .ZN(n20104) );
  INV_X1 U13028 ( .A(n20151), .ZN(n20131) );
  AND2_X1 U13029 ( .A1(n20098), .A2(n19661), .ZN(n20144) );
  INV_X1 U13030 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19955) );
  INV_X1 U13031 ( .A(n19271), .ZN(n19249) );
  NOR3_X1 U13032 ( .A1(n17838), .A2(n16945), .A3(n19062), .ZN(n19038) );
  NOR2_X1 U13033 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17081), .ZN(n17064) );
  NOR2_X1 U13034 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17152), .ZN(n17132) );
  INV_X1 U13035 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19268) );
  INV_X1 U13036 ( .A(n17318), .ZN(n17255) );
  AND2_X1 U13038 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17422), .ZN(n17409) );
  INV_X1 U13039 ( .A(n17621), .ZN(n17586) );
  NOR2_X1 U13040 ( .A1(n14088), .A2(n14102), .ZN(n16299) );
  NAND2_X1 U13041 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17654), .ZN(n17650) );
  INV_X1 U13042 ( .A(n17681), .ZN(n17677) );
  NOR2_X1 U13043 ( .A1(n17842), .A2(n17695), .ZN(n17691) );
  NAND2_X1 U13044 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17738), .ZN(n17737) );
  AND2_X1 U13045 ( .A1(n19071), .A2(n16303), .ZN(n17771) );
  INV_X1 U13046 ( .A(n17835), .ZN(n17777) );
  NOR2_X1 U13047 ( .A1(n17877), .A2(n19256), .ZN(n17885) );
  NOR2_X1 U13048 ( .A1(n19113), .A2(n18226), .ZN(n17969) );
  INV_X1 U13049 ( .A(n18040), .ZN(n18051) );
  INV_X1 U13050 ( .A(n18044), .ZN(n18115) );
  INV_X1 U13051 ( .A(n18168), .ZN(n18150) );
  NAND2_X1 U13052 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  NAND2_X1 U13053 ( .A1(n18475), .A2(n19047), .ZN(n18499) );
  NOR2_X1 U13054 ( .A1(n18450), .A2(n18592), .ZN(n18487) );
  INV_X1 U13055 ( .A(n18509), .ZN(n18489) );
  INV_X1 U13056 ( .A(n18576), .ZN(n18569) );
  NAND2_X1 U13057 ( .A1(n19102), .A2(n18608), .ZN(n18947) );
  NOR2_X1 U13058 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19206), .ZN(
        n19230) );
  OAI22_X1 U13059 ( .A1(n16744), .A2(n18304), .B1(n16743), .B2(n19041), .ZN(
        n19091) );
  NOR2_X1 U13060 ( .A1(n19105), .A2(n19268), .ZN(n19251) );
  INV_X1 U13061 ( .A(n16042), .ZN(n16040) );
  NAND2_X1 U13062 ( .A1(n16254), .A2(n12962), .ZN(n13595) );
  NAND2_X1 U13063 ( .A1(n14770), .A2(n9896), .ZN(n14765) );
  NAND2_X2 U13064 ( .A1(n11788), .A2(n11787), .ZN(n14865) );
  NAND2_X1 U13065 ( .A1(n20381), .A2(n13213), .ZN(n13368) );
  INV_X1 U13066 ( .A(n20381), .ZN(n20408) );
  INV_X1 U13067 ( .A(n20412), .ZN(n13626) );
  NAND2_X1 U13068 ( .A1(n16375), .A2(n13224), .ZN(n16370) );
  OR2_X1 U13069 ( .A1(n20302), .A2(n11448), .ZN(n16375) );
  INV_X1 U13070 ( .A(n20302), .ZN(n16349) );
  OR2_X1 U13071 ( .A1(n13667), .A2(n16481), .ZN(n16444) );
  OR2_X1 U13072 ( .A1(n12876), .A2(n12859), .ZN(n20431) );
  INV_X1 U13073 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20522) );
  INV_X1 U13074 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16486) );
  NAND2_X1 U13075 ( .A1(n20499), .A2(n20661), .ZN(n20519) );
  AOI22_X1 U13076 ( .A1(n20521), .A2(n20525), .B1(n20719), .B2(n10212), .ZN(
        n20546) );
  NAND2_X1 U13077 ( .A1(n20576), .A2(n20661), .ZN(n20629) );
  AOI22_X1 U13078 ( .A1(n20632), .A2(n20638), .B1(n10212), .B2(n20807), .ZN(
        n20660) );
  INV_X1 U13079 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U13080 ( .A1(n20662), .A2(n20661), .ZN(n20717) );
  AOI22_X1 U13081 ( .A1(n20721), .A2(n20729), .B1(n20720), .B2(n20719), .ZN(
        n20763) );
  OR2_X1 U13082 ( .A1(n20778), .A2(n20860), .ZN(n20802) );
  INV_X1 U13083 ( .A(n20912), .ZN(n20826) );
  INV_X1 U13084 ( .A(n20942), .ZN(n20850) );
  INV_X1 U13085 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U13086 ( .A1(n20902), .A2(n20861), .ZN(n20948) );
  INV_X1 U13087 ( .A(n21037), .ZN(n20964) );
  NAND2_X1 U13088 ( .A1(n16509), .A2(n16510), .ZN(n16508) );
  INV_X1 U13089 ( .A(n19448), .ZN(n19427) );
  OR2_X1 U13090 ( .A1(n16495), .A2(n16727), .ZN(n19442) );
  AND2_X1 U13091 ( .A1(n12473), .A2(n13144), .ZN(n19537) );
  INV_X1 U13092 ( .A(n16619), .ZN(n19551) );
  INV_X1 U13093 ( .A(n19558), .ZN(n19591) );
  OR2_X1 U13094 ( .A1(n12936), .A2(n16070), .ZN(n16495) );
  INV_X1 U13095 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19389) );
  OR2_X1 U13096 ( .A1(n19288), .A2(n16070), .ZN(n16664) );
  INV_X1 U13097 ( .A(n13702), .ZN(n13929) );
  INV_X1 U13098 ( .A(n19611), .ZN(n16684) );
  INV_X1 U13099 ( .A(n19693), .ZN(n19690) );
  OR2_X1 U13100 ( .A1(n20244), .A2(n19697), .ZN(n19753) );
  INV_X1 U13101 ( .A(n19760), .ZN(n19780) );
  OR2_X1 U13102 ( .A1(n19697), .A2(n19781), .ZN(n19810) );
  INV_X1 U13103 ( .A(n19817), .ZN(n19829) );
  NAND2_X1 U13104 ( .A1(n20045), .A2(n19666), .ZN(n19871) );
  AOI211_X2 U13105 ( .C1(n16061), .C2(n16064), .A(n16060), .B(n19782), .ZN(
        n19901) );
  NAND2_X1 U13106 ( .A1(n19946), .A2(n19961), .ZN(n19990) );
  INV_X1 U13107 ( .A(n20138), .ZN(n20012) );
  INV_X1 U13108 ( .A(n20040), .ZN(n20037) );
  NAND2_X1 U13109 ( .A1(n19946), .A2(n16106), .ZN(n20090) );
  NAND2_X1 U13110 ( .A1(n19946), .A2(n20045), .ZN(n20134) );
  NAND2_X1 U13111 ( .A1(n20046), .A2(n20045), .ZN(n20151) );
  INV_X1 U13112 ( .A(n20239), .ZN(n20163) );
  NOR2_X1 U13113 ( .A1(n19038), .A2(n17839), .ZN(n19271) );
  NAND2_X1 U13114 ( .A1(n19091), .A2(n19251), .ZN(n16918) );
  NOR3_X1 U13115 ( .A1(n17043), .A2(n17383), .A3(n17382), .ZN(n17381) );
  INV_X1 U13116 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17589) );
  NOR2_X2 U13117 ( .A1(n17586), .A2(n18642), .ZN(n17618) );
  INV_X1 U13118 ( .A(n17701), .ZN(n17671) );
  AND2_X1 U13119 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17722), .ZN(n17725) );
  INV_X1 U13120 ( .A(n11732), .ZN(n17752) );
  INV_X1 U13121 ( .A(n17772), .ZN(n17769) );
  NAND2_X1 U13122 ( .A1(n17837), .A2(n17776), .ZN(n17835) );
  INV_X1 U13123 ( .A(n17885), .ZN(n17880) );
  NAND2_X1 U13124 ( .A1(n17746), .A2(n18228), .ZN(n18084) );
  NAND2_X1 U13125 ( .A1(n18127), .A2(n18372), .ZN(n18040) );
  NAND2_X1 U13126 ( .A1(n16756), .A2(n18228), .ZN(n18168) );
  INV_X1 U13127 ( .A(n18248), .ZN(n18259) );
  OR2_X1 U13128 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  INV_X1 U13129 ( .A(n18575), .ZN(n18592) );
  OR3_X1 U13130 ( .A1(n19212), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18491) );
  NAND2_X1 U13131 ( .A1(n18491), .A2(n18592), .ZN(n18576) );
  INV_X1 U13132 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19206) );
  INV_X1 U13133 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19130) );
  INV_X1 U13134 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10740) );
  INV_X1 U13135 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11350) );
  OR2_X1 U13136 ( .A1(n10359), .A2(n11353), .ZN(n10228) );
  OAI211_X1 U13137 ( .C1(n10551), .C2(n11350), .A(n10229), .B(n10228), .ZN(
        n10230) );
  NAND2_X1 U13138 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10237) );
  NAND2_X1 U13139 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10236) );
  AND2_X2 U13140 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13458) );
  NAND2_X1 U13141 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10235) );
  NAND2_X4 U13142 ( .A1(n13458), .A2(n10233), .ZN(n11406) );
  NAND2_X1 U13143 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10234) );
  INV_X1 U13144 ( .A(n10283), .ZN(n10311) );
  NAND2_X1 U13145 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10240) );
  NAND2_X1 U13146 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U13147 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10247) );
  NAND2_X1 U13148 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10246) );
  AND2_X2 U13149 ( .A1(n13258), .A2(n10244), .ZN(n10382) );
  NAND2_X1 U13150 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10245) );
  NAND4_X1 U13151 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  INV_X1 U13152 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U13153 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10251) );
  OAI21_X1 U13154 ( .B1(n11176), .B2(n9671), .A(n10251), .ZN(n10259) );
  INV_X1 U13155 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U13156 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U13157 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10255) );
  NAND2_X1 U13158 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10254) );
  NAND4_X1 U13159 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10258) );
  OR2_X1 U13160 ( .A1(n11422), .A2(n11382), .ZN(n10264) );
  NAND2_X1 U13161 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U13162 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10262) );
  INV_X1 U13163 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10260) );
  OAI211_X1 U13164 ( .C1(n9657), .C2(n13440), .A(n10265), .B(n10221), .ZN(
        n10266) );
  INV_X1 U13165 ( .A(n10266), .ZN(n10272) );
  INV_X1 U13166 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U13167 ( .A1(n10311), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U13168 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10267) );
  OAI211_X1 U13169 ( .C1(n10551), .C2(n10269), .A(n10268), .B(n10267), .ZN(
        n10270) );
  INV_X1 U13170 ( .A(n10270), .ZN(n10271) );
  NAND2_X1 U13171 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10276) );
  NAND2_X1 U13172 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10275) );
  OAI211_X1 U13173 ( .C1(n9656), .C2(n13417), .A(n10276), .B(n10275), .ZN(
        n10277) );
  INV_X1 U13174 ( .A(n10277), .ZN(n10282) );
  NAND2_X1 U13175 ( .A1(n9788), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10279) );
  OR2_X1 U13176 ( .A1(n9671), .A2(n11131), .ZN(n10278) );
  OAI211_X1 U13177 ( .C1(n10551), .C2(n10617), .A(n10279), .B(n10278), .ZN(
        n10280) );
  INV_X1 U13178 ( .A(n10280), .ZN(n10281) );
  OAI22_X1 U13179 ( .A1(n11422), .A2(n11132), .B1(n11406), .B2(n11329), .ZN(
        n10284) );
  INV_X1 U13180 ( .A(n10286), .ZN(n10292) );
  NAND2_X1 U13181 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U13182 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U13183 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U13184 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10287) );
  NAND4_X1 U13185 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  OR2_X1 U13186 ( .A1(n10359), .A2(n11421), .ZN(n10296) );
  OAI21_X1 U13187 ( .B1(n11419), .B2(n9674), .A(n10298), .ZN(n10299) );
  INV_X1 U13188 ( .A(n10299), .ZN(n10318) );
  NAND2_X1 U13189 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U13190 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U13191 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10303) );
  NAND2_X1 U13192 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13193 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10301) );
  NAND4_X1 U13194 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NAND2_X1 U13195 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10310) );
  NAND2_X1 U13196 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10309) );
  NAND2_X1 U13197 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10308) );
  NAND2_X1 U13198 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10307) );
  NAND2_X1 U13199 ( .A1(n10311), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10313) );
  OAI211_X1 U13200 ( .C1(n9657), .C2(n13404), .A(n10313), .B(n10312), .ZN(
        n10314) );
  INV_X1 U13201 ( .A(n10314), .ZN(n10315) );
  NAND4_X4 U13202 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n14198) );
  NAND2_X1 U13203 ( .A1(n10319), .A2(n10424), .ZN(n10404) );
  INV_X2 U13204 ( .A(n13412), .ZN(n12856) );
  NAND2_X1 U13205 ( .A1(n9650), .A2(n12856), .ZN(n10418) );
  INV_X1 U13206 ( .A(n10418), .ZN(n12848) );
  NAND2_X1 U13207 ( .A1(n13412), .A2(n14198), .ZN(n10396) );
  OR2_X2 U13208 ( .A1(n10396), .A2(n13299), .ZN(n14218) );
  NAND2_X1 U13209 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10323) );
  NAND2_X1 U13210 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10322) );
  NAND2_X1 U13211 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10321) );
  NAND2_X1 U13212 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10325) );
  OR2_X1 U13213 ( .A1(n10359), .A2(n11246), .ZN(n10324) );
  OAI211_X1 U13214 ( .C1(n10551), .C2(n11243), .A(n10325), .B(n10324), .ZN(
        n10326) );
  INV_X1 U13215 ( .A(n10326), .ZN(n10331) );
  NAND2_X1 U13216 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10328) );
  NAND2_X1 U13217 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10327) );
  OAI211_X1 U13218 ( .C1(n9657), .C2(n13398), .A(n10328), .B(n10327), .ZN(
        n10329) );
  INV_X1 U13219 ( .A(n10329), .ZN(n10330) );
  NAND3_X1 U13220 ( .A1(n10331), .A2(n10330), .A3(n9728), .ZN(n10335) );
  OAI22_X1 U13221 ( .A1(n9672), .A2(n10508), .B1(n10495), .B2(n11256), .ZN(
        n10334) );
  INV_X1 U13222 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10332) );
  OAI22_X1 U13223 ( .A1(n11418), .A2(n10332), .B1(n11406), .B2(n11258), .ZN(
        n10333) );
  NOR2_X2 U13224 ( .A1(n10335), .A2(n10223), .ZN(n10336) );
  NAND2_X4 U13225 ( .A1(n10224), .A2(n10336), .ZN(n13635) );
  NAND2_X1 U13226 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10342) );
  NAND2_X1 U13227 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U13228 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U13229 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10339) );
  NAND4_X1 U13230 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND2_X1 U13231 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U13232 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10345) );
  NAND2_X1 U13233 ( .A1(n10518), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10344) );
  NAND2_X1 U13234 ( .A1(n10311), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10348) );
  NAND2_X1 U13235 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10347) );
  OAI211_X1 U13236 ( .C1(n9657), .C2(n13394), .A(n10348), .B(n10347), .ZN(
        n10349) );
  INV_X1 U13237 ( .A(n10349), .ZN(n10352) );
  OR2_X1 U13238 ( .A1(n10359), .A2(n11207), .ZN(n10351) );
  BUF_X4 U13239 ( .A(n10406), .Z(n13213) );
  INV_X1 U13240 ( .A(n11422), .ZN(n11394) );
  AOI22_X1 U13241 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11086), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10358) );
  INV_X1 U13242 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11274) );
  INV_X1 U13243 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11273) );
  OAI22_X1 U13244 ( .A1(n9672), .A2(n11274), .B1(n10495), .B2(n11273), .ZN(
        n10353) );
  INV_X1 U13245 ( .A(n10353), .ZN(n10357) );
  AOI22_X1 U13246 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10356) );
  INV_X1 U13247 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10354) );
  NAND4_X1 U13248 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10369) );
  AOI22_X1 U13249 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10367) );
  INV_X1 U13250 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11277) );
  INV_X1 U13251 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11276) );
  OR2_X1 U13252 ( .A1(n9674), .A2(n11276), .ZN(n10361) );
  INV_X1 U13253 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11275) );
  OR2_X1 U13254 ( .A1(n11297), .A2(n11275), .ZN(n10360) );
  OAI211_X1 U13255 ( .C1(n10551), .C2(n11277), .A(n10361), .B(n10360), .ZN(
        n10362) );
  INV_X1 U13256 ( .A(n10362), .ZN(n10366) );
  AOI22_X1 U13257 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10382), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10365) );
  INV_X1 U13258 ( .A(n10363), .ZN(n10517) );
  AOI22_X1 U13259 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10363), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10364) );
  NAND4_X1 U13260 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10368) );
  NAND2_X1 U13261 ( .A1(n13634), .A2(n13635), .ZN(n16259) );
  OAI21_X1 U13262 ( .B1(n13634), .B2(n10225), .A(n16259), .ZN(n10370) );
  INV_X1 U13263 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U13264 ( .A1(n10311), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10372) );
  NAND2_X1 U13265 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10371) );
  OAI211_X1 U13266 ( .C1(n9657), .C2(n13409), .A(n10372), .B(n10371), .ZN(
        n10378) );
  NAND2_X1 U13267 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13268 ( .A1(n10518), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10375) );
  NAND2_X1 U13269 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13270 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10373) );
  NAND4_X1 U13271 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10377) );
  INV_X1 U13272 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U13273 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10381) );
  NAND2_X1 U13274 ( .A1(n11086), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13275 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10385) );
  NAND2_X1 U13276 ( .A1(n10447), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10384) );
  NAND2_X1 U13277 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10383) );
  NAND4_X1 U13278 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  NOR2_X1 U13279 ( .A1(n10388), .A2(n10387), .ZN(n10393) );
  INV_X1 U13280 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11310) );
  INV_X1 U13281 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11309) );
  OAI22_X1 U13282 ( .A1(n10644), .A2(n11310), .B1(n11365), .B2(n11309), .ZN(
        n10390) );
  INV_X1 U13283 ( .A(n10390), .ZN(n10392) );
  NAND2_X1 U13284 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10391) );
  NAND4_X2 U13285 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n13405) );
  AND2_X4 U13286 ( .A1(n13405), .A2(n13635), .ZN(n14164) );
  INV_X1 U13287 ( .A(n13405), .ZN(n12860) );
  INV_X1 U13288 ( .A(n10810), .ZN(n10395) );
  NAND2_X2 U13289 ( .A1(n10395), .A2(n14198), .ZN(n12862) );
  NAND2_X1 U13290 ( .A1(n10397), .A2(n10421), .ZN(n10398) );
  MUX2_X1 U13291 ( .A(n10399), .B(n10398), .S(n10225), .Z(n10400) );
  NAND2_X1 U13292 ( .A1(n10225), .A2(n13405), .ZN(n12877) );
  XNOR2_X1 U13293 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12837) );
  NAND2_X1 U13294 ( .A1(n21040), .A2(n10532), .ZN(n11453) );
  INV_X1 U13295 ( .A(n11453), .ZN(n10546) );
  NAND2_X1 U13296 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10436) );
  OAI21_X1 U13297 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10436), .ZN(n20864) );
  INV_X1 U13298 ( .A(n20864), .ZN(n10410) );
  NAND2_X1 U13299 ( .A1(n16490), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20961) );
  AND2_X1 U13300 ( .A1(n20961), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10431) );
  AOI21_X1 U13301 ( .B1(n10546), .B2(n10410), .A(n10431), .ZN(n10411) );
  AND2_X1 U13302 ( .A1(n12861), .A2(n16253), .ZN(n13259) );
  NOR2_X1 U13303 ( .A1(n12862), .A2(n10397), .ZN(n10413) );
  NAND2_X1 U13304 ( .A1(n13259), .A2(n10413), .ZN(n12929) );
  NAND3_X1 U13305 ( .A1(n10412), .A2(n10414), .A3(n12929), .ZN(n10415) );
  XNOR2_X2 U13306 ( .A(n10416), .B(n10430), .ZN(n13380) );
  INV_X1 U13307 ( .A(n20961), .ZN(n16274) );
  MUX2_X1 U13308 ( .A(n16274), .B(n11453), .S(n20690), .Z(n10417) );
  NAND3_X1 U13309 ( .A1(n10418), .A2(n13635), .A3(n14218), .ZN(n10429) );
  INV_X1 U13310 ( .A(n16253), .ZN(n12871) );
  NAND3_X1 U13311 ( .A1(n12871), .A2(n13299), .A3(n13405), .ZN(n10419) );
  NAND2_X1 U13312 ( .A1(n10420), .A2(n10419), .ZN(n10428) );
  AND2_X1 U13313 ( .A1(n21040), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10423) );
  INV_X1 U13314 ( .A(n12861), .ZN(n10422) );
  OR2_X1 U13315 ( .A1(n10422), .A2(n10421), .ZN(n12873) );
  OAI211_X1 U13316 ( .C1(n10424), .C2(n16260), .A(n10423), .B(n12873), .ZN(
        n10425) );
  NOR2_X1 U13317 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  NAND3_X1 U13318 ( .A1(n10429), .A2(n10428), .A3(n10427), .ZN(n10463) );
  NAND2_X2 U13319 ( .A1(n13380), .A2(n10528), .ZN(n10531) );
  INV_X1 U13320 ( .A(n10430), .ZN(n10434) );
  INV_X1 U13321 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U13322 ( .A1(n10432), .A2(n10409), .ZN(n10433) );
  NAND2_X1 U13323 ( .A1(n10434), .A2(n10433), .ZN(n10441) );
  INV_X1 U13324 ( .A(n10436), .ZN(n10435) );
  NAND2_X1 U13325 ( .A1(n10435), .A2(n20722), .ZN(n20764) );
  NAND2_X1 U13326 ( .A1(n10436), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U13327 ( .A1(n20764), .A2(n10437), .ZN(n20464) );
  AOI22_X1 U13328 ( .A1(n10546), .A2(n20464), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20961), .ZN(n10438) );
  INV_X1 U13329 ( .A(n10439), .ZN(n10440) );
  AND2_X1 U13330 ( .A1(n10441), .A2(n10440), .ZN(n10442) );
  NAND2_X1 U13331 ( .A1(n10531), .A2(n10442), .ZN(n10443) );
  AOI22_X1 U13332 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10451) );
  INV_X1 U13334 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10913) );
  OR2_X1 U13335 ( .A1(n11365), .A2(n11274), .ZN(n10445) );
  OR2_X1 U13336 ( .A1(n10644), .A2(n11273), .ZN(n10444) );
  OAI211_X1 U13337 ( .C1(n10511), .C2(n10913), .A(n10445), .B(n10444), .ZN(
        n10446) );
  INV_X1 U13338 ( .A(n10446), .ZN(n10450) );
  INV_X1 U13339 ( .A(n10382), .ZN(n11384) );
  AOI22_X1 U13340 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10449) );
  INV_X1 U13341 ( .A(n10447), .ZN(n11225) );
  INV_X1 U13342 ( .A(n11225), .ZN(n11252) );
  AOI22_X1 U13343 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10448) );
  NAND4_X1 U13344 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10460) );
  INV_X1 U13345 ( .A(n10452), .ZN(n11424) );
  INV_X2 U13346 ( .A(n11424), .ZN(n11391) );
  AOI22_X1 U13347 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10458) );
  INV_X1 U13348 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10905) );
  INV_X1 U13349 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11278) );
  OAI22_X1 U13350 ( .A1(n9672), .A2(n10905), .B1(n11425), .B2(n11278), .ZN(
        n10453) );
  INV_X1 U13351 ( .A(n10453), .ZN(n10457) );
  OAI22_X1 U13352 ( .A1(n9664), .A2(n11277), .B1(n11406), .B2(n10354), .ZN(
        n10454) );
  INV_X1 U13353 ( .A(n10454), .ZN(n10456) );
  NAND2_X1 U13354 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10455) );
  NAND4_X1 U13355 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  OAI22_X1 U13356 ( .A1(n10549), .A2(n10598), .B1(n10789), .B2(n10913), .ZN(
        n10461) );
  INV_X1 U13357 ( .A(n10463), .ZN(n10464) );
  XNOR2_X2 U13358 ( .A(n10465), .B(n10464), .ZN(n10812) );
  INV_X1 U13359 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U13360 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10466) );
  OAI21_X1 U13361 ( .B1(n11231), .B2(n10379), .A(n10466), .ZN(n10472) );
  NAND2_X1 U13362 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13363 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13364 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13365 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10467) );
  NAND4_X1 U13366 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10471) );
  NOR2_X1 U13367 ( .A1(n10472), .A2(n10471), .ZN(n10487) );
  NAND2_X1 U13368 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10474) );
  NAND2_X1 U13369 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13370 ( .A1(n10474), .A2(n10473), .ZN(n10476) );
  OAI22_X1 U13371 ( .A1(n9664), .A2(n11407), .B1(n11406), .B2(n13404), .ZN(
        n10475) );
  NOR2_X1 U13372 ( .A1(n10476), .A2(n10475), .ZN(n10486) );
  INV_X1 U13373 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U13374 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10478) );
  NAND2_X1 U13375 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10477) );
  OAI211_X1 U13376 ( .C1(n9657), .C2(n11416), .A(n10478), .B(n10477), .ZN(
        n10479) );
  INV_X1 U13377 ( .A(n10479), .ZN(n10485) );
  INV_X1 U13378 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10482) );
  INV_X1 U13379 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11224) );
  OR2_X1 U13380 ( .A1(n11365), .A2(n11224), .ZN(n10481) );
  INV_X1 U13381 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11415) );
  OR2_X1 U13382 ( .A1(n10644), .A2(n11415), .ZN(n10480) );
  OAI211_X1 U13383 ( .C1(n10511), .C2(n10482), .A(n10481), .B(n10480), .ZN(
        n10483) );
  INV_X1 U13384 ( .A(n10483), .ZN(n10484) );
  NAND4_X1 U13385 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10712) );
  NOR2_X1 U13386 ( .A1(n10550), .A2(n10712), .ZN(n10507) );
  NAND2_X1 U13387 ( .A1(n12856), .A2(n10712), .ZN(n10505) );
  AOI22_X1 U13388 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10494) );
  INV_X1 U13389 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11215) );
  INV_X1 U13390 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11202) );
  OR2_X1 U13391 ( .A1(n11365), .A2(n11202), .ZN(n10489) );
  INV_X1 U13392 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11201) );
  OR2_X1 U13393 ( .A1(n10644), .A2(n11201), .ZN(n10488) );
  OAI211_X1 U13394 ( .C1(n10511), .C2(n11215), .A(n10489), .B(n10488), .ZN(
        n10490) );
  INV_X1 U13395 ( .A(n10490), .ZN(n10493) );
  AOI22_X1 U13396 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13397 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U13398 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10502) );
  AOI22_X1 U13399 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13400 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10499) );
  OAI22_X1 U13401 ( .A1(n9664), .A2(n11217), .B1(n11406), .B2(n13394), .ZN(
        n10496) );
  INV_X1 U13402 ( .A(n10496), .ZN(n10498) );
  NAND2_X1 U13403 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10497) );
  NAND4_X1 U13404 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10501) );
  NOR2_X1 U13405 ( .A1(n10502), .A2(n10501), .ZN(n10579) );
  MUX2_X1 U13406 ( .A(n10507), .B(n10504), .S(n10579), .Z(n10503) );
  INV_X1 U13407 ( .A(n10503), .ZN(n10573) );
  INV_X1 U13408 ( .A(n10579), .ZN(n10582) );
  AOI21_X1 U13409 ( .B1(n13634), .B2(n10582), .A(n10532), .ZN(n10506) );
  OAI211_X1 U13410 ( .C1(n10789), .C2(n11215), .A(n10506), .B(n10505), .ZN(
        n10575) );
  INV_X1 U13411 ( .A(n10507), .ZN(n10527) );
  INV_X1 U13412 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10883) );
  OR2_X1 U13413 ( .A1(n10789), .A2(n10883), .ZN(n10526) );
  AOI22_X1 U13414 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10516) );
  OR2_X1 U13415 ( .A1(n11297), .A2(n10508), .ZN(n10510) );
  OR2_X1 U13416 ( .A1(n10644), .A2(n11256), .ZN(n10509) );
  OAI211_X1 U13417 ( .C1(n10511), .C2(n10883), .A(n10510), .B(n10509), .ZN(
        n10512) );
  INV_X1 U13418 ( .A(n10512), .ZN(n10515) );
  AOI22_X1 U13419 ( .A1(n10338), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13420 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10513) );
  NAND4_X1 U13421 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10524) );
  AOI22_X1 U13422 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13423 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13424 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13425 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10519) );
  NAND4_X1 U13426 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10523) );
  NOR2_X1 U13427 ( .A1(n10524), .A2(n10523), .ZN(n10568) );
  OR2_X1 U13428 ( .A1(n10549), .A2(n10568), .ZN(n10525) );
  INV_X1 U13429 ( .A(n13380), .ZN(n10530) );
  INV_X1 U13430 ( .A(n10528), .ZN(n10529) );
  INV_X1 U13431 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10532) );
  OR2_X1 U13432 ( .A1(n10550), .A2(n10568), .ZN(n10533) );
  INV_X1 U13433 ( .A(n10803), .ZN(n10534) );
  NAND2_X1 U13434 ( .A1(n10804), .A2(n10534), .ZN(n10539) );
  INV_X1 U13435 ( .A(n10535), .ZN(n10536) );
  NAND2_X1 U13436 ( .A1(n10539), .A2(n10538), .ZN(n10593) );
  INV_X1 U13437 ( .A(n10593), .ZN(n10540) );
  INV_X1 U13438 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13439 ( .A1(n10544), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10548) );
  NAND3_X1 U13440 ( .A1(n20862), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20633) );
  INV_X1 U13441 ( .A(n20633), .ZN(n13389) );
  NAND2_X1 U13442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13389), .ZN(
        n13433) );
  NAND2_X1 U13443 ( .A1(n20862), .A2(n13433), .ZN(n10545) );
  NOR3_X1 U13444 ( .A1(n20862), .A2(n20722), .A3(n20522), .ZN(n20908) );
  NAND2_X1 U13445 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20908), .ZN(
        n20894) );
  AOI22_X1 U13446 ( .A1(n10546), .A2(n20664), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20961), .ZN(n10547) );
  INV_X1 U13447 ( .A(n11365), .ZN(n11336) );
  AOI22_X1 U13448 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10558) );
  INV_X1 U13449 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10934) );
  INV_X1 U13450 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11298) );
  OR2_X1 U13451 ( .A1(n10379), .A2(n11298), .ZN(n10553) );
  INV_X1 U13452 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11301) );
  OR2_X1 U13453 ( .A1(n10644), .A2(n11301), .ZN(n10552) );
  OAI211_X1 U13454 ( .C1(n10511), .C2(n10934), .A(n10553), .B(n10552), .ZN(
        n10554) );
  INV_X1 U13455 ( .A(n10554), .ZN(n10557) );
  INV_X1 U13456 ( .A(n10338), .ZN(n11420) );
  AOI22_X1 U13457 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13458 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10555) );
  AND4_X1 U13459 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10564) );
  AOI22_X1 U13460 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13461 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13462 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13463 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10559) );
  AND4_X1 U13464 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  NAND2_X1 U13465 ( .A1(n10564), .A2(n10563), .ZN(n10634) );
  INV_X1 U13466 ( .A(n10789), .ZN(n10792) );
  AOI22_X1 U13467 ( .A1(n10784), .A2(n10634), .B1(n10792), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U13468 ( .A1(n13635), .A2(n10397), .ZN(n10757) );
  INV_X1 U13469 ( .A(n10757), .ZN(n10711) );
  INV_X1 U13470 ( .A(n10568), .ZN(n10583) );
  NAND2_X1 U13471 ( .A1(n10583), .A2(n10582), .ZN(n10597) );
  NAND2_X1 U13472 ( .A1(n10597), .A2(n10598), .ZN(n10635) );
  INV_X1 U13473 ( .A(n10634), .ZN(n10569) );
  XNOR2_X1 U13474 ( .A(n10635), .B(n10569), .ZN(n10570) );
  INV_X1 U13475 ( .A(n16260), .ZN(n21062) );
  NAND2_X1 U13476 ( .A1(n10570), .A2(n21062), .ZN(n10571) );
  INV_X1 U13477 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10572) );
  NAND2_X1 U13478 ( .A1(n10574), .A2(n10573), .ZN(n10576) );
  OR2_X1 U13479 ( .A1(n10576), .A2(n10575), .ZN(n10578) );
  NAND2_X1 U13480 ( .A1(n10576), .A2(n10575), .ZN(n10577) );
  NAND2_X2 U13481 ( .A1(n10578), .A2(n10577), .ZN(n13551) );
  OR2_X2 U13482 ( .A1(n13551), .A2(n10757), .ZN(n10581) );
  AND2_X1 U13483 ( .A1(n13634), .A2(n13405), .ZN(n10599) );
  AOI21_X1 U13484 ( .B1(n10579), .B2(n21062), .A(n10599), .ZN(n10580) );
  OR2_X1 U13485 ( .A1(n10803), .A2(n13638), .ZN(n10587) );
  XNOR2_X1 U13486 ( .A(n10583), .B(n10582), .ZN(n10584) );
  OAI211_X1 U13487 ( .C1(n10584), .C2(n16260), .A(n9836), .B(n10397), .ZN(
        n10585) );
  INV_X1 U13488 ( .A(n10585), .ZN(n10586) );
  NAND2_X1 U13489 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13490 ( .A1(n13234), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10591) );
  INV_X1 U13491 ( .A(n10588), .ZN(n10589) );
  OR2_X1 U13492 ( .A1(n13227), .A2(n10589), .ZN(n10590) );
  INV_X1 U13493 ( .A(n10592), .ZN(n10604) );
  INV_X1 U13494 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U13495 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  OAI21_X1 U13496 ( .B1(n10598), .B2(n10597), .A(n10635), .ZN(n10600) );
  AOI21_X1 U13497 ( .B1(n10600), .B2(n21062), .A(n10599), .ZN(n10601) );
  NAND2_X1 U13498 ( .A1(n13370), .A2(n13369), .ZN(n10607) );
  NAND2_X1 U13499 ( .A1(n10605), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10606) );
  NAND2_X1 U13500 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10608) );
  OAI21_X1 U13501 ( .B1(n10379), .B2(n11329), .A(n10608), .ZN(n10614) );
  NAND2_X1 U13502 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10612) );
  NAND2_X1 U13503 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10611) );
  NAND2_X1 U13504 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10610) );
  NAND2_X1 U13505 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10609) );
  NAND4_X1 U13506 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10613) );
  NOR2_X1 U13507 ( .A1(n10614), .A2(n10613), .ZN(n10631) );
  NAND2_X1 U13508 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10616) );
  NAND2_X1 U13509 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10615) );
  NAND2_X1 U13510 ( .A1(n10616), .A2(n10615), .ZN(n10619) );
  OAI22_X1 U13511 ( .A1(n9664), .A2(n10617), .B1(n11406), .B2(n13417), .ZN(
        n10618) );
  NOR2_X1 U13512 ( .A1(n10619), .A2(n10618), .ZN(n10630) );
  INV_X1 U13513 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U13514 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13515 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10621) );
  OAI211_X1 U13516 ( .C1(n9657), .C2(n11331), .A(n10622), .B(n10621), .ZN(
        n10623) );
  INV_X1 U13517 ( .A(n10623), .ZN(n10629) );
  INV_X1 U13518 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10626) );
  OR2_X1 U13519 ( .A1(n11365), .A2(n11327), .ZN(n10625) );
  OR2_X1 U13520 ( .A1(n10644), .A2(n11326), .ZN(n10624) );
  OAI211_X1 U13521 ( .C1(n10511), .C2(n10626), .A(n10625), .B(n10624), .ZN(
        n10627) );
  INV_X1 U13522 ( .A(n10627), .ZN(n10628) );
  NAND4_X1 U13523 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10695) );
  NAND2_X1 U13524 ( .A1(n10784), .A2(n10695), .ZN(n10633) );
  NAND2_X1 U13525 ( .A1(n10792), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13526 ( .A1(n10633), .A2(n10632), .ZN(n10641) );
  XNOR2_X1 U13527 ( .A(n10642), .B(n10641), .ZN(n10842) );
  NAND2_X1 U13528 ( .A1(n10842), .A2(n10711), .ZN(n10638) );
  NAND2_X1 U13529 ( .A1(n10635), .A2(n10634), .ZN(n10698) );
  INV_X1 U13530 ( .A(n10695), .ZN(n10664) );
  XNOR2_X1 U13531 ( .A(n10698), .B(n10664), .ZN(n10636) );
  OR2_X1 U13532 ( .A1(n10636), .A2(n16260), .ZN(n10637) );
  NAND2_X1 U13533 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  INV_X1 U13534 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20425) );
  XNOR2_X1 U13535 ( .A(n10639), .B(n20425), .ZN(n13530) );
  NAND2_X1 U13536 ( .A1(n10639), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10640) );
  AOI22_X1 U13537 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10652) );
  INV_X1 U13538 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10647) );
  INV_X1 U13539 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10643) );
  OR2_X1 U13540 ( .A1(n11365), .A2(n10643), .ZN(n10646) );
  INV_X1 U13541 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11363) );
  OR2_X1 U13542 ( .A1(n10644), .A2(n11363), .ZN(n10645) );
  OAI211_X1 U13543 ( .C1(n10511), .C2(n10647), .A(n10646), .B(n10645), .ZN(
        n10648) );
  INV_X1 U13544 ( .A(n10648), .ZN(n10651) );
  AOI22_X1 U13545 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13546 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10649) );
  AND4_X1 U13547 ( .A1(n10652), .A2(n10651), .A3(n10650), .A4(n10649), .ZN(
        n10658) );
  AOI22_X1 U13548 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13549 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13550 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U13551 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10653) );
  AND4_X1 U13552 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        n10657) );
  NAND2_X1 U13553 ( .A1(n10658), .A2(n10657), .ZN(n10696) );
  NAND2_X1 U13554 ( .A1(n10784), .A2(n10696), .ZN(n10660) );
  NAND2_X1 U13555 ( .A1(n10792), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10659) );
  NAND2_X1 U13556 ( .A1(n10660), .A2(n10659), .ZN(n10661) );
  OR2_X1 U13557 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  OR2_X1 U13558 ( .A1(n10844), .A2(n10757), .ZN(n10668) );
  OR2_X1 U13559 ( .A1(n10698), .A2(n10664), .ZN(n10665) );
  XNOR2_X1 U13560 ( .A(n10665), .B(n10696), .ZN(n10666) );
  NAND2_X1 U13561 ( .A1(n10666), .A2(n21062), .ZN(n10667) );
  NAND2_X1 U13562 ( .A1(n10668), .A2(n10667), .ZN(n10670) );
  INV_X1 U13563 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10669) );
  XNOR2_X1 U13564 ( .A(n10670), .B(n10669), .ZN(n16369) );
  NAND2_X1 U13565 ( .A1(n10670), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13566 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10673) );
  NAND2_X1 U13567 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10672) );
  OAI211_X1 U13568 ( .C1(n9657), .C2(n10253), .A(n10673), .B(n10672), .ZN(
        n10679) );
  NAND2_X1 U13569 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10677) );
  NAND2_X1 U13570 ( .A1(n10518), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10676) );
  NAND2_X1 U13571 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13572 ( .A1(n11230), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10674) );
  NAND4_X1 U13573 ( .A1(n10677), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10678) );
  NOR2_X1 U13574 ( .A1(n10679), .A2(n10678), .ZN(n10692) );
  INV_X1 U13575 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10683) );
  INV_X1 U13576 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11390) );
  OR2_X1 U13577 ( .A1(n11297), .A2(n11390), .ZN(n10682) );
  INV_X1 U13578 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10680) );
  OR2_X1 U13579 ( .A1(n10644), .A2(n10680), .ZN(n10681) );
  OAI211_X1 U13580 ( .C1(n10511), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10684) );
  INV_X1 U13581 ( .A(n10684), .ZN(n10691) );
  AOI22_X1 U13582 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10690) );
  NAND2_X1 U13583 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10688) );
  NAND2_X1 U13584 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10687) );
  NAND2_X1 U13585 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10686) );
  NAND2_X1 U13586 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10685) );
  AND4_X1 U13587 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  NAND4_X1 U13588 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10700) );
  AOI22_X1 U13589 ( .A1(n10784), .A2(n10700), .B1(n10792), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13590 ( .A1(n10722), .A2(n10694), .ZN(n10856) );
  NAND2_X1 U13591 ( .A1(n10696), .A2(n10695), .ZN(n10697) );
  NOR2_X1 U13592 ( .A1(n10698), .A2(n10697), .ZN(n10699) );
  NAND2_X1 U13593 ( .A1(n10699), .A2(n10700), .ZN(n10725) );
  INV_X1 U13594 ( .A(n10699), .ZN(n10702) );
  INV_X1 U13595 ( .A(n10700), .ZN(n10701) );
  AOI21_X1 U13596 ( .B1(n10702), .B2(n10701), .A(n16260), .ZN(n10703) );
  NAND2_X1 U13597 ( .A1(n10725), .A2(n10703), .ZN(n10704) );
  NAND2_X1 U13598 ( .A1(n10705), .A2(n10704), .ZN(n10706) );
  INV_X1 U13599 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12904) );
  XNOR2_X1 U13600 ( .A(n10706), .B(n12904), .ZN(n13662) );
  NAND2_X1 U13601 ( .A1(n10706), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13602 ( .A1(n10784), .A2(n10712), .ZN(n10709) );
  NAND2_X1 U13603 ( .A1(n10792), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10708) );
  NAND2_X1 U13604 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  NAND2_X1 U13605 ( .A1(n10863), .A2(n10711), .ZN(n10716) );
  INV_X1 U13606 ( .A(n10725), .ZN(n10713) );
  INV_X1 U13607 ( .A(n10712), .ZN(n10724) );
  XNOR2_X1 U13608 ( .A(n10713), .B(n10724), .ZN(n10714) );
  NAND2_X1 U13609 ( .A1(n10714), .A2(n21062), .ZN(n10715) );
  NAND2_X1 U13610 ( .A1(n10716), .A2(n10715), .ZN(n10718) );
  INV_X1 U13611 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10717) );
  XNOR2_X1 U13612 ( .A(n10718), .B(n10717), .ZN(n13966) );
  NAND2_X1 U13613 ( .A1(n10718), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10719) );
  NOR2_X1 U13614 ( .A1(n10720), .A2(n10757), .ZN(n10721) );
  OR3_X1 U13615 ( .A1(n10725), .A2(n10724), .A3(n16260), .ZN(n10726) );
  NAND2_X1 U13616 ( .A1(n10723), .A2(n10726), .ZN(n13956) );
  AND2_X1 U13617 ( .A1(n13956), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10727) );
  NAND2_X1 U13618 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10729) );
  INV_X1 U13619 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U13620 ( .A1(n10723), .A2(n14059), .ZN(n10730) );
  INV_X1 U13621 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U13622 ( .A1(n10723), .A2(n15019), .ZN(n15001) );
  NAND2_X1 U13623 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13624 ( .A1(n10723), .A2(n10731), .ZN(n12830) );
  AND2_X1 U13625 ( .A1(n15001), .A2(n12830), .ZN(n10732) );
  XNOR2_X1 U13626 ( .A(n10723), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16334) );
  INV_X1 U13627 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13628 ( .A1(n10723), .A2(n10739), .ZN(n16331) );
  NAND2_X1 U13629 ( .A1(n16334), .A2(n16331), .ZN(n10733) );
  NOR2_X1 U13630 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10734) );
  INV_X1 U13631 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12917) );
  INV_X1 U13632 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13633 ( .A1(n12917), .A2(n10735), .ZN(n10736) );
  NAND2_X1 U13634 ( .A1(n16352), .A2(n10736), .ZN(n12832) );
  NAND2_X1 U13635 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12834) );
  NAND2_X1 U13636 ( .A1(n12832), .A2(n12834), .ZN(n15144) );
  NOR2_X1 U13637 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10737) );
  NOR2_X1 U13638 ( .A1(n10723), .A2(n10737), .ZN(n10738) );
  INV_X1 U13639 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16393) );
  INV_X1 U13640 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16398) );
  INV_X1 U13641 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U13642 ( .A1(n16352), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14962) );
  NAND2_X1 U13643 ( .A1(n10723), .A2(n16398), .ZN(n10741) );
  NAND2_X1 U13644 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15134) );
  INV_X1 U13645 ( .A(n15134), .ZN(n15032) );
  NAND2_X1 U13646 ( .A1(n15032), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15023) );
  INV_X1 U13647 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14911) );
  INV_X1 U13648 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15115) );
  INV_X1 U13649 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15106) );
  NAND3_X1 U13650 ( .A1(n14911), .A2(n15115), .A3(n15106), .ZN(n14884) );
  NAND2_X1 U13651 ( .A1(n16352), .A2(n14884), .ZN(n10742) );
  NAND2_X1 U13652 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15036) );
  NOR2_X1 U13653 ( .A1(n15036), .A2(n14911), .ZN(n10743) );
  INV_X1 U13654 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15091) );
  NAND2_X1 U13655 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15067) );
  INV_X1 U13656 ( .A(n15067), .ZN(n10746) );
  INV_X1 U13657 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15074) );
  INV_X1 U13658 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U13659 ( .A1(n15074), .A2(n14887), .ZN(n15066) );
  INV_X1 U13660 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15056) );
  NAND2_X1 U13661 ( .A1(n16352), .A2(n15056), .ZN(n14872) );
  NAND2_X1 U13662 ( .A1(n10723), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14871) );
  MUX2_X1 U13663 ( .A(n20522), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10765) );
  NAND2_X1 U13664 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20690), .ZN(
        n10767) );
  NAND2_X1 U13665 ( .A1(n10765), .A2(n10764), .ZN(n10763) );
  NAND2_X1 U13666 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20522), .ZN(
        n10752) );
  NAND2_X1 U13667 ( .A1(n10763), .A2(n10752), .ZN(n10777) );
  NAND2_X1 U13668 ( .A1(n10777), .A2(n10753), .ZN(n10755) );
  NAND2_X1 U13669 ( .A1(n20722), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10754) );
  NAND2_X1 U13670 ( .A1(n10755), .A2(n10754), .ZN(n10761) );
  XNOR2_X1 U13671 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10762) );
  INV_X1 U13672 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20451) );
  NOR2_X1 U13673 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20451), .ZN(
        n10756) );
  NAND2_X1 U13674 ( .A1(n11781), .A2(n10791), .ZN(n10800) );
  NAND2_X1 U13675 ( .A1(n11781), .A2(n10784), .ZN(n10798) );
  NAND3_X1 U13676 ( .A1(n16486), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10758), .ZN(n11779) );
  INV_X1 U13677 ( .A(n10791), .ZN(n10795) );
  INV_X1 U13678 ( .A(n10759), .ZN(n10760) );
  OAI21_X1 U13679 ( .B1(n10762), .B2(n10761), .A(n10760), .ZN(n11777) );
  OAI21_X1 U13680 ( .B1(n10765), .B2(n10764), .A(n10763), .ZN(n11776) );
  INV_X1 U13681 ( .A(n10775), .ZN(n10766) );
  NOR2_X1 U13682 ( .A1(n11776), .A2(n10766), .ZN(n10772) );
  AOI21_X1 U13683 ( .B1(n10295), .B2(n13213), .A(n13635), .ZN(n10786) );
  OAI21_X1 U13684 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20690), .A(
        n10767), .ZN(n10768) );
  AOI211_X1 U13685 ( .C1(n10399), .C2(n13213), .A(n10786), .B(n10768), .ZN(
        n10771) );
  INV_X1 U13686 ( .A(n10768), .ZN(n10769) );
  AOI21_X1 U13687 ( .B1(n10784), .B2(n10769), .A(n10791), .ZN(n10770) );
  NAND2_X1 U13688 ( .A1(n10772), .A2(n10774), .ZN(n10783) );
  NAND2_X1 U13689 ( .A1(n10775), .A2(n13635), .ZN(n10773) );
  OAI211_X1 U13690 ( .C1(n10775), .C2(n10774), .A(n11776), .B(n10773), .ZN(
        n10782) );
  INV_X1 U13691 ( .A(n10784), .ZN(n10780) );
  XNOR2_X1 U13692 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10776) );
  XNOR2_X1 U13693 ( .A(n10777), .B(n10776), .ZN(n11778) );
  NAND2_X1 U13694 ( .A1(n10792), .A2(n11778), .ZN(n10779) );
  INV_X1 U13695 ( .A(n10786), .ZN(n10778) );
  OAI211_X1 U13696 ( .C1(n10780), .C2(n11778), .A(n10779), .B(n10778), .ZN(
        n10781) );
  NAND3_X1 U13697 ( .A1(n10783), .A2(n10782), .A3(n10781), .ZN(n10788) );
  INV_X1 U13698 ( .A(n11778), .ZN(n10785) );
  NAND3_X1 U13699 ( .A1(n10786), .A2(n10785), .A3(n10784), .ZN(n10787) );
  AOI22_X1 U13700 ( .A1(n10789), .A2(n11777), .B1(n10788), .B2(n10787), .ZN(
        n10790) );
  AOI21_X1 U13701 ( .B1(n10791), .B2(n11777), .A(n10790), .ZN(n10794) );
  NOR2_X1 U13702 ( .A1(n10792), .A2(n11779), .ZN(n10793) );
  OAI22_X1 U13703 ( .A1(n11779), .A2(n10795), .B1(n10794), .B2(n10793), .ZN(
        n10796) );
  AOI21_X1 U13704 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10532), .A(
        n10796), .ZN(n10797) );
  NAND2_X1 U13705 ( .A1(n10798), .A2(n10797), .ZN(n10799) );
  NAND2_X1 U13706 ( .A1(n14218), .A2(n13634), .ZN(n10801) );
  AND2_X1 U13707 ( .A1(n10802), .A2(n10801), .ZN(n12849) );
  AND2_X1 U13708 ( .A1(n12849), .A2(n10399), .ZN(n16246) );
  AND2_X1 U13709 ( .A1(n16254), .A2(n16246), .ZN(n16264) );
  XNOR2_X2 U13710 ( .A(n10534), .B(n10804), .ZN(n13553) );
  NAND2_X1 U13711 ( .A1(n13553), .A2(n11010), .ZN(n10809) );
  AOI22_X1 U13712 ( .A1(n11192), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20769), .ZN(n10807) );
  INV_X1 U13713 ( .A(n12862), .ZN(n12843) );
  NAND2_X1 U13714 ( .A1(n12843), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10838) );
  INV_X1 U13715 ( .A(n10838), .ZN(n10805) );
  NAND2_X1 U13716 ( .A1(n10805), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10806) );
  AND2_X1 U13717 ( .A1(n10807), .A2(n10806), .ZN(n10808) );
  NAND2_X1 U13718 ( .A1(n10809), .A2(n10808), .ZN(n13233) );
  NAND2_X1 U13719 ( .A1(n13551), .A2(n10810), .ZN(n10811) );
  NAND2_X1 U13720 ( .A1(n10811), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13220) );
  NAND2_X1 U13721 ( .A1(n20769), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10814) );
  NAND2_X1 U13722 ( .A1(n11192), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10813) );
  OAI211_X1 U13723 ( .C1(n10838), .C2(n14224), .A(n10814), .B(n10813), .ZN(
        n10815) );
  AOI21_X1 U13724 ( .B1(n14221), .B2(n11010), .A(n10815), .ZN(n10816) );
  OR2_X1 U13725 ( .A1(n13220), .A2(n10816), .ZN(n13221) );
  INV_X1 U13726 ( .A(n10816), .ZN(n13222) );
  NOR2_X1 U13727 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10818) );
  OR2_X1 U13728 ( .A1(n13222), .A2(n13628), .ZN(n10817) );
  NAND2_X1 U13729 ( .A1(n13221), .A2(n10817), .ZN(n13232) );
  NAND2_X1 U13730 ( .A1(n13233), .A2(n13232), .ZN(n13231) );
  XNOR2_X1 U13731 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13674) );
  AOI21_X1 U13732 ( .B1(n10818), .B2(n13674), .A(n11443), .ZN(n10820) );
  NAND2_X1 U13733 ( .A1(n11192), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10819) );
  OAI211_X1 U13734 ( .C1(n10838), .C2(n13264), .A(n10820), .B(n10819), .ZN(
        n10821) );
  INV_X1 U13735 ( .A(n10821), .ZN(n10822) );
  NAND2_X1 U13736 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10826) );
  NAND2_X1 U13737 ( .A1(n10823), .A2(n10826), .ZN(n13330) );
  INV_X1 U13738 ( .A(n13330), .ZN(n10824) );
  INV_X1 U13739 ( .A(n10828), .ZN(n10827) );
  INV_X1 U13740 ( .A(n10839), .ZN(n10831) );
  INV_X1 U13741 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U13742 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  NAND2_X1 U13743 ( .A1(n10831), .A2(n10830), .ZN(n20362) );
  AOI22_X1 U13744 ( .A1(n20362), .A2(n11170), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13745 ( .A1(n10857), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10832) );
  OAI211_X1 U13746 ( .C1(n10838), .C2(n13461), .A(n10833), .B(n10832), .ZN(
        n10834) );
  INV_X1 U13747 ( .A(n10834), .ZN(n10835) );
  OAI21_X1 U13748 ( .B1(n20452), .B2(n11031), .A(n10835), .ZN(n13324) );
  NAND2_X1 U13749 ( .A1(n13325), .A2(n13324), .ZN(n13323) );
  NAND2_X1 U13750 ( .A1(n20769), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10837) );
  NAND2_X1 U13751 ( .A1(n11192), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10836) );
  OAI211_X1 U13752 ( .C1(n10838), .C2(n16486), .A(n10837), .B(n10836), .ZN(
        n10840) );
  OAI21_X1 U13753 ( .B1(n10839), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10846), .ZN(n20360) );
  MUX2_X1 U13754 ( .A(n10840), .B(n20360), .S(n11170), .Z(n10841) );
  INV_X1 U13755 ( .A(n10844), .ZN(n10845) );
  NAND2_X1 U13756 ( .A1(n10845), .A2(n11010), .ZN(n10851) );
  INV_X1 U13757 ( .A(n11443), .ZN(n10928) );
  AND2_X1 U13758 ( .A1(n10846), .A2(n16376), .ZN(n10847) );
  OR2_X1 U13759 ( .A1(n10847), .A2(n10852), .ZN(n20336) );
  NAND2_X1 U13760 ( .A1(n20336), .A2(n11170), .ZN(n10848) );
  OAI21_X1 U13761 ( .B1(n16376), .B2(n10928), .A(n10848), .ZN(n10849) );
  AOI21_X1 U13762 ( .B1(n11192), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10849), .ZN(
        n10850) );
  NOR2_X1 U13763 ( .A1(n10852), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10853) );
  OR2_X1 U13764 ( .A1(n10858), .A2(n10853), .ZN(n13802) );
  AOI22_X1 U13765 ( .A1(n13802), .A2(n11170), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13766 ( .A1(n10857), .A2(P1_EAX_REG_6__SCAN_IN), .ZN(n10854) );
  INV_X1 U13767 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10861) );
  NOR2_X1 U13768 ( .A1(n10858), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10859) );
  OR2_X1 U13769 ( .A1(n10882), .A2(n10859), .ZN(n16360) );
  AOI22_X1 U13770 ( .A1(n16360), .A2(n11170), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10860) );
  OAI21_X1 U13771 ( .B1(n10992), .B2(n10861), .A(n10860), .ZN(n10862) );
  AOI22_X1 U13772 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13773 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13774 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10864) );
  AND3_X1 U13775 ( .A1(n10866), .A2(n10865), .A3(n10864), .ZN(n10875) );
  AOI22_X1 U13776 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13777 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13778 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U13779 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10867) );
  AND4_X1 U13780 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(
        n10874) );
  INV_X1 U13781 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11216) );
  OAI22_X1 U13782 ( .A1(n10644), .A2(n11216), .B1(n10379), .B2(n13394), .ZN(
        n10871) );
  INV_X1 U13783 ( .A(n10871), .ZN(n10873) );
  NAND2_X1 U13784 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10872) );
  NAND4_X1 U13785 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(
        n10876) );
  NAND2_X1 U13786 ( .A1(n11010), .A2(n10876), .ZN(n10880) );
  NAND2_X1 U13787 ( .A1(n10857), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10879) );
  XNOR2_X1 U13788 ( .A(n10882), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13959) );
  NAND2_X1 U13789 ( .A1(n13959), .A2(n11170), .ZN(n10878) );
  NAND2_X1 U13790 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10877) );
  XOR2_X1 U13791 ( .A(n20322), .B(n10921), .Z(n20320) );
  INV_X1 U13792 ( .A(n20320), .ZN(n14064) );
  INV_X1 U13793 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11060) );
  OAI22_X1 U13794 ( .A1(n11425), .A2(n11060), .B1(n9664), .B2(n10883), .ZN(
        n10884) );
  INV_X1 U13795 ( .A(n10884), .ZN(n10888) );
  AOI22_X1 U13796 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13797 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13798 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10885) );
  NAND4_X1 U13799 ( .A1(n10888), .A2(n10887), .A3(n10886), .A4(n10885), .ZN(
        n10900) );
  INV_X1 U13800 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U13801 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10891) );
  INV_X1 U13802 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10889) );
  OR2_X1 U13803 ( .A1(n11297), .A2(n10889), .ZN(n10890) );
  OAI211_X1 U13804 ( .C1(n9657), .C2(n11054), .A(n10891), .B(n10890), .ZN(
        n10892) );
  INV_X1 U13805 ( .A(n10892), .ZN(n10898) );
  INV_X1 U13806 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10893) );
  OAI22_X1 U13807 ( .A1(n10644), .A2(n10893), .B1(n10379), .B2(n13398), .ZN(
        n10894) );
  INV_X1 U13808 ( .A(n10894), .ZN(n10897) );
  AOI22_X1 U13809 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13810 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10895) );
  NAND4_X1 U13811 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10899) );
  OAI21_X1 U13812 ( .B1(n10900), .B2(n10899), .A(n11010), .ZN(n10903) );
  NAND2_X1 U13813 ( .A1(n10857), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U13814 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10901) );
  NAND3_X1 U13815 ( .A1(n10903), .A2(n10902), .A3(n10901), .ZN(n10904) );
  AOI22_X1 U13816 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10912) );
  INV_X1 U13817 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11079) );
  OR2_X1 U13818 ( .A1(n10379), .A2(n10354), .ZN(n10907) );
  OR2_X1 U13819 ( .A1(n11297), .A2(n10905), .ZN(n10906) );
  OAI211_X1 U13820 ( .C1(n9657), .C2(n11079), .A(n10907), .B(n10906), .ZN(
        n10908) );
  INV_X1 U13821 ( .A(n10908), .ZN(n10911) );
  AOI22_X1 U13822 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13823 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U13824 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10920) );
  AOI22_X1 U13825 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13826 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10917) );
  INV_X1 U13827 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U13828 ( .A1(n9664), .A2(n10913), .B1(n11406), .B2(n11085), .ZN(
        n10914) );
  INV_X1 U13829 ( .A(n10914), .ZN(n10916) );
  NAND2_X1 U13830 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10915) );
  NAND4_X1 U13831 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n10919) );
  NOR2_X1 U13832 ( .A1(n10920), .A2(n10919), .ZN(n10924) );
  XNOR2_X1 U13833 ( .A(n10925), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15013) );
  NAND2_X1 U13834 ( .A1(n15013), .A2(n11170), .ZN(n10923) );
  AOI22_X1 U13835 ( .A1(n10857), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11443), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10922) );
  OAI211_X1 U13836 ( .C1(n10924), .C2(n11031), .A(n10923), .B(n10922), .ZN(
        n14067) );
  INV_X1 U13837 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10929) );
  OAI21_X1 U13838 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10926), .A(
        n10973), .ZN(n16359) );
  NAND2_X1 U13839 ( .A1(n16359), .A2(n11170), .ZN(n10927) );
  OAI21_X1 U13840 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(n10930) );
  AOI21_X1 U13841 ( .B1(n11192), .B2(P1_EAX_REG_11__SCAN_IN), .A(n10930), .ZN(
        n10931) );
  NAND2_X1 U13842 ( .A1(n10954), .A2(n10933), .ZN(n14777) );
  INV_X1 U13843 ( .A(n14777), .ZN(n10953) );
  OAI22_X1 U13844 ( .A1(n11425), .A2(n11101), .B1(n9664), .B2(n10934), .ZN(
        n10935) );
  INV_X1 U13845 ( .A(n10935), .ZN(n10939) );
  AOI22_X1 U13846 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13847 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U13848 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10936) );
  AND4_X1 U13849 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10950) );
  AOI22_X1 U13850 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10949) );
  INV_X1 U13851 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10940) );
  OAI22_X1 U13852 ( .A1(n10644), .A2(n10940), .B1(n10379), .B2(n13409), .ZN(
        n10946) );
  NAND2_X1 U13853 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10944) );
  NAND2_X1 U13854 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10943) );
  NAND2_X1 U13855 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10942) );
  NAND2_X1 U13856 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10941) );
  NAND4_X1 U13857 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10945) );
  NOR2_X1 U13858 ( .A1(n10946), .A2(n10945), .ZN(n10948) );
  NAND2_X1 U13859 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10947) );
  NAND4_X1 U13860 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(
        n10951) );
  NAND2_X1 U13861 ( .A1(n11010), .A2(n10951), .ZN(n14776) );
  INV_X1 U13862 ( .A(n14776), .ZN(n10952) );
  NAND2_X1 U13863 ( .A1(n10953), .A2(n10952), .ZN(n14779) );
  INV_X1 U13864 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14862) );
  XOR2_X1 U13865 ( .A(n14724), .B(n10973), .Z(n16345) );
  INV_X1 U13866 ( .A(n16345), .ZN(n10955) );
  AOI22_X1 U13867 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11170), .B2(n10955), .ZN(n10972) );
  AOI22_X1 U13868 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13869 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11393), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13870 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10956) );
  AND3_X1 U13871 ( .A1(n10958), .A2(n10957), .A3(n10956), .ZN(n10969) );
  AOI22_X1 U13872 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13873 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13874 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11338), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U13875 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10959) );
  AND4_X1 U13876 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(
        n10968) );
  INV_X1 U13877 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10964) );
  INV_X1 U13878 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10963) );
  OAI22_X1 U13879 ( .A1(n10964), .A2(n10644), .B1(n11365), .B2(n10963), .ZN(
        n10965) );
  INV_X1 U13880 ( .A(n10965), .ZN(n10967) );
  NAND2_X1 U13881 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10966) );
  NAND4_X1 U13882 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10970) );
  NAND2_X1 U13883 ( .A1(n11010), .A2(n10970), .ZN(n10971) );
  OAI211_X1 U13884 ( .C1(n10992), .C2(n14862), .A(n10972), .B(n10971), .ZN(
        n14721) );
  INV_X1 U13885 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14859) );
  INV_X1 U13886 ( .A(n10994), .ZN(n10974) );
  XNOR2_X1 U13887 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10974), .ZN(
        n14999) );
  AOI22_X1 U13888 ( .A1(n11170), .A2(n14999), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13889 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13890 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13891 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10975) );
  AND3_X1 U13892 ( .A1(n10977), .A2(n10976), .A3(n10975), .ZN(n10988) );
  AOI22_X1 U13893 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10982) );
  OAI22_X1 U13894 ( .A1(n9672), .A2(n13576), .B1(n11425), .B2(n11151), .ZN(
        n10978) );
  INV_X1 U13895 ( .A(n10978), .ZN(n10981) );
  AOI22_X1 U13896 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U13897 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10979) );
  AND4_X1 U13898 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10987) );
  INV_X1 U13899 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10983) );
  OAI22_X1 U13900 ( .A1(n11365), .A2(n10983), .B1(n10379), .B2(n13429), .ZN(
        n10984) );
  INV_X1 U13901 ( .A(n10984), .ZN(n10986) );
  NAND2_X1 U13902 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10985) );
  NAND4_X1 U13903 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10989) );
  NAND2_X1 U13904 ( .A1(n11010), .A2(n10989), .ZN(n10990) );
  OAI211_X1 U13905 ( .C1(n10992), .C2(n14859), .A(n10991), .B(n10990), .ZN(
        n14707) );
  XOR2_X1 U13906 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11013), .Z(
        n16340) );
  AOI22_X1 U13907 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13908 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13909 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10995) );
  AND3_X1 U13910 ( .A1(n10997), .A2(n10996), .A3(n10995), .ZN(n11008) );
  AOI22_X1 U13911 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13912 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11001) );
  OAI22_X1 U13913 ( .A1(n9664), .A2(n10683), .B1(n11406), .B2(n10253), .ZN(
        n10998) );
  INV_X1 U13914 ( .A(n10998), .ZN(n11000) );
  NAND2_X1 U13915 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10999) );
  AND4_X1 U13916 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11007) );
  INV_X1 U13917 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11003) );
  OAI22_X1 U13918 ( .A1(n10644), .A2(n11003), .B1(n10379), .B2(n13440), .ZN(
        n11004) );
  INV_X1 U13919 ( .A(n11004), .ZN(n11006) );
  NAND2_X1 U13920 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11005) );
  NAND4_X1 U13921 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n11009) );
  AOI22_X1 U13922 ( .A1(n11010), .A2(n11009), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U13923 ( .A1(n11192), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11011) );
  OAI211_X1 U13924 ( .C1(n16340), .C2(n13628), .A(n11012), .B(n11011), .ZN(
        n14698) );
  XNOR2_X1 U13925 ( .A(n11034), .B(n11033), .ZN(n16313) );
  AOI22_X1 U13926 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11020) );
  INV_X1 U13927 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11409) );
  INV_X1 U13928 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11423) );
  OR2_X1 U13929 ( .A1(n10644), .A2(n11423), .ZN(n11015) );
  INV_X1 U13930 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11417) );
  OR2_X1 U13931 ( .A1(n11297), .A2(n11417), .ZN(n11014) );
  OAI211_X1 U13932 ( .C1(n10511), .C2(n11409), .A(n11015), .B(n11014), .ZN(
        n11016) );
  INV_X1 U13933 ( .A(n11016), .ZN(n11019) );
  AOI22_X1 U13934 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U13935 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11017) );
  NAND4_X1 U13936 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11027) );
  OAI22_X1 U13937 ( .A1(n11425), .A2(n11419), .B1(n9664), .B2(n10482), .ZN(
        n11021) );
  INV_X1 U13938 ( .A(n11021), .ZN(n11025) );
  AOI22_X1 U13939 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U13940 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U13941 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11022) );
  NAND4_X1 U13942 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11026) );
  NOR2_X1 U13943 ( .A1(n11027), .A2(n11026), .ZN(n11030) );
  NAND2_X1 U13944 ( .A1(n11192), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U13945 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11028) );
  OAI211_X1 U13946 ( .C1(n11031), .C2(n11030), .A(n11029), .B(n11028), .ZN(
        n11032) );
  AOI21_X1 U13947 ( .B1(n16313), .B2(n11170), .A(n11032), .ZN(n14761) );
  OAI21_X1 U13948 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11035), .A(
        n11071), .ZN(n16339) );
  OAI22_X1 U13949 ( .A1(n10644), .A2(n11212), .B1(n11365), .B2(n13572), .ZN(
        n11036) );
  INV_X1 U13950 ( .A(n11036), .ZN(n11043) );
  NAND2_X1 U13951 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11038) );
  INV_X1 U13952 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11203) );
  OR2_X1 U13953 ( .A1(n10379), .A2(n11203), .ZN(n11037) );
  OAI211_X1 U13954 ( .C1(n9657), .C2(n11206), .A(n11038), .B(n11037), .ZN(
        n11039) );
  INV_X1 U13955 ( .A(n11039), .ZN(n11042) );
  AOI22_X1 U13956 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13957 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U13958 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n11050) );
  AOI22_X1 U13959 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13960 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11047) );
  INV_X1 U13961 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11213) );
  OAI22_X1 U13962 ( .A1(n9672), .A2(n9975), .B1(n11406), .B2(n11213), .ZN(
        n11044) );
  INV_X1 U13963 ( .A(n11044), .ZN(n11046) );
  NAND2_X1 U13964 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11045) );
  NAND4_X1 U13965 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11049) );
  NOR2_X1 U13966 ( .A1(n11050), .A2(n11049), .ZN(n11052) );
  AOI22_X1 U13967 ( .A1(n10857), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20769), .ZN(n11051) );
  OAI21_X1 U13968 ( .B1(n11438), .B2(n11052), .A(n11051), .ZN(n11053) );
  MUX2_X1 U13969 ( .A(n16339), .B(n11053), .S(n13628), .Z(n14752) );
  AOI22_X1 U13970 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U13971 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11058) );
  OAI22_X1 U13972 ( .A1(n11425), .A2(n11258), .B1(n11406), .B2(n11054), .ZN(
        n11055) );
  INV_X1 U13973 ( .A(n11055), .ZN(n11057) );
  NAND2_X1 U13974 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11056) );
  AND4_X1 U13975 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11070) );
  AOI22_X1 U13976 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11069) );
  OAI22_X1 U13977 ( .A1(n10644), .A2(n11060), .B1(n11365), .B2(n13591), .ZN(
        n11066) );
  NAND2_X1 U13978 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U13979 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U13980 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11062) );
  NAND2_X1 U13981 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11061) );
  NAND4_X1 U13982 ( .A1(n11064), .A2(n11063), .A3(n11062), .A4(n11061), .ZN(
        n11065) );
  NOR2_X1 U13983 ( .A1(n11066), .A2(n11065), .ZN(n11068) );
  NAND2_X1 U13984 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11067) );
  NAND4_X1 U13985 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11074) );
  INV_X1 U13986 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14839) );
  XNOR2_X1 U13987 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11075), .ZN(
        n14985) );
  AOI22_X1 U13988 ( .A1(n11170), .A2(n14985), .B1(n11443), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11072) );
  OAI21_X1 U13989 ( .B1(n10992), .B2(n14839), .A(n11072), .ZN(n11073) );
  AOI21_X1 U13990 ( .B1(n11402), .B2(n11074), .A(n11073), .ZN(n14686) );
  INV_X1 U13991 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14972) );
  INV_X1 U13992 ( .A(n11076), .ZN(n11077) );
  NAND2_X1 U13993 ( .A1(n14972), .A2(n11077), .ZN(n11078) );
  AND2_X1 U13994 ( .A1(n11143), .A2(n11078), .ZN(n14974) );
  AOI22_X1 U13995 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U13996 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11083) );
  INV_X1 U13997 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11279) );
  OAI22_X1 U13998 ( .A1(n11425), .A2(n11279), .B1(n11406), .B2(n11079), .ZN(
        n11080) );
  INV_X1 U13999 ( .A(n11080), .ZN(n11082) );
  NAND2_X1 U14000 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11081) );
  AND4_X1 U14001 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11096) );
  AOI22_X1 U14002 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11095) );
  INV_X1 U14003 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13560) );
  OAI22_X1 U14004 ( .A1(n11365), .A2(n13560), .B1(n10379), .B2(n11085), .ZN(
        n11092) );
  NAND2_X1 U14005 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14006 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14007 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14008 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11087) );
  NAND4_X1 U14009 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11091) );
  NOR2_X1 U14010 ( .A1(n11092), .A2(n11091), .ZN(n11094) );
  NAND2_X1 U14011 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11093) );
  NAND4_X1 U14012 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(
        n11098) );
  INV_X1 U14013 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14834) );
  OAI22_X1 U14014 ( .A1(n10992), .A2(n14834), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14972), .ZN(n11097) );
  AOI21_X1 U14015 ( .B1(n11402), .B2(n11098), .A(n11097), .ZN(n11099) );
  MUX2_X1 U14016 ( .A(n14974), .B(n11099), .S(n13628), .Z(n14672) );
  NAND2_X1 U14017 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11103) );
  OR2_X1 U14018 ( .A1(n10644), .A2(n11101), .ZN(n11102) );
  OAI211_X1 U14019 ( .C1(n9657), .C2(n11309), .A(n11103), .B(n11102), .ZN(
        n11104) );
  INV_X1 U14020 ( .A(n11104), .ZN(n11110) );
  INV_X1 U14021 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13568) );
  INV_X1 U14022 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11105) );
  OAI22_X1 U14023 ( .A1(n11365), .A2(n13568), .B1(n10379), .B2(n11105), .ZN(
        n11106) );
  INV_X1 U14024 ( .A(n11106), .ZN(n11109) );
  AOI22_X1 U14025 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14026 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11107) );
  NAND4_X1 U14027 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11118) );
  AOI22_X1 U14028 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14029 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11115) );
  INV_X1 U14030 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11111) );
  OAI22_X1 U14031 ( .A1(n11425), .A2(n11298), .B1(n11406), .B2(n11111), .ZN(
        n11112) );
  INV_X1 U14032 ( .A(n11112), .ZN(n11114) );
  NAND2_X1 U14033 ( .A1(n9976), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11113) );
  NAND4_X1 U14034 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n11117) );
  NOR2_X1 U14035 ( .A1(n11118), .A2(n11117), .ZN(n11121) );
  INV_X1 U14036 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11142) );
  AOI21_X1 U14037 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n11142), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11119) );
  AOI21_X1 U14038 ( .B1(n11192), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11119), .ZN(
        n11120) );
  OAI21_X1 U14039 ( .B1(n11438), .B2(n11121), .A(n11120), .ZN(n11123) );
  XNOR2_X1 U14040 ( .A(n11143), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14965) );
  NAND2_X1 U14041 ( .A1(n14965), .A2(n11170), .ZN(n11122) );
  NAND2_X1 U14042 ( .A1(n11123), .A2(n11122), .ZN(n14661) );
  AOI22_X1 U14043 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11130) );
  OR2_X1 U14044 ( .A1(n10379), .A2(n11331), .ZN(n11125) );
  INV_X1 U14045 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13584) );
  OR2_X1 U14046 ( .A1(n11297), .A2(n13584), .ZN(n11124) );
  OAI211_X1 U14047 ( .C1(n9657), .C2(n11330), .A(n11125), .B(n11124), .ZN(
        n11126) );
  INV_X1 U14048 ( .A(n11126), .ZN(n11129) );
  AOI22_X1 U14049 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11393), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14050 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11338), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11127) );
  AND4_X1 U14051 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11138) );
  AOI22_X1 U14052 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14053 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11230), .B1(
        n10518), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11136) );
  NOR2_X1 U14054 ( .A1(n10511), .A2(n11131), .ZN(n11134) );
  OAI22_X1 U14055 ( .A1(n9672), .A2(n11132), .B1(n11425), .B2(n11329), .ZN(
        n11133) );
  NOR2_X1 U14056 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  NAND4_X1 U14057 ( .A1(n11138), .A2(n11137), .A3(n11136), .A4(n11135), .ZN(
        n11139) );
  NAND2_X1 U14058 ( .A1(n11402), .A2(n11139), .ZN(n11150) );
  INV_X1 U14059 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21129) );
  OAI21_X1 U14060 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21129), .A(
        n20769), .ZN(n11140) );
  INV_X1 U14061 ( .A(n11140), .ZN(n11141) );
  AOI21_X1 U14062 ( .B1(n11192), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11141), .ZN(
        n11149) );
  INV_X1 U14063 ( .A(n11144), .ZN(n11146) );
  INV_X1 U14064 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14065 ( .A1(n11146), .A2(n11145), .ZN(n11147) );
  NAND2_X1 U14066 ( .A1(n11193), .A2(n11147), .ZN(n14958) );
  NOR2_X1 U14067 ( .A1(n14958), .A2(n13628), .ZN(n11148) );
  AOI21_X1 U14068 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n14647) );
  NAND2_X1 U14069 ( .A1(n10380), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11153) );
  OR2_X1 U14070 ( .A1(n10644), .A2(n11151), .ZN(n11152) );
  OAI211_X1 U14071 ( .C1(n10511), .C2(n11353), .A(n11153), .B(n11152), .ZN(
        n11154) );
  INV_X1 U14072 ( .A(n11154), .ZN(n11160) );
  INV_X1 U14073 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11155) );
  OAI22_X1 U14074 ( .A1(n11365), .A2(n13576), .B1(n10379), .B2(n11155), .ZN(
        n11156) );
  INV_X1 U14075 ( .A(n11156), .ZN(n11159) );
  AOI22_X1 U14076 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14077 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11157) );
  NAND4_X1 U14078 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(
        n11166) );
  AOI22_X1 U14079 ( .A1(n10620), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14080 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14081 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U14082 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11161) );
  NAND4_X1 U14083 ( .A1(n11164), .A2(n11163), .A3(n11162), .A4(n11161), .ZN(
        n11165) );
  NOR2_X1 U14084 ( .A1(n11166), .A2(n11165), .ZN(n11169) );
  INV_X1 U14085 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14945) );
  AOI21_X1 U14086 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14945), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11167) );
  AOI21_X1 U14087 ( .B1(n11192), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11167), .ZN(
        n11168) );
  OAI21_X1 U14088 ( .B1(n11438), .B2(n11169), .A(n11168), .ZN(n11172) );
  XNOR2_X1 U14089 ( .A(n11193), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14947) );
  NAND2_X1 U14090 ( .A1(n14947), .A2(n11170), .ZN(n11171) );
  AOI22_X1 U14091 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11181) );
  INV_X1 U14092 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13580) );
  OR2_X1 U14093 ( .A1(n11297), .A2(n13580), .ZN(n11175) );
  OR2_X1 U14094 ( .A1(n10644), .A2(n11173), .ZN(n11174) );
  OAI211_X1 U14095 ( .C1(n10511), .C2(n11176), .A(n11175), .B(n11174), .ZN(
        n11177) );
  INV_X1 U14096 ( .A(n11177), .ZN(n11180) );
  AOI22_X1 U14097 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14098 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11178) );
  AND4_X1 U14099 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11188) );
  OAI22_X1 U14100 ( .A1(n9672), .A2(n11382), .B1(n11425), .B2(n10260), .ZN(
        n11184) );
  INV_X1 U14101 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11182) );
  INV_X1 U14102 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11381) );
  OAI22_X1 U14103 ( .A1(n9664), .A2(n11182), .B1(n11406), .B2(n11381), .ZN(
        n11183) );
  NOR2_X1 U14104 ( .A1(n11184), .A2(n11183), .ZN(n11187) );
  AOI22_X1 U14105 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U14106 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11185) );
  NAND4_X1 U14107 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n11189) );
  NAND2_X1 U14108 ( .A1(n11402), .A2(n11189), .ZN(n11200) );
  OAI21_X1 U14109 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21129), .A(
        n20769), .ZN(n11190) );
  INV_X1 U14110 ( .A(n11190), .ZN(n11191) );
  AOI21_X1 U14111 ( .B1(n11192), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11191), .ZN(
        n11199) );
  INV_X1 U14112 ( .A(n11195), .ZN(n11196) );
  INV_X1 U14113 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U14114 ( .A1(n11196), .A2(n14629), .ZN(n11197) );
  NAND2_X1 U14115 ( .A1(n11265), .A2(n11197), .ZN(n14941) );
  NOR2_X1 U14116 ( .A1(n14941), .A2(n13628), .ZN(n11198) );
  OAI22_X1 U14117 ( .A1(n9657), .A2(n11202), .B1(n10511), .B2(n11201), .ZN(
        n11211) );
  INV_X1 U14118 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11204) );
  OAI22_X1 U14119 ( .A1(n11418), .A2(n11204), .B1(n11225), .B2(n11203), .ZN(
        n11210) );
  INV_X1 U14120 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11205) );
  OAI22_X1 U14121 ( .A1(n10644), .A2(n11205), .B1(n11365), .B2(n9975), .ZN(
        n11209) );
  OAI22_X1 U14122 ( .A1(n9664), .A2(n11207), .B1(n11406), .B2(n11206), .ZN(
        n11208) );
  OR4_X1 U14123 ( .A1(n11211), .A2(n11210), .A3(n11209), .A4(n11208), .ZN(
        n11223) );
  OAI22_X1 U14124 ( .A1(n11420), .A2(n11212), .B1(n11384), .B2(n13572), .ZN(
        n11221) );
  INV_X1 U14125 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11214) );
  OAI22_X1 U14126 ( .A1(n9649), .A2(n11214), .B1(n10379), .B2(n11213), .ZN(
        n11220) );
  OAI22_X1 U14127 ( .A1(n11424), .A2(n11216), .B1(n10517), .B2(n11215), .ZN(
        n11219) );
  OAI22_X1 U14128 ( .A1(n9672), .A2(n11217), .B1(n11425), .B2(n13394), .ZN(
        n11218) );
  OR4_X1 U14129 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11222) );
  NOR2_X1 U14130 ( .A1(n11223), .A2(n11222), .ZN(n11241) );
  OAI22_X1 U14131 ( .A1(n9657), .A2(n11405), .B1(n10511), .B2(n11421), .ZN(
        n11229) );
  OAI22_X1 U14132 ( .A1(n11418), .A2(n11224), .B1(n11420), .B2(n11423), .ZN(
        n11228) );
  INV_X1 U14133 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13564) );
  OAI22_X1 U14134 ( .A1(n11424), .A2(n11415), .B1(n11365), .B2(n13564), .ZN(
        n11227) );
  INV_X1 U14135 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11408) );
  OAI22_X1 U14136 ( .A1(n11225), .A2(n13404), .B1(n11406), .B2(n11408), .ZN(
        n11226) );
  OR4_X1 U14137 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11237) );
  OAI22_X1 U14138 ( .A1(n11384), .A2(n11417), .B1(n9664), .B2(n11409), .ZN(
        n11235) );
  OAI22_X1 U14139 ( .A1(n9649), .A2(n10482), .B1(n10379), .B2(n11416), .ZN(
        n11234) );
  OAI22_X1 U14140 ( .A1(n10517), .A2(n11407), .B1(n9672), .B2(n11426), .ZN(
        n11233) );
  OAI22_X1 U14141 ( .A1(n10644), .A2(n11419), .B1(n11425), .B2(n11231), .ZN(
        n11232) );
  OR4_X1 U14142 ( .A1(n11235), .A2(n11234), .A3(n11233), .A4(n11232), .ZN(
        n11236) );
  NOR2_X1 U14143 ( .A1(n11237), .A2(n11236), .ZN(n11242) );
  XOR2_X1 U14144 ( .A(n11241), .B(n11242), .Z(n11239) );
  INV_X1 U14145 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14811) );
  INV_X1 U14146 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14930) );
  OAI22_X1 U14147 ( .A1(n10992), .A2(n14811), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14930), .ZN(n11238) );
  AOI21_X1 U14148 ( .B1(n11239), .B2(n11402), .A(n11238), .ZN(n11240) );
  XNOR2_X1 U14149 ( .A(n11265), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14932) );
  MUX2_X1 U14150 ( .A(n11240), .B(n14932), .S(n11170), .Z(n14613) );
  NOR2_X1 U14151 ( .A1(n11242), .A2(n11241), .ZN(n11272) );
  AOI22_X1 U14152 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11251) );
  OAI22_X1 U14153 ( .A1(n9672), .A2(n11243), .B1(n11425), .B2(n13398), .ZN(
        n11244) );
  INV_X1 U14154 ( .A(n11244), .ZN(n11250) );
  OAI22_X1 U14155 ( .A1(n9664), .A2(n11246), .B1(n11406), .B2(n11245), .ZN(
        n11247) );
  INV_X1 U14156 ( .A(n11247), .ZN(n11249) );
  NAND2_X1 U14157 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11248) );
  NAND4_X1 U14158 ( .A1(n11251), .A2(n11250), .A3(n11249), .A4(n11248), .ZN(
        n11262) );
  AOI22_X1 U14159 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14160 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14161 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11253) );
  NAND3_X1 U14162 ( .A1(n11255), .A2(n11254), .A3(n11253), .ZN(n11261) );
  NOR2_X1 U14163 ( .A1(n10511), .A2(n11256), .ZN(n11260) );
  OAI22_X1 U14164 ( .A1(n10644), .A2(n11258), .B1(n11365), .B2(n11257), .ZN(
        n11259) );
  OR4_X1 U14165 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11271) );
  XNOR2_X1 U14166 ( .A(n11272), .B(n11271), .ZN(n11264) );
  AOI22_X1 U14167 ( .A1(n10857), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20769), .ZN(n11263) );
  OAI21_X1 U14168 ( .B1(n11264), .B2(n11438), .A(n11263), .ZN(n11270) );
  INV_X1 U14169 ( .A(n11267), .ZN(n11268) );
  INV_X1 U14170 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U14171 ( .A1(n11268), .A2(n14605), .ZN(n11269) );
  NAND2_X1 U14172 ( .A1(n11320), .A2(n11269), .ZN(n14919) );
  MUX2_X1 U14173 ( .A(n11270), .B(n14919), .S(n10818), .Z(n14602) );
  NAND2_X1 U14174 ( .A1(n14600), .A2(n14602), .ZN(n14590) );
  NAND2_X1 U14175 ( .A1(n11272), .A2(n11271), .ZN(n11294) );
  OAI22_X1 U14176 ( .A1(n9657), .A2(n11274), .B1(n10511), .B2(n11273), .ZN(
        n11283) );
  OAI22_X1 U14177 ( .A1(n11420), .A2(n11276), .B1(n11406), .B2(n11275), .ZN(
        n11282) );
  OAI22_X1 U14178 ( .A1(n11424), .A2(n11278), .B1(n9672), .B2(n11277), .ZN(
        n11281) );
  OAI22_X1 U14179 ( .A1(n10644), .A2(n11279), .B1(n11425), .B2(n10354), .ZN(
        n11280) );
  OR4_X1 U14180 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n11290) );
  AOI22_X1 U14181 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14182 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14183 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14184 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14185 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11289) );
  NOR2_X1 U14186 ( .A1(n11290), .A2(n11289), .ZN(n11295) );
  XOR2_X1 U14187 ( .A(n11294), .B(n11295), .Z(n11292) );
  INV_X1 U14188 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14801) );
  INV_X1 U14189 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14915) );
  OAI22_X1 U14190 ( .A1(n10992), .A2(n14801), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14915), .ZN(n11291) );
  AOI21_X1 U14191 ( .B1(n11292), .B2(n11402), .A(n11291), .ZN(n11293) );
  XNOR2_X1 U14192 ( .A(n11320), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14913) );
  MUX2_X1 U14193 ( .A(n11293), .B(n14913), .S(n11170), .Z(n14591) );
  NOR2_X1 U14194 ( .A1(n11295), .A2(n11294), .ZN(n11325) );
  AOI22_X1 U14195 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11306) );
  INV_X1 U14196 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11296) );
  OR2_X1 U14197 ( .A1(n11297), .A2(n11296), .ZN(n11300) );
  OR2_X1 U14198 ( .A1(n10644), .A2(n11298), .ZN(n11299) );
  OAI211_X1 U14199 ( .C1(n10511), .C2(n11301), .A(n11300), .B(n11299), .ZN(
        n11302) );
  INV_X1 U14200 ( .A(n11302), .ZN(n11305) );
  AOI22_X1 U14201 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10382), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14202 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11303) );
  AND4_X1 U14203 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n11317) );
  AOI22_X1 U14204 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11315) );
  INV_X1 U14205 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11307) );
  OAI22_X1 U14206 ( .A1(n9672), .A2(n11307), .B1(n11425), .B2(n13409), .ZN(
        n11308) );
  INV_X1 U14207 ( .A(n11308), .ZN(n11314) );
  OAI22_X1 U14208 ( .A1(n9664), .A2(n11310), .B1(n11406), .B2(n11309), .ZN(
        n11311) );
  INV_X1 U14209 ( .A(n11311), .ZN(n11313) );
  NAND2_X1 U14210 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11312) );
  AND4_X1 U14211 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n11316) );
  NAND2_X1 U14212 ( .A1(n11317), .A2(n11316), .ZN(n11324) );
  XNOR2_X1 U14213 ( .A(n11325), .B(n11324), .ZN(n11319) );
  AOI22_X1 U14214 ( .A1(n10857), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20769), .ZN(n11318) );
  OAI21_X1 U14215 ( .B1(n11319), .B2(n11438), .A(n11318), .ZN(n11323) );
  INV_X1 U14216 ( .A(n11321), .ZN(n11322) );
  INV_X1 U14217 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14580) );
  OAI21_X1 U14218 ( .B1(n11322), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11373), .ZN(n14900) );
  MUX2_X1 U14219 ( .A(n11323), .B(n14900), .S(n10818), .Z(n14577) );
  NAND2_X1 U14220 ( .A1(n11325), .A2(n11324), .ZN(n11348) );
  OAI22_X1 U14221 ( .A1(n11327), .A2(n9657), .B1(n10511), .B2(n11326), .ZN(
        n11335) );
  OAI22_X1 U14222 ( .A1(n10517), .A2(n10626), .B1(n11425), .B2(n13417), .ZN(
        n11334) );
  INV_X1 U14223 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11328) );
  OAI22_X1 U14224 ( .A1(n11329), .A2(n10644), .B1(n10379), .B2(n11328), .ZN(
        n11333) );
  OAI22_X1 U14225 ( .A1(n11225), .A2(n11331), .B1(n11406), .B2(n11330), .ZN(
        n11332) );
  OR4_X1 U14226 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11344) );
  AOI22_X1 U14227 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14228 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11393), .B1(
        n11337), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14229 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14230 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11339) );
  NAND4_X1 U14231 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11343) );
  NOR2_X1 U14232 ( .A1(n11344), .A2(n11343), .ZN(n11349) );
  XOR2_X1 U14233 ( .A(n11348), .B(n11349), .Z(n11346) );
  INV_X1 U14234 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14793) );
  INV_X1 U14235 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14896) );
  OAI22_X1 U14236 ( .A1(n10992), .A2(n14793), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14896), .ZN(n11345) );
  AOI21_X1 U14237 ( .B1(n11346), .B2(n11402), .A(n11345), .ZN(n11347) );
  XNOR2_X1 U14238 ( .A(n11373), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14894) );
  MUX2_X1 U14239 ( .A(n11347), .B(n14894), .S(n10818), .Z(n14563) );
  NOR2_X1 U14240 ( .A1(n11349), .A2(n11348), .ZN(n11380) );
  AOI22_X1 U14241 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11358) );
  OAI22_X1 U14242 ( .A1(n9672), .A2(n11350), .B1(n11425), .B2(n13429), .ZN(
        n11351) );
  INV_X1 U14243 ( .A(n11351), .ZN(n11357) );
  OAI22_X1 U14244 ( .A1(n9664), .A2(n11353), .B1(n11406), .B2(n11352), .ZN(
        n11354) );
  INV_X1 U14245 ( .A(n11354), .ZN(n11356) );
  NAND2_X1 U14246 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11355) );
  NAND4_X1 U14247 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11370) );
  AOI22_X1 U14248 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10380), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14249 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10382), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14250 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11360) );
  NAND3_X1 U14251 ( .A1(n11362), .A2(n11361), .A3(n11360), .ZN(n11369) );
  NOR2_X1 U14252 ( .A1(n10511), .A2(n11363), .ZN(n11368) );
  INV_X1 U14253 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11366) );
  INV_X1 U14254 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11364) );
  OAI22_X1 U14255 ( .A1(n10644), .A2(n11366), .B1(n11365), .B2(n11364), .ZN(
        n11367) );
  OR4_X1 U14256 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n11379) );
  XNOR2_X1 U14257 ( .A(n11380), .B(n11379), .ZN(n11372) );
  AOI22_X1 U14258 ( .A1(n10857), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20769), .ZN(n11371) );
  OAI21_X1 U14259 ( .B1(n11372), .B2(n11438), .A(n11371), .ZN(n11378) );
  INV_X1 U14260 ( .A(n11374), .ZN(n11376) );
  INV_X1 U14261 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14262 ( .A1(n11376), .A2(n11375), .ZN(n11377) );
  NAND2_X1 U14263 ( .A1(n11440), .A2(n11377), .ZN(n14881) );
  MUX2_X1 U14264 ( .A(n11378), .B(n14881), .S(n10818), .Z(n14547) );
  NAND2_X1 U14265 ( .A1(n11380), .A2(n11379), .ZN(n11433) );
  OAI22_X1 U14266 ( .A1(n11365), .A2(n11382), .B1(n10379), .B2(n11381), .ZN(
        n11386) );
  OAI22_X1 U14267 ( .A1(n11384), .A2(n13580), .B1(n11406), .B2(n11383), .ZN(
        n11385) );
  AOI211_X1 U14268 ( .C1(n9976), .C2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11386), .B(n11385), .ZN(n11389) );
  OAI22_X1 U14269 ( .A1(n10644), .A2(n10260), .B1(n11425), .B2(n13440), .ZN(
        n11387) );
  INV_X1 U14270 ( .A(n11387), .ZN(n11388) );
  OAI211_X1 U14271 ( .C1(n9657), .C2(n11390), .A(n11389), .B(n11388), .ZN(
        n11400) );
  AOI22_X1 U14272 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10447), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14273 ( .A1(n11392), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11391), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14274 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14275 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11395) );
  NAND4_X1 U14276 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11399) );
  NOR2_X1 U14277 ( .A1(n11400), .A2(n11399), .ZN(n11434) );
  XOR2_X1 U14278 ( .A(n11433), .B(n11434), .Z(n11403) );
  INV_X1 U14279 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14786) );
  INV_X1 U14280 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14877) );
  OAI22_X1 U14281 ( .A1(n10992), .A2(n14786), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14877), .ZN(n11401) );
  AOI21_X1 U14282 ( .B1(n11403), .B2(n11402), .A(n11401), .ZN(n11404) );
  XNOR2_X1 U14283 ( .A(n11440), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14875) );
  MUX2_X1 U14284 ( .A(n11404), .B(n14875), .S(n10818), .Z(n14532) );
  OAI22_X1 U14285 ( .A1(n9672), .A2(n11407), .B1(n11406), .B2(n11405), .ZN(
        n11411) );
  OAI22_X1 U14286 ( .A1(n9649), .A2(n11409), .B1(n10379), .B2(n11408), .ZN(
        n11410) );
  AOI211_X1 U14287 ( .C1(n11412), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n11411), .B(n11410), .ZN(n11414) );
  AOI22_X1 U14288 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11230), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11413) );
  OAI211_X1 U14289 ( .C1(n10511), .C2(n11415), .A(n11414), .B(n11413), .ZN(
        n11432) );
  OAI22_X1 U14290 ( .A1(n11418), .A2(n11417), .B1(n11225), .B2(n11416), .ZN(
        n11430) );
  OAI22_X1 U14291 ( .A1(n11420), .A2(n11419), .B1(n11384), .B2(n13564), .ZN(
        n11429) );
  OAI22_X1 U14292 ( .A1(n11424), .A2(n11423), .B1(n9664), .B2(n11421), .ZN(
        n11428) );
  OAI22_X1 U14293 ( .A1(n11365), .A2(n11426), .B1(n11425), .B2(n13404), .ZN(
        n11427) );
  OR4_X1 U14294 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11431) );
  NOR2_X1 U14295 ( .A1(n11432), .A2(n11431), .ZN(n11436) );
  NOR2_X1 U14296 ( .A1(n11434), .A2(n11433), .ZN(n11435) );
  XOR2_X1 U14297 ( .A(n11436), .B(n11435), .Z(n11439) );
  AOI22_X1 U14298 ( .A1(n10857), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20769), .ZN(n11437) );
  OAI21_X1 U14299 ( .B1(n11439), .B2(n11438), .A(n11437), .ZN(n11442) );
  INV_X1 U14300 ( .A(n11440), .ZN(n11441) );
  XNOR2_X1 U14301 ( .A(n11451), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14209) );
  MUX2_X1 U14302 ( .A(n11442), .B(n14209), .S(n10818), .Z(n14190) );
  AOI22_X1 U14303 ( .A1(n11192), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11443), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11444) );
  INV_X1 U14304 ( .A(n11444), .ZN(n11445) );
  XNOR2_X2 U14305 ( .A(n14189), .B(n11445), .ZN(n14168) );
  AND2_X1 U14306 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11447) );
  NOR2_X2 U14307 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20907) );
  NOR2_X1 U14308 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20901), .ZN(n11446) );
  AND2_X2 U14309 ( .A1(n11447), .A2(n11446), .ZN(n16364) );
  NAND2_X1 U14310 ( .A1(n14168), .A2(n16364), .ZN(n11457) );
  NAND2_X1 U14311 ( .A1(n11453), .A2(n20901), .ZN(n21060) );
  AND2_X1 U14312 ( .A1(n21060), .A2(n10532), .ZN(n11448) );
  NAND2_X1 U14313 ( .A1(n10532), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14314 ( .A1(n21129), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U14315 ( .A1(n11450), .A2(n11449), .ZN(n13224) );
  NAND2_X1 U14316 ( .A1(n11451), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11452) );
  INV_X1 U14317 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14179) );
  XNOR2_X1 U14318 ( .A(n11452), .B(n14179), .ZN(n13642) );
  OR2_X2 U14319 ( .A1(n11453), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20347) );
  INV_X1 U14320 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21197) );
  NOR2_X1 U14321 ( .A1(n20347), .A2(n21197), .ZN(n15027) );
  AOI21_X1 U14322 ( .B1(n16351), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15027), .ZN(n11454) );
  OAI21_X1 U14323 ( .B1(n16370), .B2(n13642), .A(n11454), .ZN(n11455) );
  INV_X1 U14324 ( .A(n11455), .ZN(n11456) );
  AOI22_X1 U14325 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11474) );
  NOR3_X2 U14326 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n19065), .ZN(n11489) );
  BUF_X4 U14327 ( .A(n11489), .Z(n17567) );
  NOR2_X2 U14328 ( .A1(n17302), .A2(n11458), .ZN(n11555) );
  AOI22_X1 U14329 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11473) );
  NOR2_X2 U14330 ( .A1(n19065), .A2(n11458), .ZN(n11512) );
  BUF_X4 U14331 ( .A(n11512), .Z(n17566) );
  INV_X2 U14332 ( .A(n17522), .ZN(n17552) );
  AOI22_X1 U14333 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11459) );
  OAI21_X1 U14334 ( .B1(n17257), .B2(n17589), .A(n11459), .ZN(n11471) );
  AOI22_X1 U14335 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14336 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11468) );
  INV_X2 U14337 ( .A(n17333), .ZN(n17553) );
  AOI22_X1 U14338 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14339 ( .A1(n9868), .A2(n19229), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U14340 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11466) );
  NAND4_X1 U14341 ( .A1(n11469), .A2(n11468), .A3(n11467), .A4(n11466), .ZN(
        n11470) );
  AOI211_X1 U14342 ( .C1(n17566), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n11471), .B(n11470), .ZN(n11472) );
  NAND3_X1 U14343 ( .A1(n11474), .A2(n11473), .A3(n11472), .ZN(n16756) );
  CLKBUF_X3 U14344 ( .A(n11553), .Z(n17573) );
  AOI22_X1 U14345 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11485) );
  INV_X1 U14346 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14347 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14348 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11475) );
  OAI211_X1 U14349 ( .C1(n16179), .C2(n11477), .A(n11476), .B(n11475), .ZN(
        n11483) );
  AOI22_X1 U14350 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14351 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14352 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14353 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14354 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11482) );
  AOI211_X1 U14355 ( .C1(n17455), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n11483), .B(n11482), .ZN(n11484) );
  NAND2_X1 U14356 ( .A1(n11485), .A2(n11484), .ZN(n11732) );
  AOI22_X1 U14357 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14358 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11497) );
  INV_X1 U14359 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U14360 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11488) );
  OAI21_X1 U14361 ( .B1(n17257), .B2(n17608), .A(n11488), .ZN(n11495) );
  AOI22_X1 U14362 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14363 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14364 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14365 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11490) );
  NAND4_X1 U14366 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11494) );
  AOI211_X1 U14367 ( .C1(n9653), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11495), .B(n11494), .ZN(n11496) );
  AOI22_X1 U14368 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14369 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14370 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14371 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14372 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11508) );
  AOI22_X1 U14373 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14374 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14375 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14376 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11503) );
  NAND4_X1 U14377 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  AOI22_X1 U14378 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11509), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9651), .ZN(n11520) );
  AOI22_X1 U14379 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11489), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11519) );
  INV_X1 U14380 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17613) );
  AOI22_X1 U14381 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11464), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11510), .ZN(n11511) );
  OAI21_X1 U14382 ( .B1(n17257), .B2(n17613), .A(n11511), .ZN(n11518) );
  AOI22_X1 U14383 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14384 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11512), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14385 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17574), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17537), .ZN(n11515) );
  AOI22_X1 U14386 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14387 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14388 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14389 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14390 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11521) );
  NAND4_X1 U14391 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11530) );
  AOI22_X1 U14392 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14393 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14394 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14395 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11525) );
  NAND4_X1 U14396 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11529) );
  AOI22_X1 U14397 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14398 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14399 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14400 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11531) );
  NAND4_X1 U14401 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11540) );
  AOI22_X1 U14402 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14403 ( .A1(n17552), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14404 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14405 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14406 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11539) );
  NAND2_X1 U14407 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18272) );
  INV_X1 U14408 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18289) );
  INV_X1 U14409 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18310) );
  NOR2_X1 U14410 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18142), .ZN(
        n18024) );
  INV_X1 U14411 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18367) );
  NAND2_X1 U14412 ( .A1(n18024), .A2(n18367), .ZN(n11541) );
  NOR2_X1 U14413 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11541), .ZN(
        n17984) );
  INV_X1 U14414 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18344) );
  NAND2_X1 U14415 ( .A1(n17984), .A2(n18344), .ZN(n17973) );
  NOR3_X1 U14416 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17973), .ZN(n11583) );
  INV_X1 U14417 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18398) );
  INV_X1 U14418 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18383) );
  NOR2_X1 U14419 ( .A1(n18398), .A2(n18383), .ZN(n18375) );
  NAND2_X1 U14420 ( .A1(n18375), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17999) );
  NAND2_X1 U14421 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18343) );
  INV_X1 U14422 ( .A(n18343), .ZN(n17986) );
  NAND2_X1 U14423 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17986), .ZN(
        n18325) );
  NOR2_X1 U14424 ( .A1(n17999), .A2(n18325), .ZN(n18334) );
  NAND2_X1 U14425 ( .A1(n18334), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17913) );
  INV_X1 U14426 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U14427 ( .A1(n17913), .A2(n17964), .ZN(n18280) );
  AOI21_X1 U14428 ( .B1(n17746), .B2(n11542), .A(n18142), .ZN(n11576) );
  XOR2_X1 U14429 ( .A(n11544), .B(n11543), .Z(n11573) );
  NAND2_X1 U14430 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11573), .ZN(
        n11574) );
  INV_X1 U14431 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18529) );
  XOR2_X1 U14432 ( .A(n17752), .B(n11545), .Z(n18195) );
  XOR2_X1 U14433 ( .A(n11547), .B(n11546), .Z(n11548) );
  NAND2_X1 U14434 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11548), .ZN(
        n11572) );
  XOR2_X1 U14435 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11548), .Z(
        n18216) );
  XNOR2_X1 U14436 ( .A(n11736), .B(n11549), .ZN(n11568) );
  INV_X1 U14437 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18567) );
  OR2_X1 U14438 ( .A1(n18567), .A2(n11566), .ZN(n11567) );
  NAND2_X1 U14439 ( .A1(n11550), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11565) );
  XNOR2_X1 U14440 ( .A(n17770), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18246) );
  AOI22_X1 U14441 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14442 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11563) );
  INV_X1 U14443 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U14444 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14445 ( .B1(n17257), .B2(n16146), .A(n11552), .ZN(n11561) );
  AOI22_X1 U14446 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14447 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9666), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14448 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14449 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11556) );
  NAND4_X1 U14450 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11560) );
  AOI211_X1 U14451 ( .C1(n17567), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n11561), .B(n11560), .ZN(n11562) );
  INV_X1 U14452 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19232) );
  NAND2_X1 U14453 ( .A1(n11565), .A2(n18245), .ZN(n18238) );
  NAND2_X1 U14454 ( .A1(n11568), .A2(n11570), .ZN(n11571) );
  XOR2_X1 U14455 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11573), .Z(
        n18183) );
  NAND2_X1 U14456 ( .A1(n11576), .A2(n11575), .ZN(n11577) );
  NOR2_X1 U14457 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18140) );
  NOR4_X1 U14458 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11578) );
  INV_X1 U14459 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18401) );
  NAND4_X1 U14460 ( .A1(n18062), .A2(n18140), .A3(n11578), .A4(n18401), .ZN(
        n11579) );
  NAND2_X1 U14461 ( .A1(n18155), .A2(n11579), .ZN(n11581) );
  INV_X1 U14462 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18426) );
  NAND2_X1 U14463 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18128) );
  INV_X1 U14464 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18436) );
  NOR2_X1 U14465 ( .A1(n18128), .A2(n18436), .ZN(n18103) );
  NAND2_X1 U14466 ( .A1(n18103), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18415) );
  INV_X1 U14467 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18420) );
  NOR2_X1 U14468 ( .A1(n18415), .A2(n18420), .ZN(n18422) );
  INV_X1 U14469 ( .A(n18422), .ZN(n18076) );
  NOR2_X1 U14470 ( .A1(n18426), .A2(n18076), .ZN(n18393) );
  NAND2_X1 U14471 ( .A1(n18393), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18048) );
  NAND2_X1 U14472 ( .A1(n18372), .A2(n18061), .ZN(n11582) );
  NAND2_X1 U14473 ( .A1(n11581), .A2(n11582), .ZN(n18049) );
  OAI221_X1 U14474 ( .B1(n11583), .B2(n18280), .C1(n11583), .C2(n18049), .A(
        n17997), .ZN(n11584) );
  INV_X1 U14475 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18018) );
  INV_X1 U14476 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18262) );
  NAND2_X1 U14477 ( .A1(n18375), .A2(n18049), .ZN(n17983) );
  NAND2_X1 U14478 ( .A1(n18155), .A2(n17949), .ZN(n11585) );
  NOR2_X1 U14479 ( .A1(n11586), .A2(n18155), .ZN(n17939) );
  NAND2_X1 U14480 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11587), .ZN(
        n11673) );
  NOR2_X2 U14481 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11587), .ZN(
        n17906) );
  INV_X1 U14482 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16211) );
  OAI22_X1 U14483 ( .A1(n16211), .A2(n18155), .B1(n18142), .B2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17890) );
  AOI22_X1 U14484 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14485 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14486 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14487 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U14488 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11597) );
  AOI22_X1 U14489 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14490 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14491 ( .A1(n17552), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14492 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14493 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  AOI22_X1 U14494 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14495 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11606) );
  INV_X1 U14496 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U14497 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11598) );
  OAI21_X1 U14498 ( .B1(n11462), .B2(n17612), .A(n11598), .ZN(n11604) );
  AOI22_X1 U14499 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14500 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14501 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14502 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U14503 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11603) );
  AOI211_X1 U14504 ( .C1(n11509), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n11604), .B(n11603), .ZN(n11605) );
  NAND3_X1 U14505 ( .A1(n11607), .A2(n11606), .A3(n11605), .ZN(n11711) );
  NOR2_X1 U14506 ( .A1(n19256), .A2(n11711), .ZN(n11694) );
  AOI22_X1 U14507 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14508 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11616) );
  INV_X1 U14509 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17593) );
  AOI22_X1 U14510 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11608) );
  OAI21_X1 U14511 ( .B1(n11462), .B2(n17593), .A(n11608), .ZN(n11614) );
  AOI22_X1 U14512 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14513 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14514 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14515 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11609) );
  NAND4_X1 U14516 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n11613) );
  AOI211_X1 U14517 ( .C1(n11509), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n11614), .B(n11613), .ZN(n11615) );
  NAND2_X1 U14518 ( .A1(n11694), .A2(n18632), .ZN(n11707) );
  AOI22_X1 U14519 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14520 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14521 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14522 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U14523 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n11627) );
  AOI22_X1 U14524 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14525 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14526 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14527 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U14528 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11626) );
  AOI22_X1 U14529 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14530 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14531 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14532 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11628) );
  NAND4_X1 U14533 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11637) );
  AOI22_X1 U14534 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14535 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14536 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14537 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11632) );
  NAND4_X1 U14538 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11636) );
  AOI22_X1 U14539 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14540 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14541 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9666), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11639) );
  OAI21_X1 U14542 ( .B1(n11462), .B2(n17589), .A(n11639), .ZN(n11646) );
  AOI22_X1 U14543 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14544 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14545 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14546 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11641) );
  NAND4_X1 U14547 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11641), .ZN(
        n11645) );
  NAND3_X2 U14548 ( .A1(n11649), .A2(n11648), .A3(n11647), .ZN(n17729) );
  AOI22_X1 U14549 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14550 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14551 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11650) );
  OAI21_X1 U14552 ( .B1(n11462), .B2(n17608), .A(n11650), .ZN(n11656) );
  AOI22_X1 U14553 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14554 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14555 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14556 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14557 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  AOI211_X1 U14558 ( .C1(n17466), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11656), .B(n11655), .ZN(n11657) );
  NAND3_X1 U14559 ( .A1(n11659), .A2(n11658), .A3(n11657), .ZN(n18619) );
  INV_X1 U14560 ( .A(n11715), .ZN(n11710) );
  AND2_X1 U14561 ( .A1(n11717), .A2(n11710), .ZN(n11671) );
  AOI22_X1 U14562 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11670) );
  INV_X1 U14563 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14564 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14565 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11660) );
  OAI211_X1 U14566 ( .C1(n16179), .C2(n11662), .A(n11661), .B(n11660), .ZN(
        n11668) );
  AOI22_X1 U14567 ( .A1(n17575), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14568 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14569 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14570 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14571 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11667) );
  NAND2_X1 U14572 ( .A1(n11712), .A2(n11714), .ZN(n11719) );
  OAI211_X1 U14573 ( .C1(n11709), .C2(n17622), .A(n11671), .B(n11719), .ZN(
        n11701) );
  NOR2_X1 U14574 ( .A1(n19041), .A2(n17746), .ZN(n18406) );
  INV_X1 U14575 ( .A(n18406), .ZN(n11672) );
  NOR2_X1 U14576 ( .A1(n17889), .A2(n11672), .ZN(n11731) );
  INV_X1 U14577 ( .A(n11673), .ZN(n17907) );
  NAND2_X1 U14578 ( .A1(n19216), .A2(n19206), .ZN(n19212) );
  AOI22_X1 U14579 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19076), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19229), .ZN(n11688) );
  INV_X1 U14580 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19081) );
  OAI21_X1 U14581 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n9868), .A(
        n11675), .ZN(n11676) );
  OAI22_X1 U14582 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19085), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11676), .ZN(n11682) );
  NOR2_X1 U14583 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19085), .ZN(
        n11677) );
  NAND2_X1 U14584 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11676), .ZN(
        n11683) );
  AOI22_X1 U14585 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11682), .B1(
        n11677), .B2(n11683), .ZN(n11692) );
  OAI21_X1 U14586 ( .B1(n11680), .B2(n11679), .A(n11692), .ZN(n11678) );
  AOI21_X1 U14587 ( .B1(n19235), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n11681), .ZN(n11687) );
  XOR2_X1 U14588 ( .A(n11688), .B(n11681), .Z(n11686) );
  AOI21_X1 U14589 ( .B1(n11683), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n11682), .ZN(n11684) );
  AOI21_X1 U14590 ( .B1(n19085), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n11684), .ZN(n11685) );
  INV_X1 U14591 ( .A(n11685), .ZN(n11689) );
  AOI21_X1 U14592 ( .B1(n11690), .B2(n11687), .A(n16915), .ZN(n19040) );
  INV_X1 U14593 ( .A(n19040), .ZN(n16743) );
  AND2_X1 U14594 ( .A1(n11688), .A2(n11687), .ZN(n11691) );
  AOI211_X1 U14595 ( .C1(n11692), .C2(n11691), .A(n11690), .B(n11689), .ZN(
        n19036) );
  NOR2_X1 U14596 ( .A1(n11712), .A2(n11711), .ZN(n11706) );
  NAND2_X1 U14597 ( .A1(n19130), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19266) );
  INV_X2 U14598 ( .A(n19266), .ZN(n19265) );
  NAND2_X1 U14599 ( .A1(n19265), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19195) );
  OAI211_X1 U14600 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19130), .B(n19189), .ZN(n19254) );
  OAI21_X1 U14601 ( .B1(n18616), .B2(n16745), .A(n19254), .ZN(n11693) );
  NAND2_X1 U14602 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19257) );
  OAI21_X1 U14603 ( .B1(n11694), .B2(n11693), .A(n19257), .ZN(n16914) );
  AOI211_X1 U14604 ( .C1(n18616), .C2(n18627), .A(n16915), .B(n16914), .ZN(
        n11705) );
  NAND2_X1 U14605 ( .A1(n18627), .A2(n18632), .ZN(n11703) );
  NAND2_X1 U14606 ( .A1(n18616), .A2(n11717), .ZN(n11697) );
  NOR2_X1 U14607 ( .A1(n11712), .A2(n18632), .ZN(n19071) );
  AOI21_X1 U14608 ( .B1(n18616), .B2(n16946), .A(n19071), .ZN(n11695) );
  AOI21_X1 U14609 ( .B1(n11714), .B2(n11703), .A(n11695), .ZN(n11696) );
  AOI21_X1 U14610 ( .B1(n11703), .B2(n11697), .A(n11696), .ZN(n11700) );
  AOI21_X1 U14611 ( .B1(n17729), .B2(n11703), .A(n11709), .ZN(n11698) );
  INV_X1 U14612 ( .A(n11698), .ZN(n11699) );
  OAI211_X1 U14613 ( .C1(n11702), .C2(n18619), .A(n11700), .B(n11699), .ZN(
        n11721) );
  NOR2_X1 U14614 ( .A1(n11701), .A2(n11721), .ZN(n11704) );
  INV_X1 U14615 ( .A(n11709), .ZN(n18623) );
  AND2_X1 U14616 ( .A1(n11711), .A2(n11723), .ZN(n11716) );
  OAI211_X1 U14617 ( .C1(n18642), .C2(n19071), .A(n19256), .B(n18610), .ZN(
        n11720) );
  OAI21_X1 U14618 ( .B1(n11704), .B2(n11716), .A(n11720), .ZN(n14101) );
  AOI211_X1 U14619 ( .C1(n19036), .C2(n11706), .A(n11705), .B(n14101), .ZN(
        n11708) );
  NAND2_X1 U14620 ( .A1(n19216), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19105) );
  INV_X1 U14621 ( .A(n19251), .ZN(n19100) );
  AOI221_X4 U14622 ( .B1(n16743), .B2(n11708), .C1(n11707), .C2(n11708), .A(
        n19100), .ZN(n18575) );
  XNOR2_X1 U14623 ( .A(n16745), .B(n18610), .ZN(n19258) );
  NOR2_X1 U14624 ( .A1(n11709), .A2(n18632), .ZN(n19054) );
  NAND3_X1 U14625 ( .A1(n11710), .A2(n19054), .A3(n18627), .ZN(n14087) );
  NOR2_X1 U14626 ( .A1(n11711), .A2(n18619), .ZN(n19053) );
  NAND3_X1 U14627 ( .A1(n11712), .A2(n19053), .A3(n18632), .ZN(n14086) );
  NOR2_X1 U14628 ( .A1(n11713), .A2(n14086), .ZN(n11718) );
  NOR2_X2 U14629 ( .A1(n17838), .A2(n11716), .ZN(n16917) );
  NAND3_X1 U14630 ( .A1(n18616), .A2(n11720), .A3(n11719), .ZN(n11722) );
  AOI21_X1 U14631 ( .B1(n18619), .B2(n11722), .A(n11721), .ZN(n11728) );
  NAND2_X1 U14632 ( .A1(n11723), .A2(n11728), .ZN(n14096) );
  INV_X1 U14633 ( .A(n11724), .ZN(n11726) );
  INV_X1 U14634 ( .A(n16945), .ZN(n11725) );
  NAND3_X1 U14635 ( .A1(n11726), .A2(n16745), .A3(n11725), .ZN(n11727) );
  NAND2_X1 U14636 ( .A1(n11728), .A2(n11727), .ZN(n19052) );
  INV_X1 U14637 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11759) );
  NAND2_X1 U14638 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18266) );
  NOR2_X1 U14639 ( .A1(n18266), .A2(n18272), .ZN(n17915) );
  INV_X1 U14640 ( .A(n17915), .ZN(n18261) );
  NOR4_X1 U14641 ( .A1(n18325), .A2(n18262), .A3(n11759), .A4(n18261), .ZN(
        n11764) );
  NOR2_X1 U14642 ( .A1(n17913), .A2(n18266), .ZN(n18292) );
  INV_X1 U14643 ( .A(n18292), .ZN(n18290) );
  NOR2_X1 U14644 ( .A1(n18290), .A2(n18272), .ZN(n17903) );
  INV_X1 U14645 ( .A(n17903), .ZN(n11760) );
  INV_X1 U14646 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18556) );
  INV_X1 U14647 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18544) );
  NOR3_X1 U14648 ( .A1(n18529), .A2(n18556), .A3(n18544), .ZN(n18369) );
  NAND3_X1 U14649 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18369), .ZN(n18493) );
  INV_X1 U14650 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18502) );
  NAND2_X1 U14651 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18498) );
  OR2_X1 U14652 ( .A1(n18502), .A2(n18498), .ZN(n18370) );
  NOR2_X1 U14653 ( .A1(n18493), .A2(n18370), .ZN(n18414) );
  NAND2_X1 U14654 ( .A1(n18372), .A2(n18414), .ZN(n18391) );
  AOI21_X1 U14655 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18536) );
  INV_X1 U14656 ( .A(n18536), .ZN(n18559) );
  NAND2_X1 U14657 ( .A1(n18369), .A2(n18559), .ZN(n18494) );
  NOR2_X1 U14658 ( .A1(n18370), .A2(n18494), .ZN(n18416) );
  NAND2_X1 U14659 ( .A1(n18372), .A2(n18416), .ZN(n18328) );
  NOR2_X1 U14660 ( .A1(n17913), .A2(n18328), .ZN(n18308) );
  AOI21_X1 U14661 ( .B1(n18308), .B2(n17915), .A(n19068), .ZN(n18271) );
  AOI221_X1 U14662 ( .B1(n11760), .B2(n18593), .C1(n18391), .C2(n18593), .A(
        n18271), .ZN(n11729) );
  INV_X1 U14663 ( .A(n17999), .ZN(n18331) );
  INV_X1 U14664 ( .A(n18391), .ZN(n18373) );
  NAND3_X1 U14665 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18331), .A3(
        n18373), .ZN(n18263) );
  NAND2_X1 U14666 ( .A1(n19070), .A2(n18263), .ZN(n18355) );
  OAI211_X1 U14667 ( .C1(n19047), .C2(n11764), .A(n11729), .B(n18355), .ZN(
        n16288) );
  INV_X1 U14668 ( .A(n16288), .ZN(n11730) );
  OAI21_X1 U14669 ( .B1(n18475), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11730), .ZN(n16214) );
  AOI211_X1 U14670 ( .C1(n11731), .C2(n16285), .A(n18569), .B(n16214), .ZN(
        n11762) );
  INV_X1 U14671 ( .A(n18304), .ZN(n19035) );
  NAND2_X1 U14672 ( .A1(n16304), .A2(n17770), .ZN(n11737) );
  NAND2_X1 U14673 ( .A1(n17765), .A2(n11737), .ZN(n11735) );
  NAND2_X1 U14674 ( .A1(n11735), .A2(n11736), .ZN(n11744) );
  NOR2_X1 U14675 ( .A1(n17756), .A2(n11744), .ZN(n11733) );
  NAND2_X1 U14676 ( .A1(n11733), .A2(n11732), .ZN(n11747) );
  NOR2_X1 U14677 ( .A1(n17749), .A2(n11747), .ZN(n11751) );
  NAND2_X1 U14678 ( .A1(n11751), .A2(n16756), .ZN(n11752) );
  XOR2_X1 U14679 ( .A(n11733), .B(n11732), .Z(n11734) );
  XOR2_X1 U14680 ( .A(n18529), .B(n11734), .Z(n18200) );
  XOR2_X1 U14681 ( .A(n11736), .B(n11735), .Z(n11742) );
  AND2_X1 U14682 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11742), .ZN(
        n11743) );
  XOR2_X1 U14683 ( .A(n17765), .B(n11737), .Z(n11740) );
  NOR2_X1 U14684 ( .A1(n11740), .A2(n18567), .ZN(n11741) );
  NOR2_X1 U14685 ( .A1(n11550), .A2(n19232), .ZN(n11739) );
  NAND3_X1 U14686 ( .A1(n18254), .A2(n11550), .A3(n19232), .ZN(n11738) );
  OAI221_X1 U14687 ( .B1(n11739), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18254), .C2(n11550), .A(n11738), .ZN(n18234) );
  XOR2_X1 U14688 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11740), .Z(
        n18233) );
  NOR2_X1 U14689 ( .A1(n18234), .A2(n18233), .ZN(n18232) );
  NOR2_X1 U14690 ( .A1(n11741), .A2(n18232), .ZN(n18224) );
  XOR2_X1 U14691 ( .A(n18556), .B(n11742), .Z(n18223) );
  NOR2_X1 U14692 ( .A1(n18224), .A2(n18223), .ZN(n18222) );
  NOR2_X1 U14693 ( .A1(n11743), .A2(n18222), .ZN(n18209) );
  XNOR2_X1 U14694 ( .A(n11744), .B(n17756), .ZN(n18210) );
  NOR2_X1 U14695 ( .A1(n18209), .A2(n18210), .ZN(n11745) );
  NAND2_X1 U14696 ( .A1(n18209), .A2(n18210), .ZN(n18208) );
  OAI21_X1 U14697 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n11745), .A(
        n18208), .ZN(n18199) );
  XNOR2_X1 U14698 ( .A(n11747), .B(n17749), .ZN(n11749) );
  NOR2_X1 U14699 ( .A1(n11748), .A2(n11749), .ZN(n11750) );
  XNOR2_X1 U14700 ( .A(n11749), .B(n11748), .ZN(n18188) );
  INV_X1 U14701 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18522) );
  NOR2_X1 U14702 ( .A1(n11750), .A2(n18187), .ZN(n11753) );
  XOR2_X1 U14703 ( .A(n11751), .B(n17746), .Z(n11754) );
  NAND2_X1 U14704 ( .A1(n11753), .A2(n11754), .ZN(n18176) );
  NAND2_X1 U14705 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18176), .ZN(
        n11756) );
  NOR2_X1 U14706 ( .A1(n11752), .A2(n11756), .ZN(n11758) );
  INV_X1 U14707 ( .A(n11752), .ZN(n11757) );
  OR2_X1 U14708 ( .A1(n11754), .A2(n11753), .ZN(n18177) );
  OAI21_X1 U14709 ( .B1(n11757), .B2(n11756), .A(n18177), .ZN(n11755) );
  AOI21_X1 U14710 ( .B1(n11757), .B2(n11756), .A(n11755), .ZN(n18163) );
  NOR3_X1 U14711 ( .A1(n11760), .A2(n11759), .A3(n16211), .ZN(n16769) );
  NAND2_X1 U14712 ( .A1(n17937), .A2(n16769), .ZN(n16774) );
  NOR2_X1 U14713 ( .A1(n19041), .A2(n16756), .ZN(n18461) );
  NAND2_X1 U14714 ( .A1(n16769), .A2(n18402), .ZN(n16216) );
  AOI22_X1 U14715 ( .A1(n19035), .A2(n16774), .B1(n18461), .B2(n16216), .ZN(
        n11761) );
  AOI211_X1 U14716 ( .C1(n11762), .C2(n11761), .A(n18581), .B(n16211), .ZN(
        n11771) );
  NOR2_X1 U14717 ( .A1(n19041), .A2(n18592), .ZN(n18590) );
  NOR2_X1 U14718 ( .A1(n18155), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16212) );
  AND3_X1 U14719 ( .A1(n18590), .A2(n16212), .A3(n17891), .ZN(n11769) );
  AND2_X1 U14720 ( .A1(n18489), .A2(n17890), .ZN(n11763) );
  NAND2_X1 U14721 ( .A1(n17906), .A2(n11763), .ZN(n11767) );
  INV_X1 U14722 ( .A(n18461), .ZN(n18438) );
  OAI22_X1 U14723 ( .A1(n18462), .A2(n18304), .B1(n18460), .B2(n18438), .ZN(
        n18371) );
  AOI21_X1 U14724 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19070), .A(
        n18593), .ZN(n18560) );
  OAI22_X1 U14725 ( .A1(n19068), .A2(n18328), .B1(n18391), .B2(n18560), .ZN(
        n18291) );
  AOI21_X1 U14726 ( .B1(n18372), .B2(n18371), .A(n18291), .ZN(n18260) );
  NOR2_X1 U14727 ( .A1(n18260), .A2(n18592), .ZN(n18279) );
  NAND2_X1 U14728 ( .A1(n18331), .A2(n18279), .ZN(n18366) );
  NAND2_X1 U14729 ( .A1(n11764), .A2(n16211), .ZN(n17905) );
  INV_X2 U14730 ( .A(n18591), .ZN(n18570) );
  NAND2_X1 U14731 ( .A1(n18570), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17897) );
  OR2_X1 U14732 ( .A1(n11771), .A2(n11770), .ZN(P3_U2834) );
  NAND2_X1 U14733 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21064) );
  INV_X1 U14734 ( .A(n21064), .ZN(n20965) );
  OR2_X1 U14735 ( .A1(n11772), .A2(n20965), .ZN(n12841) );
  AND2_X1 U14736 ( .A1(n9836), .A2(n16253), .ZN(n11773) );
  NAND2_X1 U14737 ( .A1(n13260), .A2(n11773), .ZN(n16247) );
  OAI21_X1 U14738 ( .B1(n12841), .B2(n14158), .A(n16247), .ZN(n11774) );
  NAND2_X1 U14739 ( .A1(n16254), .A2(n11774), .ZN(n11784) );
  INV_X1 U14740 ( .A(n11775), .ZN(n11782) );
  NOR3_X1 U14741 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n11780) );
  OAI21_X1 U14742 ( .B1(n11781), .B2(n11780), .A(n11779), .ZN(n16245) );
  AND2_X1 U14743 ( .A1(n21064), .A2(n16245), .ZN(n12839) );
  NAND2_X1 U14744 ( .A1(n11782), .A2(n12839), .ZN(n11783) );
  NOR2_X1 U14745 ( .A1(n13412), .A2(n20294), .ZN(n11786) );
  NOR2_X1 U14746 ( .A1(n10397), .A2(n14198), .ZN(n11785) );
  NAND4_X1 U14747 ( .A1(n12861), .A2(n11786), .A3(n11785), .A4(n10421), .ZN(
        n13282) );
  OR2_X1 U14748 ( .A1(n13282), .A2(n12871), .ZN(n11787) );
  AND2_X1 U14749 ( .A1(n14865), .A2(n9896), .ZN(n11789) );
  NAND2_X1 U14750 ( .A1(n14168), .A2(n11789), .ZN(n11805) );
  NOR4_X1 U14751 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11793) );
  NOR4_X1 U14752 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11792) );
  NOR4_X1 U14753 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11791) );
  NOR4_X1 U14754 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11790) );
  AND4_X1 U14755 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11798) );
  NOR4_X1 U14756 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11796) );
  NOR4_X1 U14757 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11795) );
  NOR4_X1 U14758 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11794) );
  INV_X1 U14759 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20983) );
  AND4_X1 U14760 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n20983), .ZN(
        n11797) );
  NAND2_X1 U14761 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  AND2_X2 U14762 ( .A1(n11799), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n13623)
         );
  AOI22_X1 U14763 ( .A1(n9632), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14847), .ZN(n11800) );
  INV_X1 U14764 ( .A(n11800), .ZN(n11803) );
  INV_X1 U14765 ( .A(n13623), .ZN(n13386) );
  NOR2_X1 U14766 ( .A1(n12862), .A2(n13386), .ZN(n11801) );
  NAND2_X1 U14767 ( .A1(n14865), .A2(n11801), .ZN(n14824) );
  INV_X1 U14768 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16808) );
  NOR2_X1 U14769 ( .A1(n14824), .A2(n16808), .ZN(n11802) );
  NOR2_X1 U14770 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  NAND2_X1 U14771 ( .A1(n11805), .A2(n11804), .ZN(P1_U2873) );
  AND2_X4 U14772 ( .A1(n15994), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12025) );
  AND3_X4 U14773 ( .A1(n12397), .A2(n16709), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U14774 ( .A1(n12025), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14775 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11806) );
  AND3_X1 U14776 ( .A1(n11807), .A2(n11806), .A3(n12026), .ZN(n11811) );
  AND2_X4 U14777 ( .A1(n15978), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12018) );
  INV_X1 U14778 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11808) );
  AND3_X2 U14779 ( .A1(n11808), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14780 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9642), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14781 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11809) );
  NAND3_X1 U14782 ( .A1(n11811), .A2(n11810), .A3(n11809), .ZN(n11818) );
  AOI22_X1 U14783 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9643), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14784 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14785 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11815) );
  NAND3_X1 U14786 ( .A1(n9726), .A2(n11816), .A3(n11815), .ZN(n11817) );
  AOI22_X1 U14787 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14788 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14789 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14790 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11819) );
  NAND4_X1 U14791 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11823) );
  AOI22_X1 U14792 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14793 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14794 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9642), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14795 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U14796 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11829) );
  NAND2_X1 U14797 ( .A1(n11844), .A2(n11830), .ZN(n11831) );
  AOI22_X1 U14798 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14799 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14800 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14801 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U14802 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11836) );
  NAND2_X1 U14803 ( .A1(n11836), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11843) );
  AOI22_X1 U14804 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14805 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14806 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9642), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14807 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9643), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11837) );
  NAND4_X1 U14808 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11841) );
  NAND2_X1 U14809 ( .A1(n11841), .A2(n12026), .ZN(n11842) );
  NAND2_X1 U14810 ( .A1(n12452), .A2(n13155), .ZN(n12451) );
  NAND2_X1 U14811 ( .A1(n11908), .A2(n19646), .ZN(n12449) );
  AOI22_X1 U14812 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9642), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14813 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14814 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14815 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12383), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14816 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  NAND2_X1 U14817 ( .A1(n11849), .A2(n12026), .ZN(n11856) );
  AOI22_X1 U14818 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14819 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14820 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11850) );
  NAND4_X1 U14821 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11854) );
  NAND2_X1 U14822 ( .A1(n11854), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11855) );
  AOI22_X1 U14823 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14824 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9661), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14825 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14826 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9643), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14827 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14828 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14829 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14830 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14831 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9661), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14832 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9641), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11867) );
  NAND2_X1 U14833 ( .A1(n11868), .A2(n11867), .ZN(n11872) );
  AOI22_X1 U14834 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14835 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U14836 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  AOI22_X1 U14837 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14838 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14839 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14840 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9638), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U14841 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  NAND2_X1 U14842 ( .A1(n11877), .A2(n12026), .ZN(n11878) );
  AOI22_X1 U14843 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14844 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11880) );
  NAND4_X1 U14845 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11884) );
  AOI22_X1 U14846 ( .A1(n12020), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14847 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14848 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14849 ( .A1(n11824), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U14850 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11889) );
  NAND2_X2 U14851 ( .A1(n11891), .A2(n11890), .ZN(n16039) );
  AOI22_X1 U14852 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14853 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14854 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11894) );
  NAND2_X1 U14855 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11897) );
  AOI22_X1 U14856 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11824), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14857 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14858 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9640), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11900) );
  NAND4_X1 U14859 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11904) );
  NAND2_X2 U14860 ( .A1(n11905), .A2(n11904), .ZN(n11915) );
  INV_X2 U14861 ( .A(n11915), .ZN(n13157) );
  NAND4_X1 U14862 ( .A1(n11906), .A2(n13157), .A3(n11919), .A4(n13155), .ZN(
        n11907) );
  INV_X1 U14863 ( .A(n11924), .ZN(n13029) );
  MUX2_X1 U14864 ( .A(n13881), .B(n11919), .S(n19646), .Z(n11909) );
  NAND3_X1 U14865 ( .A1(n11934), .A2(n11909), .A3(n10216), .ZN(n11910) );
  NAND2_X1 U14866 ( .A1(n13152), .A2(n9670), .ZN(n11912) );
  NAND2_X1 U14867 ( .A1(n11913), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11923) );
  NOR2_X1 U14868 ( .A1(n11916), .A2(n12453), .ZN(n11917) );
  NAND2_X1 U14869 ( .A1(n11920), .A2(n11917), .ZN(n16696) );
  NOR2_X1 U14870 ( .A1(n12298), .A2(n13157), .ZN(n11918) );
  NAND2_X1 U14871 ( .A1(n16696), .A2(n11918), .ZN(n11922) );
  NAND2_X1 U14872 ( .A1(n11921), .A2(n11920), .ZN(n11925) );
  NAND2_X1 U14873 ( .A1(n11922), .A2(n11925), .ZN(n12676) );
  NAND2_X1 U14874 ( .A1(n16039), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U14875 ( .A1(n11923), .A2(n11950), .ZN(n11955) );
  NAND2_X1 U14876 ( .A1(n11955), .A2(n15984), .ZN(n11932) );
  NAND2_X1 U14877 ( .A1(n11924), .A2(n9670), .ZN(n12448) );
  NAND2_X1 U14878 ( .A1(n12472), .A2(n10214), .ZN(n11929) );
  NAND2_X1 U14879 ( .A1(n20154), .A2(n16735), .ZN(n16729) );
  NOR2_X1 U14880 ( .A1(n16729), .A2(n20272), .ZN(n11930) );
  AOI21_X1 U14881 ( .B1(n15993), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11930), 
        .ZN(n11931) );
  NAND2_X1 U14882 ( .A1(n11932), .A2(n11931), .ZN(n11942) );
  INV_X1 U14883 ( .A(n11942), .ZN(n11941) );
  CLKBUF_X3 U14884 ( .A(n11830), .Z(n14328) );
  NAND2_X1 U14885 ( .A1(n12435), .A2(n13081), .ZN(n12467) );
  AND2_X1 U14886 ( .A1(n19659), .A2(n19646), .ZN(n11935) );
  NAND2_X1 U14887 ( .A1(n11971), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11939) );
  INV_X1 U14888 ( .A(n11943), .ZN(n11940) );
  NAND2_X1 U14889 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  INV_X1 U14890 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U14891 ( .A1(n13154), .A2(n13152), .ZN(n11946) );
  NAND2_X1 U14892 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  NAND2_X1 U14893 ( .A1(n11947), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14894 ( .A1(n11971), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U14895 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11948) );
  AND2_X1 U14896 ( .A1(n16729), .A2(n11948), .ZN(n11949) );
  NAND2_X1 U14897 ( .A1(n12755), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11953) );
  OAI211_X1 U14898 ( .C1(n11970), .C2(n13085), .A(n11954), .B(n11953), .ZN(
        n12006) );
  NAND2_X1 U14899 ( .A1(n12696), .A2(n16709), .ZN(n11956) );
  NAND2_X1 U14900 ( .A1(n11955), .A2(n11956), .ZN(n11963) );
  NAND2_X1 U14901 ( .A1(n11956), .A2(n13178), .ZN(n11958) );
  INV_X1 U14902 ( .A(n11957), .ZN(n14051) );
  NAND2_X1 U14903 ( .A1(n11958), .A2(n14051), .ZN(n11961) );
  NOR2_X1 U14904 ( .A1(n13156), .A2(n16735), .ZN(n11960) );
  NOR2_X1 U14905 ( .A1(n16729), .A2(n20281), .ZN(n11959) );
  AOI21_X1 U14906 ( .B1(n11961), .B2(n11960), .A(n11959), .ZN(n11962) );
  NAND2_X1 U14907 ( .A1(n11963), .A2(n11962), .ZN(n12005) );
  INV_X1 U14908 ( .A(n11968), .ZN(n11966) );
  OAI21_X1 U14909 ( .B1(n20262), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20154), 
        .ZN(n11964) );
  NAND2_X1 U14910 ( .A1(n11966), .A2(n11965), .ZN(n11969) );
  NAND2_X1 U14911 ( .A1(n11968), .A2(n11967), .ZN(n11974) );
  INV_X1 U14912 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U14913 ( .A1(n14506), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11972) );
  OAI211_X2 U14914 ( .C1(n14510), .C2(n13760), .A(n11973), .B(n11972), .ZN(
        n11990) );
  INV_X1 U14915 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13777) );
  AOI22_X1 U14916 ( .A1(n9648), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U14917 ( .A1(n14506), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11975) );
  OAI211_X1 U14918 ( .C1(n14510), .C2(n13777), .A(n11976), .B(n11975), .ZN(
        n11980) );
  NAND2_X1 U14919 ( .A1(n11955), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11978) );
  OR2_X1 U14920 ( .A1(n16729), .A2(n20254), .ZN(n11977) );
  NAND2_X1 U14921 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  NAND2_X1 U14922 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  NAND2_X1 U14923 ( .A1(n9675), .A2(n13086), .ZN(n11986) );
  NAND2_X1 U14924 ( .A1(n13881), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11982) );
  NOR2_X2 U14925 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20243) );
  NOR2_X1 U14926 ( .A1(n20262), .A2(n20272), .ZN(n20047) );
  NAND2_X1 U14927 ( .A1(n20047), .A2(n20254), .ZN(n19835) );
  INV_X1 U14928 ( .A(n19835), .ZN(n11983) );
  NAND2_X1 U14929 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20047), .ZN(
        n19624) );
  NAND2_X1 U14930 ( .A1(n19624), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U14931 ( .A1(n19873), .A2(n11984), .ZN(n19986) );
  AOI22_X1 U14932 ( .A1(n12008), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20243), .B2(n19986), .ZN(n11985) );
  NAND2_X1 U14933 ( .A1(n11987), .A2(n11844), .ZN(n13443) );
  INV_X1 U14934 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12279) );
  NOR2_X1 U14935 ( .A1(n13443), .A2(n12279), .ZN(n11988) );
  NAND2_X1 U14936 ( .A1(n12016), .A2(n11988), .ZN(n13885) );
  XNOR2_X2 U14937 ( .A(n11991), .B(n11990), .ZN(n13702) );
  NAND2_X1 U14938 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19949) );
  NAND2_X1 U14939 ( .A1(n19949), .A2(n20262), .ZN(n11992) );
  AND2_X1 U14940 ( .A1(n11992), .A2(n19624), .ZN(n16030) );
  AND2_X1 U14941 ( .A1(n16030), .A2(n20243), .ZN(n19987) );
  AOI21_X1 U14942 ( .B1(n12008), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19987), .ZN(n11993) );
  INV_X1 U14943 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12262) );
  NOR2_X1 U14944 ( .A1(n13443), .A2(n12262), .ZN(n11995) );
  INV_X1 U14945 ( .A(n11999), .ZN(n13694) );
  INV_X1 U14946 ( .A(n12007), .ZN(n12000) );
  NAND2_X1 U14947 ( .A1(n13694), .A2(n12000), .ZN(n12001) );
  NAND2_X1 U14948 ( .A1(n12008), .A2(n15984), .ZN(n12003) );
  NAND2_X1 U14949 ( .A1(n20272), .A2(n20281), .ZN(n12002) );
  AND2_X1 U14950 ( .A1(n12002), .A2(n19949), .ZN(n16029) );
  NAND2_X1 U14951 ( .A1(n16029), .A2(n20243), .ZN(n19700) );
  NAND2_X1 U14952 ( .A1(n12003), .A2(n19700), .ZN(n12004) );
  OR2_X1 U14953 ( .A1(n12006), .A2(n12005), .ZN(n13689) );
  AOI22_X1 U14954 ( .A1(n12008), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20243), .B2(n20281), .ZN(n12009) );
  INV_X1 U14955 ( .A(n13443), .ZN(n12296) );
  NAND2_X1 U14956 ( .A1(n12296), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12011) );
  XNOR2_X1 U14957 ( .A(n14054), .B(n12011), .ZN(n13097) );
  NAND2_X1 U14958 ( .A1(n13096), .A2(n13097), .ZN(n13098) );
  INV_X1 U14959 ( .A(n14054), .ZN(n12012) );
  NAND2_X1 U14960 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  NAND2_X1 U14961 ( .A1(n13098), .A2(n12013), .ZN(n13276) );
  INV_X1 U14962 ( .A(n13276), .ZN(n12014) );
  NAND2_X1 U14963 ( .A1(n12016), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12017) );
  INV_X1 U14964 ( .A(n12231), .ZN(n12349) );
  AOI22_X1 U14965 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12150), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U14966 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12023) );
  AND2_X2 U14967 ( .A1(n9645), .A2(n12026), .ZN(n12580) );
  AOI22_X1 U14968 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12580), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12022) );
  INV_X1 U14969 ( .A(n12020), .ZN(n12308) );
  AND2_X2 U14970 ( .A1(n12020), .A2(n12026), .ZN(n12581) );
  AND2_X2 U14971 ( .A1(n9661), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12115) );
  AOI22_X1 U14972 ( .A1(n12581), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U14973 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12033) );
  AOI22_X1 U14974 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12031) );
  AND2_X2 U14975 ( .A1(n9638), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12051) );
  AOI22_X1 U14976 ( .A1(n12142), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12030) );
  AND2_X2 U14977 ( .A1(n11899), .A2(n12026), .ZN(n12137) );
  AOI22_X1 U14979 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12029) );
  NAND3_X1 U14980 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15984), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13031) );
  INV_X1 U14981 ( .A(n13031), .ZN(n12027) );
  AND2_X2 U14982 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12027), .ZN(
        n12586) );
  AOI22_X1 U14983 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12586), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U14984 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12032) );
  AND2_X1 U14985 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13514) );
  NAND4_X1 U14986 ( .A1(n19479), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A4(n13514), .ZN(n12034) );
  NOR2_X1 U14987 ( .A1(n13443), .A2(n12034), .ZN(n12035) );
  AOI22_X1 U14988 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U14989 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U14990 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U14991 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12037) );
  NAND4_X1 U14992 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12046) );
  AOI22_X1 U14993 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U14994 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U14995 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U14996 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12586), .ZN(n12041) );
  NAND4_X1 U14997 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12045) );
  NOR2_X1 U14998 ( .A1(n12046), .A2(n12045), .ZN(n13485) );
  AOI22_X1 U14999 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12569), .B1(
        n12579), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15000 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15001 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15002 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15003 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12057) );
  AOI22_X1 U15004 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12073), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15005 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12137), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15006 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12072), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15007 ( .A1(n12051), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12586), .ZN(n12052) );
  NAND4_X1 U15008 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(
        n12056) );
  AOI22_X1 U15009 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15010 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15011 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15012 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12058) );
  NAND4_X1 U15013 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12058), .ZN(
        n12067) );
  AOI22_X1 U15014 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15015 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15016 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15017 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12586), .ZN(n12062) );
  NAND4_X1 U15018 ( .A1(n12065), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n12066) );
  NOR2_X1 U15019 ( .A1(n12067), .A2(n12066), .ZN(n13618) );
  AOI22_X1 U15020 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15021 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15022 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15023 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15024 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12079) );
  AOI22_X1 U15025 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12142), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15026 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15027 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12072), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15028 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12586), .ZN(n12074) );
  NAND4_X1 U15029 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12078) );
  NOR2_X1 U15030 ( .A1(n12079), .A2(n12078), .ZN(n19472) );
  AOI22_X1 U15031 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15032 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15033 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15034 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15035 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12093) );
  AOI22_X1 U15036 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12091) );
  INV_X1 U15037 ( .A(n12098), .ZN(n12086) );
  INV_X1 U15038 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12085) );
  INV_X1 U15039 ( .A(n12478), .ZN(n12084) );
  OAI22_X1 U15040 ( .A1(n12086), .A2(n12085), .B1(n12084), .B2(n12279), .ZN(
        n12087) );
  INV_X1 U15041 ( .A(n12087), .ZN(n12090) );
  AOI22_X1 U15042 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15043 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12586), .ZN(n12088) );
  NAND4_X1 U15044 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12092) );
  OR2_X1 U15045 ( .A1(n12093), .A2(n12092), .ZN(n15308) );
  AOI22_X1 U15046 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15047 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15048 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15049 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12094) );
  NAND4_X1 U15050 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12104) );
  AOI22_X1 U15051 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15052 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15053 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15054 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12586), .ZN(n12099) );
  NAND4_X1 U15055 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  OR2_X1 U15056 ( .A1(n12104), .A2(n12103), .ZN(n16597) );
  AOI22_X1 U15057 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15058 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15059 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15060 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12105) );
  NAND4_X1 U15061 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12114) );
  AOI22_X1 U15062 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15063 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15064 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15065 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12586), .ZN(n12109) );
  NAND4_X1 U15066 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(
        n12113) );
  OR2_X1 U15067 ( .A1(n12114), .A2(n12113), .ZN(n13976) );
  INV_X1 U15068 ( .A(n13976), .ZN(n12136) );
  AOI22_X1 U15069 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15070 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15071 ( .A1(n12580), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15072 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15073 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  AOI22_X1 U15074 ( .A1(n12167), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15075 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15076 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15077 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12586), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15078 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  NOR2_X1 U15079 ( .A1(n12125), .A2(n12124), .ZN(n19463) );
  AOI22_X1 U15080 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12150), .B1(
        n12579), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15081 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15082 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12580), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15083 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12581), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15084 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12135) );
  AOI22_X1 U15085 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12167), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15086 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15087 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12072), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15088 ( .A1(n12142), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12586), .ZN(n12130) );
  NAND4_X1 U15089 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12134) );
  NOR2_X1 U15090 ( .A1(n12135), .A2(n12134), .ZN(n14020) );
  OR2_X1 U15091 ( .A1(n19463), .A2(n14020), .ZN(n13972) );
  OR2_X1 U15092 ( .A1(n12136), .A2(n13972), .ZN(n12149) );
  AOI22_X1 U15093 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15094 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15095 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15096 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15097 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12148) );
  AOI22_X1 U15098 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15099 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15100 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15101 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12586), .ZN(n12143) );
  NAND4_X1 U15102 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12147) );
  NOR2_X1 U15103 ( .A1(n12148), .A2(n12147), .ZN(n13984) );
  NOR2_X1 U15104 ( .A1(n12149), .A2(n13984), .ZN(n13974) );
  AND2_X1 U15105 ( .A1(n16597), .A2(n13974), .ZN(n12161) );
  AOI22_X1 U15106 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15107 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15108 ( .A1(n12580), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15109 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U15110 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12160) );
  AOI22_X1 U15111 ( .A1(n12167), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15112 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15113 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15114 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12586), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12155) );
  NAND4_X1 U15115 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12159) );
  AND2_X1 U15116 ( .A1(n12161), .A2(n13973), .ZN(n15306) );
  AOI22_X1 U15117 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15118 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15119 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15120 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15121 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12173) );
  AOI22_X1 U15122 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15123 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15124 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15125 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12586), .ZN(n12168) );
  NAND4_X1 U15126 ( .A1(n12171), .A2(n12170), .A3(n12169), .A4(n12168), .ZN(
        n12172) );
  NOR2_X1 U15127 ( .A1(n12173), .A2(n12172), .ZN(n16591) );
  AOI22_X1 U15128 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15129 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15130 ( .A1(n12580), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15131 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15132 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12186) );
  AOI22_X1 U15133 ( .A1(n12167), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15134 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15135 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12182) );
  INV_X1 U15136 ( .A(n12586), .ZN(n12179) );
  INV_X1 U15137 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12178) );
  NOR2_X1 U15138 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  AOI21_X1 U15139 ( .B1(n12073), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n12180), .ZN(n12181) );
  NAND4_X1 U15140 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12185) );
  OR2_X1 U15141 ( .A1(n12186), .A2(n12185), .ZN(n15301) );
  AOI22_X1 U15142 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15143 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15144 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15145 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15146 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12196) );
  AOI22_X1 U15147 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15148 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15149 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15150 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12586), .ZN(n12191) );
  NAND4_X1 U15151 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  NOR2_X1 U15152 ( .A1(n12196), .A2(n12195), .ZN(n16588) );
  INV_X1 U15153 ( .A(n11899), .ZN(n12304) );
  INV_X1 U15154 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12197) );
  INV_X1 U15155 ( .A(n12383), .ZN(n12355) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16057) );
  OAI22_X1 U15157 ( .A1(n12304), .A2(n12197), .B1(n12355), .B2(n16057), .ZN(
        n12201) );
  INV_X1 U15158 ( .A(n9638), .ZN(n12361) );
  INV_X1 U15159 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12199) );
  INV_X1 U15160 ( .A(n11824), .ZN(n12359) );
  INV_X1 U15161 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12198) );
  OAI22_X1 U15162 ( .A1(n12361), .A2(n12199), .B1(n12359), .B2(n12198), .ZN(
        n12200) );
  NOR2_X1 U15163 ( .A1(n12201), .A2(n12200), .ZN(n12204) );
  AOI22_X1 U15164 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9635), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12203) );
  INV_X1 U15165 ( .A(n12308), .ZN(n16013) );
  AOI22_X1 U15166 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12202) );
  XNOR2_X1 U15167 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U15168 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12378), .ZN(
        n12213) );
  INV_X1 U15169 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16098) );
  INV_X1 U15170 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20022) );
  OAI22_X1 U15171 ( .A1(n12304), .A2(n16098), .B1(n12361), .B2(n20022), .ZN(
        n12208) );
  INV_X1 U15172 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12206) );
  INV_X1 U15173 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12205) );
  OAI22_X1 U15174 ( .A1(n12355), .A2(n12206), .B1(n12359), .B2(n12205), .ZN(
        n12207) );
  NOR2_X1 U15175 ( .A1(n12208), .A2(n12207), .ZN(n12211) );
  AOI22_X1 U15176 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9635), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15177 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15178 ( .A1(n12211), .A2(n12384), .A3(n12210), .A4(n12209), .ZN(
        n12212) );
  AND2_X1 U15179 ( .A1(n12213), .A2(n12212), .ZN(n12245) );
  NAND2_X1 U15180 ( .A1(n16070), .A2(n12245), .ZN(n12224) );
  AOI22_X1 U15181 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15182 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12580), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15183 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12581), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15184 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U15185 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12223) );
  AOI22_X1 U15186 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12478), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15187 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15188 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12072), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15189 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12586), .ZN(n12218) );
  NAND4_X1 U15190 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12222) );
  OR2_X1 U15191 ( .A1(n12223), .A2(n12222), .ZN(n12242) );
  XNOR2_X1 U15192 ( .A(n12224), .B(n12242), .ZN(n12248) );
  NAND2_X1 U15193 ( .A1(n12298), .A2(n12245), .ZN(n15295) );
  NOR2_X2 U15194 ( .A1(n15296), .A2(n15295), .ZN(n15294) );
  INV_X1 U15195 ( .A(n12018), .ZN(n12357) );
  INV_X1 U15196 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12227) );
  INV_X1 U15197 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12226) );
  OAI22_X1 U15198 ( .A1(n12357), .A2(n12227), .B1(n12359), .B2(n12226), .ZN(
        n12230) );
  INV_X1 U15199 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12228) );
  INV_X1 U15200 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13741) );
  OAI22_X1 U15201 ( .A1(n12361), .A2(n12228), .B1(n12355), .B2(n13741), .ZN(
        n12229) );
  NOR2_X1 U15202 ( .A1(n12230), .A2(n12229), .ZN(n12234) );
  AOI22_X1 U15203 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15204 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U15205 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12378), .ZN(
        n12241) );
  INV_X1 U15206 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16076) );
  INV_X1 U15207 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16089) );
  OAI22_X1 U15208 ( .A1(n12357), .A2(n16076), .B1(n12359), .B2(n16089), .ZN(
        n12236) );
  INV_X1 U15209 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13740) );
  INV_X1 U15210 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13742) );
  OAI22_X1 U15211 ( .A1(n12361), .A2(n13740), .B1(n12355), .B2(n13742), .ZN(
        n12235) );
  NOR2_X1 U15212 ( .A1(n12236), .A2(n12235), .ZN(n12239) );
  AOI22_X1 U15213 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15214 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12237) );
  NAND4_X1 U15215 ( .A1(n12239), .A2(n12384), .A3(n12238), .A4(n12237), .ZN(
        n12240) );
  NAND2_X1 U15216 ( .A1(n12241), .A2(n12240), .ZN(n12250) );
  NAND2_X1 U15217 ( .A1(n12242), .A2(n12245), .ZN(n12251) );
  XOR2_X1 U15218 ( .A(n12250), .B(n12251), .Z(n12243) );
  NAND2_X1 U15219 ( .A1(n12243), .A2(n12296), .ZN(n15281) );
  INV_X1 U15220 ( .A(n12250), .ZN(n12244) );
  NAND2_X1 U15221 ( .A1(n12298), .A2(n12244), .ZN(n15284) );
  INV_X1 U15222 ( .A(n12245), .ZN(n12246) );
  NOR2_X1 U15223 ( .A1(n15284), .A2(n12246), .ZN(n12247) );
  NOR2_X1 U15224 ( .A1(n12251), .A2(n12250), .ZN(n12272) );
  INV_X1 U15225 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12253) );
  INV_X1 U15226 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12252) );
  OAI22_X1 U15227 ( .A1(n12349), .A2(n12253), .B1(n12304), .B2(n12252), .ZN(
        n12257) );
  INV_X1 U15228 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12255) );
  INV_X1 U15229 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12254) );
  OAI22_X1 U15230 ( .A1(n12308), .A2(n12255), .B1(n9662), .B2(n12254), .ZN(
        n12256) );
  NOR2_X1 U15231 ( .A1(n12257), .A2(n12256), .ZN(n12260) );
  AOI22_X1 U15232 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15233 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15234 ( .A1(n12260), .A2(n12384), .A3(n12259), .A4(n12258), .ZN(
        n12271) );
  INV_X1 U15235 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12261) );
  OAI22_X1 U15236 ( .A1(n12357), .A2(n12262), .B1(n12359), .B2(n12261), .ZN(
        n12266) );
  INV_X1 U15237 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12264) );
  INV_X1 U15238 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12263) );
  OAI22_X1 U15239 ( .A1(n12361), .A2(n12264), .B1(n12355), .B2(n12263), .ZN(
        n12265) );
  NOR2_X1 U15240 ( .A1(n12266), .A2(n12265), .ZN(n12269) );
  AOI22_X1 U15241 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15242 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15243 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12378), .ZN(
        n12270) );
  AND2_X1 U15244 ( .A1(n12271), .A2(n12270), .ZN(n12273) );
  NAND2_X1 U15245 ( .A1(n12272), .A2(n12273), .ZN(n12325) );
  OAI211_X1 U15246 ( .C1(n12272), .C2(n12273), .A(n12296), .B(n12325), .ZN(
        n12275) );
  INV_X1 U15247 ( .A(n12273), .ZN(n12274) );
  NOR2_X1 U15248 ( .A1(n16070), .A2(n12274), .ZN(n15273) );
  NAND2_X1 U15249 ( .A1(n15274), .A2(n15273), .ZN(n15272) );
  INV_X1 U15250 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12278) );
  OAI22_X1 U15251 ( .A1(n12357), .A2(n12279), .B1(n12359), .B2(n12278), .ZN(
        n12282) );
  INV_X1 U15252 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12280) );
  INV_X1 U15253 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13711) );
  OAI22_X1 U15254 ( .A1(n12361), .A2(n12280), .B1(n12355), .B2(n13711), .ZN(
        n12281) );
  NOR2_X1 U15255 ( .A1(n12282), .A2(n12281), .ZN(n12285) );
  AOI22_X1 U15256 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15257 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12283) );
  NAND4_X1 U15258 ( .A1(n12285), .A2(n12284), .A3(n12283), .A4(n12378), .ZN(
        n12295) );
  INV_X1 U15259 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12287) );
  INV_X1 U15260 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12286) );
  OAI22_X1 U15261 ( .A1(n12357), .A2(n12287), .B1(n12359), .B2(n12286), .ZN(
        n12290) );
  INV_X1 U15262 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12288) );
  INV_X1 U15263 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13724) );
  OAI22_X1 U15264 ( .A1(n12361), .A2(n12288), .B1(n12355), .B2(n13724), .ZN(
        n12289) );
  NOR2_X1 U15265 ( .A1(n12290), .A2(n12289), .ZN(n12293) );
  AOI22_X1 U15266 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15267 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U15268 ( .A1(n12293), .A2(n12384), .A3(n12292), .A4(n12291), .ZN(
        n12294) );
  AND2_X1 U15269 ( .A1(n12295), .A2(n12294), .ZN(n12299) );
  XNOR2_X1 U15270 ( .A(n12325), .B(n12299), .ZN(n12297) );
  NAND2_X1 U15271 ( .A1(n12297), .A2(n12296), .ZN(n12301) );
  XNOR2_X1 U15272 ( .A(n12300), .B(n12301), .ZN(n15266) );
  INV_X1 U15273 ( .A(n12299), .ZN(n12324) );
  NOR2_X1 U15274 ( .A1(n16070), .A2(n12324), .ZN(n15265) );
  INV_X1 U15275 ( .A(n12300), .ZN(n12302) );
  NAND2_X1 U15276 ( .A1(n15264), .A2(n10217), .ZN(n12328) );
  INV_X1 U15277 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12305) );
  INV_X1 U15278 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12303) );
  OAI22_X1 U15279 ( .A1(n12349), .A2(n12305), .B1(n12304), .B2(n12303), .ZN(
        n12310) );
  INV_X1 U15280 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12307) );
  INV_X1 U15281 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12306) );
  OAI22_X1 U15282 ( .A1(n12308), .A2(n12307), .B1(n9662), .B2(n12306), .ZN(
        n12309) );
  NOR2_X1 U15283 ( .A1(n12310), .A2(n12309), .ZN(n12313) );
  AOI22_X1 U15284 ( .A1(n9638), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15285 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9642), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15286 ( .A1(n12313), .A2(n12384), .A3(n12312), .A4(n12311), .ZN(
        n12323) );
  INV_X1 U15287 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13442) );
  INV_X1 U15288 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12314) );
  OAI22_X1 U15289 ( .A1(n12357), .A2(n13442), .B1(n12359), .B2(n12314), .ZN(
        n12318) );
  INV_X1 U15290 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12316) );
  INV_X1 U15291 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12315) );
  OAI22_X1 U15292 ( .A1(n12361), .A2(n12316), .B1(n12355), .B2(n12315), .ZN(
        n12317) );
  NOR2_X1 U15293 ( .A1(n12318), .A2(n12317), .ZN(n12321) );
  AOI22_X1 U15294 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15295 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15296 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12378), .ZN(
        n12322) );
  NAND2_X1 U15297 ( .A1(n12323), .A2(n12322), .ZN(n12330) );
  OR2_X1 U15298 ( .A1(n12325), .A2(n12324), .ZN(n12326) );
  NOR2_X1 U15299 ( .A1(n12326), .A2(n12330), .ZN(n12369) );
  OAI21_X1 U15300 ( .B1(n12328), .B2(n12327), .A(n15253), .ZN(n12329) );
  INV_X1 U15301 ( .A(n12329), .ZN(n15261) );
  NOR2_X1 U15302 ( .A1(n16070), .A2(n12330), .ZN(n15260) );
  NAND2_X1 U15303 ( .A1(n15261), .A2(n15260), .ZN(n15259) );
  INV_X1 U15304 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13521) );
  INV_X1 U15305 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12331) );
  OAI22_X1 U15306 ( .A1(n12357), .A2(n13521), .B1(n12359), .B2(n12331), .ZN(
        n12334) );
  INV_X1 U15307 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12332) );
  INV_X1 U15308 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14247) );
  OAI22_X1 U15309 ( .A1(n12361), .A2(n12332), .B1(n12355), .B2(n14247), .ZN(
        n12333) );
  NOR2_X1 U15310 ( .A1(n12334), .A2(n12333), .ZN(n12337) );
  AOI22_X1 U15311 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15312 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12335) );
  NAND4_X1 U15313 ( .A1(n12337), .A2(n12336), .A3(n12335), .A4(n12378), .ZN(
        n12346) );
  INV_X1 U15314 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12338) );
  INV_X1 U15315 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14252) );
  OAI22_X1 U15316 ( .A1(n12357), .A2(n12338), .B1(n12359), .B2(n14252), .ZN(
        n12341) );
  INV_X1 U15317 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12339) );
  INV_X1 U15318 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14250) );
  OAI22_X1 U15319 ( .A1(n12361), .A2(n12339), .B1(n12355), .B2(n14250), .ZN(
        n12340) );
  NOR2_X1 U15320 ( .A1(n12341), .A2(n12340), .ZN(n12344) );
  AOI22_X1 U15321 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15322 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12342) );
  NAND4_X1 U15323 ( .A1(n12344), .A2(n12384), .A3(n12343), .A4(n12342), .ZN(
        n12345) );
  NAND2_X1 U15324 ( .A1(n12346), .A2(n12345), .ZN(n12370) );
  AOI21_X1 U15325 ( .B1(n15259), .B2(n15253), .A(n12370), .ZN(n15248) );
  INV_X1 U15326 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12348) );
  INV_X1 U15327 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12347) );
  OAI22_X1 U15328 ( .A1(n12349), .A2(n12348), .B1(n12359), .B2(n12347), .ZN(
        n12351) );
  INV_X1 U15329 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16113) );
  INV_X1 U15330 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14293) );
  OAI22_X1 U15331 ( .A1(n12361), .A2(n16113), .B1(n12355), .B2(n14293), .ZN(
        n12350) );
  NOR2_X1 U15332 ( .A1(n12351), .A2(n12350), .ZN(n12354) );
  AOI22_X1 U15333 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15334 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15335 ( .A1(n12354), .A2(n12384), .A3(n12353), .A4(n12352), .ZN(
        n12368) );
  INV_X1 U15336 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12356) );
  INV_X1 U15337 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14294) );
  OAI22_X1 U15338 ( .A1(n12357), .A2(n12356), .B1(n12355), .B2(n14294), .ZN(
        n12363) );
  INV_X1 U15339 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12360) );
  INV_X1 U15340 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12358) );
  OAI22_X1 U15341 ( .A1(n12361), .A2(n12360), .B1(n12359), .B2(n12358), .ZN(
        n12362) );
  NOR2_X1 U15342 ( .A1(n12363), .A2(n12362), .ZN(n12366) );
  AOI22_X1 U15343 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15344 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U15345 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12378), .ZN(
        n12367) );
  NAND2_X1 U15346 ( .A1(n12368), .A2(n12367), .ZN(n12373) );
  INV_X1 U15347 ( .A(n12369), .ZN(n15252) );
  INV_X1 U15348 ( .A(n12370), .ZN(n15254) );
  NAND2_X1 U15349 ( .A1(n16070), .A2(n15254), .ZN(n12371) );
  OR2_X1 U15350 ( .A1(n15252), .A2(n12371), .ZN(n12372) );
  NOR2_X1 U15351 ( .A1(n12372), .A2(n12373), .ZN(n12374) );
  AOI21_X1 U15352 ( .B1(n12373), .B2(n12372), .A(n12374), .ZN(n15247) );
  NAND2_X1 U15353 ( .A1(n15248), .A2(n15247), .ZN(n15249) );
  INV_X1 U15354 ( .A(n12374), .ZN(n12375) );
  NAND2_X1 U15355 ( .A1(n15249), .A2(n12375), .ZN(n12392) );
  AOI22_X1 U15356 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15357 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12376) );
  NAND2_X1 U15358 ( .A1(n12377), .A2(n12376), .ZN(n12390) );
  AOI22_X1 U15359 ( .A1(n12018), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15360 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9638), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12379) );
  NAND3_X1 U15361 ( .A1(n12380), .A2(n12379), .A3(n12378), .ZN(n12389) );
  AOI22_X1 U15362 ( .A1(n16013), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12019), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15363 ( .A1(n9658), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12381) );
  NAND2_X1 U15364 ( .A1(n12382), .A2(n12381), .ZN(n12388) );
  AOI22_X1 U15365 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15366 ( .A1(n11824), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9638), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12385) );
  NAND3_X1 U15367 ( .A1(n12386), .A2(n12385), .A3(n12384), .ZN(n12387) );
  OAI22_X1 U15368 ( .A1(n12390), .A2(n12389), .B1(n12388), .B2(n12387), .ZN(
        n12391) );
  INV_X1 U15369 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12444) );
  NAND2_X1 U15370 ( .A1(n20272), .A2(n15984), .ZN(n12394) );
  NAND2_X1 U15371 ( .A1(n11808), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12393) );
  NAND2_X1 U15372 ( .A1(n12394), .A2(n12393), .ZN(n13065) );
  NAND2_X1 U15373 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20262), .ZN(
        n12396) );
  NAND2_X1 U15374 ( .A1(n12428), .A2(n12396), .ZN(n12399) );
  NAND2_X1 U15375 ( .A1(n12397), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12398) );
  INV_X1 U15376 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16298) );
  NOR2_X1 U15377 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16298), .ZN(
        n12402) );
  NAND3_X1 U15378 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12403), .A3(
        n12444), .ZN(n12460) );
  NOR2_X1 U15379 ( .A1(n12460), .A2(n13081), .ZN(n12404) );
  OR2_X1 U15380 ( .A1(n13070), .A2(n12404), .ZN(n12442) );
  AOI22_X1 U15381 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15382 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15384 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15385 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12414) );
  AOI22_X1 U15386 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15387 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15388 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15389 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12586), .ZN(n12409) );
  NAND4_X1 U15390 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12413) );
  MUX2_X1 U15391 ( .A(n12460), .B(n14278), .S(n13178), .Z(n12804) );
  AOI22_X1 U15392 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12150), .B1(
        n12098), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15393 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15394 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12581), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15395 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12415) );
  NAND4_X1 U15396 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n12424) );
  AOI22_X1 U15397 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12167), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15398 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15399 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12072), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15400 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12586), .ZN(n12419) );
  NAND4_X1 U15401 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12423) );
  XNOR2_X1 U15402 ( .A(n12426), .B(n12425), .ZN(n12461) );
  MUX2_X1 U15403 ( .A(n12531), .B(n12461), .S(n13081), .Z(n12808) );
  NAND2_X1 U15404 ( .A1(n12804), .A2(n12808), .ZN(n13069) );
  XNOR2_X1 U15405 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12427) );
  XNOR2_X1 U15406 ( .A(n12428), .B(n12427), .ZN(n12805) );
  INV_X1 U15407 ( .A(n12805), .ZN(n12434) );
  OAI21_X1 U15408 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20281), .A(
        n12429), .ZN(n13082) );
  OAI21_X1 U15409 ( .B1(n13082), .B2(n13065), .A(n13178), .ZN(n12433) );
  INV_X1 U15410 ( .A(n13082), .ZN(n12431) );
  INV_X1 U15411 ( .A(n12429), .ZN(n12430) );
  XNOR2_X1 U15412 ( .A(n13065), .B(n12430), .ZN(n12463) );
  OAI211_X1 U15413 ( .C1(n16070), .C2(n12431), .A(n9670), .B(n12463), .ZN(
        n12432) );
  OAI211_X1 U15414 ( .C1(n12435), .C2(n12434), .A(n12433), .B(n12432), .ZN(
        n12439) );
  NAND2_X1 U15415 ( .A1(n12446), .A2(n16070), .ZN(n12436) );
  MUX2_X1 U15416 ( .A(n12436), .B(n13081), .S(n12805), .Z(n12438) );
  INV_X1 U15417 ( .A(n12461), .ZN(n12437) );
  AOI21_X1 U15418 ( .B1(n12439), .B2(n12438), .A(n12437), .ZN(n12440) );
  AOI21_X1 U15419 ( .B1(n13069), .B2(n13081), .A(n12440), .ZN(n12441) );
  NOR2_X1 U15420 ( .A1(n12442), .A2(n12441), .ZN(n12443) );
  MUX2_X1 U15421 ( .A(n12444), .B(n12443), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12445) );
  INV_X1 U15422 ( .A(n12446), .ZN(n13035) );
  NAND2_X1 U15423 ( .A1(n13070), .A2(n13035), .ZN(n12447) );
  NAND2_X1 U15424 ( .A1(n12449), .A2(n11915), .ZN(n12450) );
  NAND2_X1 U15425 ( .A1(n12448), .A2(n12450), .ZN(n12458) );
  AND2_X1 U15426 ( .A1(n12451), .A2(n13156), .ZN(n12457) );
  AND2_X1 U15427 ( .A1(n16039), .A2(n12298), .ZN(n16726) );
  OAI21_X1 U15428 ( .B1(n12452), .B2(n12453), .A(n16726), .ZN(n13165) );
  NAND2_X1 U15429 ( .A1(n12298), .A2(n19646), .ZN(n12459) );
  NAND2_X1 U15430 ( .A1(n12459), .A2(n9670), .ZN(n12454) );
  NAND2_X1 U15431 ( .A1(n12454), .A2(n19659), .ZN(n12455) );
  NAND2_X1 U15432 ( .A1(n12455), .A2(n11915), .ZN(n12456) );
  NAND4_X1 U15433 ( .A1(n12458), .A2(n12457), .A3(n13165), .A4(n12456), .ZN(
        n13019) );
  NAND2_X1 U15434 ( .A1(n16702), .A2(n15991), .ZN(n12470) );
  NAND3_X1 U15435 ( .A1(n12461), .A2(n12460), .A3(n12805), .ZN(n13073) );
  INV_X1 U15436 ( .A(n13073), .ZN(n12462) );
  NAND2_X1 U15437 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20155) );
  AND2_X1 U15438 ( .A1(n12467), .A2(n20155), .ZN(n16695) );
  NAND2_X1 U15439 ( .A1(n12466), .A2(n16695), .ZN(n12468) );
  OR2_X1 U15440 ( .A1(n16698), .A2(n12468), .ZN(n12469) );
  NAND2_X1 U15441 ( .A1(n12470), .A2(n12469), .ZN(n13016) );
  AND2_X1 U15442 ( .A1(n12472), .A2(n12471), .ZN(n13160) );
  NAND2_X1 U15443 ( .A1(n20154), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20162) );
  INV_X1 U15444 ( .A(n11908), .ZN(n12486) );
  NAND2_X1 U15445 ( .A1(n12678), .A2(n16619), .ZN(n12675) );
  AOI22_X1 U15446 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15447 ( .A1(n12581), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12586), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15448 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15449 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15450 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12484) );
  AOI22_X1 U15451 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12580), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15452 ( .A1(n12115), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15453 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15454 ( .A1(n12482), .A2(n12481), .A3(n12480), .A4(n12479), .ZN(
        n12483) );
  NOR2_X1 U15455 ( .A1(n12484), .A2(n12483), .ZN(n13105) );
  MUX2_X1 U15456 ( .A(n19659), .B(n20281), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12487) );
  AND2_X2 U15457 ( .A1(n9655), .A2(n20153), .ZN(n12595) );
  NAND2_X1 U15458 ( .A1(n12486), .A2(n12595), .ZN(n12523) );
  AND2_X1 U15459 ( .A1(n12487), .A2(n12523), .ZN(n12488) );
  INV_X1 U15460 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19303) );
  INV_X1 U15461 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13061) );
  NAND2_X1 U15462 ( .A1(n16070), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12490) );
  OAI211_X1 U15463 ( .C1(n19659), .C2(n13061), .A(n12490), .B(n20153), .ZN(
        n12491) );
  INV_X1 U15464 ( .A(n12491), .ZN(n12492) );
  INV_X1 U15465 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20184) );
  OR2_X1 U15466 ( .A1(n12648), .A2(n20184), .ZN(n12494) );
  INV_X2 U15467 ( .A(n9704), .ZN(n12649) );
  AOI22_X1 U15468 ( .A1(n12649), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15469 ( .A1(n12494), .A2(n12493), .ZN(n12508) );
  XNOR2_X1 U15470 ( .A(n12509), .B(n12508), .ZN(n13342) );
  AOI22_X1 U15471 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15472 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15473 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15474 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12504) );
  AOI22_X1 U15475 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15476 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15477 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15478 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12586), .ZN(n12499) );
  NAND4_X1 U15479 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12503) );
  INV_X1 U15480 ( .A(n13117), .ZN(n12507) );
  NAND2_X1 U15481 ( .A1(n11908), .A2(n19659), .ZN(n12505) );
  MUX2_X1 U15482 ( .A(n12505), .B(n20272), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12506) );
  OAI21_X1 U15483 ( .B1(n12507), .B2(n12619), .A(n12506), .ZN(n13341) );
  NOR2_X1 U15484 ( .A1(n13342), .A2(n13341), .ZN(n12511) );
  NOR2_X1 U15485 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  AOI22_X1 U15486 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12150), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15487 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12098), .B1(
        n12579), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15488 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12580), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15489 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12115), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12512) );
  NAND4_X1 U15490 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12521) );
  AOI22_X1 U15491 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12167), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15492 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12137), .B1(
        n12072), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15493 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n12478), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15494 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12586), .ZN(n12516) );
  NAND4_X1 U15495 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12520) );
  INV_X1 U15496 ( .A(n12806), .ZN(n13751) );
  NAND2_X1 U15497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12522) );
  OAI211_X1 U15498 ( .C1(n12619), .C2(n13751), .A(n12523), .B(n12522), .ZN(
        n12526) );
  XNOR2_X1 U15499 ( .A(n12527), .B(n12526), .ZN(n13149) );
  INV_X1 U15500 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20187) );
  OR2_X1 U15501 ( .A1(n12648), .A2(n20187), .ZN(n12525) );
  AOI22_X1 U15502 ( .A1(n12649), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U15503 ( .A1(n12525), .A2(n12524), .ZN(n13148) );
  NOR2_X1 U15504 ( .A1(n13149), .A2(n13148), .ZN(n12529) );
  NOR2_X1 U15505 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  INV_X1 U15506 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U15507 ( .A1(n12595), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12530) );
  OAI21_X1 U15508 ( .B1(n12648), .B2(n13782), .A(n12530), .ZN(n12534) );
  INV_X1 U15509 ( .A(n12531), .ZN(n13732) );
  NAND2_X1 U15510 ( .A1(n12649), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12532) );
  OAI21_X1 U15511 ( .B1(n12619), .B2(n13732), .A(n12532), .ZN(n12533) );
  INV_X1 U15512 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12535) );
  OR2_X1 U15513 ( .A1(n12648), .A2(n12535), .ZN(n12539) );
  AOI22_X1 U15514 ( .A1(n12649), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12538) );
  INV_X1 U15515 ( .A(n14278), .ZN(n12536) );
  OR2_X1 U15516 ( .A1(n12619), .A2(n12536), .ZN(n12537) );
  AOI22_X1 U15517 ( .A1(n14516), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15518 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12579), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15519 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15520 ( .A1(n12581), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15521 ( .A1(n12580), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12541) );
  NAND4_X1 U15522 ( .A1(n12544), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n12551) );
  AOI22_X1 U15523 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15524 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12072), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15525 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12167), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15526 ( .A1(n12142), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12586), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U15527 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12550) );
  INV_X1 U15528 ( .A(n14262), .ZN(n12552) );
  AOI22_X1 U15529 ( .A1(n12553), .A2(n12552), .B1(n12649), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12554) );
  NAND2_X1 U15530 ( .A1(n12555), .A2(n12554), .ZN(n15960) );
  AOI22_X1 U15531 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12137), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15532 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15533 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12580), .B1(
        n12115), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15534 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12036), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15535 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12565) );
  AOI22_X1 U15536 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12167), .B1(
        n12142), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15537 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15538 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12072), .B1(
        n12051), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15539 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12586), .ZN(n12560) );
  NAND4_X1 U15540 ( .A1(n12563), .A2(n12562), .A3(n12561), .A4(n12560), .ZN(
        n12564) );
  INV_X1 U15541 ( .A(n12810), .ZN(n14304) );
  OR2_X1 U15542 ( .A1(n12619), .A2(n14304), .ZN(n12566) );
  INV_X1 U15543 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20192) );
  OR2_X1 U15544 ( .A1(n12648), .A2(n20192), .ZN(n12568) );
  AOI22_X1 U15545 ( .A1(n12649), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U15546 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U15547 ( .A1(n12150), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U15548 ( .A1(n12137), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12571) );
  NAND2_X1 U15549 ( .A1(n12036), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12570) );
  NAND2_X1 U15550 ( .A1(n12098), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12578) );
  NAND2_X1 U15551 ( .A1(n12142), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12577) );
  NAND2_X1 U15552 ( .A1(n12167), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12576) );
  NAND2_X1 U15553 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U15554 ( .A1(n12579), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12585) );
  NAND2_X1 U15555 ( .A1(n12580), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U15556 ( .A1(n12581), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U15557 ( .A1(n12115), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U15558 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12590) );
  NAND2_X1 U15559 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12589) );
  NAND2_X1 U15560 ( .A1(n12051), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U15561 ( .A1(n12586), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12587) );
  INV_X1 U15562 ( .A(n12595), .ZN(n12629) );
  INV_X1 U15563 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16675) );
  INV_X1 U15564 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19576) );
  INV_X1 U15565 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20194) );
  OAI222_X1 U15566 ( .A1(n12629), .A2(n16675), .B1(n9704), .B2(n19576), .C1(
        n12648), .C2(n20194), .ZN(n15925) );
  INV_X1 U15567 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13870) );
  OR2_X1 U15568 ( .A1(n12648), .A2(n13870), .ZN(n12599) );
  AOI22_X1 U15569 ( .A1(n12649), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12598) );
  INV_X1 U15570 ( .A(n19479), .ZN(n12596) );
  OR2_X1 U15571 ( .A1(n12619), .A2(n12596), .ZN(n12597) );
  INV_X1 U15572 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12600) );
  OR2_X1 U15573 ( .A1(n12648), .A2(n12600), .ZN(n12602) );
  AOI22_X1 U15574 ( .A1(n12649), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12595), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12601) );
  OAI211_X1 U15575 ( .C1(n13485), .C2(n12619), .A(n12602), .B(n12601), .ZN(
        n15908) );
  INV_X1 U15576 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12603) );
  OR2_X1 U15577 ( .A1(n12648), .A2(n12603), .ZN(n12605) );
  AOI22_X1 U15578 ( .A1(n12649), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12604) );
  OAI211_X1 U15579 ( .C1(n9753), .C2(n12619), .A(n12605), .B(n12604), .ZN(
        n15895) );
  INV_X1 U15580 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12606) );
  OR2_X1 U15581 ( .A1(n12648), .A2(n12606), .ZN(n12608) );
  AOI22_X1 U15582 ( .A1(n12649), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12607) );
  OAI211_X1 U15583 ( .C1(n13618), .C2(n12619), .A(n12608), .B(n12607), .ZN(
        n15865) );
  INV_X1 U15584 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n15607) );
  OR2_X1 U15585 ( .A1(n12648), .A2(n15607), .ZN(n12611) );
  AOI22_X1 U15586 ( .A1(n12649), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12610) );
  OAI211_X1 U15587 ( .C1(n19472), .C2(n12619), .A(n12611), .B(n12610), .ZN(
        n15852) );
  INV_X1 U15588 ( .A(n13973), .ZN(n12614) );
  INV_X1 U15589 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15589) );
  OR2_X1 U15590 ( .A1(n12648), .A2(n15589), .ZN(n12613) );
  AOI22_X1 U15591 ( .A1(n12649), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12612) );
  OAI211_X1 U15592 ( .C1(n12614), .C2(n12619), .A(n12613), .B(n12612), .ZN(
        n12824) );
  INV_X1 U15593 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15576) );
  OR2_X1 U15594 ( .A1(n12648), .A2(n15576), .ZN(n12616) );
  AOI22_X1 U15595 ( .A1(n12649), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12615) );
  OAI211_X1 U15596 ( .C1(n13984), .C2(n12619), .A(n12616), .B(n12615), .ZN(
        n14009) );
  INV_X1 U15597 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20203) );
  OR2_X1 U15598 ( .A1(n12648), .A2(n20203), .ZN(n12618) );
  AOI22_X1 U15599 ( .A1(n12649), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12617) );
  OAI211_X1 U15600 ( .C1(n14020), .C2(n12619), .A(n12618), .B(n12617), .ZN(
        n15811) );
  INV_X1 U15601 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15552) );
  OR2_X1 U15602 ( .A1(n12648), .A2(n15552), .ZN(n12621) );
  AOI22_X1 U15603 ( .A1(n12649), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12620) );
  INV_X1 U15604 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20206) );
  OR2_X1 U15605 ( .A1(n12648), .A2(n20206), .ZN(n12623) );
  AOI22_X1 U15606 ( .A1(n12649), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U15607 ( .A1(n12623), .A2(n12622), .ZN(n13977) );
  NAND2_X1 U15608 ( .A1(n15236), .A2(n13977), .ZN(n15222) );
  INV_X1 U15609 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15535) );
  OR2_X1 U15610 ( .A1(n12648), .A2(n15535), .ZN(n12625) );
  AOI22_X1 U15611 ( .A1(n12649), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12624) );
  AND2_X1 U15612 ( .A1(n12625), .A2(n12624), .ZN(n15221) );
  INV_X1 U15613 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15389) );
  INV_X1 U15614 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15765) );
  OAI22_X1 U15615 ( .A1(n9704), .A2(n15389), .B1(n15765), .B2(n12629), .ZN(
        n12626) );
  AOI21_X1 U15616 ( .B1(n14516), .B2(P2_REIP_REG_19__SCAN_IN), .A(n12626), 
        .ZN(n15386) );
  NOR2_X2 U15617 ( .A1(n9708), .A2(n15386), .ZN(n15387) );
  INV_X1 U15618 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15510) );
  OR2_X1 U15619 ( .A1(n12648), .A2(n15510), .ZN(n12628) );
  AOI22_X1 U15620 ( .A1(n12649), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12627) );
  NAND2_X1 U15621 ( .A1(n12628), .A2(n12627), .ZN(n15209) );
  NAND2_X1 U15622 ( .A1(n15387), .A2(n15209), .ZN(n15380) );
  INV_X1 U15623 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15381) );
  INV_X1 U15624 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15740) );
  OAI22_X1 U15625 ( .A1(n9704), .A2(n15381), .B1(n15740), .B2(n12629), .ZN(
        n12630) );
  AOI21_X1 U15626 ( .B1(n14516), .B2(P2_REIP_REG_21__SCAN_IN), .A(n12630), 
        .ZN(n15379) );
  INV_X1 U15627 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15482) );
  OR2_X1 U15628 ( .A1(n12648), .A2(n15482), .ZN(n12632) );
  AOI22_X1 U15629 ( .A1(n12649), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12631) );
  AND2_X1 U15630 ( .A1(n12632), .A2(n12631), .ZN(n15722) );
  INV_X1 U15631 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20215) );
  OR2_X1 U15632 ( .A1(n12648), .A2(n20215), .ZN(n12634) );
  AOI22_X1 U15633 ( .A1(n12649), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12633) );
  AND2_X1 U15634 ( .A1(n12634), .A2(n12633), .ZN(n15371) );
  INV_X1 U15635 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20217) );
  OR2_X1 U15636 ( .A1(n12648), .A2(n20217), .ZN(n12636) );
  AOI22_X1 U15637 ( .A1(n12649), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15638 ( .A1(n12636), .A2(n12635), .ZN(n15363) );
  INV_X1 U15639 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20219) );
  OR2_X1 U15640 ( .A1(n12648), .A2(n20219), .ZN(n12638) );
  AOI22_X1 U15641 ( .A1(n12649), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U15642 ( .A1(n12638), .A2(n12637), .ZN(n15357) );
  INV_X1 U15643 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20221) );
  OR2_X1 U15644 ( .A1(n12648), .A2(n20221), .ZN(n12640) );
  AOI22_X1 U15645 ( .A1(n12649), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12639) );
  AND2_X1 U15646 ( .A1(n12640), .A2(n12639), .ZN(n15347) );
  INV_X1 U15647 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20224) );
  OR2_X1 U15648 ( .A1(n12648), .A2(n20224), .ZN(n12642) );
  AOI22_X1 U15649 ( .A1(n12649), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12641) );
  AND2_X1 U15650 ( .A1(n12642), .A2(n12641), .ZN(n14475) );
  NOR2_X2 U15651 ( .A1(n9707), .A2(n14475), .ZN(n14476) );
  INV_X1 U15652 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n14444) );
  OR2_X1 U15653 ( .A1(n12648), .A2(n14444), .ZN(n12644) );
  AOI22_X1 U15654 ( .A1(n12649), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U15655 ( .A1(n12644), .A2(n12643), .ZN(n14460) );
  NAND2_X1 U15656 ( .A1(n14476), .A2(n14460), .ZN(n15323) );
  INV_X1 U15657 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20226) );
  OR2_X1 U15658 ( .A1(n12648), .A2(n20226), .ZN(n12646) );
  AOI22_X1 U15659 ( .A1(n12649), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12645) );
  AND2_X1 U15660 ( .A1(n12646), .A2(n12645), .ZN(n15322) );
  INV_X1 U15661 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12647) );
  OR2_X1 U15662 ( .A1(n12648), .A2(n12647), .ZN(n12651) );
  AOI22_X1 U15663 ( .A1(n12649), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12650) );
  AND2_X1 U15664 ( .A1(n12651), .A2(n12650), .ZN(n12654) );
  INV_X1 U15665 ( .A(n12654), .ZN(n12652) );
  INV_X1 U15666 ( .A(n12653), .ZN(n15325) );
  NAND2_X1 U15667 ( .A1(n15325), .A2(n12654), .ZN(n12655) );
  NAND2_X1 U15668 ( .A1(n14518), .A2(n12655), .ZN(n16506) );
  NAND2_X1 U15669 ( .A1(n19537), .A2(n12453), .ZN(n19538) );
  NOR2_X1 U15670 ( .A1(n12453), .A2(n11844), .ZN(n12656) );
  NOR4_X1 U15671 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12660) );
  NOR4_X1 U15672 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12659) );
  NOR4_X1 U15673 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12658) );
  NOR4_X1 U15674 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12657) );
  NAND4_X1 U15675 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12665) );
  NOR4_X1 U15676 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12663) );
  NOR4_X1 U15677 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12662) );
  NOR4_X1 U15678 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12661) );
  INV_X1 U15679 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20188) );
  NAND4_X1 U15680 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n20188), .ZN(
        n12664) );
  INV_X1 U15681 ( .A(n19497), .ZN(n15356) );
  INV_X1 U15682 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n12670) );
  NAND2_X1 U15683 ( .A1(n12968), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12668) );
  INV_X1 U15684 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16841) );
  OR2_X1 U15685 ( .A1(n12968), .A2(n16841), .ZN(n12667) );
  NAND2_X1 U15686 ( .A1(n12668), .A2(n12667), .ZN(n19507) );
  AOI22_X1 U15687 ( .A1(n19495), .A2(n19507), .B1(n19546), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n12669) );
  OAI21_X1 U15688 ( .B1(n15356), .B2(n12670), .A(n12669), .ZN(n12671) );
  AOI21_X1 U15689 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n19496), .A(n12671), .ZN(
        n12672) );
  NAND2_X1 U15690 ( .A1(n12675), .A2(n12674), .ZN(P2_U2889) );
  NAND2_X1 U15691 ( .A1(n11957), .A2(n12676), .ZN(n15990) );
  OR2_X1 U15692 ( .A1(n16702), .A2(n15990), .ZN(n13023) );
  INV_X1 U15693 ( .A(n13170), .ZN(n15995) );
  NAND2_X1 U15694 ( .A1(n13023), .A2(n15995), .ZN(n12677) );
  NAND2_X1 U15695 ( .A1(n12678), .A2(n19487), .ZN(n12771) );
  INV_X1 U15696 ( .A(n12679), .ZN(n12680) );
  INV_X1 U15697 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15965) );
  AOI22_X1 U15698 ( .A1(n9648), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12683) );
  NAND2_X1 U15699 ( .A1(n14506), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12682) );
  OAI211_X1 U15700 ( .C1(n14510), .C2(n15965), .A(n12683), .B(n12682), .ZN(
        n13893) );
  NAND2_X1 U15701 ( .A1(n14506), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15702 ( .A1(n9648), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12684) );
  OAI211_X1 U15703 ( .C1(n20154), .C2(n12686), .A(n12685), .B(n12684), .ZN(
        n12687) );
  AOI21_X1 U15704 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12687), .ZN(n13445) );
  NOR2_X2 U15705 ( .A1(n13895), .A2(n13445), .ZN(n13524) );
  INV_X1 U15706 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15940) );
  AOI22_X1 U15707 ( .A1(n9648), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12689) );
  NAND2_X1 U15708 ( .A1(n14506), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12688) );
  OAI211_X1 U15709 ( .C1(n14510), .C2(n15940), .A(n12689), .B(n12688), .ZN(
        n13525) );
  NAND2_X1 U15710 ( .A1(n14506), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U15711 ( .A1(n9648), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12690) );
  OAI211_X1 U15712 ( .C1(n20154), .C2(n12692), .A(n12691), .B(n12690), .ZN(
        n12693) );
  AOI21_X1 U15713 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12693), .ZN(n13516) );
  INV_X1 U15714 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16689) );
  AOI22_X1 U15715 ( .A1(n9648), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12695) );
  NAND2_X1 U15716 ( .A1(n14506), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12694) );
  OAI211_X1 U15717 ( .C1(n14510), .C2(n16689), .A(n12695), .B(n12694), .ZN(
        n13872) );
  NAND2_X1 U15718 ( .A1(n12760), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12701) );
  INV_X1 U15719 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U15720 ( .A1(n9648), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U15721 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12697) );
  OAI211_X1 U15722 ( .C1(n13493), .C2(n12696), .A(n12698), .B(n12697), .ZN(
        n12699) );
  INV_X1 U15723 ( .A(n12699), .ZN(n12700) );
  NAND2_X1 U15724 ( .A1(n12701), .A2(n12700), .ZN(n13489) );
  INV_X1 U15725 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15726 ( .A1(n9648), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U15727 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12702) );
  OAI211_X1 U15728 ( .C1(n12704), .C2(n12696), .A(n12703), .B(n12702), .ZN(
        n12705) );
  AOI21_X1 U15729 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12705), .ZN(n15889) );
  INV_X1 U15730 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12708) );
  NAND2_X1 U15731 ( .A1(n9648), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U15732 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12706) );
  OAI211_X1 U15733 ( .C1(n12708), .C2(n12696), .A(n12707), .B(n12706), .ZN(
        n12709) );
  AOI21_X1 U15734 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12709), .ZN(n13619) );
  NOR2_X2 U15735 ( .A1(n15892), .A2(n13619), .ZN(n15604) );
  INV_X1 U15736 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15858) );
  AOI22_X1 U15737 ( .A1(n9648), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12711) );
  NAND2_X1 U15738 ( .A1(n14506), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12710) );
  OAI211_X1 U15739 ( .C1(n14510), .C2(n15858), .A(n12711), .B(n12710), .ZN(
        n15603) );
  INV_X1 U15740 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U15741 ( .A1(n9648), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U15742 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12712) );
  OAI211_X1 U15743 ( .C1(n12812), .C2(n12696), .A(n12713), .B(n12712), .ZN(
        n12714) );
  AOI21_X1 U15744 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12714), .ZN(n12818) );
  INV_X1 U15745 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U15746 ( .A1(n9648), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U15747 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12715) );
  OAI211_X1 U15748 ( .C1(n14002), .C2(n12696), .A(n12716), .B(n12715), .ZN(
        n12717) );
  AOI21_X1 U15749 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12717), .ZN(n13986) );
  INV_X1 U15750 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U15751 ( .A1(n9648), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12719) );
  NAND2_X1 U15752 ( .A1(n14506), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12718) );
  OAI211_X1 U15753 ( .C1(n14510), .C2(n15784), .A(n12719), .B(n12718), .ZN(
        n14018) );
  INV_X1 U15754 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U15755 ( .A1(n9648), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12721) );
  NAND2_X1 U15756 ( .A1(n14506), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12720) );
  OAI211_X1 U15757 ( .C1(n14510), .C2(n15800), .A(n12721), .B(n12720), .ZN(
        n15232) );
  INV_X1 U15758 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n14228) );
  NAND2_X1 U15759 ( .A1(n9648), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15760 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12722) );
  OAI211_X1 U15761 ( .C1(n14228), .C2(n12696), .A(n12723), .B(n12722), .ZN(
        n12724) );
  AOI21_X1 U15762 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12724), .ZN(n15318) );
  INV_X1 U15763 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U15764 ( .A1(n9648), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U15765 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12725) );
  OAI211_X1 U15766 ( .C1(n14229), .C2(n12696), .A(n12726), .B(n12725), .ZN(
        n12727) );
  AOI21_X1 U15767 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12727), .ZN(n15225) );
  INV_X1 U15768 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n14230) );
  NAND2_X1 U15769 ( .A1(n9648), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15770 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12728) );
  OAI211_X1 U15771 ( .C1(n14230), .C2(n12696), .A(n12729), .B(n12728), .ZN(
        n12730) );
  AOI21_X1 U15772 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12730), .ZN(n15310) );
  INV_X1 U15773 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U15774 ( .A1(n9648), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12732) );
  NAND2_X1 U15775 ( .A1(n14506), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12731) );
  OAI211_X1 U15776 ( .C1(n14510), .C2(n15748), .A(n12732), .B(n12731), .ZN(
        n15206) );
  INV_X1 U15777 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U15778 ( .A1(n9648), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U15779 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12733) );
  OAI211_X1 U15780 ( .C1(n14367), .C2(n12696), .A(n12734), .B(n12733), .ZN(
        n12735) );
  AOI21_X1 U15781 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12735), .ZN(n15302) );
  INV_X1 U15782 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12738) );
  NAND2_X1 U15783 ( .A1(n9648), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U15784 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12736) );
  OAI211_X1 U15785 ( .C1(n12738), .C2(n12696), .A(n12737), .B(n12736), .ZN(
        n12739) );
  AOI21_X1 U15786 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12739), .ZN(n15478) );
  INV_X1 U15787 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U15788 ( .A1(n9648), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12741) );
  NAND2_X1 U15789 ( .A1(n14506), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12740) );
  OAI211_X1 U15790 ( .C1(n14510), .C2(n15713), .A(n12741), .B(n12740), .ZN(
        n15291) );
  INV_X1 U15791 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15288) );
  NAND2_X1 U15792 ( .A1(n9648), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15793 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12742) );
  OAI211_X1 U15794 ( .C1(n15288), .C2(n12696), .A(n12743), .B(n12742), .ZN(
        n12744) );
  AOI21_X1 U15795 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12744), .ZN(n15287) );
  INV_X1 U15796 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U15797 ( .A1(n9648), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15798 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12745) );
  OAI211_X1 U15799 ( .C1(n15278), .C2(n12696), .A(n12746), .B(n12745), .ZN(
        n12747) );
  AOI21_X1 U15800 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12747), .ZN(n15275) );
  INV_X1 U15801 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U15802 ( .A1(n9648), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12749) );
  NAND2_X1 U15803 ( .A1(n14506), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12748) );
  OAI211_X1 U15804 ( .C1(n14510), .C2(n15677), .A(n12749), .B(n12748), .ZN(
        n15267) );
  INV_X1 U15805 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U15806 ( .A1(n9648), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12751) );
  NAND2_X1 U15807 ( .A1(n14506), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12750) );
  OAI211_X1 U15808 ( .C1(n14510), .C2(n14486), .A(n12751), .B(n12750), .ZN(
        n14473) );
  INV_X1 U15809 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U15810 ( .A1(n9648), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U15811 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12752) );
  OAI211_X1 U15812 ( .C1(n14413), .C2(n12696), .A(n12753), .B(n12752), .ZN(
        n12754) );
  AOI21_X1 U15813 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12754), .ZN(n14442) );
  INV_X1 U15814 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12758) );
  NAND2_X1 U15815 ( .A1(n9648), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U15816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12756) );
  OAI211_X1 U15817 ( .C1(n12696), .C2(n12758), .A(n12757), .B(n12756), .ZN(
        n12759) );
  AOI21_X1 U15818 ( .B1(n12760), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12759), .ZN(n15246) );
  NOR2_X2 U15819 ( .A1(n9706), .A2(n15246), .ZN(n12763) );
  INV_X1 U15820 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U15821 ( .A1(n9648), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12762) );
  NAND2_X1 U15822 ( .A1(n14506), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12761) );
  OAI211_X1 U15823 ( .C1(n14510), .C2(n15647), .A(n12762), .B(n12761), .ZN(
        n12764) );
  NAND2_X1 U15824 ( .A1(n12763), .A2(n12764), .ZN(n14511) );
  INV_X1 U15825 ( .A(n12763), .ZN(n12766) );
  INV_X1 U15826 ( .A(n12764), .ZN(n12765) );
  NAND2_X1 U15827 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U15828 ( .A1(n14511), .A2(n12767), .ZN(n15644) );
  INV_X2 U15829 ( .A(n19490), .ZN(n19484) );
  NAND2_X1 U15830 ( .A1(n19484), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12768) );
  OAI21_X1 U15831 ( .B1(n15644), .B2(n19484), .A(n12768), .ZN(n12769) );
  INV_X1 U15832 ( .A(n12769), .ZN(n12770) );
  NAND2_X1 U15833 ( .A1(n12771), .A2(n12770), .ZN(P2_U2857) );
  NOR2_X1 U15834 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12773) );
  NOR4_X1 U15835 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12772) );
  NAND4_X1 U15836 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12773), .A4(n12772), .ZN(n12776) );
  NOR2_X1 U15837 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12776), .ZN(n16896)
         );
  INV_X1 U15838 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21055) );
  NOR3_X1 U15839 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21055), .ZN(n12775) );
  NOR4_X1 U15840 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12774)
         );
  NAND4_X1 U15841 ( .A1(n13623), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12775), .A4(
        n12774), .ZN(U214) );
  NOR2_X1 U15842 ( .A1(n16040), .A2(n12776), .ZN(n16807) );
  NAND2_X1 U15843 ( .A1(n16807), .A2(U214), .ZN(U212) );
  INV_X1 U15844 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15590) );
  NAND2_X1 U15845 ( .A1(n12790), .A2(n15590), .ZN(n12777) );
  AND2_X1 U15846 ( .A1(n14005), .A2(n12777), .ZN(n15592) );
  AND2_X1 U15847 ( .A1(n12787), .A2(n15624), .ZN(n12778) );
  NOR2_X1 U15848 ( .A1(n9748), .A2(n12778), .ZN(n19373) );
  AOI21_X1 U15849 ( .B1(n19389), .B2(n12785), .A(n12788), .ZN(n19396) );
  AOI21_X1 U15850 ( .B1(n12692), .B2(n12784), .A(n12786), .ZN(n19402) );
  AOI21_X1 U15851 ( .B1(n12686), .B2(n12782), .A(n9678), .ZN(n19435) );
  AOI21_X1 U15852 ( .B1(n14040), .B2(n12781), .A(n12783), .ZN(n14038) );
  OAI22_X1 U15853 ( .A1(n16735), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n12779) );
  INV_X1 U15854 ( .A(n12779), .ZN(n14049) );
  INV_X1 U15855 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U15856 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12780), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16735), .ZN(n14027) );
  NOR2_X1 U15857 ( .A1(n14049), .A2(n14027), .ZN(n14026) );
  OAI21_X1 U15858 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12781), .ZN(n13921) );
  NAND2_X1 U15859 ( .A1(n14026), .A2(n13921), .ZN(n14036) );
  NOR2_X1 U15860 ( .A1(n14038), .A2(n14036), .ZN(n13889) );
  OAI21_X1 U15861 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12783), .A(
        n12782), .ZN(n19602) );
  NAND2_X1 U15862 ( .A1(n13889), .A2(n19602), .ZN(n19432) );
  NOR2_X1 U15863 ( .A1(n19435), .A2(n19432), .ZN(n19415) );
  OAI21_X1 U15864 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9678), .A(
        n12784), .ZN(n19417) );
  NAND2_X1 U15865 ( .A1(n19415), .A2(n19417), .ZN(n19401) );
  NOR2_X1 U15866 ( .A1(n19402), .A2(n19401), .ZN(n13866) );
  OAI21_X1 U15867 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12786), .A(
        n12785), .ZN(n16653) );
  NAND2_X1 U15868 ( .A1(n13866), .A2(n16653), .ZN(n19394) );
  NOR2_X1 U15869 ( .A1(n19396), .A2(n19394), .ZN(n19379) );
  OAI21_X1 U15870 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12788), .A(
        n12787), .ZN(n19381) );
  NAND2_X1 U15871 ( .A1(n19379), .A2(n19381), .ZN(n19372) );
  NOR2_X1 U15872 ( .A1(n19373), .A2(n19372), .ZN(n19358) );
  OR2_X1 U15873 ( .A1(n9748), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12789) );
  NAND2_X1 U15874 ( .A1(n12790), .A2(n12789), .ZN(n19359) );
  NAND2_X1 U15875 ( .A1(n19358), .A2(n19359), .ZN(n12793) );
  NOR2_X1 U15876 ( .A1(n15592), .A2(n12793), .ZN(n15175) );
  INV_X1 U15877 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20049) );
  NAND4_X1 U15878 ( .A1(n20049), .A2(n19955), .A3(n16735), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20159) );
  INV_X1 U15879 ( .A(n20159), .ZN(n19420) );
  INV_X1 U15880 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14004) );
  INV_X1 U15881 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19335) );
  INV_X1 U15882 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15180) );
  INV_X1 U15883 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19322) );
  INV_X1 U15884 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15467) );
  INV_X1 U15885 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15451) );
  INV_X1 U15886 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15169) );
  INV_X1 U15887 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15431) );
  INV_X1 U15888 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12792) );
  INV_X1 U15889 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14509) );
  NAND2_X1 U15890 ( .A1(n19420), .A2(n9647), .ZN(n16504) );
  AOI211_X1 U15891 ( .C1(n15592), .C2(n12793), .A(n15175), .B(n16504), .ZN(
        n12828) );
  INV_X1 U15892 ( .A(n12794), .ZN(n12795) );
  INV_X1 U15893 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19279) );
  INV_X1 U15894 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20183) );
  NOR2_X1 U15895 ( .A1(n19279), .A2(n20183), .ZN(n20174) );
  NOR2_X1 U15896 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20176) );
  NOR3_X1 U15897 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20174), .A3(n20176), 
        .ZN(n20168) );
  NAND2_X1 U15898 ( .A1(n20155), .A2(n20168), .ZN(n13017) );
  INV_X1 U15899 ( .A(n13017), .ZN(n16694) );
  NAND2_X1 U15900 ( .A1(n20049), .A2(n16694), .ZN(n16727) );
  INV_X1 U15901 ( .A(n16727), .ZN(n16494) );
  OR2_X1 U15902 ( .A1(n16495), .A2(n16494), .ZN(n12797) );
  INV_X1 U15903 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16586) );
  INV_X1 U15904 ( .A(n12936), .ZN(n12937) );
  INV_X1 U15905 ( .A(n20155), .ZN(n20175) );
  OR2_X1 U15906 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20175), .ZN(n12819) );
  NAND3_X1 U15907 ( .A1(n16586), .A2(n12937), .A3(n12819), .ZN(n12796) );
  INV_X1 U15908 ( .A(n19443), .ZN(n19429) );
  INV_X1 U15909 ( .A(n12448), .ZN(n12798) );
  NAND2_X1 U15910 ( .A1(n12799), .A2(n12798), .ZN(n19277) );
  NAND2_X1 U15911 ( .A1(n12936), .A2(n19277), .ZN(n19282) );
  INV_X1 U15912 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20153) );
  NAND2_X1 U15913 ( .A1(n20154), .A2(n20153), .ZN(n19283) );
  NOR2_X1 U15914 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19283), .ZN(n12800) );
  AND2_X1 U15915 ( .A1(n12800), .A2(n16735), .ZN(n16662) );
  NOR3_X1 U15916 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20162), .A3(n20153), 
        .ZN(n16724) );
  INV_X1 U15917 ( .A(n16724), .ZN(n12801) );
  NAND2_X1 U15918 ( .A1(n20159), .A2(n12801), .ZN(n12802) );
  NAND2_X1 U15919 ( .A1(n19425), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19390) );
  OAI22_X1 U15920 ( .A1(n19429), .A2(n12812), .B1(n15590), .B2(n19390), .ZN(
        n12827) );
  INV_X1 U15921 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12803) );
  MUX2_X1 U15922 ( .A(n12804), .B(n12803), .S(n14328), .Z(n13897) );
  MUX2_X1 U15923 ( .A(n12806), .B(n12805), .S(n13081), .Z(n13067) );
  INV_X1 U15924 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13924) );
  MUX2_X1 U15925 ( .A(n13067), .B(n13924), .S(n14328), .Z(n13126) );
  NOR2_X1 U15926 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12807) );
  MUX2_X1 U15927 ( .A(n13117), .B(n12807), .S(n14328), .Z(n13127) );
  INV_X1 U15928 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14044) );
  MUX2_X1 U15929 ( .A(n12808), .B(n14044), .S(n14328), .Z(n12809) );
  MUX2_X1 U15931 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n14262), .S(n19650), .Z(
        n14267) );
  INV_X1 U15932 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19412) );
  MUX2_X1 U15933 ( .A(n12810), .B(n19412), .S(n14328), .Z(n14309) );
  INV_X1 U15934 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12811) );
  MUX2_X1 U15935 ( .A(n12811), .B(n14497), .S(n19650), .Z(n14313) );
  NAND2_X1 U15936 ( .A1(n14328), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U15938 ( .A1(n14328), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14342) );
  NOR2_X1 U15939 ( .A1(n19650), .A2(n12812), .ZN(n14000) );
  INV_X1 U15940 ( .A(n14000), .ZN(n12813) );
  XNOR2_X1 U15941 ( .A(n14344), .B(n12813), .ZN(n14346) );
  NAND2_X1 U15942 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12819), .ZN(n12814) );
  NOR2_X1 U15943 ( .A1(n13081), .A2(n12814), .ZN(n12815) );
  NOR2_X1 U15944 ( .A1(n9647), .A2(n20159), .ZN(n19458) );
  AOI22_X1 U15945 ( .A1(n14346), .A2(n19448), .B1(n19458), .B2(n15592), .ZN(
        n12816) );
  INV_X2 U15946 ( .A(n16662), .ZN(n19424) );
  OAI211_X1 U15947 ( .C1(n15589), .C2(n19425), .A(n12816), .B(n19424), .ZN(
        n12826) );
  INV_X1 U15948 ( .A(n13987), .ZN(n12817) );
  AOI21_X1 U15949 ( .B1(n12818), .B2(n15606), .A(n12817), .ZN(n15841) );
  INV_X1 U15950 ( .A(n15841), .ZN(n15594) );
  NOR2_X1 U15951 ( .A1(n13081), .A2(n12819), .ZN(n12820) );
  NAND2_X1 U15952 ( .A1(n19282), .A2(n12820), .ZN(n19453) );
  INV_X1 U15953 ( .A(n12822), .ZN(n12823) );
  OAI21_X1 U15954 ( .B1(n12821), .B2(n12824), .A(n12823), .ZN(n19511) );
  OAI22_X1 U15955 ( .A1(n15594), .A2(n19453), .B1(n19511), .B2(n19442), .ZN(
        n12825) );
  OR4_X1 U15956 ( .A1(n12828), .A2(n12827), .A3(n12826), .A4(n12825), .ZN(
        P2_U2842) );
  INV_X1 U15957 ( .A(n12830), .ZN(n12831) );
  NOR2_X1 U15958 ( .A1(n12829), .A2(n12831), .ZN(n15002) );
  INV_X1 U15959 ( .A(n12832), .ZN(n12833) );
  NOR2_X1 U15960 ( .A1(n15002), .A2(n12833), .ZN(n12836) );
  NAND2_X1 U15961 ( .A1(n12834), .A2(n15001), .ZN(n12835) );
  XNOR2_X1 U15962 ( .A(n12836), .B(n12835), .ZN(n16350) );
  INV_X1 U15963 ( .A(n12837), .ZN(n12838) );
  NAND2_X1 U15964 ( .A1(n12838), .A2(n20971), .ZN(n21061) );
  NAND2_X1 U15965 ( .A1(n13635), .A2(n21061), .ZN(n12840) );
  NAND2_X1 U15966 ( .A1(n12840), .A2(n12839), .ZN(n12845) );
  AOI22_X1 U15967 ( .A1(n12841), .A2(n13213), .B1(n21062), .B2(n21061), .ZN(
        n12842) );
  OAI21_X1 U15968 ( .B1(n12843), .B2(n12842), .A(n16254), .ZN(n12844) );
  MUX2_X1 U15969 ( .A(n12845), .B(n12844), .S(n10225), .Z(n12854) );
  OR2_X1 U15970 ( .A1(n13299), .A2(n13638), .ZN(n12851) );
  NAND2_X1 U15971 ( .A1(n12851), .A2(n13213), .ZN(n12847) );
  OR2_X1 U15972 ( .A1(n12848), .A2(n12847), .ZN(n12869) );
  NAND2_X1 U15973 ( .A1(n12849), .A2(n12869), .ZN(n12850) );
  NAND2_X1 U15974 ( .A1(n10137), .A2(n12850), .ZN(n13250) );
  OAI21_X1 U15975 ( .B1(n16254), .B2(n12851), .A(n13250), .ZN(n12852) );
  INV_X1 U15976 ( .A(n12852), .ZN(n12853) );
  NAND2_X1 U15977 ( .A1(n12854), .A2(n12853), .ZN(n12855) );
  INV_X1 U15978 ( .A(n12931), .ZN(n12876) );
  OAI21_X1 U15979 ( .B1(n12929), .B2(n12856), .A(n16247), .ZN(n12857) );
  NOR2_X1 U15980 ( .A1(n16246), .A2(n12857), .ZN(n12858) );
  AND2_X1 U15981 ( .A1(n10412), .A2(n12858), .ZN(n12859) );
  NOR2_X1 U15982 ( .A1(n16350), .A2(n20431), .ZN(n12934) );
  INV_X1 U15983 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13311) );
  NOR2_X1 U15984 ( .A1(n13314), .A2(n13311), .ZN(n13374) );
  AND2_X1 U15985 ( .A1(n12846), .A2(n13635), .ZN(n16232) );
  NAND2_X2 U15986 ( .A1(n12860), .A2(n13213), .ZN(n14150) );
  NAND2_X1 U15987 ( .A1(n12861), .A2(n13635), .ZN(n12864) );
  INV_X1 U15988 ( .A(n10225), .ZN(n13418) );
  OAI21_X1 U15989 ( .B1(n12862), .B2(n13213), .A(n13418), .ZN(n12863) );
  OAI211_X1 U15990 ( .C1(n10399), .C2(n16259), .A(n12864), .B(n12863), .ZN(
        n12865) );
  INV_X1 U15991 ( .A(n12865), .ZN(n12867) );
  NAND2_X1 U15992 ( .A1(n10404), .A2(n14164), .ZN(n12866) );
  OAI211_X1 U15993 ( .C1(n14121), .C2(n9836), .A(n12867), .B(n12866), .ZN(
        n12868) );
  INV_X1 U15994 ( .A(n12868), .ZN(n12870) );
  OAI211_X1 U15995 ( .C1(n12872), .C2(n12871), .A(n12870), .B(n12869), .ZN(
        n13239) );
  OAI21_X1 U15996 ( .B1(n13240), .B2(n13213), .A(n12873), .ZN(n12874) );
  NOR2_X1 U15997 ( .A1(n13239), .A2(n12874), .ZN(n12875) );
  NOR2_X1 U15998 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20447), .ZN(
        n13292) );
  NOR2_X1 U15999 ( .A1(n12877), .A2(n14158), .ZN(n12878) );
  NAND2_X1 U16000 ( .A1(n13260), .A2(n12878), .ZN(n13261) );
  INV_X1 U16001 ( .A(n13261), .ZN(n16249) );
  AOI21_X1 U16002 ( .B1(n13374), .B2(n15022), .A(n15151), .ZN(n13371) );
  AOI21_X1 U16003 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13372) );
  NOR2_X1 U16004 ( .A1(n20425), .A2(n10572), .ZN(n20436) );
  NAND2_X1 U16005 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20436), .ZN(
        n13667) );
  NOR2_X1 U16006 ( .A1(n13372), .A2(n13667), .ZN(n16446) );
  NAND3_X1 U16007 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16451) );
  NOR3_X1 U16008 ( .A1(n12917), .A2(n14059), .A3(n16451), .ZN(n12879) );
  NAND3_X1 U16009 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16446), .A3(
        n12879), .ZN(n15018) );
  NOR2_X1 U16010 ( .A1(n13371), .A2(n15018), .ZN(n12886) );
  NAND2_X1 U16011 ( .A1(n12879), .A2(n10735), .ZN(n16443) );
  INV_X1 U16012 ( .A(n16443), .ZN(n12883) );
  NOR3_X1 U16013 ( .A1(n13314), .A2(n13311), .A3(n13667), .ZN(n16448) );
  AND2_X1 U16014 ( .A1(n12879), .A2(n16448), .ZN(n15020) );
  NAND2_X1 U16015 ( .A1(n15151), .A2(n15018), .ZN(n12882) );
  INV_X1 U16016 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20443) );
  NAND2_X1 U16017 ( .A1(n20441), .A2(n20443), .ZN(n12881) );
  INV_X2 U16018 ( .A(n20347), .ZN(n20334) );
  OR2_X1 U16019 ( .A1(n12931), .A2(n20334), .ZN(n12880) );
  OAI211_X1 U16020 ( .C1(n16447), .C2(n15020), .A(n12882), .B(n16445), .ZN(
        n16439) );
  AOI21_X1 U16021 ( .B1(n15022), .B2(n12883), .A(n16439), .ZN(n12884) );
  INV_X1 U16022 ( .A(n12884), .ZN(n12885) );
  MUX2_X1 U16023 ( .A(n12886), .B(n12885), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n12933) );
  NAND2_X1 U16024 ( .A1(n14150), .A2(n13311), .ZN(n12887) );
  NAND2_X1 U16025 ( .A1(n14150), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12890) );
  OAI21_X1 U16026 ( .B1(n14164), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12890), .ZN(
        n13296) );
  XNOR2_X1 U16027 ( .A(n12891), .B(n13296), .ZN(n13286) );
  NAND2_X1 U16028 ( .A1(n13285), .A2(n12891), .ZN(n13317) );
  OR2_X1 U16029 ( .A1(n14163), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U16030 ( .A1(n14150), .A2(n13314), .ZN(n12892) );
  OAI211_X1 U16031 ( .C1(n14158), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12892), .B(
        n14204), .ZN(n12893) );
  AND2_X1 U16032 ( .A1(n12894), .A2(n12893), .ZN(n13316) );
  MUX2_X1 U16033 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12896) );
  NAND2_X1 U16034 ( .A1(n10572), .A2(n14121), .ZN(n12895) );
  AND2_X1 U16035 ( .A1(n12896), .A2(n12895), .ZN(n13337) );
  OR2_X1 U16036 ( .A1(n14163), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n12899) );
  OAI21_X1 U16037 ( .B1(n14164), .B2(n20425), .A(n14150), .ZN(n12897) );
  OAI21_X1 U16038 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n14158), .A(n12897), .ZN(
        n12898) );
  INV_X1 U16039 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U16040 ( .A1(n14113), .A2(n12900), .ZN(n12903) );
  OAI211_X1 U16041 ( .C1(n14164), .C2(n10669), .A(n12901), .B(n14150), .ZN(
        n12902) );
  NAND2_X1 U16042 ( .A1(n12903), .A2(n12902), .ZN(n13543) );
  OR2_X1 U16043 ( .A1(n14163), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12907) );
  OAI21_X1 U16044 ( .B1(n14164), .B2(n12904), .A(n14150), .ZN(n12905) );
  OAI21_X1 U16045 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n14158), .A(n12905), .ZN(
        n12906) );
  INV_X1 U16046 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U16047 ( .A1(n14113), .A2(n13817), .ZN(n12910) );
  OAI211_X1 U16048 ( .C1(n14164), .C2(n10717), .A(n12908), .B(n14150), .ZN(
        n12909) );
  INV_X1 U16049 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16472) );
  OAI21_X1 U16050 ( .B1(n14164), .B2(n16472), .A(n14150), .ZN(n12911) );
  OAI21_X1 U16051 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n14158), .A(n12911), .ZN(
        n12913) );
  OR2_X1 U16052 ( .A1(n14163), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12912) );
  NAND2_X1 U16053 ( .A1(n12913), .A2(n12912), .ZN(n13911) );
  INV_X1 U16054 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20323) );
  NAND2_X1 U16055 ( .A1(n14113), .A2(n20323), .ZN(n12916) );
  OAI211_X1 U16056 ( .C1(n14164), .C2(n14059), .A(n12914), .B(n14150), .ZN(
        n12915) );
  NAND2_X1 U16057 ( .A1(n12916), .A2(n12915), .ZN(n13994) );
  OR2_X1 U16058 ( .A1(n14163), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U16059 ( .A1(n14150), .A2(n12917), .ZN(n12918) );
  OAI211_X1 U16060 ( .C1(n14158), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12918), .B(
        n14204), .ZN(n12919) );
  MUX2_X1 U16061 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12922) );
  OR2_X1 U16062 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U16063 ( .A1(n12922), .A2(n12921), .ZN(n14782) );
  OR2_X1 U16064 ( .A1(n14163), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U16065 ( .A1(n14150), .A2(n15019), .ZN(n12923) );
  OAI211_X1 U16066 ( .C1(n14158), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12923), .B(
        n14204), .ZN(n12924) );
  NAND2_X1 U16067 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  OR2_X1 U16068 ( .A1(n14780), .A2(n12926), .ZN(n12927) );
  NAND2_X1 U16069 ( .A1(n14710), .A2(n12927), .ZN(n14772) );
  OR2_X1 U16070 ( .A1(n12928), .A2(n13635), .ZN(n16276) );
  OAI21_X1 U16071 ( .B1(n12929), .B2(n13412), .A(n16276), .ZN(n12930) );
  INV_X1 U16072 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21001) );
  OAI22_X1 U16073 ( .A1(n14772), .A2(n16466), .B1(n21001), .B2(n20347), .ZN(
        n12932) );
  OR3_X1 U16074 ( .A1(n12934), .A2(n12933), .A3(n12932), .ZN(P1_U3019) );
  INV_X1 U16075 ( .A(n12467), .ZN(n13159) );
  INV_X1 U16076 ( .A(n19277), .ZN(n19457) );
  INV_X1 U16077 ( .A(n20243), .ZN(n20245) );
  OAI21_X1 U16078 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n20245), .A(n12936), 
        .ZN(n19276) );
  NOR3_X1 U16079 ( .A1(n19457), .A2(P2_READREQUEST_REG_SCAN_IN), .A3(n19276), 
        .ZN(n12935) );
  AOI21_X1 U16080 ( .B1(n13159), .B2(n19282), .A(n12935), .ZN(P2_U3612) );
  INV_X1 U16081 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19561) );
  NAND2_X1 U16082 ( .A1(n9779), .A2(n19507), .ZN(n12943) );
  OAI21_X1 U16083 ( .B1(n12298), .B2(n20155), .A(n12937), .ZN(n12956) );
  NAND2_X1 U16084 ( .A1(n12956), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12938) );
  OAI211_X1 U16085 ( .C1(n19561), .C2(n16495), .A(n12943), .B(n12938), .ZN(
        P2_U2981) );
  INV_X1 U16086 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19574) );
  NAND2_X1 U16087 ( .A1(n12968), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12940) );
  INV_X1 U16088 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16852) );
  OR2_X1 U16089 ( .A1(n12968), .A2(n16852), .ZN(n12939) );
  NAND2_X1 U16090 ( .A1(n12940), .A2(n12939), .ZN(n19523) );
  NAND2_X1 U16091 ( .A1(n9779), .A2(n19523), .ZN(n12953) );
  NAND2_X1 U16092 ( .A1(n12956), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12941) );
  OAI211_X1 U16093 ( .C1(n19574), .C2(n16495), .A(n12953), .B(n12941), .ZN(
        P2_U2975) );
  INV_X1 U16094 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13208) );
  NAND2_X1 U16095 ( .A1(n12956), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12942) );
  OAI211_X1 U16096 ( .C1(n13208), .C2(n16495), .A(n12943), .B(n12942), .ZN(
        P2_U2966) );
  INV_X1 U16097 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19569) );
  NAND2_X1 U16098 ( .A1(n12968), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12945) );
  INV_X1 U16099 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16849) );
  OR2_X1 U16100 ( .A1(n16040), .A2(n16849), .ZN(n12944) );
  NAND2_X1 U16101 ( .A1(n12945), .A2(n12944), .ZN(n19517) );
  NAND2_X1 U16102 ( .A1(n9779), .A2(n19517), .ZN(n12948) );
  NAND2_X1 U16103 ( .A1(n12956), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12946) );
  OAI211_X1 U16104 ( .C1(n19569), .C2(n16495), .A(n12948), .B(n12946), .ZN(
        P2_U2977) );
  INV_X1 U16105 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U16106 ( .A1(n12956), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12947) );
  OAI211_X1 U16107 ( .C1(n13205), .C2(n16495), .A(n12948), .B(n12947), .ZN(
        P2_U2962) );
  INV_X1 U16108 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19565) );
  NAND2_X1 U16109 ( .A1(n12968), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12950) );
  INV_X1 U16110 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16845) );
  OR2_X1 U16111 ( .A1(n12968), .A2(n16845), .ZN(n12949) );
  NAND2_X1 U16112 ( .A1(n12950), .A2(n12949), .ZN(n19512) );
  NAND2_X1 U16113 ( .A1(n9779), .A2(n19512), .ZN(n12955) );
  NAND2_X1 U16114 ( .A1(n12956), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12951) );
  OAI211_X1 U16115 ( .C1(n19565), .C2(n16495), .A(n12955), .B(n12951), .ZN(
        P2_U2979) );
  INV_X1 U16116 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U16117 ( .A1(n12956), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12952) );
  OAI211_X1 U16118 ( .C1(n13043), .C2(n16495), .A(n12953), .B(n12952), .ZN(
        P2_U2960) );
  INV_X1 U16119 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U16120 ( .A1(n12956), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12954) );
  OAI211_X1 U16121 ( .C1(n13046), .C2(n16495), .A(n12955), .B(n12954), .ZN(
        P2_U2964) );
  INV_X1 U16122 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12958) );
  INV_X1 U16123 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12957) );
  INV_X1 U16124 ( .A(n12956), .ZN(n12978) );
  INV_X1 U16125 ( .A(n9779), .ZN(n12961) );
  AOI22_X1 U16126 ( .A1(n16042), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16040), .ZN(n19505) );
  OAI222_X1 U16127 ( .A1(n16495), .A2(n12958), .B1(n12957), .B2(n12978), .C1(
        n12961), .C2(n19505), .ZN(P2_U2982) );
  INV_X1 U16128 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12959) );
  OAI22_X1 U16129 ( .A1(n16040), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16042), .ZN(n16037) );
  OAI222_X1 U16130 ( .A1(n13061), .A2(n16495), .B1(n12959), .B2(n12978), .C1(
        n12961), .C2(n16037), .ZN(P2_U2967) );
  INV_X1 U16131 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13200) );
  INV_X1 U16132 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12960) );
  OAI222_X1 U16133 ( .A1(n12961), .A2(n16037), .B1(n16495), .B2(n13200), .C1(
        n12960), .C2(n12978), .ZN(P2_U2952) );
  AND2_X1 U16134 ( .A1(n16245), .A2(n12846), .ZN(n16255) );
  NAND2_X1 U16135 ( .A1(n16255), .A2(n20300), .ZN(n13013) );
  INV_X1 U16136 ( .A(n13013), .ZN(n12963) );
  INV_X1 U16137 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21167) );
  NOR2_X1 U16138 ( .A1(n12928), .A2(n20294), .ZN(n12962) );
  NAND2_X1 U16139 ( .A1(n20907), .A2(n16490), .ZN(n13012) );
  OAI211_X1 U16140 ( .C1(n12963), .C2(n21167), .A(n13595), .B(n13012), .ZN(
        P1_U2801) );
  INV_X1 U16141 ( .A(n12978), .ZN(n13009) );
  AOI22_X1 U16142 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16143 ( .A1(n16042), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16040), .ZN(n19651) );
  INV_X1 U16144 ( .A(n19651), .ZN(n12964) );
  NAND2_X1 U16145 ( .A1(n9779), .A2(n12964), .ZN(n12986) );
  NAND2_X1 U16146 ( .A1(n12965), .A2(n12986), .ZN(P2_U2957) );
  AOI22_X1 U16147 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16148 ( .A1(n16042), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16040), .ZN(n19643) );
  INV_X1 U16149 ( .A(n19643), .ZN(n12966) );
  NAND2_X1 U16150 ( .A1(n9779), .A2(n12966), .ZN(n12998) );
  NAND2_X1 U16151 ( .A1(n12967), .A2(n12998), .ZN(P2_U2955) );
  AOI22_X1 U16152 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12972) );
  INV_X1 U16153 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16843) );
  OR2_X1 U16154 ( .A1(n16040), .A2(n16843), .ZN(n12970) );
  NAND2_X1 U16155 ( .A1(n12968), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12969) );
  AND2_X1 U16156 ( .A1(n12970), .A2(n12969), .ZN(n19510) );
  INV_X1 U16157 ( .A(n19510), .ZN(n12971) );
  NAND2_X1 U16158 ( .A1(n9779), .A2(n12971), .ZN(n13006) );
  NAND2_X1 U16159 ( .A1(n12972), .A2(n13006), .ZN(P2_U2965) );
  AOI22_X1 U16160 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16161 ( .A1(n16042), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16040), .ZN(n19556) );
  INV_X1 U16162 ( .A(n19556), .ZN(n13979) );
  NAND2_X1 U16163 ( .A1(n9779), .A2(n13979), .ZN(n13000) );
  NAND2_X1 U16164 ( .A1(n12973), .A2(n13000), .ZN(P2_U2968) );
  AOI22_X1 U16165 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12977) );
  INV_X1 U16166 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12974) );
  OR2_X1 U16167 ( .A1(n16040), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U16168 ( .A1(n16040), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12975) );
  AND2_X1 U16169 ( .A1(n12976), .A2(n12975), .ZN(n19520) );
  INV_X1 U16170 ( .A(n19520), .ZN(n15353) );
  NAND2_X1 U16171 ( .A1(n9779), .A2(n15353), .ZN(n13002) );
  NAND2_X1 U16172 ( .A1(n12977), .A2(n13002), .ZN(P2_U2961) );
  AOI22_X1 U16173 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12979) );
  OAI22_X1 U16174 ( .A1(n16040), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16042), .ZN(n19638) );
  INV_X1 U16175 ( .A(n19638), .ZN(n16617) );
  NAND2_X1 U16176 ( .A1(n9779), .A2(n16617), .ZN(n12996) );
  NAND2_X1 U16177 ( .A1(n12979), .A2(n12996), .ZN(P2_U2954) );
  AOI22_X1 U16178 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12956), .B1(n13008), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12980) );
  OAI22_X1 U16179 ( .A1(n16040), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16042), .ZN(n19647) );
  INV_X1 U16180 ( .A(n19647), .ZN(n16610) );
  NAND2_X1 U16181 ( .A1(n9779), .A2(n16610), .ZN(n13010) );
  NAND2_X1 U16182 ( .A1(n12980), .A2(n13010), .ZN(P2_U2971) );
  AOI22_X1 U16183 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12981) );
  OAI22_X1 U16184 ( .A1(n16040), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16042), .ZN(n19528) );
  INV_X1 U16185 ( .A(n19528), .ZN(n16603) );
  NAND2_X1 U16186 ( .A1(n9779), .A2(n16603), .ZN(n12988) );
  NAND2_X1 U16187 ( .A1(n12981), .A2(n12988), .ZN(P2_U2958) );
  AOI22_X1 U16188 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12985) );
  INV_X1 U16189 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n12982) );
  OR2_X1 U16190 ( .A1(n16040), .A2(n12982), .ZN(n12984) );
  NAND2_X1 U16191 ( .A1(n16040), .A2(BUF2_REG_7__SCAN_IN), .ZN(n12983) );
  AND2_X1 U16192 ( .A1(n12984), .A2(n12983), .ZN(n19526) );
  INV_X1 U16193 ( .A(n19526), .ZN(n19661) );
  NAND2_X1 U16194 ( .A1(n9779), .A2(n19661), .ZN(n12990) );
  NAND2_X1 U16195 ( .A1(n12985), .A2(n12990), .ZN(P2_U2959) );
  AOI22_X1 U16196 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12956), .B1(n13008), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U16197 ( .A1(n12987), .A2(n12986), .ZN(P2_U2972) );
  AOI22_X1 U16198 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U16199 ( .A1(n12989), .A2(n12988), .ZN(P2_U2973) );
  AOI22_X1 U16200 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U16201 ( .A1(n12991), .A2(n12990), .ZN(P2_U2974) );
  AOI22_X1 U16202 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12995) );
  INV_X1 U16203 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16847) );
  OR2_X1 U16204 ( .A1(n16040), .A2(n16847), .ZN(n12993) );
  NAND2_X1 U16205 ( .A1(n16040), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12992) );
  AND2_X1 U16206 ( .A1(n12993), .A2(n12992), .ZN(n19515) );
  INV_X1 U16207 ( .A(n19515), .ZN(n15339) );
  NAND2_X1 U16208 ( .A1(n9779), .A2(n15339), .ZN(n13004) );
  NAND2_X1 U16209 ( .A1(n12995), .A2(n13004), .ZN(P2_U2963) );
  AOI22_X1 U16210 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12997) );
  NAND2_X1 U16211 ( .A1(n12997), .A2(n12996), .ZN(P2_U2969) );
  AOI22_X1 U16212 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16213 ( .A1(n12999), .A2(n12998), .ZN(P2_U2970) );
  AOI22_X1 U16214 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13001) );
  NAND2_X1 U16215 ( .A1(n13001), .A2(n13000), .ZN(P2_U2953) );
  AOI22_X1 U16216 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U16217 ( .A1(n13003), .A2(n13002), .ZN(P2_U2976) );
  AOI22_X1 U16218 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16219 ( .A1(n13005), .A2(n13004), .ZN(P2_U2978) );
  AOI22_X1 U16220 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13007) );
  NAND2_X1 U16221 ( .A1(n13007), .A2(n13006), .ZN(P2_U2980) );
  AOI22_X1 U16222 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13009), .B1(n13008), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U16223 ( .A1(n13011), .A2(n13010), .ZN(P2_U2956) );
  INV_X1 U16224 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21187) );
  AND2_X1 U16225 ( .A1(n21187), .A2(n13012), .ZN(n13015) );
  OAI21_X1 U16226 ( .B1(n14164), .B2(n16253), .A(n21059), .ZN(n13014) );
  OAI21_X1 U16227 ( .B1(n13015), .B2(n21059), .A(n13014), .ZN(P1_U3487) );
  NAND2_X1 U16228 ( .A1(n16702), .A2(n16070), .ZN(n13143) );
  OR2_X1 U16229 ( .A1(n12448), .A2(n13017), .ZN(n13026) );
  INV_X1 U16230 ( .A(n13016), .ZN(n13025) );
  OR2_X1 U16231 ( .A1(n11925), .A2(n13017), .ZN(n13018) );
  OR2_X1 U16232 ( .A1(n16698), .A2(n13018), .ZN(n13021) );
  INV_X1 U16233 ( .A(n13019), .ZN(n13020) );
  NAND2_X1 U16234 ( .A1(n13021), .A2(n13020), .ZN(n13138) );
  INV_X1 U16235 ( .A(n13138), .ZN(n13022) );
  AND2_X1 U16236 ( .A1(n13023), .A2(n13022), .ZN(n13024) );
  OAI211_X1 U16237 ( .C1(n13143), .C2(n13026), .A(n13025), .B(n13024), .ZN(
        n16715) );
  NAND2_X1 U16238 ( .A1(n16715), .A2(n13144), .ZN(n13028) );
  NAND2_X1 U16239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16025) );
  NOR2_X1 U16240 ( .A1(n16735), .A2(n16025), .ZN(n16740) );
  AOI22_X1 U16241 ( .A1(n16735), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16740), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n13027) );
  AND2_X1 U16242 ( .A1(n13028), .A2(n13027), .ZN(n15986) );
  INV_X1 U16243 ( .A(n15986), .ZN(n16022) );
  NAND2_X1 U16244 ( .A1(n12444), .A2(n13031), .ZN(n13075) );
  NAND2_X1 U16245 ( .A1(n13030), .A2(n13075), .ZN(n16697) );
  OR4_X1 U16246 ( .A1(n15986), .A2(n19283), .A3(n13029), .A4(n16697), .ZN(
        n13032) );
  OAI21_X1 U16247 ( .B1(n12444), .B2(n16022), .A(n13032), .ZN(P2_U3595) );
  INV_X1 U16248 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13037) );
  OR2_X1 U16249 ( .A1(n12448), .A2(n19286), .ZN(n13033) );
  OAI21_X1 U16250 ( .B1(n13143), .B2(n13033), .A(n16495), .ZN(n13034) );
  AND2_X1 U16251 ( .A1(n13034), .A2(n20168), .ZN(n19558) );
  NAND2_X1 U16252 ( .A1(n19558), .A2(n13035), .ZN(n13207) );
  NOR2_X1 U16253 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16025), .ZN(n19589) );
  AOI22_X1 U16254 ( .A1(n19572), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13036) );
  OAI21_X1 U16255 ( .B1(n13037), .B2(n13207), .A(n13036), .ZN(P2_U2933) );
  INV_X1 U16256 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16257 ( .A1(n19572), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16258 ( .B1(n13039), .B2(n13207), .A(n13038), .ZN(P2_U2931) );
  INV_X1 U16259 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16260 ( .A1(n19572), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13040) );
  OAI21_X1 U16261 ( .B1(n13041), .B2(n13207), .A(n13040), .ZN(P2_U2926) );
  AOI22_X1 U16262 ( .A1(n19572), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13042) );
  OAI21_X1 U16263 ( .B1(n13043), .B2(n13207), .A(n13042), .ZN(P2_U2927) );
  AOI22_X1 U16264 ( .A1(n19572), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13044) );
  OAI21_X1 U16265 ( .B1(n15389), .B2(n13207), .A(n13044), .ZN(P2_U2932) );
  AOI22_X1 U16266 ( .A1(n19572), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13045) );
  OAI21_X1 U16267 ( .B1(n13046), .B2(n13207), .A(n13045), .ZN(P2_U2923) );
  INV_X1 U16268 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U16269 ( .A1(n19572), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U16270 ( .B1(n13048), .B2(n13207), .A(n13047), .ZN(P2_U2928) );
  INV_X1 U16271 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16272 ( .A1(n19572), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13049) );
  OAI21_X1 U16273 ( .B1(n13050), .B2(n13207), .A(n13049), .ZN(P2_U2929) );
  INV_X1 U16274 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16275 ( .A1(n19572), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13051) );
  OAI21_X1 U16276 ( .B1(n13052), .B2(n13207), .A(n13051), .ZN(P2_U2924) );
  AOI22_X1 U16277 ( .A1(n19572), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19557), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13053) );
  OAI21_X1 U16278 ( .B1(n15381), .B2(n13207), .A(n13053), .ZN(P2_U2930) );
  NAND2_X1 U16279 ( .A1(n16070), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13054) );
  AND4_X1 U16280 ( .A1(n11844), .A2(n13054), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20153), .ZN(n13055) );
  AOI21_X1 U16281 ( .B1(n16619), .B2(n20276), .A(n19547), .ZN(n13064) );
  XNOR2_X1 U16282 ( .A(n13057), .B(n13056), .ZN(n19445) );
  INV_X1 U16283 ( .A(n16037), .ZN(n19494) );
  INV_X1 U16284 ( .A(n13058), .ZN(n13059) );
  NAND3_X1 U16285 ( .A1(n16619), .A2(n19456), .A3(n19445), .ZN(n13060) );
  OAI21_X1 U16286 ( .B1(n19537), .B2(n13061), .A(n13060), .ZN(n13062) );
  AOI21_X1 U16287 ( .B1(n19494), .B2(n19522), .A(n13062), .ZN(n13063) );
  OAI21_X1 U16288 ( .B1(n13064), .B2(n19445), .A(n13063), .ZN(P2_U2919) );
  INV_X1 U16289 ( .A(n14053), .ZN(n19454) );
  NOR2_X1 U16290 ( .A1(n13065), .A2(n13082), .ZN(n13066) );
  NOR2_X1 U16291 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NOR2_X1 U16292 ( .A1(n13069), .A2(n13068), .ZN(n13071) );
  OR2_X1 U16293 ( .A1(n13071), .A2(n13070), .ZN(n20288) );
  INV_X1 U16294 ( .A(n16696), .ZN(n13179) );
  NAND2_X1 U16295 ( .A1(n13179), .A2(n16726), .ZN(n13172) );
  INV_X1 U16296 ( .A(n16698), .ZN(n13072) );
  OAI21_X1 U16297 ( .B1(n13082), .B2(n13073), .A(n13072), .ZN(n13074) );
  INV_X1 U16298 ( .A(n13074), .ZN(n13077) );
  INV_X1 U16299 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19289) );
  OAI21_X1 U16300 ( .B1(n12478), .B2(n13075), .A(n19289), .ZN(n20273) );
  MUX2_X1 U16301 ( .A(n13077), .B(n20273), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20284) );
  NAND3_X1 U16302 ( .A1(n13179), .A2(n16070), .A3(n20284), .ZN(n13078) );
  OAI21_X1 U16303 ( .B1(n20288), .B2(n13172), .A(n13078), .ZN(n13137) );
  AND2_X1 U16304 ( .A1(n16039), .A2(n13144), .ZN(n13079) );
  NAND2_X1 U16305 ( .A1(n13137), .A2(n13079), .ZN(n19288) );
  INV_X1 U16306 ( .A(n19283), .ZN(n20246) );
  OR2_X1 U16307 ( .A1(n20243), .A2(n20246), .ZN(n20263) );
  NAND2_X1 U16308 ( .A1(n20263), .A2(n16735), .ZN(n13080) );
  NOR2_X1 U16309 ( .A1(n20049), .A2(n20154), .ZN(n20264) );
  MUX2_X1 U16310 ( .A(n13105), .B(n13082), .S(n13081), .Z(n13083) );
  INV_X1 U16311 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U16312 ( .A(n13083), .B(n13094), .S(n14328), .Z(n19446) );
  OR2_X1 U16313 ( .A1(n19446), .A2(n13085), .ZN(n13123) );
  NAND2_X1 U16314 ( .A1(n19446), .A2(n13085), .ZN(n13084) );
  NAND2_X1 U16315 ( .A1(n13123), .A2(n13084), .ZN(n13190) );
  INV_X1 U16316 ( .A(n13190), .ZN(n13092) );
  NOR2_X1 U16317 ( .A1(n9709), .A2(n13085), .ZN(n13114) );
  AOI21_X1 U16318 ( .B1(n9709), .B2(n13085), .A(n13114), .ZN(n13194) );
  INV_X1 U16319 ( .A(n13194), .ZN(n13090) );
  INV_X1 U16320 ( .A(n13086), .ZN(n13088) );
  NAND2_X1 U16321 ( .A1(n20049), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13087) );
  NAND2_X1 U16322 ( .A1(n13088), .A2(n13087), .ZN(n13108) );
  OAI21_X1 U16323 ( .B1(n19593), .B2(n13108), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13089) );
  NAND2_X1 U16324 ( .A1(n19592), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13191) );
  OAI211_X1 U16325 ( .C1(n13090), .C2(n16664), .A(n13089), .B(n13191), .ZN(
        n13091) );
  AOI21_X1 U16326 ( .B1(n19598), .B2(n13092), .A(n13091), .ZN(n13093) );
  OAI21_X1 U16327 ( .B1(n19454), .B2(n15640), .A(n13093), .ZN(P2_U3014) );
  MUX2_X1 U16328 ( .A(n13094), .B(n19454), .S(n19490), .Z(n13095) );
  OAI21_X1 U16329 ( .B1(n19481), .B2(n20276), .A(n13095), .ZN(P2_U2887) );
  OR2_X1 U16330 ( .A1(n13097), .A2(n13096), .ZN(n13099) );
  NOR2_X1 U16331 ( .A1(n19484), .A2(n14031), .ZN(n13100) );
  AOI21_X1 U16332 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n19484), .A(n13100), .ZN(
        n13101) );
  OAI21_X1 U16333 ( .B1(n20265), .B2(n19481), .A(n13101), .ZN(P2_U2886) );
  INV_X1 U16334 ( .A(n13127), .ZN(n13103) );
  NAND3_X1 U16335 ( .A1(n14328), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n13102) );
  NAND2_X1 U16336 ( .A1(n13103), .A2(n13102), .ZN(n14030) );
  NAND2_X1 U16337 ( .A1(n13123), .A2(n14030), .ZN(n13124) );
  OAI21_X1 U16338 ( .B1(n14030), .B2(n13123), .A(n13124), .ZN(n13104) );
  XNOR2_X1 U16339 ( .A(n13104), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19605) );
  XNOR2_X1 U16340 ( .A(n13105), .B(n13117), .ZN(n13113) );
  XOR2_X1 U16341 ( .A(n13113), .B(n13114), .Z(n13106) );
  NAND2_X1 U16342 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13106), .ZN(
        n13115) );
  OAI21_X1 U16343 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13106), .A(
        n13115), .ZN(n19609) );
  AND2_X1 U16344 ( .A1(n19592), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19607) );
  INV_X1 U16345 ( .A(n19607), .ZN(n13107) );
  OAI21_X1 U16346 ( .B1(n16664), .B2(n19609), .A(n13107), .ZN(n13111) );
  INV_X1 U16347 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13109) );
  MUX2_X1 U16348 ( .A(n19593), .B(n16661), .S(n13109), .Z(n13110) );
  AOI211_X1 U16349 ( .C1(n19605), .C2(n19598), .A(n13111), .B(n13110), .ZN(
        n13112) );
  OAI21_X1 U16350 ( .B1(n14031), .B2(n15640), .A(n13112), .ZN(P2_U3013) );
  NAND2_X1 U16351 ( .A1(n13114), .A2(n13113), .ZN(n13116) );
  NAND2_X1 U16352 ( .A1(n13116), .A2(n13115), .ZN(n13762) );
  XNOR2_X1 U16353 ( .A(n13760), .B(n13762), .ZN(n13119) );
  NAND2_X1 U16354 ( .A1(n9709), .A2(n13117), .ZN(n13752) );
  XNOR2_X1 U16355 ( .A(n13751), .B(n13752), .ZN(n13118) );
  NAND2_X1 U16356 ( .A1(n13119), .A2(n13118), .ZN(n13764) );
  OAI21_X1 U16357 ( .B1(n13119), .B2(n13118), .A(n13764), .ZN(n13120) );
  INV_X1 U16358 ( .A(n13120), .ZN(n13177) );
  NAND2_X1 U16359 ( .A1(n19592), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U16360 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13121) );
  OAI211_X1 U16361 ( .C1(n19603), .C2(n13921), .A(n13175), .B(n13121), .ZN(
        n13122) );
  AOI21_X1 U16362 ( .B1(n19595), .B2(n13177), .A(n13122), .ZN(n13131) );
  NOR2_X1 U16363 ( .A1(n13123), .A2(n14030), .ZN(n13125) );
  OAI21_X1 U16364 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13125), .A(
        n13124), .ZN(n13129) );
  OAI21_X1 U16365 ( .B1(n13127), .B2(n13126), .A(n13756), .ZN(n13925) );
  XNOR2_X1 U16366 ( .A(n13925), .B(n13760), .ZN(n13128) );
  OR2_X1 U16367 ( .A1(n13129), .A2(n13128), .ZN(n13759) );
  NAND2_X1 U16368 ( .A1(n13129), .A2(n13128), .ZN(n13180) );
  NAND3_X1 U16369 ( .A1(n13759), .A2(n13180), .A3(n19598), .ZN(n13130) );
  OAI211_X1 U16370 ( .C1(n13929), .C2(n15640), .A(n13131), .B(n13130), .ZN(
        P2_U3012) );
  NAND2_X1 U16371 ( .A1(n13157), .A2(n16694), .ZN(n13142) );
  AOI21_X1 U16372 ( .B1(n13132), .B2(n9670), .A(n13155), .ZN(n13133) );
  NAND2_X1 U16373 ( .A1(n13143), .A2(n13133), .ZN(n13141) );
  MUX2_X1 U16374 ( .A(n11926), .B(n13157), .S(n12298), .Z(n13134) );
  NAND2_X1 U16375 ( .A1(n13134), .A2(n20155), .ZN(n13135) );
  NOR2_X1 U16376 ( .A1(n16698), .A2(n13135), .ZN(n13136) );
  OR2_X1 U16377 ( .A1(n13137), .A2(n13136), .ZN(n13139) );
  NOR2_X1 U16378 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  OAI211_X1 U16379 ( .C1(n13143), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        n13145) );
  NAND2_X1 U16380 ( .A1(n12466), .A2(n16070), .ZN(n13146) );
  AND2_X1 U16381 ( .A1(n13146), .A2(n15990), .ZN(n13147) );
  XNOR2_X1 U16382 ( .A(n13149), .B(n13148), .ZN(n20256) );
  INV_X1 U16383 ( .A(n20256), .ZN(n15397) );
  INV_X1 U16384 ( .A(n13181), .ZN(n13173) );
  AND2_X1 U16385 ( .A1(n13150), .A2(n13173), .ZN(n19613) );
  AND2_X1 U16386 ( .A1(n13152), .A2(n13151), .ZN(n13153) );
  NAND2_X1 U16387 ( .A1(n13154), .A2(n13153), .ZN(n13169) );
  NAND2_X1 U16388 ( .A1(n13156), .A2(n13155), .ZN(n13158) );
  AOI22_X1 U16389 ( .A1(n13159), .A2(n13158), .B1(n16039), .B2(n13157), .ZN(
        n13162) );
  INV_X1 U16390 ( .A(n13160), .ZN(n13161) );
  AND3_X1 U16391 ( .A1(n13163), .A2(n13162), .A3(n13161), .ZN(n13168) );
  NAND2_X1 U16392 ( .A1(n13164), .A2(n16070), .ZN(n14050) );
  NAND2_X1 U16393 ( .A1(n14050), .A2(n13165), .ZN(n13166) );
  NAND2_X1 U16394 ( .A1(n13166), .A2(n11914), .ZN(n13167) );
  NAND3_X1 U16395 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(n16006) );
  NOR2_X1 U16396 ( .A1(n16006), .A2(n13170), .ZN(n13171) );
  NOR2_X1 U16397 ( .A1(n13181), .A2(n13171), .ZN(n15785) );
  NAND2_X1 U16398 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19618) );
  AND2_X1 U16399 ( .A1(n13181), .A2(n19424), .ZN(n19608) );
  AOI21_X1 U16400 ( .B1(n15785), .B2(n19618), .A(n19608), .ZN(n13774) );
  INV_X1 U16401 ( .A(n13172), .ZN(n20289) );
  NAND2_X1 U16402 ( .A1(n15785), .A2(n13760), .ZN(n13770) );
  OR2_X1 U16403 ( .A1(n13770), .A2(n19618), .ZN(n13174) );
  NAND2_X1 U16404 ( .A1(n13175), .A2(n13174), .ZN(n13176) );
  AOI21_X1 U16405 ( .B1(n19611), .B2(n13177), .A(n13176), .ZN(n13187) );
  NAND2_X1 U16406 ( .A1(n13179), .A2(n13178), .ZN(n20285) );
  OR2_X2 U16407 ( .A1(n13181), .A2(n20285), .ZN(n15974) );
  NAND2_X1 U16408 ( .A1(n13759), .A2(n13180), .ZN(n13184) );
  INV_X1 U16409 ( .A(n15991), .ZN(n16701) );
  INV_X1 U16410 ( .A(n19618), .ZN(n13182) );
  NOR2_X1 U16411 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13182), .ZN(
        n13768) );
  INV_X1 U16412 ( .A(n13768), .ZN(n13771) );
  NAND2_X1 U16413 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13182), .ZN(
        n13769) );
  AND2_X1 U16414 ( .A1(n13771), .A2(n13769), .ZN(n13183) );
  OAI22_X1 U16415 ( .A1(n15974), .A2(n13184), .B1(n15782), .B2(n13183), .ZN(
        n13185) );
  INV_X1 U16416 ( .A(n13185), .ZN(n13186) );
  OAI211_X1 U16417 ( .C1(n13774), .C2(n13760), .A(n13187), .B(n13186), .ZN(
        n13188) );
  AOI21_X1 U16418 ( .B1(n19613), .B2(n13702), .A(n13188), .ZN(n13189) );
  OAI21_X1 U16419 ( .B1(n16677), .B2(n15397), .A(n13189), .ZN(P2_U3044) );
  OAI22_X1 U16420 ( .A1(n15974), .A2(n13190), .B1(n16677), .B2(n19445), .ZN(
        n13193) );
  OAI21_X1 U16421 ( .B1(n15927), .B2(n19454), .A(n13191), .ZN(n13192) );
  AOI211_X1 U16422 ( .C1(n19611), .C2(n13194), .A(n13193), .B(n13192), .ZN(
        n13198) );
  INV_X1 U16423 ( .A(n15782), .ZN(n13195) );
  INV_X1 U16424 ( .A(n19608), .ZN(n13196) );
  MUX2_X1 U16425 ( .A(n15786), .B(n13196), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13197) );
  NAND2_X1 U16426 ( .A1(n13198), .A2(n13197), .ZN(P2_U3046) );
  AOI22_X1 U16427 ( .A1(n19589), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13199) );
  OAI21_X1 U16428 ( .B1(n13200), .B2(n13207), .A(n13199), .ZN(P2_U2935) );
  INV_X1 U16429 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U16430 ( .A1(n19589), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13201) );
  OAI21_X1 U16431 ( .B1(n13202), .B2(n13207), .A(n13201), .ZN(P2_U2934) );
  INV_X1 U16432 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15327) );
  AOI22_X1 U16433 ( .A1(n19572), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13203) );
  OAI21_X1 U16434 ( .B1(n15327), .B2(n13207), .A(n13203), .ZN(P2_U2922) );
  AOI22_X1 U16435 ( .A1(n19572), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13204) );
  OAI21_X1 U16436 ( .B1(n13205), .B2(n13207), .A(n13204), .ZN(P2_U2925) );
  AOI22_X1 U16437 ( .A1(n19572), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n19588), .ZN(n13206) );
  OAI21_X1 U16438 ( .B1(n13208), .B2(n13207), .A(n13206), .ZN(P2_U2921) );
  INV_X1 U16439 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13598) );
  INV_X1 U16440 ( .A(n16232), .ZN(n13468) );
  NAND2_X1 U16441 ( .A1(n13468), .A2(n16276), .ZN(n13212) );
  INV_X1 U16442 ( .A(n16254), .ZN(n13209) );
  INV_X1 U16443 ( .A(n16271), .ZN(n13210) );
  NOR2_X1 U16444 ( .A1(n20294), .A2(n13210), .ZN(n13211) );
  NOR2_X1 U16445 ( .A1(n20769), .A2(n16490), .ZN(n13383) );
  NAND2_X1 U16446 ( .A1(n10532), .A2(n13383), .ZN(n20380) );
  INV_X2 U16447 ( .A(n20380), .ZN(n20394) );
  NOR2_X4 U16448 ( .A1(n20381), .A2(n20394), .ZN(n20391) );
  AOI22_X1 U16449 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20391), .B1(n20394), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13214) );
  OAI21_X1 U16450 ( .B1(n13598), .B2(n13368), .A(n13214), .ZN(P1_U2906) );
  INV_X1 U16451 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U16452 ( .A1(n20394), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13215) );
  OAI21_X1 U16453 ( .B1(n13604), .B2(n13368), .A(n13215), .ZN(P1_U2912) );
  AOI22_X1 U16454 ( .A1(n20394), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13216) );
  OAI21_X1 U16455 ( .B1(n14811), .B2(n13368), .A(n13216), .ZN(P1_U2913) );
  AOI22_X1 U16456 ( .A1(n20394), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13217) );
  OAI21_X1 U16457 ( .B1(n14793), .B2(n13368), .A(n13217), .ZN(P1_U2909) );
  AOI22_X1 U16458 ( .A1(n20394), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13218) );
  OAI21_X1 U16459 ( .B1(n14801), .B2(n13368), .A(n13218), .ZN(P1_U2911) );
  INV_X1 U16460 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13601) );
  AOI22_X1 U16461 ( .A1(n20394), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13219) );
  OAI21_X1 U16462 ( .B1(n13601), .B2(n13368), .A(n13219), .ZN(P1_U2908) );
  INV_X1 U16463 ( .A(n13220), .ZN(n13223) );
  OAI21_X1 U16464 ( .B1(n13223), .B2(n13222), .A(n13221), .ZN(n13654) );
  INV_X1 U16465 ( .A(n16364), .ZN(n16371) );
  OR2_X1 U16466 ( .A1(n16351), .A2(n13224), .ZN(n13225) );
  AOI22_X1 U16467 ( .A1(n13225), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n13230) );
  OR2_X1 U16468 ( .A1(n13226), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13228) );
  AND2_X1 U16469 ( .A1(n13228), .A2(n13227), .ZN(n20440) );
  NAND2_X1 U16470 ( .A1(n20440), .A2(n20302), .ZN(n13229) );
  OAI211_X1 U16471 ( .C1(n13654), .C2(n16371), .A(n13230), .B(n13229), .ZN(
        P1_U2999) );
  OAI21_X1 U16472 ( .B1(n13233), .B2(n13232), .A(n13231), .ZN(n13688) );
  XNOR2_X1 U16473 ( .A(n13234), .B(n13311), .ZN(n13288) );
  INV_X1 U16474 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21047) );
  NOR2_X1 U16475 ( .A1(n20347), .A2(n21047), .ZN(n13291) );
  AOI21_X1 U16476 ( .B1(n16351), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13291), .ZN(n13235) );
  OAI21_X1 U16477 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16370), .A(
        n13235), .ZN(n13236) );
  AOI21_X1 U16478 ( .B1(n13288), .B2(n20302), .A(n13236), .ZN(n13237) );
  OAI21_X1 U16479 ( .B1(n13688), .B2(n16371), .A(n13237), .ZN(P1_U2998) );
  INV_X1 U16480 ( .A(n13239), .ZN(n13241) );
  NAND4_X1 U16481 ( .A1(n13241), .A2(n10397), .A3(n11775), .A4(n13240), .ZN(
        n14220) );
  INV_X1 U16482 ( .A(n14220), .ZN(n13242) );
  OR2_X1 U16483 ( .A1(n9669), .A2(n13242), .ZN(n13246) );
  NOR2_X1 U16484 ( .A1(n13243), .A2(n13263), .ZN(n13244) );
  AOI22_X1 U16485 ( .A1(n16232), .A2(n10409), .B1(n13244), .B2(n13260), .ZN(
        n13245) );
  NAND2_X1 U16486 ( .A1(n13246), .A2(n13245), .ZN(n16231) );
  AOI22_X1 U16487 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13311), .B2(n10751), .ZN(
        n13273) );
  NOR2_X1 U16488 ( .A1(n16490), .A2(n20443), .ZN(n13272) );
  INV_X1 U16489 ( .A(n13272), .ZN(n14222) );
  NOR2_X1 U16490 ( .A1(n13273), .A2(n14222), .ZN(n13248) );
  NOR3_X1 U16491 ( .A1(n13243), .A2(n13263), .A3(n13382), .ZN(n13247) );
  AOI211_X1 U16492 ( .C1(n16231), .C2(n21040), .A(n13248), .B(n13247), .ZN(
        n13256) );
  INV_X1 U16493 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20811) );
  OR2_X1 U16494 ( .A1(n16254), .A2(n13261), .ZN(n13281) );
  INV_X1 U16495 ( .A(n13281), .ZN(n13254) );
  INV_X1 U16496 ( .A(n11772), .ZN(n13249) );
  OAI211_X1 U16497 ( .C1(n16232), .C2(n13249), .A(n21064), .B(n16271), .ZN(
        n13251) );
  OAI211_X1 U16498 ( .C1(n16259), .C2(n13418), .A(n13251), .B(n13250), .ZN(
        n13252) );
  INV_X1 U16499 ( .A(n13383), .ZN(n16491) );
  NOR2_X1 U16500 ( .A1(n10532), .A2(n16491), .ZN(n13479) );
  AOI22_X1 U16501 ( .A1(n16230), .A2(n20300), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13479), .ZN(n16482) );
  OAI21_X1 U16502 ( .B1(n20811), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n16482), 
        .ZN(n21045) );
  NAND2_X1 U16503 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21043), .ZN(
        n13255) );
  OAI21_X1 U16504 ( .B1(n13256), .B2(n21043), .A(n13255), .ZN(P1_U3473) );
  INV_X1 U16505 ( .A(n13257), .ZN(n20459) );
  NOR3_X1 U16506 ( .A1(n13468), .A2(n13458), .A3(n13258), .ZN(n13268) );
  AND2_X1 U16507 ( .A1(n13260), .A2(n13259), .ZN(n13462) );
  NAND2_X1 U16508 ( .A1(n16247), .A2(n13261), .ZN(n13464) );
  INV_X1 U16509 ( .A(n13262), .ZN(n13266) );
  INV_X1 U16510 ( .A(n13263), .ZN(n13265) );
  NAND2_X1 U16511 ( .A1(n13265), .A2(n13264), .ZN(n13459) );
  NAND2_X1 U16512 ( .A1(n13266), .A2(n13459), .ZN(n13270) );
  MUX2_X1 U16513 ( .A(n13462), .B(n13464), .S(n13270), .Z(n13267) );
  AOI211_X1 U16514 ( .C1(n20459), .C2(n14220), .A(n13268), .B(n13267), .ZN(
        n13269) );
  INV_X1 U16515 ( .A(n13269), .ZN(n13457) );
  INV_X1 U16516 ( .A(n13382), .ZN(n21038) );
  INV_X1 U16517 ( .A(n13270), .ZN(n13271) );
  AOI222_X1 U16518 ( .A1(n13457), .A2(n21040), .B1(n13273), .B2(n13272), .C1(
        n21038), .C2(n13271), .ZN(n13275) );
  NAND2_X1 U16519 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21043), .ZN(
        n13274) );
  OAI21_X1 U16520 ( .B1(n13275), .B2(n21043), .A(n13274), .ZN(P1_U3472) );
  NAND2_X1 U16521 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  INV_X1 U16522 ( .A(n20258), .ZN(n16002) );
  MUX2_X1 U16523 ( .A(n13924), .B(n13929), .S(n19490), .Z(n13280) );
  OAI21_X1 U16524 ( .B1(n16002), .B2(n19481), .A(n13280), .ZN(P2_U2885) );
  AOI22_X1 U16525 ( .A1(n14784), .A2(n13686), .B1(n14783), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13287) );
  OAI21_X1 U16526 ( .B1(n13688), .B2(n14769), .A(n13287), .ZN(P1_U2871) );
  INV_X1 U16527 ( .A(n13288), .ZN(n13295) );
  OAI21_X1 U16528 ( .B1(n20442), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16445), .ZN(n20446) );
  INV_X1 U16529 ( .A(n20446), .ZN(n13289) );
  NOR2_X1 U16530 ( .A1(n13289), .A2(n13311), .ZN(n13290) );
  AOI211_X1 U16531 ( .C1(n20438), .C2(n13686), .A(n13291), .B(n13290), .ZN(
        n13294) );
  INV_X1 U16532 ( .A(n16416), .ZN(n15041) );
  OR3_X1 U16533 ( .A1(n15041), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13292), .ZN(n13293) );
  OAI211_X1 U16534 ( .C1(n13295), .C2(n20431), .A(n13294), .B(n13293), .ZN(
        P1_U3030) );
  NAND2_X1 U16535 ( .A1(n14121), .A2(n20443), .ZN(n13297) );
  AND2_X1 U16536 ( .A1(n13297), .A2(n13296), .ZN(n20437) );
  INV_X1 U16537 ( .A(n20437), .ZN(n13298) );
  INV_X1 U16538 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13647) );
  OAI222_X1 U16539 ( .A1(n13298), .A2(n14765), .B1(n14770), .B2(n13647), .C1(
        n13654), .C2(n14769), .ZN(P1_U2872) );
  NAND2_X1 U16540 ( .A1(n13299), .A2(n14198), .ZN(n13300) );
  NAND2_X1 U16541 ( .A1(n13386), .A2(DATAI_0_), .ZN(n13302) );
  NAND2_X1 U16542 ( .A1(n13623), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13301) );
  AND2_X1 U16543 ( .A1(n13302), .A2(n13301), .ZN(n13826) );
  INV_X1 U16544 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20409) );
  OAI222_X1 U16545 ( .A1(n13654), .A2(n14869), .B1(n14868), .B2(n13826), .C1(
        n14865), .C2(n20409), .ZN(P1_U2904) );
  NAND2_X1 U16546 ( .A1(n13386), .A2(DATAI_1_), .ZN(n13304) );
  NAND2_X1 U16547 ( .A1(n13623), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13303) );
  AND2_X1 U16548 ( .A1(n13304), .A2(n13303), .ZN(n14841) );
  INV_X1 U16549 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20406) );
  OAI222_X1 U16550 ( .A1(n13688), .A2(n14869), .B1(n14868), .B2(n14841), .C1(
        n14865), .C2(n20406), .ZN(P1_U2903) );
  NOR2_X1 U16551 ( .A1(n13785), .A2(n19484), .ZN(n13308) );
  AOI21_X1 U16552 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19484), .A(n13308), .ZN(
        n13309) );
  OAI21_X1 U16553 ( .B1(n20248), .B2(n19481), .A(n13309), .ZN(P2_U2884) );
  NOR2_X1 U16554 ( .A1(n20443), .A2(n13311), .ZN(n13312) );
  AOI22_X1 U16555 ( .A1(n13312), .A2(n15151), .B1(n13311), .B2(n15154), .ZN(
        n13313) );
  AOI21_X1 U16556 ( .B1(n16445), .B2(n13313), .A(n13314), .ZN(n13321) );
  AND3_X1 U16557 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15022), .A3(
        n13314), .ZN(n13320) );
  INV_X1 U16558 ( .A(n13372), .ZN(n13315) );
  NOR2_X1 U16559 ( .A1(n20442), .A2(n13315), .ZN(n13375) );
  AND2_X1 U16560 ( .A1(n13317), .A2(n13316), .ZN(n13318) );
  OR2_X1 U16561 ( .A1(n13338), .A2(n13318), .ZN(n13676) );
  INV_X1 U16562 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20981) );
  OAI22_X1 U16563 ( .A1(n16466), .A2(n13676), .B1(n20981), .B2(n20347), .ZN(
        n13319) );
  NOR4_X1 U16564 ( .A1(n13321), .A2(n13320), .A3(n13375), .A4(n13319), .ZN(
        n13322) );
  OAI21_X1 U16565 ( .B1(n20431), .B2(n13336), .A(n13322), .ZN(P1_U3029) );
  OAI21_X1 U16566 ( .B1(n13325), .B2(n13324), .A(n13323), .ZN(n13451) );
  NAND2_X1 U16567 ( .A1(n13386), .A2(DATAI_3_), .ZN(n13327) );
  NAND2_X1 U16568 ( .A1(n13623), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13326) );
  AND2_X1 U16569 ( .A1(n13327), .A2(n13326), .ZN(n13822) );
  INV_X1 U16570 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20402) );
  OAI222_X1 U16571 ( .A1(n13451), .A2(n14869), .B1(n14868), .B2(n13822), .C1(
        n14865), .C2(n20402), .ZN(P1_U2901) );
  INV_X1 U16572 ( .A(n13328), .ZN(n13329) );
  AOI21_X1 U16573 ( .B1(n13330), .B2(n13231), .A(n13329), .ZN(n13671) );
  INV_X1 U16574 ( .A(n13671), .ZN(n13353) );
  INV_X1 U16575 ( .A(n13676), .ZN(n13331) );
  AOI22_X1 U16576 ( .A1(n14784), .A2(n13331), .B1(n14783), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13332) );
  OAI21_X1 U16577 ( .B1(n13353), .B2(n14769), .A(n13332), .ZN(P1_U2870) );
  AOI22_X1 U16578 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16579 ( .B1(n13674), .B2(n16370), .A(n13333), .ZN(n13334) );
  AOI21_X1 U16580 ( .B1(n13671), .B2(n16364), .A(n13334), .ZN(n13335) );
  OAI21_X1 U16581 ( .B1(n16349), .B2(n13336), .A(n13335), .ZN(P1_U2997) );
  OR2_X1 U16582 ( .A1(n13338), .A2(n13337), .ZN(n13339) );
  NAND2_X1 U16583 ( .A1(n13545), .A2(n13339), .ZN(n20376) );
  INV_X1 U16584 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13340) );
  OAI222_X1 U16585 ( .A1(n20376), .A2(n14765), .B1(n14770), .B2(n13340), .C1(
        n14769), .C2(n13451), .ZN(P1_U2869) );
  XNOR2_X1 U16586 ( .A(n13342), .B(n13341), .ZN(n20270) );
  INV_X1 U16587 ( .A(n20270), .ZN(n13343) );
  NAND2_X1 U16588 ( .A1(n20265), .A2(n13343), .ZN(n13344) );
  OAI21_X1 U16589 ( .B1(n20265), .B2(n13343), .A(n13344), .ZN(n19549) );
  NOR2_X1 U16590 ( .A1(n20276), .A2(n19445), .ZN(n19550) );
  NOR2_X1 U16591 ( .A1(n19549), .A2(n19550), .ZN(n19548) );
  INV_X1 U16592 ( .A(n13344), .ZN(n13345) );
  NOR2_X1 U16593 ( .A1(n19548), .A2(n13345), .ZN(n13347) );
  XNOR2_X1 U16594 ( .A(n20258), .B(n20256), .ZN(n13346) );
  NOR2_X1 U16595 ( .A1(n13346), .A2(n13347), .ZN(n15396) );
  AOI21_X1 U16596 ( .B1(n13347), .B2(n13346), .A(n15396), .ZN(n13350) );
  AOI22_X1 U16597 ( .A1(n19522), .A2(n16617), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19546), .ZN(n13349) );
  NAND2_X1 U16598 ( .A1(n20256), .A2(n19547), .ZN(n13348) );
  OAI211_X1 U16599 ( .C1(n13350), .C2(n19551), .A(n13349), .B(n13348), .ZN(
        P2_U2917) );
  NAND2_X1 U16600 ( .A1(n13386), .A2(DATAI_2_), .ZN(n13352) );
  NAND2_X1 U16601 ( .A1(n13623), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13351) );
  AND2_X1 U16602 ( .A1(n13352), .A2(n13351), .ZN(n14835) );
  INV_X1 U16603 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20404) );
  OAI222_X1 U16604 ( .A1(n13353), .A2(n14869), .B1(n14868), .B2(n14835), .C1(
        n14865), .C2(n20404), .ZN(P1_U2902) );
  INV_X1 U16605 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U16606 ( .A1(n20394), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13354) );
  OAI21_X1 U16607 ( .B1(n13355), .B2(n13368), .A(n13354), .ZN(P1_U2915) );
  INV_X1 U16608 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13357) );
  AOI22_X1 U16609 ( .A1(n20394), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16610 ( .B1(n13357), .B2(n13368), .A(n13356), .ZN(P1_U2916) );
  INV_X1 U16611 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U16612 ( .A1(n20394), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13358) );
  OAI21_X1 U16613 ( .B1(n13359), .B2(n13368), .A(n13358), .ZN(P1_U2917) );
  INV_X1 U16614 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U16615 ( .A1(n20394), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13360) );
  OAI21_X1 U16616 ( .B1(n13361), .B2(n13368), .A(n13360), .ZN(P1_U2920) );
  INV_X1 U16617 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U16618 ( .A1(n20394), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13362) );
  OAI21_X1 U16619 ( .B1(n13363), .B2(n13368), .A(n13362), .ZN(P1_U2914) );
  AOI22_X1 U16620 ( .A1(n20394), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13364) );
  OAI21_X1 U16621 ( .B1(n14786), .B2(n13368), .A(n13364), .ZN(P1_U2907) );
  INV_X1 U16622 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U16623 ( .A1(n20394), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U16624 ( .B1(n13617), .B2(n13368), .A(n13365), .ZN(P1_U2910) );
  AOI22_X1 U16625 ( .A1(n20394), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13366) );
  OAI21_X1 U16626 ( .B1(n14839), .B2(n13368), .A(n13366), .ZN(P1_U2919) );
  AOI22_X1 U16627 ( .A1(n20394), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13367) );
  OAI21_X1 U16628 ( .B1(n14834), .B2(n13368), .A(n13367), .ZN(P1_U2918) );
  XNOR2_X1 U16629 ( .A(n13370), .B(n13369), .ZN(n13456) );
  NOR2_X1 U16630 ( .A1(n13372), .A2(n13371), .ZN(n20424) );
  INV_X1 U16631 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13373) );
  OR2_X1 U16632 ( .A1(n20347), .A2(n13373), .ZN(n13453) );
  OAI21_X1 U16633 ( .B1(n16466), .B2(n20376), .A(n13453), .ZN(n13377) );
  OAI21_X1 U16634 ( .B1(n16447), .B2(n13374), .A(n16445), .ZN(n13665) );
  NOR2_X1 U16635 ( .A1(n13665), .A2(n13375), .ZN(n20426) );
  NOR2_X1 U16636 ( .A1(n20426), .A2(n10572), .ZN(n13376) );
  AOI211_X1 U16637 ( .C1(n20424), .C2(n10572), .A(n13377), .B(n13376), .ZN(
        n13378) );
  OAI21_X1 U16638 ( .B1(n20431), .B2(n13456), .A(n13378), .ZN(P1_U3028) );
  OR2_X1 U16639 ( .A1(n13553), .A2(n20901), .ZN(n13379) );
  NAND2_X1 U16640 ( .A1(n21129), .A2(n20907), .ZN(n13496) );
  NAND2_X1 U16641 ( .A1(n13379), .A2(n13496), .ZN(n20771) );
  INV_X1 U16642 ( .A(n20771), .ZN(n20900) );
  OAI21_X1 U16643 ( .B1(n20576), .B2(n20901), .A(n20900), .ZN(n13385) );
  OR2_X1 U16644 ( .A1(n13257), .A2(n13475), .ZN(n20631) );
  NAND2_X1 U16645 ( .A1(n14221), .A2(n13380), .ZN(n20767) );
  INV_X1 U16646 ( .A(n20767), .ZN(n20895) );
  INV_X1 U16647 ( .A(n13433), .ZN(n13381) );
  AOI21_X1 U16648 ( .B1(n20604), .B2(n20895), .A(n13381), .ZN(n13388) );
  NOR2_X1 U16649 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21068) );
  OAI21_X1 U16650 ( .B1(n20907), .B2(n13389), .A(n20906), .ZN(n13384) );
  NOR2_X2 U16651 ( .A1(n20609), .A2(n20860), .ZN(n20656) );
  INV_X1 U16652 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16822) );
  INV_X1 U16653 ( .A(DATAI_24_), .ZN(n21195) );
  OAI22_X1 U16654 ( .A1(n16822), .A2(n13436), .B1(n21195), .B2(n13437), .ZN(
        n20909) );
  NAND2_X1 U16655 ( .A1(n13432), .A2(n13213), .ZN(n20723) );
  INV_X1 U16656 ( .A(n13388), .ZN(n13390) );
  AOI22_X1 U16657 ( .A1(n13390), .A2(n20907), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13389), .ZN(n13434) );
  INV_X1 U16658 ( .A(n20898), .ZN(n20819) );
  OAI22_X1 U16659 ( .A1(n20723), .A2(n13433), .B1(n13434), .B2(n20819), .ZN(
        n13391) );
  AOI21_X1 U16660 ( .B1(n20656), .B2(n20909), .A(n13391), .ZN(n13393) );
  NOR2_X2 U16661 ( .A1(n20609), .A2(n20777), .ZN(n20686) );
  INV_X1 U16662 ( .A(DATAI_16_), .ZN(n21171) );
  INV_X1 U16663 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16838) );
  OAI22_X1 U16664 ( .A1(n21171), .A2(n13437), .B1(n16838), .B2(n13436), .ZN(
        n20810) );
  NAND2_X1 U16665 ( .A1(n20686), .A2(n9778), .ZN(n13392) );
  OAI211_X1 U16666 ( .C1(n13441), .C2(n13394), .A(n13393), .B(n13392), .ZN(
        P1_U3089) );
  INV_X1 U16667 ( .A(DATAI_25_), .ZN(n21210) );
  INV_X1 U16668 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16820) );
  OAI22_X1 U16669 ( .A1(n21210), .A2(n13437), .B1(n16820), .B2(n13436), .ZN(
        n20914) );
  NAND2_X1 U16670 ( .A1(n13432), .A2(n13635), .ZN(n20820) );
  OAI22_X1 U16671 ( .A1(n20820), .A2(n13433), .B1(n13434), .B2(n20826), .ZN(
        n13395) );
  AOI21_X1 U16672 ( .B1(n20656), .B2(n20914), .A(n13395), .ZN(n13397) );
  INV_X1 U16673 ( .A(DATAI_17_), .ZN(n21147) );
  INV_X1 U16674 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16836) );
  OAI22_X1 U16675 ( .A1(n21147), .A2(n13437), .B1(n16836), .B2(n13436), .ZN(
        n20823) );
  NAND2_X1 U16676 ( .A1(n20686), .A2(n20823), .ZN(n13396) );
  OAI211_X1 U16677 ( .C1(n13441), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        P1_U3090) );
  INV_X1 U16678 ( .A(DATAI_31_), .ZN(n21151) );
  OAI22_X1 U16679 ( .A1(n16808), .A2(n13436), .B1(n21151), .B2(n13437), .ZN(
        n20954) );
  INV_X1 U16680 ( .A(DATAI_7_), .ZN(n13400) );
  NAND2_X1 U16681 ( .A1(n13623), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13399) );
  OAI21_X1 U16682 ( .B1(n13623), .B2(n13400), .A(n13399), .ZN(n14813) );
  INV_X1 U16683 ( .A(n14813), .ZN(n13812) );
  INV_X1 U16684 ( .A(n20951), .ZN(n20858) );
  NAND2_X1 U16685 ( .A1(n13432), .A2(n14198), .ZN(n20756) );
  OAI22_X1 U16686 ( .A1(n20858), .A2(n13434), .B1(n13433), .B2(n20756), .ZN(
        n13401) );
  AOI21_X1 U16687 ( .B1(n20954), .B2(n20656), .A(n13401), .ZN(n13403) );
  INV_X1 U16688 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16824) );
  INV_X1 U16689 ( .A(DATAI_23_), .ZN(n21218) );
  NAND2_X1 U16690 ( .A1(n20686), .A2(n20852), .ZN(n13402) );
  OAI211_X1 U16691 ( .C1(n13441), .C2(n13404), .A(n13403), .B(n13402), .ZN(
        P1_U3096) );
  INV_X1 U16692 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16816) );
  INV_X1 U16693 ( .A(DATAI_27_), .ZN(n21149) );
  OAI22_X1 U16694 ( .A1(n16816), .A2(n13436), .B1(n21149), .B2(n13437), .ZN(
        n20926) );
  NAND2_X1 U16695 ( .A1(n13432), .A2(n13405), .ZN(n20739) );
  INV_X1 U16696 ( .A(n20924), .ZN(n20835) );
  OAI22_X1 U16697 ( .A1(n20739), .A2(n13433), .B1(n13434), .B2(n20835), .ZN(
        n13406) );
  AOI21_X1 U16698 ( .B1(n20656), .B2(n20926), .A(n13406), .ZN(n13408) );
  INV_X1 U16699 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16832) );
  INV_X1 U16700 ( .A(DATAI_19_), .ZN(n21214) );
  OAI22_X1 U16701 ( .A1(n16832), .A2(n13436), .B1(n21214), .B2(n13437), .ZN(
        n20832) );
  NAND2_X1 U16702 ( .A1(n20832), .A2(n20686), .ZN(n13407) );
  OAI211_X1 U16703 ( .C1(n13441), .C2(n13409), .A(n13408), .B(n13407), .ZN(
        P1_U3092) );
  INV_X1 U16704 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16814) );
  INV_X1 U16705 ( .A(DATAI_28_), .ZN(n21119) );
  OAI22_X1 U16706 ( .A1(n16814), .A2(n13436), .B1(n21119), .B2(n13437), .ZN(
        n20932) );
  INV_X1 U16707 ( .A(DATAI_4_), .ZN(n13411) );
  INV_X1 U16708 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13410) );
  MUX2_X1 U16709 ( .A(n13411), .B(n13410), .S(n13623), .Z(n14825) );
  INV_X1 U16710 ( .A(n20930), .ZN(n20839) );
  NAND2_X1 U16711 ( .A1(n13432), .A2(n13412), .ZN(n20743) );
  OAI22_X1 U16712 ( .A1(n20839), .A2(n13434), .B1(n13433), .B2(n20743), .ZN(
        n13413) );
  AOI21_X1 U16713 ( .B1(n20932), .B2(n20656), .A(n13413), .ZN(n13416) );
  INV_X1 U16714 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16830) );
  INV_X1 U16715 ( .A(DATAI_20_), .ZN(n13414) );
  NAND2_X1 U16716 ( .A1(n20686), .A2(n20836), .ZN(n13415) );
  OAI211_X1 U16717 ( .C1(n13441), .C2(n13417), .A(n13416), .B(n13415), .ZN(
        P1_U3093) );
  INV_X1 U16718 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16818) );
  INV_X1 U16719 ( .A(DATAI_26_), .ZN(n21237) );
  OAI22_X1 U16720 ( .A1(n16818), .A2(n13436), .B1(n21237), .B2(n13437), .ZN(
        n20876) );
  NAND2_X1 U16721 ( .A1(n13432), .A2(n13418), .ZN(n20827) );
  INV_X1 U16722 ( .A(n20918), .ZN(n20831) );
  OAI22_X1 U16723 ( .A1(n20827), .A2(n13433), .B1(n13434), .B2(n20831), .ZN(
        n13419) );
  AOI21_X1 U16724 ( .B1(n20656), .B2(n20876), .A(n13419), .ZN(n13422) );
  INV_X1 U16725 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16834) );
  INV_X1 U16726 ( .A(DATAI_18_), .ZN(n13420) );
  OAI22_X1 U16727 ( .A1(n16834), .A2(n13436), .B1(n13420), .B2(n13437), .ZN(
        n20920) );
  NAND2_X1 U16728 ( .A1(n20686), .A2(n9774), .ZN(n13421) );
  OAI211_X1 U16729 ( .C1(n13441), .C2(n10354), .A(n13422), .B(n13421), .ZN(
        P1_U3091) );
  INV_X1 U16730 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16812) );
  INV_X1 U16731 ( .A(DATAI_29_), .ZN(n21170) );
  OAI22_X1 U16732 ( .A1(n16812), .A2(n13436), .B1(n21170), .B2(n13437), .ZN(
        n20938) );
  INV_X1 U16733 ( .A(DATAI_5_), .ZN(n13424) );
  INV_X1 U16734 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13423) );
  MUX2_X1 U16735 ( .A(n13424), .B(n13423), .S(n13623), .Z(n14820) );
  INV_X1 U16736 ( .A(n20936), .ZN(n20843) );
  NAND2_X1 U16737 ( .A1(n13432), .A2(n10397), .ZN(n20747) );
  OAI22_X1 U16738 ( .A1(n20843), .A2(n13434), .B1(n13433), .B2(n20747), .ZN(
        n13425) );
  AOI21_X1 U16739 ( .B1(n20938), .B2(n20656), .A(n13425), .ZN(n13428) );
  INV_X1 U16740 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16828) );
  INV_X1 U16741 ( .A(DATAI_21_), .ZN(n13426) );
  NAND2_X1 U16742 ( .A1(n20840), .A2(n20686), .ZN(n13427) );
  OAI211_X1 U16743 ( .C1(n13441), .C2(n13429), .A(n13428), .B(n13427), .ZN(
        P1_U3094) );
  INV_X1 U16744 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16810) );
  INV_X1 U16745 ( .A(DATAI_30_), .ZN(n21115) );
  OAI22_X1 U16746 ( .A1(n16810), .A2(n13436), .B1(n21115), .B2(n13437), .ZN(
        n20885) );
  INV_X1 U16747 ( .A(DATAI_6_), .ZN(n13431) );
  NAND2_X1 U16748 ( .A1(n13623), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U16749 ( .B1(n13623), .B2(n13431), .A(n13430), .ZN(n14817) );
  INV_X1 U16750 ( .A(n14817), .ZN(n13657) );
  NAND2_X1 U16751 ( .A1(n13432), .A2(n10421), .ZN(n20845) );
  OAI22_X1 U16752 ( .A1(n20850), .A2(n13434), .B1(n13433), .B2(n20845), .ZN(
        n13435) );
  AOI21_X1 U16753 ( .B1(n20885), .B2(n20656), .A(n13435), .ZN(n13439) );
  INV_X1 U16754 ( .A(DATAI_22_), .ZN(n21217) );
  INV_X1 U16755 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16826) );
  OAI22_X1 U16756 ( .A1(n21217), .A2(n13437), .B1(n16826), .B2(n13436), .ZN(
        n20944) );
  NAND2_X1 U16757 ( .A1(n20686), .A2(n9776), .ZN(n13438) );
  OAI211_X1 U16758 ( .C1(n13441), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        P1_U3095) );
  NOR2_X1 U16759 ( .A1(n13443), .A2(n13442), .ZN(n13883) );
  NAND2_X1 U16760 ( .A1(n13444), .A2(n13883), .ZN(n13888) );
  XOR2_X1 U16761 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13888), .Z(n13450)
         );
  NAND2_X1 U16762 ( .A1(n13445), .A2(n13895), .ZN(n13447) );
  INV_X1 U16763 ( .A(n13524), .ZN(n13446) );
  AND2_X1 U16764 ( .A1(n13447), .A2(n13446), .ZN(n19436) );
  INV_X1 U16765 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19428) );
  NOR2_X1 U16766 ( .A1(n19490), .A2(n19428), .ZN(n13448) );
  AOI21_X1 U16767 ( .B1(n19436), .B2(n19490), .A(n13448), .ZN(n13449) );
  OAI21_X1 U16768 ( .B1(n13450), .B2(n19481), .A(n13449), .ZN(P2_U2882) );
  INV_X1 U16769 ( .A(n13451), .ZN(n20373) );
  NAND2_X1 U16770 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13452) );
  OAI211_X1 U16771 ( .C1(n16370), .C2(n20362), .A(n13453), .B(n13452), .ZN(
        n13454) );
  AOI21_X1 U16772 ( .B1(n20373), .B2(n16364), .A(n13454), .ZN(n13455) );
  OAI21_X1 U16773 ( .B1(n16349), .B2(n13456), .A(n13455), .ZN(P1_U2996) );
  NOR2_X1 U16774 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16490), .ZN(n13472) );
  MUX2_X1 U16775 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13457), .S(
        n16230), .Z(n16239) );
  AOI22_X1 U16776 ( .A1(n13472), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16490), .B2(n16239), .ZN(n13474) );
  XNOR2_X1 U16777 ( .A(n13458), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13467) );
  NAND2_X1 U16778 ( .A1(n20663), .A2(n14220), .ZN(n13466) );
  XNOR2_X1 U16779 ( .A(n13459), .B(n13461), .ZN(n13463) );
  OAI21_X1 U16780 ( .B1(n13262), .B2(n13461), .A(n9657), .ZN(n21039) );
  AOI22_X1 U16781 ( .A1(n13464), .A2(n13463), .B1(n13462), .B2(n21039), .ZN(
        n13465) );
  OAI211_X1 U16782 ( .C1(n13468), .C2(n13467), .A(n13466), .B(n13465), .ZN(
        n21041) );
  NAND2_X1 U16783 ( .A1(n21041), .A2(n16230), .ZN(n13471) );
  INV_X1 U16784 ( .A(n16230), .ZN(n13469) );
  NAND2_X1 U16785 ( .A1(n13469), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13470) );
  NAND2_X1 U16786 ( .A1(n13471), .A2(n13470), .ZN(n16240) );
  AOI22_X1 U16787 ( .A1(n16240), .A2(n16490), .B1(n13472), .B2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13473) );
  NOR2_X1 U16788 ( .A1(n10542), .A2(n9826), .ZN(n13476) );
  XOR2_X1 U16789 ( .A(n16486), .B(n13476), .Z(n20350) );
  NOR2_X1 U16790 ( .A1(n20350), .A2(n11775), .ZN(n16484) );
  NAND2_X1 U16791 ( .A1(n16230), .A2(n16490), .ZN(n13478) );
  OAI21_X1 U16792 ( .B1(n16486), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13478), .ZN(
        n13477) );
  OAI21_X1 U16793 ( .B1(n16484), .B2(n13478), .A(n13477), .ZN(n16267) );
  OAI21_X1 U16794 ( .B1(n16244), .B2(n13243), .A(n16267), .ZN(n13509) );
  OAI21_X1 U16795 ( .B1(n13509), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13479), .ZN(
        n13480) );
  NAND2_X1 U16796 ( .A1(n13480), .A2(n20582), .ZN(n20450) );
  NAND2_X1 U16797 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20811), .ZN(n13497) );
  INV_X1 U16798 ( .A(n13497), .ZN(n13510) );
  OAI21_X1 U16799 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13553), .A(n20771), 
        .ZN(n13481) );
  OAI21_X1 U16800 ( .B1(n13510), .B2(n9669), .A(n13481), .ZN(n13482) );
  NAND2_X1 U16801 ( .A1(n20450), .A2(n13482), .ZN(n13483) );
  OAI21_X1 U16802 ( .B1(n20450), .B2(n20522), .A(n13483), .ZN(P1_U3477) );
  INV_X1 U16803 ( .A(n13485), .ZN(n13488) );
  INV_X1 U16804 ( .A(n13486), .ZN(n13487) );
  OAI211_X1 U16805 ( .C1(n10051), .C2(n13488), .A(n13487), .B(n19487), .ZN(
        n13492) );
  OR2_X1 U16806 ( .A1(n13489), .A2(n13873), .ZN(n13490) );
  AND2_X1 U16807 ( .A1(n13490), .A2(n15890), .ZN(n19397) );
  NAND2_X1 U16808 ( .A1(n19490), .A2(n19397), .ZN(n13491) );
  OAI211_X1 U16809 ( .C1(n19490), .C2(n13493), .A(n13492), .B(n13491), .ZN(
        P2_U2878) );
  INV_X1 U16810 ( .A(n13553), .ZN(n13504) );
  MUX2_X1 U16811 ( .A(n20609), .B(n13554), .S(n13504), .Z(n13495) );
  NAND2_X1 U16812 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20907), .ZN(n13503) );
  AOI21_X1 U16813 ( .B1(n20778), .B2(n13495), .A(n13503), .ZN(n13501) );
  INV_X1 U16814 ( .A(n13496), .ZN(n20804) );
  AOI22_X1 U16815 ( .A1(n13498), .A2(n20804), .B1(n13497), .B2(n20663), .ZN(
        n13499) );
  INV_X1 U16816 ( .A(n13499), .ZN(n13500) );
  OAI21_X1 U16817 ( .B1(n13501), .B2(n13500), .A(n20450), .ZN(n13502) );
  OAI21_X1 U16818 ( .B1(n20450), .B2(n20862), .A(n13502), .ZN(P1_U3475) );
  NOR2_X1 U16819 ( .A1(n13257), .A2(n13510), .ZN(n13507) );
  NOR2_X1 U16820 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  MUX2_X1 U16821 ( .A(n20771), .B(n13505), .S(n20453), .Z(n13506) );
  OAI21_X1 U16822 ( .B1(n13507), .B2(n13506), .A(n20450), .ZN(n13508) );
  OAI21_X1 U16823 ( .B1(n20450), .B2(n20722), .A(n13508), .ZN(P1_U3476) );
  NOR2_X1 U16824 ( .A1(n13509), .A2(n16491), .ZN(n16281) );
  INV_X1 U16825 ( .A(n14221), .ZN(n13511) );
  OAI22_X1 U16826 ( .A1(n13551), .A2(n20901), .B1(n13511), .B2(n13510), .ZN(
        n13512) );
  OAI21_X1 U16827 ( .B1(n16281), .B2(n13512), .A(n20450), .ZN(n13513) );
  OAI21_X1 U16828 ( .B1(n20450), .B2(n20690), .A(n13513), .ZN(P1_U3478) );
  INV_X1 U16829 ( .A(n13514), .ZN(n13515) );
  NOR2_X1 U16830 ( .A1(n13888), .A2(n13515), .ZN(n19480) );
  XNOR2_X1 U16831 ( .A(n19480), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13520) );
  NAND2_X1 U16832 ( .A1(n13516), .A2(n13526), .ZN(n13518) );
  INV_X1 U16833 ( .A(n13871), .ZN(n13517) );
  NAND2_X1 U16834 ( .A1(n13518), .A2(n13517), .ZN(n19406) );
  MUX2_X1 U16835 ( .A(n12811), .B(n19406), .S(n19490), .Z(n13519) );
  OAI21_X1 U16836 ( .B1(n13520), .B2(n19481), .A(n13519), .ZN(P2_U2880) );
  NOR2_X1 U16837 ( .A1(n13888), .A2(n13521), .ZN(n13523) );
  INV_X1 U16838 ( .A(n19480), .ZN(n13522) );
  OAI211_X1 U16839 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13523), .A(
        n13522), .B(n19487), .ZN(n13529) );
  OR2_X1 U16840 ( .A1(n13525), .A2(n13524), .ZN(n13527) );
  AND2_X1 U16841 ( .A1(n13527), .A2(n13526), .ZN(n19419) );
  NAND2_X1 U16842 ( .A1(n19490), .A2(n19419), .ZN(n13528) );
  OAI211_X1 U16843 ( .C1(n19490), .C2(n19412), .A(n13529), .B(n13528), .ZN(
        P2_U2881) );
  XNOR2_X1 U16844 ( .A(n13531), .B(n13530), .ZN(n20432) );
  AOI21_X1 U16845 ( .B1(n13533), .B2(n13323), .A(n9800), .ZN(n13537) );
  INV_X1 U16846 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20984) );
  NOR2_X1 U16847 ( .A1(n20347), .A2(n20984), .ZN(n20427) );
  AOI21_X1 U16848 ( .B1(n16351), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20427), .ZN(n13534) );
  OAI21_X1 U16849 ( .B1(n20360), .B2(n16370), .A(n13534), .ZN(n13535) );
  AOI21_X1 U16850 ( .B1(n13537), .B2(n16364), .A(n13535), .ZN(n13536) );
  OAI21_X1 U16851 ( .B1(n16349), .B2(n20432), .A(n13536), .ZN(P1_U2995) );
  INV_X1 U16852 ( .A(n13537), .ZN(n20355) );
  INV_X1 U16853 ( .A(n13544), .ZN(n13538) );
  XNOR2_X1 U16854 ( .A(n13545), .B(n13538), .ZN(n20428) );
  AOI22_X1 U16855 ( .A1(n14784), .A2(n20428), .B1(n14783), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U16856 ( .B1(n20355), .B2(n14769), .A(n13539), .ZN(P1_U2868) );
  INV_X1 U16857 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20400) );
  OAI222_X1 U16858 ( .A1(n20355), .A2(n14869), .B1(n14868), .B2(n14825), .C1(
        n14865), .C2(n20400), .ZN(P1_U2900) );
  AND2_X1 U16859 ( .A1(n13532), .A2(n13541), .ZN(n13542) );
  OR2_X1 U16860 ( .A1(n13540), .A2(n13542), .ZN(n20332) );
  OAI21_X1 U16861 ( .B1(n13545), .B2(n13544), .A(n13543), .ZN(n13546) );
  AND2_X1 U16862 ( .A1(n13546), .A2(n13659), .ZN(n20333) );
  AOI22_X1 U16863 ( .A1(n14784), .A2(n20333), .B1(n14783), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U16864 ( .B1(n20332), .B2(n14769), .A(n13547), .ZN(P1_U2867) );
  OR3_X1 U16865 ( .A1(n20722), .A2(n20862), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20809) );
  INV_X1 U16866 ( .A(n20906), .ZN(n20772) );
  OR2_X1 U16867 ( .A1(n13257), .A2(n9826), .ZN(n20865) );
  NOR2_X1 U16868 ( .A1(n20690), .A2(n20809), .ZN(n13586) );
  INV_X1 U16869 ( .A(n13586), .ZN(n13549) );
  OAI21_X1 U16870 ( .B1(n20865), .B2(n13548), .A(n13549), .ZN(n13555) );
  AOI211_X1 U16871 ( .C1(n20902), .C2(P1_STATEBS16_REG_SCAN_IN), .A(n20901), 
        .B(n13555), .ZN(n13550) );
  AOI211_X2 U16872 ( .C1(n20901), .C2(n20809), .A(n20772), .B(n13550), .ZN(
        n13592) );
  NOR2_X2 U16873 ( .A1(n13554), .A2(n20697), .ZN(n20890) );
  INV_X1 U16874 ( .A(n20853), .ZN(n13588) );
  INV_X1 U16875 ( .A(n20876), .ZN(n20923) );
  INV_X1 U16876 ( .A(n13555), .ZN(n13556) );
  INV_X1 U16877 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20769) );
  OAI22_X1 U16878 ( .A1(n13556), .A2(n20901), .B1(n20809), .B2(n20769), .ZN(
        n13585) );
  AOI22_X1 U16879 ( .A1(n20919), .A2(n13586), .B1(n20918), .B2(n13585), .ZN(
        n13557) );
  OAI21_X1 U16880 ( .B1(n13588), .B2(n20923), .A(n13557), .ZN(n13558) );
  AOI21_X1 U16881 ( .B1(n20890), .B2(n9774), .A(n13558), .ZN(n13559) );
  OAI21_X1 U16882 ( .B1(n13592), .B2(n13560), .A(n13559), .ZN(P1_U3139) );
  INV_X1 U16883 ( .A(n20954), .ZN(n20803) );
  AOI22_X1 U16884 ( .A1(n20953), .A2(n13586), .B1(n20951), .B2(n13585), .ZN(
        n13561) );
  OAI21_X1 U16885 ( .B1(n13588), .B2(n20803), .A(n13561), .ZN(n13562) );
  AOI21_X1 U16886 ( .B1(n20890), .B2(n20852), .A(n13562), .ZN(n13563) );
  OAI21_X1 U16887 ( .B1(n13592), .B2(n13564), .A(n13563), .ZN(P1_U3144) );
  INV_X1 U16888 ( .A(n20926), .ZN(n20788) );
  AOI22_X1 U16889 ( .A1(n20925), .A2(n13586), .B1(n20924), .B2(n13585), .ZN(
        n13565) );
  OAI21_X1 U16890 ( .B1(n13588), .B2(n20788), .A(n13565), .ZN(n13566) );
  AOI21_X1 U16891 ( .B1(n20890), .B2(n20832), .A(n13566), .ZN(n13567) );
  OAI21_X1 U16892 ( .B1(n13592), .B2(n13568), .A(n13567), .ZN(P1_U3140) );
  INV_X1 U16893 ( .A(n20909), .ZN(n20781) );
  AOI22_X1 U16894 ( .A1(n20899), .A2(n13586), .B1(n20898), .B2(n13585), .ZN(
        n13569) );
  OAI21_X1 U16895 ( .B1(n13588), .B2(n20781), .A(n13569), .ZN(n13570) );
  AOI21_X1 U16896 ( .B1(n20890), .B2(n9778), .A(n13570), .ZN(n13571) );
  OAI21_X1 U16897 ( .B1(n13592), .B2(n13572), .A(n13571), .ZN(P1_U3137) );
  INV_X1 U16898 ( .A(n20938), .ZN(n20794) );
  AOI22_X1 U16899 ( .A1(n20937), .A2(n13586), .B1(n20936), .B2(n13585), .ZN(
        n13573) );
  OAI21_X1 U16900 ( .B1(n13588), .B2(n20794), .A(n13573), .ZN(n13574) );
  AOI21_X1 U16901 ( .B1(n20890), .B2(n20840), .A(n13574), .ZN(n13575) );
  OAI21_X1 U16902 ( .B1(n13592), .B2(n13576), .A(n13575), .ZN(P1_U3142) );
  INV_X1 U16903 ( .A(n20885), .ZN(n20949) );
  AOI22_X1 U16904 ( .A1(n20943), .A2(n13586), .B1(n20942), .B2(n13585), .ZN(
        n13577) );
  OAI21_X1 U16905 ( .B1(n13588), .B2(n20949), .A(n13577), .ZN(n13578) );
  AOI21_X1 U16906 ( .B1(n20890), .B2(n9776), .A(n13578), .ZN(n13579) );
  OAI21_X1 U16907 ( .B1(n13592), .B2(n13580), .A(n13579), .ZN(P1_U3143) );
  INV_X1 U16908 ( .A(n20932), .ZN(n20791) );
  AOI22_X1 U16909 ( .A1(n20931), .A2(n13586), .B1(n20930), .B2(n13585), .ZN(
        n13581) );
  OAI21_X1 U16910 ( .B1(n13588), .B2(n20791), .A(n13581), .ZN(n13582) );
  AOI21_X1 U16911 ( .B1(n20890), .B2(n20836), .A(n13582), .ZN(n13583) );
  OAI21_X1 U16912 ( .B1(n13592), .B2(n13584), .A(n13583), .ZN(P1_U3141) );
  INV_X1 U16913 ( .A(n20914), .ZN(n20821) );
  AOI22_X1 U16914 ( .A1(n20913), .A2(n13586), .B1(n20912), .B2(n13585), .ZN(
        n13587) );
  OAI21_X1 U16915 ( .B1(n13588), .B2(n20821), .A(n13587), .ZN(n13589) );
  AOI21_X1 U16916 ( .B1(n20890), .B2(n20823), .A(n13589), .ZN(n13590) );
  OAI21_X1 U16917 ( .B1(n13592), .B2(n13591), .A(n13590), .ZN(P1_U3138) );
  INV_X1 U16918 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13593) );
  OAI222_X1 U16919 ( .A1(n20332), .A2(n14869), .B1(n14868), .B2(n14820), .C1(
        n13593), .C2(n14865), .ZN(P1_U2899) );
  AND2_X1 U16920 ( .A1(n16260), .A2(n20965), .ZN(n13594) );
  OR2_X2 U16921 ( .A1(n13595), .A2(n13594), .ZN(n20412) );
  NAND2_X1 U16922 ( .A1(n13626), .A2(n13635), .ZN(n13627) );
  INV_X1 U16923 ( .A(DATAI_14_), .ZN(n21180) );
  MUX2_X1 U16924 ( .A(n21180), .B(n16841), .S(n13623), .Z(n14857) );
  INV_X1 U16925 ( .A(n14857), .ZN(n13596) );
  NAND2_X1 U16926 ( .A1(n13846), .A2(n13596), .ZN(n20422) );
  NAND2_X1 U16927 ( .A1(n20412), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13597) );
  OAI211_X1 U16928 ( .C1(n13598), .C2(n13820), .A(n20422), .B(n13597), .ZN(
        P1_U2951) );
  INV_X1 U16929 ( .A(DATAI_12_), .ZN(n21203) );
  NAND2_X1 U16930 ( .A1(n13623), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U16931 ( .B1(n13623), .B2(n21203), .A(n13599), .ZN(n14861) );
  NAND2_X1 U16932 ( .A1(n13846), .A2(n14861), .ZN(n20417) );
  NAND2_X1 U16933 ( .A1(n20412), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13600) );
  OAI211_X1 U16934 ( .C1(n13601), .C2(n13820), .A(n20417), .B(n13600), .ZN(
        P1_U2949) );
  INV_X1 U16935 ( .A(DATAI_8_), .ZN(n21198) );
  MUX2_X1 U16936 ( .A(n21198), .B(n16852), .S(n13623), .Z(n14807) );
  INV_X1 U16937 ( .A(n14807), .ZN(n13602) );
  NAND2_X1 U16938 ( .A1(n13846), .A2(n13602), .ZN(n13613) );
  NAND2_X1 U16939 ( .A1(n20412), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13603) );
  OAI211_X1 U16940 ( .C1(n13604), .C2(n13820), .A(n13613), .B(n13603), .ZN(
        P1_U2945) );
  INV_X1 U16941 ( .A(DATAI_13_), .ZN(n21200) );
  MUX2_X1 U16942 ( .A(n21200), .B(n16843), .S(n13623), .Z(n14860) );
  INV_X1 U16943 ( .A(n14860), .ZN(n13605) );
  NAND2_X1 U16944 ( .A1(n13846), .A2(n13605), .ZN(n20419) );
  NAND2_X1 U16945 ( .A1(n20412), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13606) );
  OAI211_X1 U16946 ( .C1(n14786), .C2(n13820), .A(n20419), .B(n13606), .ZN(
        P1_U2950) );
  INV_X1 U16947 ( .A(DATAI_9_), .ZN(n13608) );
  NAND2_X1 U16948 ( .A1(n13623), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13607) );
  OAI21_X1 U16949 ( .B1(n13623), .B2(n13608), .A(n13607), .ZN(n14803) );
  NAND2_X1 U16950 ( .A1(n13846), .A2(n14803), .ZN(n20410) );
  NAND2_X1 U16951 ( .A1(n20412), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13609) );
  OAI211_X1 U16952 ( .C1(n14801), .C2(n13820), .A(n20410), .B(n13609), .ZN(
        P1_U2946) );
  INV_X1 U16953 ( .A(DATAI_11_), .ZN(n21212) );
  MUX2_X1 U16954 ( .A(n21212), .B(n16847), .S(n13623), .Z(n14867) );
  INV_X1 U16955 ( .A(n14867), .ZN(n13610) );
  NAND2_X1 U16956 ( .A1(n13846), .A2(n13610), .ZN(n20415) );
  NAND2_X1 U16957 ( .A1(n20412), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13611) );
  OAI211_X1 U16958 ( .C1(n14793), .C2(n13820), .A(n20415), .B(n13611), .ZN(
        P1_U2948) );
  INV_X1 U16959 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20393) );
  NAND2_X1 U16960 ( .A1(n20412), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13612) );
  OAI211_X1 U16961 ( .C1(n20393), .C2(n13820), .A(n13613), .B(n13612), .ZN(
        P1_U2960) );
  INV_X1 U16962 ( .A(DATAI_10_), .ZN(n13615) );
  NAND2_X1 U16963 ( .A1(n13623), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13614) );
  OAI21_X1 U16964 ( .B1(n13623), .B2(n13615), .A(n13614), .ZN(n14798) );
  NAND2_X1 U16965 ( .A1(n13846), .A2(n14798), .ZN(n20413) );
  NAND2_X1 U16966 ( .A1(n20412), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13616) );
  OAI211_X1 U16967 ( .C1(n13617), .C2(n13820), .A(n20413), .B(n13616), .ZN(
        P1_U2947) );
  OAI211_X1 U16968 ( .C1(n9765), .C2(n10050), .A(n19487), .B(n19471), .ZN(
        n13622) );
  AND2_X1 U16969 ( .A1(n15892), .A2(n13619), .ZN(n13620) );
  OR2_X1 U16970 ( .A1(n13620), .A2(n15604), .ZN(n15627) );
  INV_X1 U16971 ( .A(n15627), .ZN(n19375) );
  NAND2_X1 U16972 ( .A1(n19375), .A2(n19490), .ZN(n13621) );
  OAI211_X1 U16973 ( .C1(n19490), .C2(n12708), .A(n13622), .B(n13621), .ZN(
        P2_U2876) );
  INV_X1 U16974 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14855) );
  INV_X1 U16975 ( .A(DATAI_15_), .ZN(n13625) );
  INV_X1 U16976 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13624) );
  MUX2_X1 U16977 ( .A(n13625), .B(n13624), .S(n13623), .Z(n14856) );
  INV_X1 U16978 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20379) );
  OAI222_X1 U16979 ( .A1(n13820), .A2(n14855), .B1(n13627), .B2(n14856), .C1(
        n13626), .C2(n20379), .ZN(P1_U2967) );
  NAND2_X1 U16980 ( .A1(n21059), .A2(n16253), .ZN(n13633) );
  NAND2_X1 U16981 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21068), .ZN(n16278) );
  NOR2_X1 U16982 ( .A1(n16278), .A2(n10532), .ZN(n13631) );
  NAND2_X1 U16983 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10532), .ZN(n13629) );
  OAI21_X1 U16984 ( .B1(n13629), .B2(n13628), .A(n20347), .ZN(n13630) );
  NOR2_X1 U16985 ( .A1(n13642), .A2(n16490), .ZN(n13632) );
  NAND2_X1 U16986 ( .A1(n13633), .A2(n14732), .ZN(n20372) );
  INV_X1 U16987 ( .A(n20372), .ZN(n20354) );
  NOR2_X1 U16988 ( .A1(n13644), .A2(n13634), .ZN(n13650) );
  NAND2_X1 U16989 ( .A1(n13635), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13639) );
  AND2_X1 U16990 ( .A1(n21064), .A2(n21129), .ZN(n16272) );
  NOR2_X1 U16991 ( .A1(n13639), .A2(n16272), .ZN(n13636) );
  INV_X1 U16992 ( .A(n16272), .ZN(n13637) );
  AOI21_X1 U16993 ( .B1(n13638), .B2(n21061), .A(n13637), .ZN(n13649) );
  INV_X1 U16994 ( .A(n13639), .ZN(n13640) );
  NOR2_X1 U16995 ( .A1(n13649), .A2(n13640), .ZN(n13641) );
  NAND2_X1 U16996 ( .A1(n13650), .A2(n13641), .ZN(n20363) );
  AND2_X1 U16997 ( .A1(n13642), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13643) );
  OAI21_X1 U16998 ( .B1(n20365), .B2(n20319), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13646) );
  NOR2_X1 U16999 ( .A1(n13644), .A2(n16259), .ZN(n20367) );
  NAND2_X1 U17000 ( .A1(n20367), .A2(n14221), .ZN(n13645) );
  OAI211_X1 U17001 ( .C1(n20363), .C2(n13647), .A(n13646), .B(n13645), .ZN(
        n13648) );
  AOI21_X1 U17002 ( .B1(n20345), .B2(n20437), .A(n13648), .ZN(n13653) );
  NAND2_X1 U17003 ( .A1(n20352), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13652) );
  OAI211_X1 U17004 ( .C1(n13654), .C2(n20354), .A(n13653), .B(n13652), .ZN(
        P1_U2840) );
  OAI21_X1 U17005 ( .B1(n13540), .B2(n13656), .A(n13655), .ZN(n13799) );
  INV_X1 U17006 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20397) );
  OAI222_X1 U17007 ( .A1(n13799), .A2(n14869), .B1(n14868), .B2(n13657), .C1(
        n14865), .C2(n20397), .ZN(P1_U2898) );
  AND2_X1 U17008 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  OR2_X1 U17009 ( .A1(n13660), .A2(n13815), .ZN(n13794) );
  INV_X1 U17010 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13661) );
  OAI222_X1 U17011 ( .A1(n13794), .A2(n14765), .B1(n14770), .B2(n13661), .C1(
        n14769), .C2(n13799), .ZN(P1_U2866) );
  XNOR2_X1 U17012 ( .A(n13663), .B(n13662), .ZN(n13806) );
  INV_X1 U17013 ( .A(n15022), .ZN(n13666) );
  NAND2_X1 U17014 ( .A1(n20436), .A2(n10669), .ZN(n16480) );
  OAI22_X1 U17015 ( .A1(n16447), .A2(n20436), .B1(n16446), .B2(n20442), .ZN(
        n13664) );
  NOR2_X1 U17016 ( .A1(n13665), .A2(n13664), .ZN(n16476) );
  OAI21_X1 U17017 ( .B1(n13666), .B2(n16480), .A(n16476), .ZN(n13964) );
  NAND2_X1 U17018 ( .A1(n20334), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17019 ( .B1(n16466), .B2(n13794), .A(n13801), .ZN(n13669) );
  INV_X1 U17020 ( .A(n20424), .ZN(n16481) );
  NOR2_X1 U17021 ( .A1(n16444), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13668) );
  AOI211_X1 U17022 ( .C1(n13964), .C2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13669), .B(n13668), .ZN(n13670) );
  OAI21_X1 U17023 ( .B1(n20431), .B2(n13806), .A(n13670), .ZN(P1_U3025) );
  NAND2_X1 U17024 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13792) );
  AOI21_X1 U17025 ( .B1(n13683), .B2(n13792), .A(n13791), .ZN(n20370) );
  NAND2_X1 U17026 ( .A1(n13671), .A2(n20372), .ZN(n13680) );
  AND2_X1 U17027 ( .A1(n13792), .A2(n13683), .ZN(n13672) );
  AOI22_X1 U17028 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n13672), .ZN(n13673) );
  OAI21_X1 U17029 ( .B1(n20361), .B2(n13674), .A(n13673), .ZN(n13678) );
  INV_X1 U17030 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13675) );
  OAI22_X1 U17031 ( .A1(n20377), .A2(n13676), .B1(n13675), .B2(n20363), .ZN(
        n13677) );
  AOI211_X1 U17032 ( .C1(n20459), .C2(n20367), .A(n13678), .B(n13677), .ZN(
        n13679) );
  OAI211_X1 U17033 ( .C1(n20981), .C2(n20370), .A(n13680), .B(n13679), .ZN(
        P1_U2838) );
  INV_X1 U17034 ( .A(n9669), .ZN(n20866) );
  NAND2_X1 U17035 ( .A1(n20367), .A2(n20866), .ZN(n13682) );
  AOI22_X1 U17036 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13791), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13681) );
  OAI211_X1 U17037 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20361), .A(
        n13682), .B(n13681), .ZN(n13685) );
  OAI22_X1 U17038 ( .A1(n13790), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n9979), .B2(
        n20363), .ZN(n13684) );
  AOI211_X1 U17039 ( .C1(n20345), .C2(n13686), .A(n13685), .B(n13684), .ZN(
        n13687) );
  OAI21_X1 U17040 ( .B1(n13688), .B2(n20354), .A(n13687), .ZN(P1_U2839) );
  NAND2_X1 U17041 ( .A1(n14292), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13698) );
  INV_X1 U17042 ( .A(n13689), .ZN(n13690) );
  NOR2_X1 U17043 ( .A1(n11998), .A2(n13690), .ZN(n13699) );
  INV_X1 U17044 ( .A(n13699), .ZN(n13691) );
  OR2_X1 U17045 ( .A1(n9667), .A2(n13691), .ZN(n13692) );
  NOR2_X1 U17046 ( .A1(n9676), .A2(n13692), .ZN(n14234) );
  AND2_X1 U17047 ( .A1(n13694), .A2(n14053), .ZN(n13701) );
  INV_X1 U17048 ( .A(n13701), .ZN(n13695) );
  OR2_X1 U17049 ( .A1(n9668), .A2(n13695), .ZN(n13696) );
  NOR2_X1 U17050 ( .A1(n13696), .A2(n9676), .ZN(n14235) );
  AOI22_X1 U17051 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14234), .B1(
        n14235), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13697) );
  NAND2_X1 U17052 ( .A1(n13698), .A2(n13697), .ZN(n13708) );
  AND2_X1 U17053 ( .A1(n9676), .A2(n13699), .ZN(n13717) );
  INV_X1 U17054 ( .A(n14296), .ZN(n14241) );
  NAND2_X1 U17055 ( .A1(n13702), .A2(n13699), .ZN(n13700) );
  INV_X1 U17056 ( .A(n14237), .ZN(n13704) );
  NAND2_X1 U17057 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  NOR2_X1 U17058 ( .A1(n9676), .A2(n13703), .ZN(n14236) );
  NAND2_X1 U17059 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  NOR2_X1 U17060 ( .A1(n13708), .A2(n13707), .ZN(n13731) );
  NOR2_X1 U17061 ( .A1(n13746), .A2(n13709), .ZN(n13714) );
  INV_X1 U17062 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13712) );
  NOR2_X1 U17063 ( .A1(n16001), .A2(n14031), .ZN(n13721) );
  NAND2_X1 U17064 ( .A1(n13710), .A2(n13721), .ZN(n19698) );
  AND2_X1 U17065 ( .A1(n16001), .A2(n19612), .ZN(n13722) );
  NAND2_X1 U17066 ( .A1(n13710), .A2(n13722), .ZN(n16049) );
  OAI22_X1 U17067 ( .A1(n13712), .A2(n19698), .B1(n16049), .B2(n13711), .ZN(
        n13713) );
  NOR2_X1 U17068 ( .A1(n13714), .A2(n13713), .ZN(n13730) );
  AOI22_X1 U17069 ( .A1(n19628), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13729) );
  INV_X1 U17070 ( .A(n13719), .ZN(n13727) );
  INV_X1 U17071 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U17072 ( .A1(n13723), .A2(n13721), .ZN(n14283) );
  OAI22_X1 U17073 ( .A1(n13725), .A2(n14283), .B1(n20055), .B2(n13724), .ZN(
        n13726) );
  NOR2_X1 U17074 ( .A1(n13727), .A2(n13726), .ZN(n13728) );
  NAND2_X1 U17075 ( .A1(n13732), .A2(n12298), .ZN(n13940) );
  NAND2_X1 U17076 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13733) );
  INV_X1 U17077 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n19928) );
  INV_X1 U17078 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13735) );
  OAI21_X1 U17079 ( .B1(n14237), .B2(n13735), .A(n16070), .ZN(n13736) );
  INV_X1 U17080 ( .A(n13736), .ZN(n13738) );
  NAND2_X1 U17081 ( .A1(n14236), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13737) );
  OAI211_X1 U17082 ( .C1(n14283), .C2(n19928), .A(n13738), .B(n13737), .ZN(
        n13739) );
  OAI22_X1 U17083 ( .A1(n16049), .A2(n13741), .B1(n14296), .B2(n13740), .ZN(
        n13745) );
  INV_X1 U17084 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13743) );
  OAI22_X1 U17085 ( .A1(n19698), .A2(n13743), .B1(n20055), .B2(n13742), .ZN(
        n13744) );
  NOR2_X1 U17086 ( .A1(n13745), .A2(n13744), .ZN(n13749) );
  AOI22_X1 U17087 ( .A1(n19628), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13748) );
  INV_X1 U17088 ( .A(n13746), .ZN(n14282) );
  AOI22_X1 U17089 ( .A1(n14282), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13747) );
  NAND4_X1 U17090 ( .A1(n13750), .A2(n13749), .A3(n13748), .A4(n13747), .ZN(
        n13754) );
  NAND2_X1 U17091 ( .A1(n13752), .A2(n13751), .ZN(n13753) );
  INV_X1 U17092 ( .A(n13898), .ZN(n13758) );
  NAND2_X1 U17093 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  NAND2_X1 U17094 ( .A1(n13758), .A2(n13757), .ZN(n14043) );
  OAI21_X1 U17095 ( .B1(n13925), .B2(n13760), .A(n13759), .ZN(n13933) );
  XOR2_X1 U17096 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13933), .Z(
        n13761) );
  XNOR2_X1 U17097 ( .A(n13934), .B(n13761), .ZN(n13789) );
  NAND2_X1 U17098 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13762), .ZN(
        n13763) );
  NAND2_X1 U17099 ( .A1(n13764), .A2(n13763), .ZN(n13938) );
  XNOR2_X1 U17100 ( .A(n13938), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13937) );
  OR2_X1 U17101 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  NAND2_X1 U17102 ( .A1(n13767), .A2(n13900), .ZN(n20240) );
  OAI21_X1 U17103 ( .B1(n15782), .B2(n13771), .A(n13770), .ZN(n13772) );
  INV_X1 U17104 ( .A(n13772), .ZN(n13773) );
  INV_X1 U17105 ( .A(n14456), .ZN(n13776) );
  NOR2_X1 U17106 ( .A1(n13782), .A2(n19424), .ZN(n13775) );
  AOI221_X1 U17107 ( .B1(n15941), .B2(n13777), .C1(n13776), .C2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13775), .ZN(n13779) );
  NAND2_X1 U17108 ( .A1(n9675), .A2(n19613), .ZN(n13778) );
  OAI211_X1 U17109 ( .C1(n16677), .C2(n20240), .A(n13779), .B(n13778), .ZN(
        n13780) );
  AOI21_X1 U17110 ( .B1(n13787), .B2(n19611), .A(n13780), .ZN(n13781) );
  OAI21_X1 U17111 ( .B1(n15974), .B2(n13789), .A(n13781), .ZN(P2_U3043) );
  OAI22_X1 U17112 ( .A1(n16670), .A2(n14040), .B1(n13782), .B2(n19424), .ZN(
        n13783) );
  AOI21_X1 U17113 ( .B1(n16661), .B2(n14038), .A(n13783), .ZN(n13784) );
  OAI21_X1 U17114 ( .B1(n13785), .B2(n15640), .A(n13784), .ZN(n13786) );
  AOI21_X1 U17115 ( .B1(n13787), .B2(n19595), .A(n13786), .ZN(n13788) );
  OAI21_X1 U17116 ( .B1(n16665), .B2(n13789), .A(n13788), .ZN(P2_U3011) );
  NAND3_X1 U17117 ( .A1(n20366), .A2(P1_REIP_REG_4__SCAN_IN), .A3(
        P1_REIP_REG_3__SCAN_IN), .ZN(n20344) );
  NOR2_X1 U17118 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20344), .ZN(n13797) );
  INV_X1 U17119 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20989) );
  NAND2_X1 U17120 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13858) );
  OAI21_X1 U17121 ( .B1(n13858), .B2(n20351), .A(n20352), .ZN(n13856) );
  OAI22_X1 U17122 ( .A1(n13802), .A2(n20361), .B1(n20989), .B2(n13856), .ZN(
        n13796) );
  AOI22_X1 U17123 ( .A1(n20346), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20365), .ZN(n13793) );
  OAI211_X1 U17124 ( .C1(n20377), .C2(n13794), .A(n13793), .B(n20347), .ZN(
        n13795) );
  AOI211_X1 U17125 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n13797), .A(n13796), .B(
        n13795), .ZN(n13798) );
  OAI21_X1 U17126 ( .B1(n14732), .B2(n13799), .A(n13798), .ZN(P1_U2834) );
  INV_X1 U17127 ( .A(n13799), .ZN(n13804) );
  NAND2_X1 U17128 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13800) );
  OAI211_X1 U17129 ( .C1(n16370), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n13803) );
  AOI21_X1 U17130 ( .B1(n13804), .B2(n16364), .A(n13803), .ZN(n13805) );
  OAI21_X1 U17131 ( .B1(n13806), .B2(n16349), .A(n13805), .ZN(P1_U2993) );
  NAND2_X1 U17132 ( .A1(n15307), .A2(n13973), .ZN(n13985) );
  OAI211_X1 U17133 ( .C1(n15307), .C2(n13973), .A(n13985), .B(n19487), .ZN(
        n13808) );
  NAND2_X1 U17134 ( .A1(n15841), .A2(n19490), .ZN(n13807) );
  OAI211_X1 U17135 ( .C1(n19490), .C2(n12812), .A(n13808), .B(n13807), .ZN(
        P2_U2874) );
  INV_X1 U17136 ( .A(n13809), .ZN(n13908) );
  NAND2_X1 U17137 ( .A1(n13655), .A2(n13810), .ZN(n13811) );
  AND2_X1 U17138 ( .A1(n13908), .A2(n13811), .ZN(n16363) );
  INV_X1 U17139 ( .A(n16363), .ZN(n13813) );
  OAI222_X1 U17140 ( .A1(n13813), .A2(n14869), .B1(n14868), .B2(n13812), .C1(
        n14865), .C2(n10861), .ZN(P1_U2897) );
  INV_X1 U17141 ( .A(n14769), .ZN(n14774) );
  NOR2_X1 U17142 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  OR2_X1 U17143 ( .A1(n13912), .A2(n13816), .ZN(n13967) );
  OAI22_X1 U17144 ( .A1(n13967), .A2(n14765), .B1(n13817), .B2(n14770), .ZN(
        n13818) );
  AOI21_X1 U17145 ( .B1(n16363), .B2(n14774), .A(n13818), .ZN(n13819) );
  INV_X1 U17146 ( .A(n13819), .ZN(P1_U2865) );
  AOI22_X1 U17147 ( .A1(n20421), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20412), .ZN(n13821) );
  NAND2_X1 U17148 ( .A1(n13846), .A2(n14817), .ZN(n13829) );
  NAND2_X1 U17149 ( .A1(n13821), .A2(n13829), .ZN(P1_U2943) );
  AOI22_X1 U17150 ( .A1(n20421), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20412), .ZN(n13823) );
  INV_X1 U17151 ( .A(n13822), .ZN(n14830) );
  NAND2_X1 U17152 ( .A1(n13846), .A2(n14830), .ZN(n13850) );
  NAND2_X1 U17153 ( .A1(n13823), .A2(n13850), .ZN(P1_U2955) );
  AOI22_X1 U17154 ( .A1(n20421), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20412), .ZN(n13825) );
  INV_X1 U17155 ( .A(n14841), .ZN(n13824) );
  NAND2_X1 U17156 ( .A1(n13846), .A2(n13824), .ZN(n13833) );
  NAND2_X1 U17157 ( .A1(n13825), .A2(n13833), .ZN(P1_U2938) );
  AOI22_X1 U17158 ( .A1(n20421), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20412), .ZN(n13827) );
  INV_X1 U17159 ( .A(n13826), .ZN(n14849) );
  NAND2_X1 U17160 ( .A1(n13846), .A2(n14849), .ZN(n13835) );
  NAND2_X1 U17161 ( .A1(n13827), .A2(n13835), .ZN(P1_U2937) );
  AOI22_X1 U17162 ( .A1(n20421), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20412), .ZN(n13828) );
  NAND2_X1 U17163 ( .A1(n13846), .A2(n14813), .ZN(n13839) );
  NAND2_X1 U17164 ( .A1(n13828), .A2(n13839), .ZN(P1_U2944) );
  AOI22_X1 U17165 ( .A1(n20421), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20412), .ZN(n13830) );
  NAND2_X1 U17166 ( .A1(n13830), .A2(n13829), .ZN(P1_U2958) );
  AOI22_X1 U17167 ( .A1(n20421), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20412), .ZN(n13832) );
  INV_X1 U17168 ( .A(n14825), .ZN(n13831) );
  NAND2_X1 U17169 ( .A1(n13846), .A2(n13831), .ZN(n13843) );
  NAND2_X1 U17170 ( .A1(n13832), .A2(n13843), .ZN(P1_U2941) );
  AOI22_X1 U17171 ( .A1(n20421), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20412), .ZN(n13834) );
  NAND2_X1 U17172 ( .A1(n13834), .A2(n13833), .ZN(P1_U2953) );
  AOI22_X1 U17173 ( .A1(n20421), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20412), .ZN(n13836) );
  NAND2_X1 U17174 ( .A1(n13836), .A2(n13835), .ZN(P1_U2952) );
  AOI22_X1 U17175 ( .A1(n20421), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20412), .ZN(n13838) );
  INV_X1 U17176 ( .A(n14835), .ZN(n13837) );
  NAND2_X1 U17177 ( .A1(n13846), .A2(n13837), .ZN(n13841) );
  NAND2_X1 U17178 ( .A1(n13838), .A2(n13841), .ZN(P1_U2939) );
  AOI22_X1 U17179 ( .A1(n20421), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20412), .ZN(n13840) );
  NAND2_X1 U17180 ( .A1(n13840), .A2(n13839), .ZN(P1_U2959) );
  AOI22_X1 U17181 ( .A1(n20421), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20412), .ZN(n13842) );
  NAND2_X1 U17182 ( .A1(n13842), .A2(n13841), .ZN(P1_U2954) );
  AOI22_X1 U17183 ( .A1(n20421), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20412), .ZN(n13844) );
  NAND2_X1 U17184 ( .A1(n13844), .A2(n13843), .ZN(P1_U2956) );
  AOI22_X1 U17185 ( .A1(n20421), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20412), .ZN(n13847) );
  INV_X1 U17186 ( .A(n14820), .ZN(n13845) );
  NAND2_X1 U17187 ( .A1(n13846), .A2(n13845), .ZN(n13848) );
  NAND2_X1 U17188 ( .A1(n13847), .A2(n13848), .ZN(P1_U2942) );
  AOI22_X1 U17189 ( .A1(n20421), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20412), .ZN(n13849) );
  NAND2_X1 U17190 ( .A1(n13849), .A2(n13848), .ZN(P1_U2957) );
  AOI22_X1 U17191 ( .A1(n20421), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20412), .ZN(n13851) );
  NAND2_X1 U17192 ( .A1(n13851), .A2(n13850), .ZN(P1_U2940) );
  INV_X1 U17193 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20991) );
  AOI21_X1 U17194 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20334), .ZN(n13852) );
  OAI21_X1 U17195 ( .B1(n16360), .B2(n20361), .A(n13852), .ZN(n13854) );
  NOR2_X1 U17196 ( .A1(n20377), .A2(n13967), .ZN(n13853) );
  AOI211_X1 U17197 ( .C1(n20346), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13854), .B(
        n13853), .ZN(n13855) );
  OAI21_X1 U17198 ( .B1(n13856), .B2(n20991), .A(n13855), .ZN(n13857) );
  AOI21_X1 U17199 ( .B1(n16363), .B2(n20327), .A(n13857), .ZN(n13862) );
  INV_X1 U17200 ( .A(n20344), .ZN(n13860) );
  INV_X1 U17201 ( .A(n13858), .ZN(n13859) );
  NAND3_X1 U17202 ( .A1(n13860), .A2(n20991), .A3(n13859), .ZN(n13861) );
  NAND2_X1 U17203 ( .A1(n13862), .A2(n13861), .ZN(P1_U2833) );
  INV_X1 U17204 ( .A(n14320), .ZN(n13863) );
  OAI21_X1 U17205 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n14319) );
  NOR2_X1 U17206 ( .A1(n19416), .A2(n13866), .ZN(n13867) );
  XNOR2_X1 U17207 ( .A(n13867), .B(n16653), .ZN(n13868) );
  INV_X1 U17208 ( .A(n20159), .ZN(n19438) );
  NAND2_X1 U17209 ( .A1(n13868), .A2(n19438), .ZN(n13880) );
  AOI21_X1 U17210 ( .B1(n13869), .B2(n15924), .A(n9745), .ZN(n19524) );
  INV_X1 U17211 ( .A(n19524), .ZN(n16676) );
  OAI22_X1 U17212 ( .A1(n19442), .A2(n16676), .B1(n19425), .B2(n13870), .ZN(
        n13878) );
  OR2_X1 U17213 ( .A1(n13872), .A2(n13871), .ZN(n13875) );
  NAND2_X1 U17214 ( .A1(n13875), .A2(n13874), .ZN(n19486) );
  AOI22_X1 U17215 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19459), .ZN(n13876) );
  OAI211_X1 U17216 ( .C1(n19453), .C2(n19486), .A(n13876), .B(n19424), .ZN(
        n13877) );
  NOR2_X1 U17217 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  OAI211_X1 U17218 ( .C1(n19427), .C2(n14319), .A(n13880), .B(n13879), .ZN(
        P2_U2847) );
  NAND2_X1 U17219 ( .A1(n13881), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13882) );
  AND2_X1 U17220 ( .A1(n13305), .A2(n13882), .ZN(n13886) );
  INV_X1 U17221 ( .A(n13883), .ZN(n13884) );
  NAND3_X1 U17222 ( .A1(n13886), .A2(n13885), .A3(n13884), .ZN(n13887) );
  NAND2_X1 U17223 ( .A1(n13888), .A2(n13887), .ZN(n15398) );
  INV_X1 U17224 ( .A(n19602), .ZN(n13892) );
  NOR2_X1 U17225 ( .A1(n19416), .A2(n13889), .ZN(n13891) );
  AOI21_X1 U17226 ( .B1(n13892), .B2(n13891), .A(n20159), .ZN(n13890) );
  OAI21_X1 U17227 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(n13905) );
  OR2_X1 U17228 ( .A1(n13894), .A2(n13893), .ZN(n13896) );
  AND2_X1 U17229 ( .A1(n13896), .A2(n13895), .ZN(n19596) );
  OAI21_X1 U17230 ( .B1(n13898), .B2(n13897), .A(n14268), .ZN(n14272) );
  AOI22_X1 U17231 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19459), .ZN(n13899) );
  OAI211_X1 U17232 ( .C1(n19427), .C2(n14272), .A(n13899), .B(n19424), .ZN(
        n13903) );
  XNOR2_X1 U17233 ( .A(n13901), .B(n13900), .ZN(n15399) );
  OAI22_X1 U17234 ( .A1(n19442), .A2(n15399), .B1(n19425), .B2(n12535), .ZN(
        n13902) );
  AOI211_X1 U17235 ( .C1(n19596), .C2(n19437), .A(n13903), .B(n13902), .ZN(
        n13904) );
  OAI211_X1 U17236 ( .C1(n19277), .C2(n15398), .A(n13905), .B(n13904), .ZN(
        P2_U2851) );
  INV_X1 U17237 ( .A(n13906), .ZN(n13907) );
  AOI21_X1 U17238 ( .B1(n13909), .B2(n13908), .A(n13907), .ZN(n13961) );
  NAND3_X1 U17239 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13910) );
  NOR3_X1 U17240 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20344), .A3(n13910), .ZN(
        n13916) );
  OR2_X1 U17241 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  NAND2_X1 U17242 ( .A1(n13995), .A2(n13913), .ZN(n16465) );
  AOI22_X1 U17243 ( .A1(n20346), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20365), .ZN(n13914) );
  OAI211_X1 U17244 ( .C1(n20377), .C2(n16465), .A(n13914), .B(n20347), .ZN(
        n13915) );
  NOR2_X1 U17245 ( .A1(n13916), .A2(n13915), .ZN(n13918) );
  INV_X1 U17246 ( .A(n20352), .ZN(n14717) );
  NAND4_X1 U17247 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14077)
         );
  NOR2_X1 U17248 ( .A1(n14077), .A2(n20351), .ZN(n14079) );
  NOR2_X1 U17249 ( .A1(n14717), .A2(n14079), .ZN(n20318) );
  NAND2_X1 U17250 ( .A1(n20318), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U17251 ( .C1(n20361), .C2(n13959), .A(n13918), .B(n13917), .ZN(
        n13919) );
  AOI21_X1 U17252 ( .B1(n13961), .B2(n20327), .A(n13919), .ZN(n13920) );
  INV_X1 U17253 ( .A(n13920), .ZN(P1_U2832) );
  NOR2_X1 U17254 ( .A1(n19416), .A2(n14026), .ZN(n13922) );
  XNOR2_X1 U17255 ( .A(n13922), .B(n13921), .ZN(n13923) );
  NAND2_X1 U17256 ( .A1(n13923), .A2(n19420), .ZN(n13932) );
  INV_X1 U17257 ( .A(n19442), .ZN(n19450) );
  OAI22_X1 U17258 ( .A1(n19429), .A2(n13924), .B1(n20187), .B2(n19425), .ZN(
        n13927) );
  NOR2_X1 U17259 ( .A1(n19427), .A2(n13925), .ZN(n13926) );
  AOI211_X1 U17260 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19459), .A(
        n13927), .B(n13926), .ZN(n13928) );
  OAI21_X1 U17261 ( .B1(n13929), .B2(n19453), .A(n13928), .ZN(n13930) );
  AOI21_X1 U17262 ( .B1(n20256), .B2(n19450), .A(n13930), .ZN(n13931) );
  OAI211_X1 U17263 ( .C1(n16002), .C2(n19277), .A(n13932), .B(n13931), .ZN(
        P2_U2853) );
  INV_X1 U17264 ( .A(n13961), .ZN(n13998) );
  OAI222_X1 U17265 ( .A1(n13998), .A2(n14869), .B1(n14868), .B2(n14807), .C1(
        n20393), .C2(n14865), .ZN(P1_U2896) );
  XNOR2_X1 U17266 ( .A(n14272), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14274) );
  NAND2_X1 U17267 ( .A1(n13936), .A2(n13935), .ZN(n14275) );
  XOR2_X1 U17268 ( .A(n14274), .B(n14275), .Z(n19599) );
  INV_X1 U17269 ( .A(n19599), .ZN(n13954) );
  NAND2_X1 U17270 ( .A1(n13938), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13939) );
  INV_X1 U17271 ( .A(n13946), .ZN(n13944) );
  XNOR2_X1 U17272 ( .A(n13942), .B(n14278), .ZN(n13945) );
  INV_X1 U17273 ( .A(n13945), .ZN(n13943) );
  NAND2_X1 U17274 ( .A1(n13944), .A2(n13943), .ZN(n14420) );
  NAND2_X1 U17275 ( .A1(n13946), .A2(n13945), .ZN(n14419) );
  NAND2_X1 U17276 ( .A1(n14420), .A2(n14419), .ZN(n13947) );
  XNOR2_X1 U17277 ( .A(n13947), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19594) );
  NAND2_X1 U17278 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15941), .ZN(
        n15962) );
  OAI21_X1 U17279 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15786), .A(
        n14456), .ZN(n15968) );
  NOR2_X1 U17280 ( .A1(n12535), .A2(n19424), .ZN(n13948) );
  AOI21_X1 U17281 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15968), .A(
        n13948), .ZN(n13949) );
  OAI21_X1 U17282 ( .B1(n16677), .B2(n15399), .A(n13949), .ZN(n13950) );
  AOI21_X1 U17283 ( .B1(n19596), .B2(n19613), .A(n13950), .ZN(n13951) );
  OAI21_X1 U17284 ( .B1(n15962), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13951), .ZN(n13952) );
  AOI21_X1 U17285 ( .B1(n19594), .B2(n19611), .A(n13952), .ZN(n13953) );
  OAI21_X1 U17286 ( .B1(n13954), .B2(n15974), .A(n13953), .ZN(P2_U3042) );
  XNOR2_X1 U17287 ( .A(n13956), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13957) );
  XNOR2_X1 U17288 ( .A(n13955), .B(n13957), .ZN(n16468) );
  INV_X1 U17289 ( .A(n16468), .ZN(n13963) );
  AOI22_X1 U17290 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13958) );
  OAI21_X1 U17291 ( .B1(n13959), .B2(n16370), .A(n13958), .ZN(n13960) );
  AOI21_X1 U17292 ( .B1(n13961), .B2(n16364), .A(n13960), .ZN(n13962) );
  OAI21_X1 U17293 ( .B1(n13963), .B2(n16349), .A(n13962), .ZN(P1_U2991) );
  AOI21_X1 U17294 ( .B1(n12904), .B2(n16416), .A(n13964), .ZN(n16473) );
  XOR2_X1 U17295 ( .A(n13966), .B(n13965), .Z(n16365) );
  NAND2_X1 U17296 ( .A1(n16365), .A2(n20439), .ZN(n13971) );
  NOR2_X1 U17297 ( .A1(n12904), .A2(n16444), .ZN(n16469) );
  NAND2_X1 U17298 ( .A1(n20334), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n16366) );
  INV_X1 U17299 ( .A(n16366), .ZN(n13969) );
  NOR2_X1 U17300 ( .A1(n16466), .A2(n13967), .ZN(n13968) );
  AOI211_X1 U17301 ( .C1(n10717), .C2(n16469), .A(n13969), .B(n13968), .ZN(
        n13970) );
  OAI211_X1 U17302 ( .C1(n10717), .C2(n16473), .A(n13971), .B(n13970), .ZN(
        P1_U3024) );
  NOR2_X1 U17303 ( .A1(n14021), .A2(n13972), .ZN(n19465) );
  AND2_X1 U17304 ( .A1(n15307), .A2(n13973), .ZN(n13975) );
  NAND2_X1 U17305 ( .A1(n13975), .A2(n13974), .ZN(n16599) );
  OAI21_X1 U17306 ( .B1(n19465), .B2(n13976), .A(n16599), .ZN(n15321) );
  OR2_X1 U17307 ( .A1(n15236), .A2(n13977), .ZN(n13978) );
  NAND2_X1 U17308 ( .A1(n15222), .A2(n13978), .ZN(n19346) );
  AOI22_X1 U17309 ( .A1(n19496), .A2(BUF1_REG_17__SCAN_IN), .B1(n19497), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U17310 ( .A1(n19495), .A2(n13979), .B1(n19546), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13980) );
  OAI211_X1 U17311 ( .C1(n19538), .C2(n19346), .A(n13981), .B(n13980), .ZN(
        n13982) );
  INV_X1 U17312 ( .A(n13982), .ZN(n13983) );
  OAI21_X1 U17313 ( .B1(n15321), .B2(n19551), .A(n13983), .ZN(P2_U2902) );
  XNOR2_X1 U17314 ( .A(n13985), .B(n13984), .ZN(n13990) );
  AND2_X1 U17315 ( .A1(n13987), .A2(n13986), .ZN(n13988) );
  OR2_X1 U17316 ( .A1(n13988), .A2(n9750), .ZN(n15832) );
  MUX2_X1 U17317 ( .A(n15832), .B(n14002), .S(n19484), .Z(n13989) );
  OAI21_X1 U17318 ( .B1(n13990), .B2(n19481), .A(n13989), .ZN(P2_U2873) );
  AND2_X1 U17319 ( .A1(n13906), .A2(n13991), .ZN(n13993) );
  OR2_X1 U17320 ( .A1(n13993), .A2(n13992), .ZN(n14062) );
  AOI21_X1 U17321 ( .B1(n13995), .B2(n13994), .A(n10093), .ZN(n20325) );
  AOI22_X1 U17322 ( .A1(n20325), .A2(n14784), .B1(n14783), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13996) );
  OAI21_X1 U17323 ( .B1(n14062), .B2(n14769), .A(n13996), .ZN(P1_U2863) );
  INV_X1 U17324 ( .A(n14868), .ZN(n14068) );
  AOI22_X1 U17325 ( .A1(n14068), .A2(n14803), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14847), .ZN(n13997) );
  OAI21_X1 U17326 ( .B1(n14062), .B2(n14869), .A(n13997), .ZN(P1_U2895) );
  INV_X1 U17327 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13999) );
  OAI222_X1 U17328 ( .A1(n16465), .A2(n14765), .B1(n14770), .B2(n13999), .C1(
        n14769), .C2(n13998), .ZN(P1_U2864) );
  NAND2_X1 U17329 ( .A1(n14328), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14001) );
  MUX2_X1 U17330 ( .A(n14001), .B(n14328), .S(n9713), .Z(n14003) );
  NAND2_X1 U17331 ( .A1(n9713), .A2(n14002), .ZN(n14361) );
  NAND2_X1 U17332 ( .A1(n14003), .A2(n14361), .ZN(n14380) );
  NOR2_X1 U17333 ( .A1(n19416), .A2(n15175), .ZN(n14007) );
  AND2_X1 U17334 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  OR2_X1 U17335 ( .A1(n14006), .A2(n15173), .ZN(n15578) );
  XNOR2_X1 U17336 ( .A(n14007), .B(n15578), .ZN(n14008) );
  NAND2_X1 U17337 ( .A1(n14008), .A2(n19420), .ZN(n14016) );
  INV_X1 U17338 ( .A(n15832), .ZN(n15580) );
  NOR2_X1 U17339 ( .A1(n19425), .A2(n15576), .ZN(n14014) );
  NOR2_X1 U17340 ( .A1(n12822), .A2(n14009), .ZN(n14010) );
  NOR2_X1 U17341 ( .A1(n15812), .A2(n14010), .ZN(n19508) );
  INV_X1 U17342 ( .A(n19508), .ZN(n14012) );
  AOI22_X1 U17343 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19459), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19443), .ZN(n14011) );
  OAI211_X1 U17344 ( .C1(n14012), .C2(n19442), .A(n14011), .B(n19424), .ZN(
        n14013) );
  AOI211_X1 U17345 ( .C1(n15580), .C2(n19437), .A(n14014), .B(n14013), .ZN(
        n14015) );
  OAI211_X1 U17346 ( .C1(n19427), .C2(n14380), .A(n14016), .B(n14015), .ZN(
        P2_U2841) );
  NOR2_X1 U17347 ( .A1(n9750), .A2(n14018), .ZN(n14019) );
  OR2_X1 U17348 ( .A1(n14017), .A2(n14019), .ZN(n15809) );
  INV_X1 U17349 ( .A(n14021), .ZN(n14023) );
  INV_X1 U17350 ( .A(n14020), .ZN(n14022) );
  OR2_X1 U17351 ( .A1(n14021), .A2(n14020), .ZN(n19464) );
  OAI211_X1 U17352 ( .C1(n14023), .C2(n14022), .A(n19487), .B(n19464), .ZN(
        n14025) );
  NAND2_X1 U17353 ( .A1(n19484), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14024) );
  OAI211_X1 U17354 ( .C1(n15809), .C2(n19484), .A(n14025), .B(n14024), .ZN(
        P2_U2872) );
  AOI211_X1 U17355 ( .C1(n14049), .C2(n14027), .A(n19416), .B(n14026), .ZN(
        n15975) );
  AOI22_X1 U17356 ( .A1(n15975), .A2(n19420), .B1(n19458), .B2(n13109), .ZN(
        n14035) );
  AOI22_X1 U17357 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19459), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19443), .ZN(n14029) );
  NAND2_X1 U17358 ( .A1(n19444), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14028) );
  OAI211_X1 U17359 ( .C1(n19427), .C2(n14030), .A(n14029), .B(n14028), .ZN(
        n14033) );
  NOR2_X1 U17360 ( .A1(n14031), .A2(n19453), .ZN(n14032) );
  AOI211_X1 U17361 ( .C1(n20270), .C2(n19450), .A(n14033), .B(n14032), .ZN(
        n14034) );
  OAI211_X1 U17362 ( .C1(n20265), .C2(n19277), .A(n14035), .B(n14034), .ZN(
        P2_U2854) );
  NAND2_X1 U17363 ( .A1(n9647), .A2(n14036), .ZN(n14037) );
  XNOR2_X1 U17364 ( .A(n14038), .B(n14037), .ZN(n14039) );
  NAND2_X1 U17365 ( .A1(n14039), .A2(n19420), .ZN(n14048) );
  OAI22_X1 U17366 ( .A1(n14040), .A2(n19390), .B1(n19442), .B2(n20240), .ZN(
        n14041) );
  INV_X1 U17367 ( .A(n14041), .ZN(n14042) );
  OAI21_X1 U17368 ( .B1(n19427), .B2(n14043), .A(n14042), .ZN(n14046) );
  OAI22_X1 U17369 ( .A1(n19429), .A2(n14044), .B1(n13782), .B2(n19425), .ZN(
        n14045) );
  AOI211_X1 U17370 ( .C1(n9676), .C2(n19437), .A(n14046), .B(n14045), .ZN(
        n14047) );
  OAI211_X1 U17371 ( .C1(n20248), .C2(n19277), .A(n14048), .B(n14047), .ZN(
        P2_U2852) );
  NAND2_X1 U17372 ( .A1(n9647), .A2(n14049), .ZN(n19462) );
  OAI21_X1 U17373 ( .B1(n9647), .B2(n13085), .A(n19462), .ZN(n15976) );
  INV_X1 U17374 ( .A(n15976), .ZN(n14056) );
  AND2_X1 U17375 ( .A1(n14051), .A2(n14050), .ZN(n15979) );
  NOR2_X1 U17376 ( .A1(n15979), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14052) );
  AOI21_X1 U17377 ( .B1(n14053), .B2(n16006), .A(n14052), .ZN(n16708) );
  INV_X1 U17378 ( .A(n16732), .ZN(n16021) );
  OAI22_X1 U17379 ( .A1(n19283), .A2(n16708), .B1(n16021), .B2(n14054), .ZN(
        n14055) );
  AOI21_X1 U17380 ( .B1(n14056), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n14055), 
        .ZN(n14058) );
  AOI21_X1 U17381 ( .B1(n15993), .B2(n20246), .A(n15986), .ZN(n14057) );
  OAI22_X1 U17382 ( .A1(n14058), .A2(n15986), .B1(n14057), .B2(n16709), .ZN(
        P2_U3601) );
  XNOR2_X1 U17383 ( .A(n10723), .B(n14059), .ZN(n14060) );
  XNOR2_X1 U17384 ( .A(n14061), .B(n14060), .ZN(n16460) );
  INV_X1 U17385 ( .A(n14062), .ZN(n20328) );
  AOI22_X1 U17386 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14063) );
  OAI21_X1 U17387 ( .B1(n14064), .B2(n16370), .A(n14063), .ZN(n14065) );
  AOI21_X1 U17388 ( .B1(n20328), .B2(n16364), .A(n14065), .ZN(n14066) );
  OAI21_X1 U17389 ( .B1(n16460), .B2(n16349), .A(n14066), .ZN(P1_U2990) );
  XOR2_X1 U17390 ( .A(n14067), .B(n13992), .Z(n15015) );
  INV_X1 U17391 ( .A(n15015), .ZN(n14070) );
  AOI22_X1 U17392 ( .A1(n14068), .A2(n14798), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14847), .ZN(n14069) );
  OAI21_X1 U17393 ( .B1(n14070), .B2(n14869), .A(n14069), .ZN(P1_U2894) );
  NAND2_X1 U17394 ( .A1(n14072), .A2(n14071), .ZN(n14073) );
  NAND2_X1 U17395 ( .A1(n14781), .A2(n14073), .ZN(n16455) );
  INV_X1 U17396 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14074) );
  OAI22_X1 U17397 ( .A1(n16455), .A2(n14765), .B1(n14074), .B2(n14770), .ZN(
        n14075) );
  AOI21_X1 U17398 ( .B1(n15015), .B2(n14774), .A(n14075), .ZN(n14076) );
  INV_X1 U17399 ( .A(n14076), .ZN(P1_U2862) );
  NOR2_X2 U17400 ( .A1(n20344), .A2(n14077), .ZN(n20326) );
  INV_X1 U17401 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20996) );
  NAND3_X1 U17402 ( .A1(n20326), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n20996), 
        .ZN(n14083) );
  AOI22_X1 U17403 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20365), .B1(
        n20346), .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n14078) );
  OAI211_X1 U17404 ( .C1(n20377), .C2(n16455), .A(n14078), .B(n20347), .ZN(
        n14081) );
  NAND3_X1 U17405 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n14079), .ZN(n14169) );
  NAND2_X1 U17406 ( .A1(n20352), .A2(n14169), .ZN(n16326) );
  NOR2_X1 U17407 ( .A1(n20996), .A2(n16326), .ZN(n14080) );
  NOR2_X1 U17408 ( .A1(n14081), .A2(n14080), .ZN(n14082) );
  OAI211_X1 U17409 ( .C1(n20361), .C2(n15013), .A(n14083), .B(n14082), .ZN(
        n14084) );
  AOI21_X1 U17410 ( .B1(n15015), .B2(n20327), .A(n14084), .ZN(n14085) );
  INV_X1 U17411 ( .A(n14085), .ZN(P1_U2830) );
  INV_X1 U17412 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17351) );
  NAND2_X1 U17413 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .ZN(n14092) );
  INV_X1 U17414 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17424) );
  NOR3_X1 U17415 ( .A1(n14086), .A2(n18623), .A3(n17729), .ZN(n14088) );
  INV_X1 U17416 ( .A(n19036), .ZN(n16744) );
  NOR4_X2 U17417 ( .A1(n19256), .A2(n16946), .A3(n16299), .A4(n19100), .ZN(
        n17621) );
  INV_X1 U17418 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17479) );
  NAND2_X1 U17419 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .ZN(n16204) );
  NAND4_X1 U17420 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n14090) );
  INV_X1 U17421 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17601) );
  INV_X1 U17422 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17281) );
  NAND3_X1 U17423 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17600) );
  NOR3_X1 U17424 ( .A1(n17601), .A2(n17281), .A3(n17600), .ZN(n17585) );
  INV_X1 U17425 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17216) );
  INV_X1 U17426 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17587) );
  INV_X1 U17427 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17252) );
  NOR3_X1 U17428 ( .A1(n17216), .A2(n17587), .A3(n17252), .ZN(n16203) );
  NAND4_X1 U17429 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17585), .A4(n16203), .ZN(n14089) );
  NOR4_X1 U17430 ( .A1(n17479), .A2(n16204), .A3(n14090), .A4(n14089), .ZN(
        n17463) );
  NAND2_X1 U17431 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17463), .ZN(n17462) );
  NOR2_X1 U17432 ( .A1(n17586), .A2(n17462), .ZN(n17449) );
  NAND2_X1 U17433 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17449), .ZN(n17448) );
  NAND2_X1 U17434 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17437), .ZN(n17407) );
  INV_X1 U17435 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17366) );
  INV_X1 U17436 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17362) );
  NOR2_X1 U17437 ( .A1(n17366), .A2(n17362), .ZN(n16114) );
  AND2_X1 U17438 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17352) );
  NAND4_X1 U17439 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16114), .A4(n17352), .ZN(n14091) );
  NOR4_X1 U17440 ( .A1(n17351), .A2(n14092), .A3(n17407), .A4(n14091), .ZN(
        n17344) );
  NAND2_X1 U17441 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17344), .ZN(n14093) );
  NOR2_X1 U17442 ( .A1(n17729), .A2(n14093), .ZN(n14095) );
  NAND2_X1 U17443 ( .A1(n17596), .A2(n14093), .ZN(n17345) );
  INV_X1 U17444 ( .A(n17345), .ZN(n14094) );
  MUX2_X1 U17445 ( .A(n14095), .B(n14094), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NOR2_X1 U17446 ( .A1(n9868), .A2(n19229), .ZN(n19056) );
  AOI21_X1 U17447 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19056), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14107) );
  OR2_X1 U17448 ( .A1(n14097), .A2(n14107), .ZN(n19043) );
  NOR2_X1 U17449 ( .A1(n19212), .A2(n19043), .ZN(n14106) );
  AOI21_X1 U17450 ( .B1(n16745), .B2(n17838), .A(n19062), .ZN(n14098) );
  INV_X1 U17451 ( .A(n14098), .ZN(n16300) );
  NAND2_X1 U17452 ( .A1(n19256), .A2(n17838), .ZN(n19094) );
  INV_X1 U17453 ( .A(n19094), .ZN(n14099) );
  NOR2_X1 U17454 ( .A1(n16945), .A2(n14099), .ZN(n14100) );
  INV_X1 U17455 ( .A(n19257), .ZN(n19122) );
  NOR2_X1 U17456 ( .A1(n19122), .A2(n16915), .ZN(n16301) );
  OAI21_X1 U17457 ( .B1(n16300), .B2(n17776), .A(n16301), .ZN(n14104) );
  NOR2_X1 U17458 ( .A1(n14102), .A2(n14101), .ZN(n14103) );
  NAND2_X1 U17459 ( .A1(n14104), .A2(n14103), .ZN(n19069) );
  NOR2_X1 U17460 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19206), .ZN(n18609) );
  INV_X1 U17461 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18598) );
  NAND3_X1 U17462 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19204)
         );
  NOR2_X1 U17463 ( .A1(n18598), .A2(n19204), .ZN(n14105) );
  MUX2_X1 U17464 ( .A(n14106), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19236), .Z(P3_U3284) );
  NAND2_X1 U17465 ( .A1(n14107), .A2(n10220), .ZN(n18597) );
  NOR2_X1 U17466 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18597), .ZN(n14108) );
  INV_X1 U17467 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19102) );
  NOR2_X1 U17468 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19260) );
  AOI21_X1 U17469 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19260), .ZN(n19110) );
  OAI21_X1 U17470 ( .B1(n14108), .B2(n19204), .A(n18947), .ZN(n18603) );
  INV_X1 U17471 ( .A(n18603), .ZN(n14109) );
  NAND2_X1 U17472 ( .A1(n19268), .A2(n19206), .ZN(n16911) );
  AND2_X1 U17473 ( .A1(n19212), .A2(n16911), .ZN(n19250) );
  INV_X1 U17474 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19255) );
  NOR2_X1 U17475 ( .A1(n19216), .A2(n19255), .ZN(n18156) );
  NOR2_X1 U17476 ( .A1(n19250), .A2(n18156), .ZN(n16208) );
  AOI21_X1 U17477 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n16208), .ZN(n16209) );
  NOR2_X1 U17478 ( .A1(n14109), .A2(n16209), .ZN(n14111) );
  NAND3_X1 U17479 ( .A1(n19268), .A2(n19206), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18847) );
  INV_X1 U17480 ( .A(n18847), .ZN(n18897) );
  NOR2_X1 U17481 ( .A1(n19206), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18646) );
  OR2_X1 U17482 ( .A1(n18646), .A2(n14109), .ZN(n16207) );
  OR2_X1 U17483 ( .A1(n18897), .A2(n16207), .ZN(n14110) );
  MUX2_X1 U17484 ( .A(n14111), .B(n14110), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17485 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14112) );
  AOI21_X1 U17486 ( .B1(n14165), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14112), .ZN(
        n14205) );
  INV_X1 U17487 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U17488 ( .A1(n14113), .A2(n14114), .ZN(n14117) );
  INV_X1 U17489 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15021) );
  OAI211_X1 U17490 ( .C1(n14164), .C2(n15021), .A(n14115), .B(n14150), .ZN(
        n14116) );
  NAND2_X1 U17491 ( .A1(n14117), .A2(n14116), .ZN(n14711) );
  OR2_X1 U17492 ( .A1(n14163), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U17493 ( .A1(n14150), .A2(n16417), .ZN(n14118) );
  OAI211_X1 U17494 ( .C1(n14158), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14118), .B(
        n14204), .ZN(n14119) );
  MUX2_X1 U17495 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14123) );
  NAND2_X1 U17496 ( .A1(n10739), .A2(n14121), .ZN(n14122) );
  OR2_X1 U17497 ( .A1(n14163), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14126) );
  INV_X1 U17498 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16424) );
  NAND2_X1 U17499 ( .A1(n14150), .A2(n16424), .ZN(n14124) );
  OAI211_X1 U17500 ( .C1(n14158), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14124), .B(
        n14204), .ZN(n14125) );
  NAND2_X1 U17501 ( .A1(n14126), .A2(n14125), .ZN(n14753) );
  MUX2_X1 U17502 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14128) );
  OR2_X1 U17503 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14127) );
  NAND2_X1 U17504 ( .A1(n14128), .A2(n14127), .ZN(n14683) );
  OR2_X1 U17505 ( .A1(n14163), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17506 ( .A1(n14150), .A2(n16398), .ZN(n14129) );
  OAI211_X1 U17507 ( .C1(n14158), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14129), .B(
        n14204), .ZN(n14130) );
  MUX2_X1 U17508 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14133) );
  OR2_X1 U17509 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14132) );
  AND2_X1 U17510 ( .A1(n14133), .A2(n14132), .ZN(n14662) );
  INV_X1 U17511 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15137) );
  OAI21_X1 U17512 ( .B1(n14164), .B2(n15137), .A(n14150), .ZN(n14134) );
  OAI21_X1 U17513 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n14158), .A(n14134), .ZN(
        n14136) );
  OR2_X1 U17514 ( .A1(n14163), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n14135) );
  NAND2_X1 U17515 ( .A1(n14136), .A2(n14135), .ZN(n14650) );
  OR2_X1 U17516 ( .A1(n14154), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14139) );
  OR2_X1 U17517 ( .A1(n14158), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14137) );
  OAI211_X1 U17518 ( .C1(n14164), .C2(n15133), .A(n14137), .B(n14150), .ZN(
        n14138) );
  NAND2_X1 U17519 ( .A1(n14139), .A2(n14138), .ZN(n14638) );
  OR2_X1 U17520 ( .A1(n14163), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14142) );
  INV_X1 U17521 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U17522 ( .A1(n14150), .A2(n14937), .ZN(n14140) );
  OAI211_X1 U17523 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n14158), .A(n14140), .B(
        n14204), .ZN(n14141) );
  AND2_X1 U17524 ( .A1(n14142), .A2(n14141), .ZN(n14626) );
  MUX2_X1 U17525 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14144) );
  OR2_X1 U17526 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14143) );
  NAND2_X1 U17527 ( .A1(n14144), .A2(n14143), .ZN(n14615) );
  OAI21_X1 U17528 ( .B1(n14164), .B2(n15106), .A(n14150), .ZN(n14145) );
  OAI21_X1 U17529 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n14158), .A(n14145), .ZN(
        n14147) );
  OR2_X1 U17530 ( .A1(n14163), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U17531 ( .A1(n14147), .A2(n14146), .ZN(n14604) );
  MUX2_X1 U17532 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14149) );
  OR2_X1 U17533 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14148) );
  NAND2_X1 U17534 ( .A1(n14149), .A2(n14148), .ZN(n14593) );
  OR2_X1 U17535 ( .A1(n14163), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U17536 ( .A1(n14150), .A2(n15091), .ZN(n14151) );
  OAI211_X1 U17537 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n14158), .A(n14151), .B(
        n14204), .ZN(n14152) );
  AND2_X1 U17538 ( .A1(n14153), .A2(n14152), .ZN(n14579) );
  MUX2_X1 U17539 ( .A(n14154), .B(n14204), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14156) );
  OR2_X1 U17540 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14155) );
  AND2_X1 U17541 ( .A1(n14156), .A2(n14155), .ZN(n14564) );
  OR2_X1 U17542 ( .A1(n14163), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U17543 ( .A1(n14150), .A2(n14887), .ZN(n14157) );
  OAI211_X1 U17544 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n14158), .A(n14157), .B(
        n14204), .ZN(n14159) );
  NAND2_X1 U17545 ( .A1(n14160), .A2(n14159), .ZN(n14548) );
  OR2_X1 U17546 ( .A1(n14165), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14162) );
  OR2_X1 U17547 ( .A1(n14158), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U17548 ( .A1(n14162), .A2(n14161), .ZN(n14202) );
  OAI22_X1 U17549 ( .A1(n14202), .A2(n14164), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14163), .ZN(n14535) );
  MUX2_X1 U17550 ( .A(n14204), .B(n14205), .S(n14537), .Z(n14167) );
  AOI22_X1 U17551 ( .A1(n14165), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14158), .ZN(n14166) );
  NAND2_X1 U17552 ( .A1(n14168), .A2(n20327), .ZN(n14188) );
  INV_X1 U17553 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21182) );
  INV_X1 U17554 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21201) );
  NOR2_X1 U17555 ( .A1(n21182), .A2(n21201), .ZN(n14178) );
  NAND2_X1 U17556 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14180) );
  NOR2_X1 U17557 ( .A1(n14180), .A2(n14169), .ZN(n14716) );
  NAND3_X1 U17558 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14716), .ZN(n14702) );
  NAND3_X1 U17559 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14170) );
  OAI21_X1 U17560 ( .B1(n14702), .B2(n14170), .A(n20352), .ZN(n14687) );
  AND3_X1 U17561 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14181) );
  INV_X1 U17562 ( .A(n14181), .ZN(n14171) );
  NAND2_X1 U17563 ( .A1(n20352), .A2(n14171), .ZN(n14172) );
  NAND2_X1 U17564 ( .A1(n14687), .A2(n14172), .ZN(n14656) );
  AND3_X1 U17565 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_23__SCAN_IN), .ZN(n14182) );
  INV_X1 U17566 ( .A(n14182), .ZN(n14173) );
  AND2_X1 U17567 ( .A1(n20352), .A2(n14173), .ZN(n14174) );
  NAND2_X1 U17568 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14585) );
  INV_X1 U17569 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21173) );
  NOR2_X1 U17570 ( .A1(n14585), .A2(n21173), .ZN(n14183) );
  INV_X1 U17571 ( .A(n14183), .ZN(n14175) );
  AND2_X1 U17572 ( .A1(n20352), .A2(n14175), .ZN(n14176) );
  NAND2_X1 U17573 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14184) );
  AND2_X1 U17574 ( .A1(n20352), .A2(n14184), .ZN(n14177) );
  NOR2_X1 U17575 ( .A1(n14588), .A2(n14177), .ZN(n14554) );
  OAI21_X1 U17576 ( .B1(n14178), .B2(n14717), .A(n14554), .ZN(n14213) );
  INV_X1 U17577 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14733) );
  OAI22_X1 U17578 ( .A1(n20363), .A2(n14733), .B1(n14179), .B2(n20321), .ZN(
        n14186) );
  INV_X1 U17579 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21004) );
  NAND3_X1 U17580 ( .A1(n20326), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16329) );
  NAND2_X1 U17581 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14715), .ZN(n14703) );
  NOR2_X2 U17582 ( .A1(n21004), .A2(n14703), .ZN(n16317) );
  NAND3_X1 U17583 ( .A1(n16317), .A2(P1_REIP_REG_16__SCAN_IN), .A3(
        P1_REIP_REG_15__SCAN_IN), .ZN(n14688) );
  INV_X1 U17584 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21010) );
  NAND2_X1 U17585 ( .A1(n14584), .A2(n14183), .ZN(n14572) );
  AOI211_X1 U17586 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14213), .A(n14186), 
        .B(n14185), .ZN(n14187) );
  OAI211_X1 U17587 ( .C1(n15017), .C2(n20377), .A(n14188), .B(n14187), .ZN(
        P1_U2809) );
  NOR2_X1 U17588 ( .A1(n20347), .A2(n21201), .ZN(n15047) );
  NOR2_X1 U17589 ( .A1(n16370), .A2(n14209), .ZN(n14191) );
  AOI211_X1 U17590 ( .C1(n16351), .C2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15047), .B(n14191), .ZN(n14197) );
  NAND2_X1 U17591 ( .A1(n15045), .A2(n20302), .ZN(n14196) );
  OAI211_X1 U17592 ( .C1(n14217), .C2(n16371), .A(n14197), .B(n14196), .ZN(
        P1_U2969) );
  NOR2_X1 U17593 ( .A1(n14824), .A2(n16810), .ZN(n14200) );
  NAND3_X1 U17595 ( .A1(n14865), .A2(n10295), .A3(n14198), .ZN(n14840) );
  OAI22_X1 U17596 ( .A1(n21270), .A2(n21115), .B1(n14857), .B2(n14840), .ZN(
        n14199) );
  AOI211_X1 U17597 ( .C1(n14847), .C2(P1_EAX_REG_30__SCAN_IN), .A(n14200), .B(
        n14199), .ZN(n14201) );
  OAI21_X1 U17598 ( .B1(n14217), .B2(n14869), .A(n14201), .ZN(P1_U2874) );
  INV_X1 U17599 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14208) );
  INV_X1 U17600 ( .A(n14550), .ZN(n14203) );
  OAI22_X1 U17601 ( .A1(n14537), .A2(n14204), .B1(n14203), .B2(n14202), .ZN(
        n14207) );
  INV_X1 U17602 ( .A(n14205), .ZN(n14206) );
  INV_X1 U17603 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14210) );
  OAI22_X1 U17604 ( .A1(n14210), .A2(n20321), .B1(n20361), .B2(n14209), .ZN(
        n14212) );
  NOR2_X1 U17605 ( .A1(n14543), .A2(n21182), .ZN(n14214) );
  OAI21_X1 U17606 ( .B1(n14214), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14213), 
        .ZN(n14215) );
  OAI211_X1 U17607 ( .C1(n14217), .C2(n14732), .A(n14216), .B(n14215), .ZN(
        P1_U2810) );
  NOR2_X1 U17608 ( .A1(n14218), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14219) );
  AOI21_X1 U17609 ( .B1(n14221), .B2(n14220), .A(n14219), .ZN(n16234) );
  OAI21_X1 U17610 ( .B1(n16234), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16490), 
        .ZN(n14223) );
  AOI22_X1 U17611 ( .A1(n14223), .A2(n14222), .B1(n14224), .B2(n21038), .ZN(
        n14226) );
  AOI21_X1 U17612 ( .B1(n16232), .B2(n21040), .A(n21043), .ZN(n14225) );
  OAI22_X1 U17613 ( .A1(n14226), .A2(n21043), .B1(n14225), .B2(n14224), .ZN(
        P1_U3474) );
  OAI21_X1 U17614 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n14328), .ZN(n14227) );
  INV_X1 U17615 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19467) );
  NOR2_X1 U17616 ( .A1(n19650), .A2(n14228), .ZN(n14354) );
  OR2_X2 U17617 ( .A1(n14355), .A2(n14354), .ZN(n14357) );
  NOR2_X1 U17618 ( .A1(n19650), .A2(n14229), .ZN(n14349) );
  OR2_X2 U17619 ( .A1(n14357), .A2(n14349), .ZN(n14351) );
  NOR2_X1 U17620 ( .A1(n19650), .A2(n14230), .ZN(n14347) );
  INV_X1 U17621 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U17623 ( .A1(n14328), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14388) );
  NAND2_X2 U17624 ( .A1(n14371), .A2(n14388), .ZN(n14393) );
  INV_X1 U17625 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16574) );
  NOR2_X1 U17626 ( .A1(n19650), .A2(n16574), .ZN(n14392) );
  NAND2_X1 U17627 ( .A1(n14328), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14231) );
  NAND2_X1 U17628 ( .A1(n10184), .A2(n9710), .ZN(n14232) );
  NAND2_X1 U17629 ( .A1(n14414), .A2(n14232), .ZN(n16526) );
  NAND2_X1 U17630 ( .A1(n14281), .A2(n14278), .ZN(n14266) );
  AOI22_X1 U17631 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14234), .B1(
        n14235), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14240) );
  NAND3_X1 U17632 ( .A1(n14240), .A2(n14239), .A3(n14238), .ZN(n14245) );
  AOI22_X1 U17633 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n14295), .B1(
        n14241), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U17634 ( .A1(n14292), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14242) );
  NOR2_X1 U17635 ( .A1(n14245), .A2(n14244), .ZN(n14261) );
  INV_X1 U17636 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14246) );
  NOR2_X1 U17637 ( .A1(n13746), .A2(n14246), .ZN(n14249) );
  OAI22_X1 U17638 ( .A1(n12178), .A2(n19698), .B1(n16049), .B2(n14247), .ZN(
        n14248) );
  AOI22_X1 U17639 ( .A1(n19628), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14259) );
  INV_X1 U17640 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14251) );
  OAI22_X1 U17641 ( .A1(n14251), .A2(n14283), .B1(n20055), .B2(n14250), .ZN(
        n14257) );
  INV_X1 U17642 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14255) );
  INV_X1 U17643 ( .A(n19953), .ZN(n14254) );
  INV_X1 U17644 ( .A(n16083), .ZN(n14253) );
  OAI22_X1 U17645 ( .A1(n14255), .A2(n14254), .B1(n14253), .B2(n14252), .ZN(
        n14256) );
  NOR2_X1 U17646 ( .A1(n14257), .A2(n14256), .ZN(n14258) );
  NAND4_X1 U17647 ( .A1(n14261), .A2(n14260), .A3(n14259), .A4(n14258), .ZN(
        n14264) );
  NAND2_X1 U17648 ( .A1(n14262), .A2(n12298), .ZN(n14263) );
  NAND2_X1 U17649 ( .A1(n14264), .A2(n14263), .ZN(n14279) );
  NAND2_X1 U17650 ( .A1(n14418), .A2(n14233), .ZN(n14271) );
  INV_X1 U17651 ( .A(n14310), .ZN(n14270) );
  NAND2_X1 U17652 ( .A1(n14268), .A2(n14267), .ZN(n14269) );
  NAND2_X1 U17653 ( .A1(n14270), .A2(n14269), .ZN(n19426) );
  NAND2_X1 U17654 ( .A1(n14271), .A2(n19426), .ZN(n14276) );
  XNOR2_X1 U17655 ( .A(n14276), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15952) );
  NOR2_X1 U17656 ( .A1(n14272), .A2(n15965), .ZN(n14273) );
  AOI21_X1 U17657 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n15951) );
  NAND2_X1 U17658 ( .A1(n14276), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14277) );
  NOR2_X1 U17659 ( .A1(n14279), .A2(n12536), .ZN(n14280) );
  INV_X1 U17660 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14285) );
  INV_X1 U17661 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14284) );
  OAI22_X1 U17662 ( .A1(n19698), .A2(n14285), .B1(n14283), .B2(n14284), .ZN(
        n14286) );
  AOI21_X1 U17663 ( .B1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n14282), .A(
        n14286), .ZN(n14303) );
  AOI22_X1 U17664 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19953), .B1(
        n16083), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U17665 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n14290) );
  AOI22_X1 U17666 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13704), .B1(
        n14235), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U17667 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14234), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17668 ( .A1(n19628), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14292), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14301) );
  OAI22_X1 U17669 ( .A1(n16049), .A2(n14294), .B1(n20055), .B2(n14293), .ZN(
        n14299) );
  INV_X1 U17670 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14297) );
  OAI22_X1 U17671 ( .A1(n20096), .A2(n14297), .B1(n14296), .B2(n16113), .ZN(
        n14298) );
  NOR2_X1 U17672 ( .A1(n14299), .A2(n14298), .ZN(n14300) );
  NAND4_X1 U17673 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14300), .ZN(
        n14306) );
  NAND2_X1 U17674 ( .A1(n14304), .A2(n12298), .ZN(n14305) );
  NOR2_X1 U17675 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  OR2_X1 U17676 ( .A1(n14315), .A2(n14311), .ZN(n19411) );
  INV_X1 U17677 ( .A(n14313), .ZN(n14314) );
  XNOR2_X1 U17678 ( .A(n14315), .B(n14314), .ZN(n19404) );
  AND2_X1 U17679 ( .A1(n19404), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15636) );
  INV_X1 U17680 ( .A(n15636), .ZN(n14317) );
  NAND2_X1 U17681 ( .A1(n14316), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15634) );
  OR2_X1 U17682 ( .A1(n14319), .A2(n14233), .ZN(n14324) );
  NOR2_X1 U17683 ( .A1(n14324), .A2(n16689), .ZN(n16645) );
  INV_X1 U17684 ( .A(n14326), .ZN(n14323) );
  NAND2_X1 U17685 ( .A1(n14328), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14321) );
  MUX2_X1 U17686 ( .A(n14321), .B(n14328), .S(n14320), .Z(n14322) );
  AND2_X1 U17687 ( .A1(n14323), .A2(n14322), .ZN(n19388) );
  NAND2_X1 U17688 ( .A1(n19388), .A2(n14497), .ZN(n14337) );
  INV_X1 U17689 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15921) );
  NAND2_X1 U17690 ( .A1(n14337), .A2(n15921), .ZN(n15616) );
  NAND2_X1 U17691 ( .A1(n14324), .A2(n16689), .ZN(n16643) );
  INV_X1 U17692 ( .A(n19404), .ZN(n14325) );
  NAND2_X1 U17693 ( .A1(n14325), .A2(n16675), .ZN(n16641) );
  AND2_X1 U17694 ( .A1(n16643), .A2(n16641), .ZN(n15613) );
  NOR2_X1 U17695 ( .A1(n14326), .A2(n12704), .ZN(n14327) );
  NAND2_X1 U17696 ( .A1(n14328), .A2(n14327), .ZN(n14329) );
  AND2_X1 U17697 ( .A1(n14406), .A2(n14329), .ZN(n14330) );
  NAND2_X1 U17698 ( .A1(n14332), .A2(n14330), .ZN(n14340) );
  OR2_X1 U17699 ( .A1(n14340), .A2(n14233), .ZN(n14331) );
  INV_X1 U17700 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15885) );
  NAND2_X1 U17701 ( .A1(n14331), .A2(n15885), .ZN(n15882) );
  NAND2_X1 U17702 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n14332), .ZN(n14333) );
  NOR2_X1 U17703 ( .A1(n19650), .A2(n14333), .ZN(n14334) );
  OR2_X1 U17704 ( .A1(n14335), .A2(n14334), .ZN(n19370) );
  INV_X1 U17705 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15875) );
  OAI21_X1 U17706 ( .B1(n19370), .B2(n14233), .A(n15875), .ZN(n15618) );
  NAND4_X1 U17707 ( .A1(n15616), .A2(n15613), .A3(n15882), .A4(n15618), .ZN(
        n14336) );
  INV_X1 U17708 ( .A(n14337), .ZN(n14338) );
  NAND2_X1 U17709 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14339) );
  NOR2_X1 U17710 ( .A1(n19370), .A2(n14339), .ZN(n15617) );
  INV_X1 U17711 ( .A(n14340), .ZN(n19382) );
  AND2_X1 U17712 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14341) );
  NAND2_X1 U17713 ( .A1(n10182), .A2(n9633), .ZN(n14343) );
  NAND2_X1 U17714 ( .A1(n14344), .A2(n14343), .ZN(n19362) );
  INV_X1 U17715 ( .A(n15597), .ZN(n14345) );
  OAI21_X1 U17716 ( .B1(n19362), .B2(n14233), .A(n15858), .ZN(n15598) );
  AND2_X1 U17717 ( .A1(n14346), .A2(n14497), .ZN(n14381) );
  NOR2_X1 U17718 ( .A1(n14381), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15586) );
  AND2_X1 U17719 ( .A1(n14351), .A2(n14347), .ZN(n14348) );
  NOR2_X1 U17720 ( .A1(n14373), .A2(n14348), .ZN(n19321) );
  AOI21_X1 U17721 ( .B1(n19321), .B2(n14497), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U17722 ( .A1(n14357), .A2(n14349), .ZN(n14350) );
  AND2_X1 U17723 ( .A1(n14351), .A2(n14350), .ZN(n15218) );
  NAND2_X1 U17724 ( .A1(n15218), .A2(n14497), .ZN(n14378) );
  INV_X1 U17725 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15534) );
  AND2_X1 U17726 ( .A1(n14378), .A2(n15534), .ZN(n15530) );
  NAND3_X1 U17727 ( .A1(n14362), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n14328), 
        .ZN(n14352) );
  OAI211_X1 U17728 ( .C1(n14362), .C2(P2_EBX_REG_16__SCAN_IN), .A(n14352), .B(
        n14406), .ZN(n15245) );
  OAI21_X1 U17729 ( .B1(n15245), .B2(n14233), .A(n15800), .ZN(n14353) );
  NAND2_X1 U17730 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  NAND2_X1 U17731 ( .A1(n14357), .A2(n14356), .ZN(n19336) );
  OR2_X1 U17732 ( .A1(n19336), .A2(n14233), .ZN(n14358) );
  INV_X1 U17733 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15790) );
  NAND2_X1 U17734 ( .A1(n14358), .A2(n15790), .ZN(n15492) );
  INV_X1 U17735 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14359) );
  NOR2_X1 U17736 ( .A1(n19650), .A2(n14359), .ZN(n14360) );
  NAND2_X1 U17737 ( .A1(n14361), .A2(n14360), .ZN(n14363) );
  NAND2_X1 U17738 ( .A1(n14363), .A2(n14362), .ZN(n19352) );
  OR2_X1 U17739 ( .A1(n19352), .A2(n14233), .ZN(n14364) );
  NAND2_X1 U17740 ( .A1(n14364), .A2(n15784), .ZN(n15562) );
  OR2_X1 U17741 ( .A1(n14380), .A2(n14233), .ZN(n14365) );
  INV_X1 U17742 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15827) );
  NAND2_X1 U17743 ( .A1(n14365), .A2(n15827), .ZN(n15572) );
  NAND4_X1 U17744 ( .A1(n15550), .A2(n15492), .A3(n15562), .A4(n15572), .ZN(
        n14366) );
  NOR3_X1 U17745 ( .A1(n15494), .A2(n15530), .A3(n14366), .ZN(n14374) );
  NOR2_X1 U17746 ( .A1(n19650), .A2(n14367), .ZN(n14368) );
  AND2_X1 U17747 ( .A1(n14369), .A2(n14368), .ZN(n14370) );
  NOR2_X1 U17748 ( .A1(n14371), .A2(n14370), .ZN(n19311) );
  NAND2_X1 U17749 ( .A1(n19311), .A2(n14497), .ZN(n14375) );
  NAND2_X1 U17750 ( .A1(n14375), .A2(n15740), .ZN(n15497) );
  NOR2_X1 U17751 ( .A1(n19650), .A2(n15208), .ZN(n14372) );
  XNOR2_X1 U17752 ( .A(n14373), .B(n14372), .ZN(n15202) );
  NAND2_X1 U17753 ( .A1(n15202), .A2(n14497), .ZN(n14376) );
  NAND2_X1 U17754 ( .A1(n14376), .A2(n15748), .ZN(n15506) );
  NAND4_X1 U17755 ( .A1(n15560), .A2(n14374), .A3(n15497), .A4(n15506), .ZN(
        n14387) );
  OR2_X1 U17756 ( .A1(n14375), .A2(n15740), .ZN(n15498) );
  AND2_X1 U17757 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14377) );
  NAND2_X1 U17758 ( .A1(n19321), .A2(n14377), .ZN(n15518) );
  INV_X1 U17759 ( .A(n14378), .ZN(n14379) );
  NAND2_X1 U17760 ( .A1(n14379), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15516) );
  NAND2_X1 U17761 ( .A1(n15518), .A2(n15516), .ZN(n15495) );
  OR3_X1 U17762 ( .A1(n14380), .A2(n14233), .A3(n15827), .ZN(n15571) );
  OR3_X1 U17763 ( .A1(n19352), .A2(n14233), .A3(n15784), .ZN(n15561) );
  INV_X1 U17764 ( .A(n14381), .ZN(n14383) );
  INV_X1 U17765 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14382) );
  AND3_X1 U17766 ( .A1(n15571), .A2(n15561), .A3(n15584), .ZN(n15488) );
  NAND2_X1 U17767 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14384) );
  NAND3_X1 U17768 ( .A1(n15488), .A2(n15490), .A3(n15493), .ZN(n14385) );
  NOR2_X1 U17769 ( .A1(n15495), .A2(n14385), .ZN(n14386) );
  INV_X1 U17770 ( .A(n14388), .ZN(n14389) );
  NAND2_X1 U17771 ( .A1(n14390), .A2(n14389), .ZN(n14391) );
  NAND2_X1 U17772 ( .A1(n14393), .A2(n14391), .ZN(n16220) );
  INV_X1 U17773 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15729) );
  OAI21_X1 U17774 ( .B1(n16220), .B2(n14233), .A(n15729), .ZN(n15476) );
  AND2_X1 U17775 ( .A1(n14393), .A2(n14392), .ZN(n14394) );
  OR2_X1 U17776 ( .A1(n14394), .A2(n14397), .ZN(n16578) );
  NOR2_X1 U17777 ( .A1(n16578), .A2(n14233), .ZN(n14395) );
  XNOR2_X1 U17778 ( .A(n14395), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15464) );
  INV_X1 U17779 ( .A(n16578), .ZN(n14396) );
  INV_X1 U17780 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15698) );
  NAND2_X1 U17781 ( .A1(n14328), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14398) );
  MUX2_X1 U17782 ( .A(n14398), .B(P2_EBX_REG_24__SCAN_IN), .S(n14397), .Z(
        n14399) );
  NAND2_X1 U17783 ( .A1(n14399), .A2(n14406), .ZN(n16561) );
  NOR2_X1 U17784 ( .A1(n16561), .A2(n14233), .ZN(n15457) );
  NAND2_X1 U17785 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n9724), .ZN(n14400) );
  NOR2_X1 U17786 ( .A1(n19650), .A2(n14400), .ZN(n14401) );
  OAI21_X1 U17787 ( .B1(n16537), .B2(n14233), .A(n15677), .ZN(n14403) );
  NAND2_X1 U17788 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14402) );
  NOR2_X1 U17789 ( .A1(n14408), .A2(n15278), .ZN(n14404) );
  NAND2_X1 U17790 ( .A1(n14328), .A2(n14404), .ZN(n14405) );
  NAND2_X1 U17791 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  AOI21_X1 U17792 ( .B1(n14408), .B2(n15278), .A(n14407), .ZN(n16549) );
  AND2_X1 U17793 ( .A1(n16549), .A2(n14497), .ZN(n14409) );
  NAND3_X1 U17794 ( .A1(n15450), .A2(n15440), .A3(n15446), .ZN(n14484) );
  INV_X1 U17795 ( .A(n14409), .ZN(n14410) );
  INV_X1 U17796 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15690) );
  INV_X1 U17797 ( .A(n14411), .ZN(n14412) );
  NOR2_X1 U17798 ( .A1(n15447), .A2(n14412), .ZN(n14489) );
  NOR2_X1 U17799 ( .A1(n19650), .A2(n14413), .ZN(n14415) );
  AOI21_X1 U17800 ( .B1(n14415), .B2(n14414), .A(n14490), .ZN(n15199) );
  NAND2_X1 U17801 ( .A1(n15199), .A2(n14497), .ZN(n14487) );
  XNOR2_X1 U17802 ( .A(n14487), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14416) );
  INV_X1 U17803 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U17804 ( .A1(n14419), .A2(n15965), .ZN(n14421) );
  AND2_X2 U17805 ( .A1(n14421), .A2(n14420), .ZN(n15956) );
  INV_X1 U17806 ( .A(n14418), .ZN(n14422) );
  INV_X1 U17807 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15964) );
  NAND2_X1 U17808 ( .A1(n14422), .A2(n15964), .ZN(n15953) );
  NAND2_X1 U17809 ( .A1(n15956), .A2(n15953), .ZN(n15958) );
  NAND2_X1 U17810 ( .A1(n15958), .A2(n15954), .ZN(n14425) );
  NAND2_X1 U17811 ( .A1(n14425), .A2(n14417), .ZN(n14426) );
  NAND2_X1 U17812 ( .A1(n15632), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14430) );
  NAND2_X1 U17813 ( .A1(n14427), .A2(n14233), .ZN(n14429) );
  NAND2_X1 U17814 ( .A1(n14434), .A2(n14429), .ZN(n15630) );
  INV_X1 U17815 ( .A(n15632), .ZN(n14431) );
  XNOR2_X1 U17816 ( .A(n14434), .B(n16689), .ZN(n16637) );
  INV_X1 U17817 ( .A(n14434), .ZN(n14435) );
  NAND2_X1 U17818 ( .A1(n14435), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14436) );
  AND2_X1 U17819 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15872) );
  AND2_X1 U17820 ( .A1(n15872), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15825) );
  NAND2_X1 U17821 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15826) );
  NOR2_X1 U17822 ( .A1(n15826), .A2(n15827), .ZN(n14437) );
  NAND2_X1 U17823 ( .A1(n15825), .A2(n14437), .ZN(n15461) );
  AND2_X1 U17824 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15791) );
  NAND2_X1 U17825 ( .A1(n15791), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14438) );
  NOR2_X1 U17826 ( .A1(n15461), .A2(n14438), .ZN(n15770) );
  NAND2_X1 U17827 ( .A1(n15770), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15710) );
  NAND2_X1 U17828 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15712) );
  AND2_X1 U17829 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15699) );
  AND2_X1 U17830 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14439) );
  NAND2_X1 U17831 ( .A1(n15699), .A2(n14439), .ZN(n14451) );
  OR3_X1 U17832 ( .A1(n15710), .A2(n15712), .A3(n14451), .ZN(n14457) );
  INV_X1 U17833 ( .A(n14457), .ZN(n14440) );
  NAND2_X1 U17834 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14458) );
  AOI21_X1 U17835 ( .B1(n15662), .B2(n14471), .A(n15419), .ZN(n14468) );
  NAND2_X1 U17836 ( .A1(n14441), .A2(n14442), .ZN(n14443) );
  NAND2_X1 U17837 ( .A1(n9706), .A2(n14443), .ZN(n15256) );
  NOR2_X1 U17838 ( .A1(n19424), .A2(n14444), .ZN(n14463) );
  NOR2_X1 U17839 ( .A1(n15190), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14446) );
  OR2_X1 U17840 ( .A1(n14445), .A2(n14446), .ZN(n15192) );
  NOR2_X1 U17841 ( .A1(n19603), .A2(n15192), .ZN(n14447) );
  AOI211_X1 U17842 ( .C1(n19593), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14463), .B(n14447), .ZN(n14448) );
  OAI21_X1 U17843 ( .B1(n15256), .B2(n15640), .A(n14448), .ZN(n14449) );
  AOI21_X1 U17844 ( .B1(n14468), .B2(n19595), .A(n14449), .ZN(n14450) );
  OAI21_X1 U17845 ( .B1(n14470), .B2(n16665), .A(n14450), .ZN(P2_U2986) );
  NOR2_X1 U17846 ( .A1(n15965), .A2(n15964), .ZN(n15963) );
  AND3_X1 U17847 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n15963), .ZN(n14452) );
  NAND2_X1 U17848 ( .A1(n14452), .A2(n15941), .ZN(n16673) );
  NAND2_X1 U17849 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16672) );
  INV_X1 U17850 ( .A(n15710), .ZN(n15749) );
  NAND2_X1 U17851 ( .A1(n15922), .A2(n15749), .ZN(n15747) );
  NOR2_X1 U17852 ( .A1(n15741), .A2(n14451), .ZN(n15691) );
  NAND2_X1 U17853 ( .A1(n15691), .A2(n9895), .ZN(n15660) );
  NOR2_X1 U17854 ( .A1(n15660), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14480) );
  INV_X1 U17855 ( .A(n14452), .ZN(n14453) );
  NAND2_X1 U17856 ( .A1(n19617), .A2(n14453), .ZN(n14454) );
  NAND2_X1 U17857 ( .A1(n14456), .A2(n14454), .ZN(n16671) );
  AND2_X1 U17858 ( .A1(n19617), .A2(n16672), .ZN(n14455) );
  OR2_X1 U17859 ( .A1(n16671), .A2(n14455), .ZN(n15780) );
  NAND2_X1 U17860 ( .A1(n14456), .A2(n15786), .ZN(n15893) );
  OAI21_X1 U17861 ( .B1(n15780), .B2(n14457), .A(n15893), .ZN(n15697) );
  NAND2_X1 U17862 ( .A1(n15893), .A2(n14458), .ZN(n14459) );
  AND2_X1 U17863 ( .A1(n15697), .A2(n14459), .ZN(n14521) );
  INV_X1 U17864 ( .A(n14521), .ZN(n14478) );
  NOR2_X1 U17865 ( .A1(n14480), .A2(n14478), .ZN(n15659) );
  INV_X1 U17866 ( .A(n15256), .ZN(n14464) );
  OR2_X1 U17867 ( .A1(n14476), .A2(n14460), .ZN(n14461) );
  NAND2_X1 U17868 ( .A1(n15323), .A2(n14461), .ZN(n15334) );
  NOR2_X1 U17869 ( .A1(n15334), .A2(n16677), .ZN(n14462) );
  AOI211_X1 U17870 ( .C1(n14464), .C2(n19613), .A(n14463), .B(n14462), .ZN(
        n14466) );
  NOR2_X1 U17871 ( .A1(n15660), .A2(n14486), .ZN(n14525) );
  NAND2_X1 U17872 ( .A1(n14525), .A2(n15662), .ZN(n14465) );
  OAI211_X1 U17873 ( .C1(n15659), .C2(n15662), .A(n14466), .B(n14465), .ZN(
        n14467) );
  AOI21_X1 U17874 ( .B1(n14468), .B2(n19611), .A(n14467), .ZN(n14469) );
  OAI21_X1 U17875 ( .B1(n9717), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14471), .ZN(n15438) );
  XNOR2_X1 U17876 ( .A(n14472), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15429) );
  INV_X1 U17877 ( .A(n15974), .ZN(n19606) );
  NAND2_X1 U17878 ( .A1(n15429), .A2(n19606), .ZN(n14483) );
  OR2_X1 U17879 ( .A1(n15269), .A2(n14473), .ZN(n14474) );
  NAND2_X1 U17880 ( .A1(n14441), .A2(n14474), .ZN(n15432) );
  INV_X1 U17881 ( .A(n15432), .ZN(n16530) );
  AND2_X1 U17882 ( .A1(n9707), .A2(n14475), .ZN(n14477) );
  OR2_X1 U17883 ( .A1(n14477), .A2(n14476), .ZN(n16536) );
  NAND2_X1 U17884 ( .A1(n14478), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14479) );
  NAND2_X1 U17885 ( .A1(n19592), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15430) );
  OAI211_X1 U17886 ( .C1(n16536), .C2(n16677), .A(n14479), .B(n15430), .ZN(
        n14481) );
  AOI211_X1 U17887 ( .C1(n19613), .C2(n16530), .A(n14481), .B(n14480), .ZN(
        n14482) );
  OAI211_X1 U17888 ( .C1(n15438), .C2(n16684), .A(n14483), .B(n14482), .ZN(
        P2_U3019) );
  AOI21_X1 U17889 ( .B1(n15662), .B2(n14486), .A(n14487), .ZN(n14488) );
  NAND2_X1 U17890 ( .A1(n14328), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14491) );
  XNOR2_X1 U17891 ( .A(n14490), .B(n14491), .ZN(n14496) );
  INV_X1 U17892 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U17893 ( .B1(n14496), .B2(n14233), .A(n15663), .ZN(n15416) );
  INV_X1 U17894 ( .A(n14491), .ZN(n14492) );
  NAND2_X1 U17895 ( .A1(n14328), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14494) );
  XNOR2_X1 U17896 ( .A(n14498), .B(n14494), .ZN(n16505) );
  AOI21_X1 U17897 ( .B1(n16505), .B2(n14497), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15408) );
  AND2_X1 U17898 ( .A1(n14497), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14495) );
  NAND2_X1 U17899 ( .A1(n16505), .A2(n14495), .ZN(n15406) );
  INV_X1 U17900 ( .A(n14496), .ZN(n16515) );
  NAND3_X1 U17901 ( .A1(n16515), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14497), .ZN(n15415) );
  OAI211_X1 U17902 ( .C1(n15405), .C2(n15408), .A(n15406), .B(n15415), .ZN(
        n14505) );
  INV_X1 U17903 ( .A(n14498), .ZN(n14500) );
  INV_X1 U17904 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U17905 ( .A1(n14500), .A2(n14499), .ZN(n14501) );
  MUX2_X1 U17906 ( .A(n14502), .B(n14501), .S(n14328), .Z(n16498) );
  NOR2_X1 U17907 ( .A1(n16498), .A2(n14233), .ZN(n14503) );
  XNOR2_X1 U17908 ( .A(n14505), .B(n14504), .ZN(n14530) );
  NAND2_X1 U17909 ( .A1(n15419), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15420) );
  AOI22_X1 U17910 ( .A1(n9648), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14508) );
  NAND2_X1 U17911 ( .A1(n14506), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14507) );
  OAI211_X1 U17912 ( .C1(n14510), .C2(n14509), .A(n14508), .B(n14507), .ZN(
        n14512) );
  NAND2_X1 U17913 ( .A1(n19592), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U17914 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14513) );
  OAI211_X1 U17915 ( .C1(n19603), .C2(n14514), .A(n14524), .B(n14513), .ZN(
        n14515) );
  INV_X1 U17916 ( .A(n16587), .ZN(n16501) );
  AOI222_X1 U17917 ( .A1(n14516), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12595), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12649), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n14517) );
  NAND3_X1 U17918 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U17919 ( .A1(n19617), .A2(n14519), .ZN(n14520) );
  AND2_X1 U17920 ( .A1(n14521), .A2(n14520), .ZN(n15648) );
  OAI21_X1 U17921 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15786), .A(
        n15648), .ZN(n14522) );
  NAND2_X1 U17922 ( .A1(n14522), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14523) );
  NAND3_X1 U17923 ( .A1(n14525), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15649) );
  NOR3_X1 U17924 ( .A1(n15649), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15647), .ZN(n14526) );
  NAND2_X1 U17925 ( .A1(n14527), .A2(n19611), .ZN(n14528) );
  OAI211_X1 U17926 ( .C1(n14530), .C2(n15974), .A(n14529), .B(n14528), .ZN(
        P2_U3015) );
  INV_X1 U17927 ( .A(n14531), .ZN(n14534) );
  NOR2_X1 U17928 ( .A1(n14550), .A2(n14535), .ZN(n14536) );
  INV_X1 U17929 ( .A(n15059), .ZN(n14540) );
  INV_X1 U17930 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U17931 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14875), .ZN(n14538) );
  OAI21_X1 U17932 ( .B1(n20363), .B2(n14734), .A(n14538), .ZN(n14539) );
  AOI21_X1 U17933 ( .B1(n14540), .B2(n20345), .A(n14539), .ZN(n14542) );
  OR2_X1 U17934 ( .A1(n14554), .A2(n21182), .ZN(n14541) );
  OAI211_X1 U17935 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14543), .A(n14542), 
        .B(n14541), .ZN(n14544) );
  AOI21_X1 U17936 ( .B1(n14879), .B2(n20327), .A(n14544), .ZN(n14545) );
  INV_X1 U17937 ( .A(n14545), .ZN(P1_U2811) );
  INV_X1 U17938 ( .A(n14572), .ZN(n14559) );
  INV_X1 U17939 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21185) );
  NOR2_X1 U17940 ( .A1(n21185), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14558) );
  NOR2_X1 U17941 ( .A1(n14566), .A2(n14548), .ZN(n14549) );
  INV_X1 U17942 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14735) );
  INV_X1 U17943 ( .A(n14881), .ZN(n14551) );
  AOI22_X1 U17944 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14551), .ZN(n14552) );
  OAI21_X1 U17945 ( .B1(n20363), .B2(n14735), .A(n14552), .ZN(n14553) );
  INV_X1 U17946 ( .A(n14553), .ZN(n14556) );
  INV_X1 U17947 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21138) );
  OR2_X1 U17948 ( .A1(n14554), .A2(n21138), .ZN(n14555) );
  OAI211_X1 U17949 ( .C1(n15070), .C2(n20377), .A(n14556), .B(n14555), .ZN(
        n14557) );
  AOI21_X1 U17950 ( .B1(n14559), .B2(n14558), .A(n14557), .ZN(n14560) );
  OAI21_X1 U17951 ( .B1(n14891), .B2(n14732), .A(n14560), .ZN(P1_U2812) );
  NOR2_X1 U17952 ( .A1(n14578), .A2(n14564), .ZN(n14565) );
  OR2_X1 U17953 ( .A1(n14566), .A2(n14565), .ZN(n15078) );
  INV_X1 U17954 ( .A(n15078), .ZN(n14569) );
  INV_X1 U17955 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U17956 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14894), .ZN(n14567) );
  OAI21_X1 U17957 ( .B1(n20363), .B2(n14736), .A(n14567), .ZN(n14568) );
  AOI21_X1 U17958 ( .B1(n14569), .B2(n20345), .A(n14568), .ZN(n14571) );
  NAND2_X1 U17959 ( .A1(n14588), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14570) );
  OAI211_X1 U17960 ( .C1(n14572), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14571), 
        .B(n14570), .ZN(n14573) );
  AOI21_X1 U17961 ( .B1(n14898), .B2(n20327), .A(n14573), .ZN(n14574) );
  INV_X1 U17962 ( .A(n14574), .ZN(P1_U2813) );
  AOI21_X1 U17963 ( .B1(n14579), .B2(n9718), .A(n14578), .ZN(n15088) );
  INV_X1 U17964 ( .A(n15088), .ZN(n14583) );
  OAI22_X1 U17965 ( .A1(n14580), .A2(n20321), .B1(n20361), .B2(n14900), .ZN(
        n14581) );
  AOI21_X1 U17966 ( .B1(n20346), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14581), .ZN(
        n14582) );
  OAI21_X1 U17967 ( .B1(n14583), .B2(n20377), .A(n14582), .ZN(n14587) );
  INV_X1 U17968 ( .A(n14584), .ZN(n14608) );
  NOR3_X1 U17969 ( .A1(n14608), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14585), 
        .ZN(n14586) );
  AOI211_X1 U17970 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n14588), .A(n14587), 
        .B(n14586), .ZN(n14589) );
  OAI21_X1 U17971 ( .B1(n14906), .B2(n14732), .A(n14589), .ZN(P1_U2814) );
  XNOR2_X1 U17972 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14599) );
  AOI21_X1 U17973 ( .B1(n14591), .B2(n14601), .A(n14576), .ZN(n14917) );
  NAND2_X1 U17974 ( .A1(n14917), .A2(n20327), .ZN(n14598) );
  INV_X1 U17975 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14738) );
  AOI22_X1 U17976 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14913), .ZN(n14592) );
  OAI21_X1 U17977 ( .B1(n20363), .B2(n14738), .A(n14592), .ZN(n14596) );
  NAND2_X1 U17978 ( .A1(n14603), .A2(n14593), .ZN(n14594) );
  NAND2_X1 U17979 ( .A1(n9718), .A2(n14594), .ZN(n15095) );
  NOR2_X1 U17980 ( .A1(n15095), .A2(n20377), .ZN(n14595) );
  AOI211_X1 U17981 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14620), .A(n14596), 
        .B(n14595), .ZN(n14597) );
  OAI211_X1 U17982 ( .C1(n14608), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        P1_U2815) );
  OAI21_X1 U17983 ( .B1(n14600), .B2(n14602), .A(n14601), .ZN(n14927) );
  OAI21_X1 U17984 ( .B1(n14614), .B2(n14604), .A(n14603), .ZN(n15102) );
  OAI22_X1 U17985 ( .A1(n14605), .A2(n20321), .B1(n20361), .B2(n14919), .ZN(
        n14606) );
  AOI21_X1 U17986 ( .B1(n20346), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14606), .ZN(
        n14607) );
  OAI21_X1 U17987 ( .B1(n15102), .B2(n20377), .A(n14607), .ZN(n14610) );
  NOR2_X1 U17988 ( .A1(n14608), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14609) );
  AOI211_X1 U17989 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14620), .A(n14610), 
        .B(n14609), .ZN(n14611) );
  OAI21_X1 U17990 ( .B1(n14927), .B2(n14732), .A(n14611), .ZN(P1_U2816) );
  AOI21_X1 U17991 ( .B1(n14613), .B2(n14624), .A(n14600), .ZN(n14929) );
  INV_X1 U17992 ( .A(n14929), .ZN(n14816) );
  INV_X1 U17993 ( .A(n14614), .ZN(n14617) );
  NAND2_X1 U17994 ( .A1(n14628), .A2(n14615), .ZN(n14616) );
  NAND2_X1 U17995 ( .A1(n14617), .A2(n14616), .ZN(n14741) );
  INV_X1 U17996 ( .A(n14741), .ZN(n15118) );
  INV_X1 U17997 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U17998 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14932), .ZN(n14618) );
  OAI21_X1 U17999 ( .B1(n20363), .B2(n14740), .A(n14618), .ZN(n14619) );
  AOI21_X1 U18000 ( .B1(n15118), .B2(n20345), .A(n14619), .ZN(n14623) );
  INV_X1 U18001 ( .A(n14635), .ZN(n14643) );
  INV_X1 U18002 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21131) );
  INV_X1 U18003 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21168) );
  NOR3_X1 U18004 ( .A1(n14643), .A2(n21131), .A3(n21168), .ZN(n14621) );
  OAI21_X1 U18005 ( .B1(n14621), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14620), 
        .ZN(n14622) );
  OAI211_X1 U18006 ( .C1(n14816), .C2(n14732), .A(n14623), .B(n14622), .ZN(
        P1_U2817) );
  OAI21_X1 U18007 ( .B1(n9721), .B2(n14625), .A(n14624), .ZN(n14939) );
  XOR2_X1 U18008 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .Z(n14634) );
  NAND2_X1 U18009 ( .A1(n14640), .A2(n14626), .ZN(n14627) );
  NAND2_X1 U18010 ( .A1(n14628), .A2(n14627), .ZN(n16379) );
  NAND2_X1 U18011 ( .A1(n14656), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14632) );
  OAI22_X1 U18012 ( .A1(n14629), .A2(n20321), .B1(n20361), .B2(n14941), .ZN(
        n14630) );
  AOI21_X1 U18013 ( .B1(n20346), .B2(P1_EBX_REG_22__SCAN_IN), .A(n14630), .ZN(
        n14631) );
  OAI211_X1 U18014 ( .C1(n16379), .C2(n20377), .A(n14632), .B(n14631), .ZN(
        n14633) );
  AOI21_X1 U18015 ( .B1(n14635), .B2(n14634), .A(n14633), .ZN(n14636) );
  OAI21_X1 U18016 ( .B1(n14939), .B2(n14732), .A(n14636), .ZN(P1_U2818) );
  XNOR2_X1 U18017 ( .A(n9712), .B(n14637), .ZN(n14954) );
  NAND2_X1 U18018 ( .A1(n14652), .A2(n14638), .ZN(n14639) );
  NAND2_X1 U18019 ( .A1(n14640), .A2(n14639), .ZN(n15129) );
  AOI22_X1 U18020 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14947), .ZN(n14642) );
  NAND2_X1 U18021 ( .A1(n20346), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14641) );
  OAI211_X1 U18022 ( .C1(n15129), .C2(n20377), .A(n14642), .B(n14641), .ZN(
        n14645) );
  NOR2_X1 U18023 ( .A1(n14643), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14644) );
  AOI211_X1 U18024 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n14656), .A(n14645), 
        .B(n14644), .ZN(n14646) );
  OAI21_X1 U18025 ( .B1(n14954), .B2(n14732), .A(n14646), .ZN(P1_U2819) );
  INV_X1 U18026 ( .A(n14647), .ZN(n14649) );
  INV_X1 U18027 ( .A(n9743), .ZN(n14648) );
  AOI21_X1 U18028 ( .B1(n14649), .B2(n14648), .A(n9712), .ZN(n14960) );
  INV_X1 U18029 ( .A(n14960), .ZN(n14829) );
  OR2_X1 U18030 ( .A1(n14664), .A2(n14650), .ZN(n14651) );
  NAND2_X1 U18031 ( .A1(n14652), .A2(n14651), .ZN(n14745) );
  INV_X1 U18032 ( .A(n14745), .ZN(n15141) );
  INV_X1 U18033 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14744) );
  INV_X1 U18034 ( .A(n14958), .ZN(n14653) );
  AOI22_X1 U18035 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20365), .B1(
        n20319), .B2(n14653), .ZN(n14654) );
  OAI21_X1 U18036 ( .B1(n20363), .B2(n14744), .A(n14654), .ZN(n14655) );
  AOI21_X1 U18037 ( .B1(n15141), .B2(n20345), .A(n14655), .ZN(n14659) );
  AND3_X1 U18038 ( .A1(n14681), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14657) );
  OAI21_X1 U18039 ( .B1(n14657), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14656), 
        .ZN(n14658) );
  OAI211_X1 U18040 ( .C1(n14829), .C2(n14732), .A(n14659), .B(n14658), .ZN(
        P1_U2820) );
  AOI21_X1 U18041 ( .B1(n14661), .B2(n14660), .A(n9743), .ZN(n14969) );
  INV_X1 U18042 ( .A(n14969), .ZN(n14833) );
  NOR2_X1 U18043 ( .A1(n14677), .A2(n14662), .ZN(n14663) );
  OR2_X1 U18044 ( .A1(n14664), .A2(n14663), .ZN(n14747) );
  INV_X1 U18045 ( .A(n14747), .ZN(n16388) );
  INV_X1 U18046 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21014) );
  AOI21_X1 U18047 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20334), .ZN(n14666) );
  AOI22_X1 U18048 ( .A1(n20346), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n14965), 
        .B2(n20319), .ZN(n14665) );
  OAI211_X1 U18049 ( .C1(n21014), .C2(n14687), .A(n14666), .B(n14665), .ZN(
        n14670) );
  INV_X1 U18050 ( .A(n14681), .ZN(n14668) );
  XNOR2_X1 U18051 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14667) );
  NOR2_X1 U18052 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  AOI211_X1 U18053 ( .C1(n16388), .C2(n20345), .A(n14670), .B(n14669), .ZN(
        n14671) );
  OAI21_X1 U18054 ( .B1(n14833), .B2(n14732), .A(n14671), .ZN(P1_U2821) );
  OAI21_X1 U18055 ( .B1(n9715), .B2(n11100), .A(n14660), .ZN(n14979) );
  INV_X1 U18056 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14971) );
  INV_X1 U18057 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14748) );
  INV_X1 U18058 ( .A(n14974), .ZN(n14673) );
  OAI22_X1 U18059 ( .A1(n14748), .A2(n20363), .B1(n14673), .B2(n20361), .ZN(
        n14674) );
  AOI211_X1 U18060 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20334), .B(n14674), .ZN(n14679) );
  AND2_X1 U18061 ( .A1(n9705), .A2(n14675), .ZN(n14676) );
  NOR2_X1 U18062 ( .A1(n14677), .A2(n14676), .ZN(n16402) );
  NAND2_X1 U18063 ( .A1(n16402), .A2(n20345), .ZN(n14678) );
  OAI211_X1 U18064 ( .C1(n14687), .C2(n14971), .A(n14679), .B(n14678), .ZN(
        n14680) );
  AOI21_X1 U18065 ( .B1(n14681), .B2(n14971), .A(n14680), .ZN(n14682) );
  OAI21_X1 U18066 ( .B1(n14979), .B2(n14732), .A(n14682), .ZN(P1_U2822) );
  NAND2_X1 U18067 ( .A1(n9752), .A2(n14683), .ZN(n14684) );
  NAND2_X1 U18068 ( .A1(n9705), .A2(n14684), .ZN(n16409) );
  AOI21_X1 U18069 ( .B1(n14686), .B2(n14685), .A(n9715), .ZN(n14987) );
  NAND2_X1 U18070 ( .A1(n14987), .A2(n20327), .ZN(n14695) );
  AOI21_X1 U18071 ( .B1(n21010), .B2(n14688), .A(n14687), .ZN(n14693) );
  INV_X1 U18072 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14691) );
  INV_X1 U18073 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14751) );
  OAI22_X1 U18074 ( .A1(n20363), .A2(n14751), .B1(n14985), .B2(n20361), .ZN(
        n14689) );
  INV_X1 U18075 ( .A(n14689), .ZN(n14690) );
  OAI211_X1 U18076 ( .C1(n20321), .C2(n14691), .A(n14690), .B(n20347), .ZN(
        n14692) );
  NOR2_X1 U18077 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  OAI211_X1 U18078 ( .C1(n16409), .C2(n20377), .A(n14695), .B(n14694), .ZN(
        P1_U2823) );
  OAI21_X1 U18079 ( .B1(n14696), .B2(n14698), .A(n14697), .ZN(n14858) );
  AND2_X1 U18080 ( .A1(n14708), .A2(n14699), .ZN(n14700) );
  OR2_X1 U18081 ( .A1(n14700), .A2(n14758), .ZN(n15158) );
  AOI22_X1 U18082 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20365), .B1(
        n20346), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n14701) );
  OAI211_X1 U18083 ( .C1(n20377), .C2(n15158), .A(n14701), .B(n20347), .ZN(
        n14705) );
  NAND2_X1 U18084 ( .A1(n20352), .A2(n14702), .ZN(n16321) );
  AOI21_X1 U18085 ( .B1(n21004), .B2(n14703), .A(n16321), .ZN(n14704) );
  AOI211_X1 U18086 ( .C1(n16340), .C2(n20319), .A(n14705), .B(n14704), .ZN(
        n14706) );
  OAI21_X1 U18087 ( .B1(n14858), .B2(n14732), .A(n14706), .ZN(P1_U2826) );
  OAI21_X1 U18088 ( .B1(n9686), .B2(n14707), .A(n10161), .ZN(n15007) );
  INV_X1 U18089 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21003) );
  INV_X1 U18090 ( .A(n14708), .ZN(n14709) );
  AOI21_X1 U18091 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n16432) );
  AOI22_X1 U18092 ( .A1(n16432), .A2(n20345), .B1(n20346), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14712) );
  OAI211_X1 U18093 ( .C1(n20321), .C2(n14713), .A(n14712), .B(n20347), .ZN(
        n14714) );
  AOI21_X1 U18094 ( .B1(n14715), .B2(n21003), .A(n14714), .ZN(n14720) );
  NOR2_X1 U18095 ( .A1(n14717), .A2(n14716), .ZN(n14730) );
  INV_X1 U18096 ( .A(n14999), .ZN(n14718) );
  AOI22_X1 U18097 ( .A1(n14730), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n20319), 
        .B2(n14718), .ZN(n14719) );
  OAI211_X1 U18098 ( .C1(n15007), .C2(n14732), .A(n14720), .B(n14719), .ZN(
        P1_U2827) );
  NOR2_X1 U18099 ( .A1(n14722), .A2(n14721), .ZN(n14723) );
  NOR2_X1 U18100 ( .A1(n9686), .A2(n14723), .ZN(n16346) );
  INV_X1 U18101 ( .A(n16346), .ZN(n14864) );
  INV_X1 U18102 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20999) );
  OAI21_X1 U18103 ( .B1(n16329), .B2(n20999), .A(n21001), .ZN(n14729) );
  NOR2_X1 U18104 ( .A1(n14772), .A2(n20377), .ZN(n14728) );
  INV_X1 U18105 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14771) );
  NOR2_X1 U18106 ( .A1(n20321), .A2(n14724), .ZN(n14725) );
  AOI211_X1 U18107 ( .C1(n16345), .C2(n20319), .A(n20334), .B(n14725), .ZN(
        n14726) );
  OAI21_X1 U18108 ( .B1(n14771), .B2(n20363), .A(n14726), .ZN(n14727) );
  AOI211_X1 U18109 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14731) );
  OAI21_X1 U18110 ( .B1(n14864), .B2(n14732), .A(n14731), .ZN(P1_U2828) );
  OAI22_X1 U18111 ( .A1(n15017), .A2(n14765), .B1(n14733), .B2(n14770), .ZN(
        P1_U2841) );
  INV_X1 U18112 ( .A(n14879), .ZN(n14790) );
  OAI222_X1 U18113 ( .A1(n14734), .A2(n14770), .B1(n14765), .B2(n15059), .C1(
        n14790), .C2(n14769), .ZN(P1_U2843) );
  OAI222_X1 U18114 ( .A1(n15070), .A2(n14765), .B1(n14735), .B2(n14770), .C1(
        n14891), .C2(n14769), .ZN(P1_U2844) );
  INV_X1 U18115 ( .A(n14898), .ZN(n14797) );
  AOI22_X1 U18116 ( .A1(n15088), .A2(n14784), .B1(n14783), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14737) );
  OAI21_X1 U18117 ( .B1(n14906), .B2(n14769), .A(n14737), .ZN(P1_U2846) );
  INV_X1 U18118 ( .A(n14917), .ZN(n14806) );
  OAI222_X1 U18119 ( .A1(n15095), .A2(n14765), .B1(n14738), .B2(n14770), .C1(
        n14806), .C2(n14769), .ZN(P1_U2847) );
  INV_X1 U18120 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14739) );
  OAI222_X1 U18121 ( .A1(n15102), .A2(n14765), .B1(n14739), .B2(n14770), .C1(
        n14927), .C2(n14769), .ZN(P1_U2848) );
  OAI222_X1 U18122 ( .A1(n14741), .A2(n14765), .B1(n14740), .B2(n14770), .C1(
        n14816), .C2(n14769), .ZN(P1_U2849) );
  INV_X1 U18123 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14742) );
  OAI222_X1 U18124 ( .A1(n16379), .A2(n14765), .B1(n14742), .B2(n14770), .C1(
        n14939), .C2(n14769), .ZN(P1_U2850) );
  INV_X1 U18125 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14743) );
  OAI222_X1 U18126 ( .A1(n15129), .A2(n14765), .B1(n14743), .B2(n14770), .C1(
        n14954), .C2(n14769), .ZN(P1_U2851) );
  OAI222_X1 U18127 ( .A1(n14745), .A2(n14765), .B1(n14744), .B2(n14770), .C1(
        n14829), .C2(n14769), .ZN(P1_U2852) );
  INV_X1 U18128 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14746) );
  OAI222_X1 U18129 ( .A1(n14747), .A2(n14765), .B1(n14746), .B2(n14770), .C1(
        n14833), .C2(n14769), .ZN(P1_U2853) );
  NOR2_X1 U18130 ( .A1(n14770), .A2(n14748), .ZN(n14749) );
  AOI21_X1 U18131 ( .B1(n16402), .B2(n14784), .A(n14749), .ZN(n14750) );
  OAI21_X1 U18132 ( .B1(n14979), .B2(n14769), .A(n14750), .ZN(P1_U2854) );
  INV_X1 U18133 ( .A(n14987), .ZN(n14846) );
  OAI222_X1 U18134 ( .A1(n16409), .A2(n14765), .B1(n14751), .B2(n14770), .C1(
        n14846), .C2(n14769), .ZN(P1_U2855) );
  OAI21_X1 U18135 ( .B1(n9677), .B2(n14752), .A(n14685), .ZN(n14854) );
  INV_X1 U18136 ( .A(n14854), .ZN(n16336) );
  OR2_X1 U18137 ( .A1(n14760), .A2(n14753), .ZN(n14754) );
  NAND2_X1 U18138 ( .A1(n9752), .A2(n14754), .ZN(n16419) );
  INV_X1 U18139 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16307) );
  OAI22_X1 U18140 ( .A1(n16419), .A2(n14765), .B1(n16307), .B2(n14770), .ZN(
        n14755) );
  AOI21_X1 U18141 ( .B1(n16336), .B2(n14774), .A(n14755), .ZN(n14756) );
  INV_X1 U18142 ( .A(n14756), .ZN(P1_U2856) );
  NOR2_X1 U18143 ( .A1(n14758), .A2(n14757), .ZN(n14759) );
  OR2_X1 U18144 ( .A1(n14760), .A2(n14759), .ZN(n16426) );
  INV_X1 U18145 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14763) );
  AND2_X1 U18146 ( .A1(n14697), .A2(n14761), .ZN(n14762) );
  OR2_X1 U18147 ( .A1(n14762), .A2(n9677), .ZN(n14995) );
  OAI222_X1 U18148 ( .A1(n16426), .A2(n14765), .B1(n14770), .B2(n14763), .C1(
        n14769), .C2(n14995), .ZN(P1_U2857) );
  INV_X1 U18149 ( .A(n14858), .ZN(n16341) );
  INV_X1 U18150 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14764) );
  OAI22_X1 U18151 ( .A1(n15158), .A2(n14765), .B1(n14764), .B2(n14770), .ZN(
        n14766) );
  AOI21_X1 U18152 ( .B1(n16341), .B2(n14774), .A(n14766), .ZN(n14767) );
  INV_X1 U18153 ( .A(n14767), .ZN(P1_U2858) );
  AOI22_X1 U18154 ( .A1(n16432), .A2(n14784), .B1(n14783), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14768) );
  OAI21_X1 U18155 ( .B1(n15007), .B2(n14769), .A(n14768), .ZN(P1_U2859) );
  OAI22_X1 U18156 ( .A1(n14772), .A2(n14765), .B1(n14771), .B2(n14770), .ZN(
        n14773) );
  AOI21_X1 U18157 ( .B1(n16346), .B2(n14774), .A(n14773), .ZN(n14775) );
  INV_X1 U18158 ( .A(n14775), .ZN(P1_U2860) );
  NAND2_X1 U18159 ( .A1(n14777), .A2(n14776), .ZN(n14778) );
  AND2_X1 U18160 ( .A1(n14779), .A2(n14778), .ZN(n16356) );
  INV_X1 U18161 ( .A(n16356), .ZN(n14870) );
  AOI21_X1 U18162 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n16438) );
  AOI22_X1 U18163 ( .A1(n16438), .A2(n14784), .B1(n14783), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U18164 ( .B1(n14870), .B2(n14769), .A(n14785), .ZN(P1_U2861) );
  OAI22_X1 U18165 ( .A1(n14824), .A2(n16812), .B1(n14786), .B2(n14865), .ZN(
        n14788) );
  NOR2_X1 U18166 ( .A1(n14840), .A2(n14860), .ZN(n14787) );
  AOI211_X1 U18167 ( .C1(n9632), .C2(DATAI_29_), .A(n14788), .B(n14787), .ZN(
        n14789) );
  OAI21_X1 U18168 ( .B1(n14790), .B2(n14869), .A(n14789), .ZN(P1_U2875) );
  AOI22_X1 U18169 ( .A1(n14848), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14847), .ZN(n14792) );
  AOI22_X1 U18170 ( .A1(n9632), .A2(DATAI_28_), .B1(n14850), .B2(n14861), .ZN(
        n14791) );
  OAI211_X1 U18171 ( .C1(n14891), .C2(n14869), .A(n14792), .B(n14791), .ZN(
        P1_U2876) );
  NOR2_X1 U18172 ( .A1(n14865), .A2(n14793), .ZN(n14795) );
  OAI22_X1 U18173 ( .A1(n21270), .A2(n21149), .B1(n14867), .B2(n14840), .ZN(
        n14794) );
  AOI211_X1 U18174 ( .C1(n14848), .C2(BUF1_REG_27__SCAN_IN), .A(n14795), .B(
        n14794), .ZN(n14796) );
  OAI21_X1 U18175 ( .B1(n14797), .B2(n14869), .A(n14796), .ZN(P1_U2877) );
  AOI22_X1 U18176 ( .A1(n14848), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14847), .ZN(n14800) );
  AOI22_X1 U18177 ( .A1(n9632), .A2(DATAI_26_), .B1(n14850), .B2(n14798), .ZN(
        n14799) );
  OAI211_X1 U18178 ( .C1(n14906), .C2(n14869), .A(n14800), .B(n14799), .ZN(
        P1_U2878) );
  OAI22_X1 U18179 ( .A1(n14824), .A2(n16820), .B1(n14801), .B2(n14865), .ZN(
        n14802) );
  INV_X1 U18180 ( .A(n14802), .ZN(n14805) );
  AOI22_X1 U18181 ( .A1(n9632), .A2(DATAI_25_), .B1(n14850), .B2(n14803), .ZN(
        n14804) );
  OAI211_X1 U18182 ( .C1(n14806), .C2(n14869), .A(n14805), .B(n14804), .ZN(
        P1_U2879) );
  OAI22_X1 U18183 ( .A1(n14824), .A2(n16822), .B1(n13604), .B2(n14865), .ZN(
        n14809) );
  NOR2_X1 U18184 ( .A1(n14840), .A2(n14807), .ZN(n14808) );
  AOI211_X1 U18185 ( .C1(n9632), .C2(DATAI_24_), .A(n14809), .B(n14808), .ZN(
        n14810) );
  OAI21_X1 U18186 ( .B1(n14927), .B2(n14869), .A(n14810), .ZN(P1_U2880) );
  OAI22_X1 U18187 ( .A1(n14824), .A2(n16824), .B1(n14811), .B2(n14865), .ZN(
        n14812) );
  INV_X1 U18188 ( .A(n14812), .ZN(n14815) );
  AOI22_X1 U18189 ( .A1(n9632), .A2(DATAI_23_), .B1(n14850), .B2(n14813), .ZN(
        n14814) );
  OAI211_X1 U18190 ( .C1(n14816), .C2(n14869), .A(n14815), .B(n14814), .ZN(
        P1_U2881) );
  AOI22_X1 U18191 ( .A1(n14848), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14847), .ZN(n14819) );
  AOI22_X1 U18192 ( .A1(n9632), .A2(DATAI_22_), .B1(n14850), .B2(n14817), .ZN(
        n14818) );
  OAI211_X1 U18193 ( .C1(n14939), .C2(n14869), .A(n14819), .B(n14818), .ZN(
        P1_U2882) );
  NOR2_X1 U18194 ( .A1(n14824), .A2(n16828), .ZN(n14822) );
  OAI22_X1 U18195 ( .A1(n21270), .A2(n13426), .B1(n14820), .B2(n14840), .ZN(
        n14821) );
  AOI211_X1 U18196 ( .C1(n14847), .C2(P1_EAX_REG_21__SCAN_IN), .A(n14822), .B(
        n14821), .ZN(n14823) );
  OAI21_X1 U18197 ( .B1(n14954), .B2(n14869), .A(n14823), .ZN(P1_U2883) );
  NOR2_X1 U18198 ( .A1(n14824), .A2(n16830), .ZN(n14827) );
  OAI22_X1 U18199 ( .A1(n21270), .A2(n13414), .B1(n14825), .B2(n14840), .ZN(
        n14826) );
  AOI211_X1 U18200 ( .C1(n14847), .C2(P1_EAX_REG_20__SCAN_IN), .A(n14827), .B(
        n14826), .ZN(n14828) );
  OAI21_X1 U18201 ( .B1(n14829), .B2(n14869), .A(n14828), .ZN(P1_U2884) );
  AOI22_X1 U18202 ( .A1(n14848), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14847), .ZN(n14832) );
  AOI22_X1 U18203 ( .A1(n9632), .A2(DATAI_19_), .B1(n14850), .B2(n14830), .ZN(
        n14831) );
  OAI211_X1 U18204 ( .C1(n14833), .C2(n14869), .A(n14832), .B(n14831), .ZN(
        P1_U2885) );
  NOR2_X1 U18205 ( .A1(n14865), .A2(n14834), .ZN(n14837) );
  OAI22_X1 U18206 ( .A1(n21270), .A2(n13420), .B1(n14835), .B2(n14840), .ZN(
        n14836) );
  AOI211_X1 U18207 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n14848), .A(n14837), .B(
        n14836), .ZN(n14838) );
  OAI21_X1 U18208 ( .B1(n14979), .B2(n14869), .A(n14838), .ZN(P1_U2886) );
  NOR2_X1 U18209 ( .A1(n14865), .A2(n14839), .ZN(n14844) );
  OAI22_X1 U18210 ( .A1(n21270), .A2(n21147), .B1(n14841), .B2(n14840), .ZN(
        n14843) );
  AOI211_X1 U18211 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n14848), .A(n14844), .B(
        n14843), .ZN(n14845) );
  OAI21_X1 U18212 ( .B1(n14846), .B2(n14869), .A(n14845), .ZN(P1_U2887) );
  AOI22_X1 U18213 ( .A1(n14848), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14847), .ZN(n14853) );
  AOI22_X1 U18214 ( .A1(n9632), .A2(DATAI_16_), .B1(n14850), .B2(n14849), .ZN(
        n14852) );
  OAI211_X1 U18215 ( .C1(n14854), .C2(n14869), .A(n14853), .B(n14852), .ZN(
        P1_U2888) );
  OAI222_X1 U18216 ( .A1(n14995), .A2(n14869), .B1(n14868), .B2(n14856), .C1(
        n14865), .C2(n14855), .ZN(P1_U2889) );
  OAI222_X1 U18217 ( .A1(n14858), .A2(n14869), .B1(n14868), .B2(n14857), .C1(
        n20383), .C2(n14865), .ZN(P1_U2890) );
  OAI222_X1 U18218 ( .A1(n15007), .A2(n14869), .B1(n14868), .B2(n14860), .C1(
        n14859), .C2(n14865), .ZN(P1_U2891) );
  INV_X1 U18219 ( .A(n14861), .ZN(n14863) );
  OAI222_X1 U18220 ( .A1(n14864), .A2(n14869), .B1(n14868), .B2(n14863), .C1(
        n14862), .C2(n14865), .ZN(P1_U2892) );
  INV_X1 U18221 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14866) );
  OAI222_X1 U18222 ( .A1(n14870), .A2(n14869), .B1(n14868), .B2(n14867), .C1(
        n14866), .C2(n14865), .ZN(P1_U2893) );
  NAND2_X1 U18223 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  XNOR2_X1 U18224 ( .A(n14874), .B(n14873), .ZN(n15063) );
  NAND2_X1 U18225 ( .A1(n16361), .A2(n14875), .ZN(n14876) );
  NAND2_X1 U18226 ( .A1(n20334), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15058) );
  OAI211_X1 U18227 ( .C1(n16375), .C2(n14877), .A(n14876), .B(n15058), .ZN(
        n14878) );
  AOI21_X1 U18228 ( .B1(n14879), .B2(n16364), .A(n14878), .ZN(n14880) );
  OAI21_X1 U18229 ( .B1(n16349), .B2(n15063), .A(n14880), .ZN(P1_U2970) );
  NOR2_X1 U18230 ( .A1(n20347), .A2(n21138), .ZN(n15065) );
  NOR2_X1 U18231 ( .A1(n16370), .A2(n14881), .ZN(n14882) );
  AOI211_X1 U18232 ( .C1(n16351), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15065), .B(n14882), .ZN(n14890) );
  NOR2_X1 U18233 ( .A1(n10723), .A2(n15074), .ZN(n14886) );
  NOR3_X1 U18234 ( .A1(n10723), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14884), .ZN(n14885) );
  XNOR2_X1 U18235 ( .A(n14888), .B(n14887), .ZN(n15064) );
  NAND2_X1 U18236 ( .A1(n15064), .A2(n20302), .ZN(n14889) );
  OAI211_X1 U18237 ( .C1(n14891), .C2(n16371), .A(n14890), .B(n14889), .ZN(
        P1_U2971) );
  NOR2_X1 U18238 ( .A1(n14892), .A2(n14903), .ZN(n14893) );
  XNOR2_X1 U18239 ( .A(n14893), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15082) );
  NAND2_X1 U18240 ( .A1(n16361), .A2(n14894), .ZN(n14895) );
  NAND2_X1 U18241 ( .A1(n20334), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15077) );
  OAI211_X1 U18242 ( .C1(n16375), .C2(n14896), .A(n14895), .B(n15077), .ZN(
        n14897) );
  AOI21_X1 U18243 ( .B1(n14898), .B2(n16364), .A(n14897), .ZN(n14899) );
  OAI21_X1 U18244 ( .B1(n16349), .B2(n15082), .A(n14899), .ZN(P1_U2972) );
  NOR2_X1 U18245 ( .A1(n20347), .A2(n21173), .ZN(n15087) );
  NOR2_X1 U18246 ( .A1(n16370), .A2(n14900), .ZN(n14901) );
  AOI211_X1 U18247 ( .C1(n16351), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15087), .B(n14901), .ZN(n14905) );
  INV_X1 U18248 ( .A(n14902), .ZN(n15084) );
  NAND2_X1 U18249 ( .A1(n14903), .A2(n15091), .ZN(n15083) );
  NAND3_X1 U18250 ( .A1(n15084), .A2(n20302), .A3(n15083), .ZN(n14904) );
  OAI211_X1 U18251 ( .C1(n14906), .C2(n16371), .A(n14905), .B(n14904), .ZN(
        P1_U2973) );
  AOI21_X1 U18252 ( .B1(n14907), .B2(n10723), .A(n15115), .ZN(n14922) );
  MUX2_X1 U18253 ( .A(n16352), .B(n14922), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n14910) );
  OR2_X1 U18254 ( .A1(n10723), .A2(n15115), .ZN(n14908) );
  NAND3_X1 U18255 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n14912) );
  XNOR2_X1 U18256 ( .A(n14912), .B(n14911), .ZN(n15100) );
  NAND2_X1 U18257 ( .A1(n16361), .A2(n14913), .ZN(n14914) );
  NAND2_X1 U18258 ( .A1(n20334), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15094) );
  OAI211_X1 U18259 ( .C1(n16375), .C2(n14915), .A(n14914), .B(n15094), .ZN(
        n14916) );
  AOI21_X1 U18260 ( .B1(n14917), .B2(n16364), .A(n14916), .ZN(n14918) );
  OAI21_X1 U18261 ( .B1(n16349), .B2(n15100), .A(n14918), .ZN(P1_U2974) );
  INV_X1 U18262 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21095) );
  NOR2_X1 U18263 ( .A1(n20347), .A2(n21095), .ZN(n15103) );
  NOR2_X1 U18264 ( .A1(n16370), .A2(n14919), .ZN(n14920) );
  AOI211_X1 U18265 ( .C1(n16351), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15103), .B(n14920), .ZN(n14926) );
  NOR2_X1 U18266 ( .A1(n14922), .A2(n14921), .ZN(n14923) );
  MUX2_X1 U18267 ( .A(n14923), .B(n14922), .S(n10723), .Z(n14924) );
  XNOR2_X1 U18268 ( .A(n14924), .B(n15106), .ZN(n15101) );
  NAND2_X1 U18269 ( .A1(n15101), .A2(n20302), .ZN(n14925) );
  OAI211_X1 U18270 ( .C1(n14927), .C2(n16371), .A(n14926), .B(n14925), .ZN(
        P1_U2975) );
  XNOR2_X1 U18271 ( .A(n10723), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14928) );
  XNOR2_X1 U18272 ( .A(n14921), .B(n14928), .ZN(n15120) );
  NAND2_X1 U18273 ( .A1(n14929), .A2(n16364), .ZN(n14934) );
  INV_X1 U18274 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21018) );
  OAI22_X1 U18275 ( .A1(n16375), .A2(n14930), .B1(n20347), .B2(n21018), .ZN(
        n14931) );
  AOI21_X1 U18276 ( .B1(n16361), .B2(n14932), .A(n14931), .ZN(n14933) );
  OAI211_X1 U18277 ( .C1(n15120), .C2(n16349), .A(n14934), .B(n14933), .ZN(
        P1_U2976) );
  NAND2_X1 U18278 ( .A1(n14936), .A2(n14935), .ZN(n14938) );
  XNOR2_X1 U18279 ( .A(n14938), .B(n14937), .ZN(n16377) );
  INV_X1 U18280 ( .A(n14939), .ZN(n14943) );
  AOI22_X1 U18281 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14940) );
  OAI21_X1 U18282 ( .B1(n14941), .B2(n16370), .A(n14940), .ZN(n14942) );
  AOI21_X1 U18283 ( .B1(n14943), .B2(n16364), .A(n14942), .ZN(n14944) );
  OAI21_X1 U18284 ( .B1(n16349), .B2(n16377), .A(n14944), .ZN(P1_U2977) );
  NOR2_X1 U18285 ( .A1(n20347), .A2(n21131), .ZN(n15127) );
  NOR2_X1 U18286 ( .A1(n16375), .A2(n14945), .ZN(n14946) );
  AOI211_X1 U18287 ( .C1(n16361), .C2(n14947), .A(n15127), .B(n14946), .ZN(
        n14953) );
  NOR2_X1 U18288 ( .A1(n14948), .A2(n15134), .ZN(n14949) );
  MUX2_X1 U18289 ( .A(n14950), .B(n14949), .S(n10723), .Z(n14951) );
  XNOR2_X1 U18290 ( .A(n14951), .B(n15133), .ZN(n15121) );
  NAND2_X1 U18291 ( .A1(n15121), .A2(n20302), .ZN(n14952) );
  OAI211_X1 U18292 ( .C1(n14954), .C2(n16371), .A(n14953), .B(n14952), .ZN(
        P1_U2978) );
  NOR2_X1 U18293 ( .A1(n14948), .A2(n16393), .ZN(n14955) );
  MUX2_X1 U18294 ( .A(n9739), .B(n14955), .S(n10723), .Z(n14956) );
  XNOR2_X1 U18295 ( .A(n14956), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15143) );
  INV_X1 U18296 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21164) );
  NOR2_X1 U18297 ( .A1(n20347), .A2(n21164), .ZN(n15140) );
  AOI21_X1 U18298 ( .B1(n16351), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15140), .ZN(n14957) );
  OAI21_X1 U18299 ( .B1(n14958), .B2(n16370), .A(n14957), .ZN(n14959) );
  AOI21_X1 U18300 ( .B1(n14960), .B2(n16364), .A(n14959), .ZN(n14961) );
  OAI21_X1 U18301 ( .B1(n16349), .B2(n15143), .A(n14961), .ZN(P1_U2979) );
  NAND2_X1 U18302 ( .A1(n14948), .A2(n14962), .ZN(n14964) );
  XNOR2_X1 U18303 ( .A(n10723), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14963) );
  XNOR2_X1 U18304 ( .A(n14964), .B(n14963), .ZN(n16387) );
  INV_X1 U18305 ( .A(n14965), .ZN(n14967) );
  AOI22_X1 U18306 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14966) );
  OAI21_X1 U18307 ( .B1(n14967), .B2(n16370), .A(n14966), .ZN(n14968) );
  AOI21_X1 U18308 ( .B1(n14969), .B2(n16364), .A(n14968), .ZN(n14970) );
  OAI21_X1 U18309 ( .B1(n16387), .B2(n16349), .A(n14970), .ZN(P1_U2980) );
  OAI22_X1 U18310 ( .A1(n16375), .A2(n14972), .B1(n20347), .B2(n14971), .ZN(
        n14973) );
  AOI21_X1 U18311 ( .B1(n16361), .B2(n14974), .A(n14973), .ZN(n14978) );
  OR2_X1 U18312 ( .A1(n14976), .A2(n14975), .ZN(n16399) );
  NAND3_X1 U18313 ( .A1(n16399), .A2(n14948), .A3(n20302), .ZN(n14977) );
  OAI211_X1 U18314 ( .C1(n14979), .C2(n16371), .A(n14978), .B(n14977), .ZN(
        P1_U2981) );
  NOR2_X1 U18315 ( .A1(n10723), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14982) );
  NAND2_X1 U18316 ( .A1(n14980), .A2(n16330), .ZN(n14981) );
  MUX2_X1 U18317 ( .A(n14982), .B(n10723), .S(n14981), .Z(n14983) );
  XNOR2_X1 U18318 ( .A(n14983), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16408) );
  AOI22_X1 U18319 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14984) );
  OAI21_X1 U18320 ( .B1(n14985), .B2(n16370), .A(n14984), .ZN(n14986) );
  AOI21_X1 U18321 ( .B1(n14987), .B2(n16364), .A(n14986), .ZN(n14988) );
  OAI21_X1 U18322 ( .B1(n16408), .B2(n16349), .A(n14988), .ZN(P1_U2982) );
  INV_X1 U18323 ( .A(n16331), .ZN(n14989) );
  NOR2_X1 U18324 ( .A1(n14990), .A2(n14989), .ZN(n14994) );
  NOR2_X1 U18325 ( .A1(n12829), .A2(n14991), .ZN(n16333) );
  NOR2_X1 U18326 ( .A1(n16333), .A2(n14992), .ZN(n14993) );
  XOR2_X1 U18327 ( .A(n14994), .B(n14993), .Z(n16425) );
  INV_X1 U18328 ( .A(n14995), .ZN(n16318) );
  AOI22_X1 U18329 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14996) );
  OAI21_X1 U18330 ( .B1(n16313), .B2(n16370), .A(n14996), .ZN(n14997) );
  AOI21_X1 U18331 ( .B1(n16318), .B2(n16364), .A(n14997), .ZN(n14998) );
  OAI21_X1 U18332 ( .B1(n16425), .B2(n16349), .A(n14998), .ZN(P1_U2984) );
  NOR2_X1 U18333 ( .A1(n20347), .A2(n21003), .ZN(n16431) );
  NOR2_X1 U18334 ( .A1(n16370), .A2(n14999), .ZN(n15000) );
  AOI211_X1 U18335 ( .C1(n16351), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16431), .B(n15000), .ZN(n15006) );
  OAI21_X1 U18336 ( .B1(n15002), .B2(n15144), .A(n15001), .ZN(n15004) );
  XNOR2_X1 U18337 ( .A(n15004), .B(n15003), .ZN(n16434) );
  NAND2_X1 U18338 ( .A1(n16434), .A2(n20302), .ZN(n15005) );
  OAI211_X1 U18339 ( .C1(n15007), .C2(n16371), .A(n15006), .B(n15005), .ZN(
        P1_U2986) );
  AND2_X1 U18340 ( .A1(n15008), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15010) );
  XNOR2_X1 U18341 ( .A(n12829), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15009) );
  MUX2_X1 U18342 ( .A(n15010), .B(n15009), .S(n10723), .Z(n15011) );
  NOR3_X1 U18343 ( .A1(n15008), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10723), .ZN(n16353) );
  NOR2_X1 U18344 ( .A1(n15011), .A2(n16353), .ZN(n16452) );
  AOI22_X1 U18345 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15012) );
  OAI21_X1 U18346 ( .B1(n15013), .B2(n16370), .A(n15012), .ZN(n15014) );
  AOI21_X1 U18347 ( .B1(n15015), .B2(n16364), .A(n15014), .ZN(n15016) );
  OAI21_X1 U18348 ( .B1(n16452), .B2(n16349), .A(n15016), .ZN(P1_U2989) );
  INV_X1 U18349 ( .A(n15017), .ZN(n15028) );
  OR2_X1 U18350 ( .A1(n15019), .A2(n15018), .ZN(n15124) );
  NOR2_X1 U18351 ( .A1(n15021), .A2(n15124), .ZN(n15030) );
  INV_X1 U18352 ( .A(n15030), .ZN(n15150) );
  NAND3_X1 U18353 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n15020), .ZN(n15123) );
  NOR2_X1 U18354 ( .A1(n15021), .A2(n15123), .ZN(n15152) );
  NAND2_X1 U18355 ( .A1(n15022), .A2(n15152), .ZN(n15105) );
  INV_X1 U18356 ( .A(n15023), .ZN(n15024) );
  NAND4_X1 U18357 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16406) );
  NOR2_X1 U18358 ( .A1(n16398), .A2(n16406), .ZN(n15029) );
  NAND4_X1 U18359 ( .A1(n16418), .A2(n15024), .A3(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n15029), .ZN(n15116) );
  NAND2_X1 U18360 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15038) );
  NOR2_X1 U18361 ( .A1(n15093), .A2(n15038), .ZN(n15075) );
  NAND3_X1 U18362 ( .A1(n15075), .A2(n10746), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15049) );
  INV_X1 U18363 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15025) );
  NOR3_X1 U18364 ( .A1(n15049), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15025), .ZN(n15026) );
  AOI211_X1 U18365 ( .C1(n15028), .C2(n20438), .A(n15027), .B(n15026), .ZN(
        n15043) );
  NAND2_X1 U18366 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15029), .ZN(
        n15126) );
  OAI221_X1 U18367 ( .B1(n20442), .B2(n15030), .C1(n20442), .C2(n15029), .A(
        n16445), .ZN(n15031) );
  AOI221_X1 U18368 ( .B1(n15123), .B2(n15154), .C1(n15126), .C2(n15154), .A(
        n15031), .ZN(n16390) );
  NAND2_X1 U18369 ( .A1(n16390), .A2(n15032), .ZN(n15033) );
  NAND2_X1 U18370 ( .A1(n15041), .A2(n16445), .ZN(n16449) );
  NAND2_X1 U18371 ( .A1(n15033), .A2(n16449), .ZN(n16378) );
  NAND2_X1 U18372 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U18373 ( .A1(n16416), .A2(n16383), .ZN(n15034) );
  AND2_X1 U18374 ( .A1(n16378), .A2(n15034), .ZN(n15114) );
  OR2_X1 U18375 ( .A1(n20442), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15035) );
  NAND2_X1 U18376 ( .A1(n15114), .A2(n15035), .ZN(n15109) );
  AND2_X1 U18377 ( .A1(n16416), .A2(n15036), .ZN(n15037) );
  AND2_X1 U18378 ( .A1(n16416), .A2(n15038), .ZN(n15039) );
  AND2_X1 U18379 ( .A1(n16416), .A2(n15067), .ZN(n15040) );
  NOR2_X1 U18380 ( .A1(n15080), .A2(n15040), .ZN(n15055) );
  OAI211_X1 U18381 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15041), .A(
        n15055), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15050) );
  NAND3_X1 U18382 ( .A1(n15050), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16449), .ZN(n15042) );
  INV_X1 U18383 ( .A(n15045), .ZN(n15054) );
  INV_X1 U18384 ( .A(n15046), .ZN(n15048) );
  AOI21_X1 U18385 ( .B1(n15048), .B2(n20438), .A(n15047), .ZN(n15053) );
  INV_X1 U18386 ( .A(n15049), .ZN(n15051) );
  OAI21_X1 U18387 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15051), .A(
        n15050), .ZN(n15052) );
  OAI211_X1 U18388 ( .C1(n15054), .C2(n20431), .A(n15053), .B(n15052), .ZN(
        P1_U3001) );
  INV_X1 U18389 ( .A(n15055), .ZN(n15061) );
  NAND3_X1 U18390 ( .A1(n15075), .A2(n10746), .A3(n15056), .ZN(n15057) );
  OAI211_X1 U18391 ( .C1(n15059), .C2(n16466), .A(n15058), .B(n15057), .ZN(
        n15060) );
  AOI21_X1 U18392 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15061), .A(
        n15060), .ZN(n15062) );
  OAI21_X1 U18393 ( .B1(n15063), .B2(n20431), .A(n15062), .ZN(P1_U3002) );
  INV_X1 U18394 ( .A(n15064), .ZN(n15073) );
  INV_X1 U18395 ( .A(n15065), .ZN(n15069) );
  NAND3_X1 U18396 ( .A1(n15075), .A2(n15067), .A3(n15066), .ZN(n15068) );
  OAI211_X1 U18397 ( .C1(n15070), .C2(n16466), .A(n15069), .B(n15068), .ZN(
        n15071) );
  AOI21_X1 U18398 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15080), .A(
        n15071), .ZN(n15072) );
  OAI21_X1 U18399 ( .B1(n15073), .B2(n20431), .A(n15072), .ZN(P1_U3003) );
  NAND2_X1 U18400 ( .A1(n15075), .A2(n15074), .ZN(n15076) );
  OAI211_X1 U18401 ( .C1(n15078), .C2(n16466), .A(n15077), .B(n15076), .ZN(
        n15079) );
  AOI21_X1 U18402 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15080), .A(
        n15079), .ZN(n15081) );
  OAI21_X1 U18403 ( .B1(n15082), .B2(n20431), .A(n15081), .ZN(P1_U3004) );
  INV_X1 U18404 ( .A(n15098), .ZN(n15092) );
  NAND3_X1 U18405 ( .A1(n15084), .A2(n20439), .A3(n15083), .ZN(n15090) );
  XNOR2_X1 U18406 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15085) );
  NOR2_X1 U18407 ( .A1(n15093), .A2(n15085), .ZN(n15086) );
  AOI211_X1 U18408 ( .C1(n15088), .C2(n20438), .A(n15087), .B(n15086), .ZN(
        n15089) );
  OAI211_X1 U18409 ( .C1(n15092), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        P1_U3005) );
  NOR2_X1 U18410 ( .A1(n15093), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15097) );
  OAI21_X1 U18411 ( .B1(n15095), .B2(n16466), .A(n15094), .ZN(n15096) );
  AOI211_X1 U18412 ( .C1(n15098), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15097), .B(n15096), .ZN(n15099) );
  OAI21_X1 U18413 ( .B1(n15100), .B2(n20431), .A(n15099), .ZN(P1_U3006) );
  INV_X1 U18414 ( .A(n15101), .ZN(n15112) );
  INV_X1 U18415 ( .A(n15102), .ZN(n15104) );
  AOI21_X1 U18416 ( .B1(n15104), .B2(n20438), .A(n15103), .ZN(n15111) );
  OAI21_X1 U18417 ( .B1(n15105), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15108) );
  OAI21_X1 U18418 ( .B1(n15115), .B2(n15116), .A(n15106), .ZN(n15107) );
  OAI21_X1 U18419 ( .B1(n15109), .B2(n15108), .A(n15107), .ZN(n15110) );
  OAI211_X1 U18420 ( .C1(n15112), .C2(n20431), .A(n15111), .B(n15110), .ZN(
        P1_U3007) );
  NAND2_X1 U18421 ( .A1(n20334), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15113) );
  OAI221_X1 U18422 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15116), 
        .C1(n15115), .C2(n15114), .A(n15113), .ZN(n15117) );
  AOI21_X1 U18423 ( .B1(n15118), .B2(n20438), .A(n15117), .ZN(n15119) );
  OAI21_X1 U18424 ( .B1(n15120), .B2(n20431), .A(n15119), .ZN(P1_U3008) );
  NAND2_X1 U18425 ( .A1(n15121), .A2(n20439), .ZN(n15132) );
  INV_X1 U18426 ( .A(n15123), .ZN(n15125) );
  NAND2_X1 U18427 ( .A1(n20441), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15122) );
  OAI22_X1 U18428 ( .A1(n20442), .A2(n15124), .B1(n15123), .B2(n15122), .ZN(
        n15135) );
  AOI21_X1 U18429 ( .B1(n20447), .B2(n15125), .A(n15135), .ZN(n16437) );
  NOR2_X1 U18430 ( .A1(n16437), .A2(n15126), .ZN(n16394) );
  NAND2_X1 U18431 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16394), .ZN(
        n15136) );
  NOR2_X1 U18432 ( .A1(n15137), .A2(n15136), .ZN(n16384) );
  INV_X1 U18433 ( .A(n15127), .ZN(n15128) );
  OAI21_X1 U18434 ( .B1(n15129), .B2(n16466), .A(n15128), .ZN(n15130) );
  AOI21_X1 U18435 ( .B1(n16384), .B2(n15133), .A(n15130), .ZN(n15131) );
  OAI211_X1 U18436 ( .C1(n16378), .C2(n15133), .A(n15132), .B(n15131), .ZN(
        P1_U3010) );
  OAI21_X1 U18437 ( .B1(n20447), .B2(n15135), .A(n15134), .ZN(n15138) );
  AOI22_X1 U18438 ( .A1(n16390), .A2(n15138), .B1(n15137), .B2(n15136), .ZN(
        n15139) );
  AOI211_X1 U18439 ( .C1(n20438), .C2(n15141), .A(n15140), .B(n15139), .ZN(
        n15142) );
  OAI21_X1 U18440 ( .B1(n15143), .B2(n20431), .A(n15142), .ZN(P1_U3011) );
  INV_X1 U18441 ( .A(n15144), .ZN(n15146) );
  AOI21_X1 U18442 ( .B1(n12829), .B2(n15146), .A(n15145), .ZN(n15147) );
  AOI21_X1 U18443 ( .B1(n16352), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15147), .ZN(n15149) );
  INV_X1 U18444 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16417) );
  MUX2_X1 U18445 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n16417), .S(
        n10723), .Z(n15148) );
  XNOR2_X1 U18446 ( .A(n15149), .B(n15148), .ZN(n16344) );
  NAND2_X1 U18447 ( .A1(n15151), .A2(n15150), .ZN(n15157) );
  INV_X1 U18448 ( .A(n15152), .ZN(n15153) );
  NAND2_X1 U18449 ( .A1(n15154), .A2(n15153), .ZN(n15155) );
  AND2_X1 U18450 ( .A1(n16445), .A2(n15155), .ZN(n15156) );
  NAND2_X1 U18451 ( .A1(n15157), .A2(n15156), .ZN(n16433) );
  OAI22_X1 U18452 ( .A1(n15158), .A2(n16466), .B1(n21004), .B2(n20347), .ZN(
        n15159) );
  AOI21_X1 U18453 ( .B1(n16433), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15159), .ZN(n15161) );
  NAND2_X1 U18454 ( .A1(n16418), .A2(n16417), .ZN(n15160) );
  OAI211_X1 U18455 ( .C1(n16344), .C2(n20431), .A(n15161), .B(n15160), .ZN(
        P1_U3017) );
  NAND2_X1 U18456 ( .A1(n20168), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n15163) );
  NOR3_X1 U18457 ( .A1(n12298), .A2(n16039), .A3(n20168), .ZN(n15162) );
  AOI21_X1 U18458 ( .B1(n16726), .B2(n15163), .A(n15162), .ZN(n15165) );
  NAND2_X1 U18459 ( .A1(n20154), .A2(n19955), .ZN(n16026) );
  INV_X1 U18460 ( .A(n16026), .ZN(n16733) );
  OAI22_X1 U18461 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16733), .B1(n20175), 
        .B2(n19955), .ZN(n15164) );
  OAI21_X1 U18462 ( .B1(n15165), .B2(n16735), .A(n15164), .ZN(n15168) );
  AOI21_X1 U18463 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16729), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15166) );
  AOI211_X1 U18464 ( .C1(n19572), .C2(n20155), .A(n15166), .B(n19282), .ZN(
        n15167) );
  MUX2_X1 U18465 ( .A(n15168), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15167), 
        .Z(P2_U3610) );
  NAND2_X1 U18466 ( .A1(n15187), .A2(n15169), .ZN(n15170) );
  NAND2_X1 U18467 ( .A1(n15191), .A2(n15170), .ZN(n16544) );
  OR2_X1 U18468 ( .A1(n9766), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15171) );
  NAND2_X1 U18469 ( .A1(n15189), .A2(n15171), .ZN(n16568) );
  OAI21_X1 U18470 ( .B1(n15185), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15186), .ZN(n16225) );
  OAI21_X1 U18471 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15183), .A(
        n15172), .ZN(n15511) );
  NOR2_X1 U18472 ( .A1(n15173), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15174) );
  OR2_X1 U18473 ( .A1(n15177), .A2(n15174), .ZN(n15566) );
  INV_X1 U18474 ( .A(n15566), .ZN(n19354) );
  NAND2_X1 U18475 ( .A1(n15175), .A2(n15578), .ZN(n19348) );
  NOR2_X1 U18476 ( .A1(n19354), .A2(n19348), .ZN(n15237) );
  OR2_X1 U18477 ( .A1(n15177), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15178) );
  NAND2_X1 U18478 ( .A1(n15176), .A2(n15178), .ZN(n15554) );
  NAND2_X1 U18479 ( .A1(n15237), .A2(n15554), .ZN(n19339) );
  NAND2_X1 U18480 ( .A1(n15176), .A2(n19335), .ZN(n15179) );
  AND2_X1 U18481 ( .A1(n15181), .A2(n15179), .ZN(n15543) );
  NAND2_X1 U18482 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  NAND2_X1 U18483 ( .A1(n15184), .A2(n15182), .ZN(n15536) );
  NAND2_X1 U18484 ( .A1(n9647), .A2(n15219), .ZN(n19330) );
  AOI21_X1 U18485 ( .B1(n19322), .B2(n15184), .A(n15183), .ZN(n15526) );
  INV_X1 U18486 ( .A(n15526), .ZN(n19331) );
  NAND2_X1 U18487 ( .A1(n9647), .A2(n19329), .ZN(n15204) );
  NAND2_X1 U18488 ( .A1(n15511), .A2(n15204), .ZN(n15203) );
  NAND2_X1 U18489 ( .A1(n15203), .A2(n9647), .ZN(n19315) );
  AOI21_X1 U18490 ( .B1(n15172), .B2(n12791), .A(n15185), .ZN(n15503) );
  INV_X1 U18491 ( .A(n15503), .ZN(n19316) );
  NAND2_X1 U18492 ( .A1(n9647), .A2(n19314), .ZN(n16224) );
  NAND2_X1 U18493 ( .A1(n16225), .A2(n16224), .ZN(n16223) );
  NAND2_X1 U18494 ( .A1(n16223), .A2(n9647), .ZN(n16581) );
  AOI21_X1 U18495 ( .B1(n15467), .B2(n15186), .A(n9766), .ZN(n15470) );
  INV_X1 U18496 ( .A(n15470), .ZN(n16582) );
  NAND2_X1 U18497 ( .A1(n9647), .A2(n16580), .ZN(n16567) );
  NAND2_X1 U18498 ( .A1(n16568), .A2(n16567), .ZN(n16566) );
  NAND2_X1 U18499 ( .A1(n16566), .A2(n9647), .ZN(n16555) );
  INV_X1 U18500 ( .A(n15187), .ZN(n15188) );
  AOI21_X1 U18501 ( .B1(n15451), .B2(n15189), .A(n15188), .ZN(n15454) );
  INV_X1 U18502 ( .A(n15454), .ZN(n16556) );
  NAND2_X1 U18503 ( .A1(n9647), .A2(n16554), .ZN(n16543) );
  NAND2_X1 U18504 ( .A1(n16544), .A2(n16543), .ZN(n16542) );
  NAND2_X1 U18505 ( .A1(n16542), .A2(n9647), .ZN(n16532) );
  AOI21_X1 U18506 ( .B1(n15431), .B2(n15191), .A(n15190), .ZN(n15435) );
  INV_X1 U18507 ( .A(n15435), .ZN(n16533) );
  NAND2_X1 U18508 ( .A1(n9647), .A2(n16531), .ZN(n15193) );
  NAND2_X1 U18509 ( .A1(n15192), .A2(n15193), .ZN(n16492) );
  OAI211_X1 U18510 ( .C1(n15193), .C2(n15192), .A(n19420), .B(n16492), .ZN(
        n15201) );
  AOI22_X1 U18511 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19459), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19444), .ZN(n15194) );
  INV_X1 U18512 ( .A(n15194), .ZN(n15196) );
  NOR2_X1 U18513 ( .A1(n19429), .A2(n14413), .ZN(n15195) );
  NOR2_X1 U18514 ( .A1(n15196), .A2(n15195), .ZN(n15197) );
  OAI21_X1 U18515 ( .B1(n15334), .B2(n19442), .A(n15197), .ZN(n15198) );
  AOI21_X1 U18516 ( .B1(n15199), .B2(n19448), .A(n15198), .ZN(n15200) );
  OAI211_X1 U18517 ( .C1(n15256), .C2(n19453), .A(n15201), .B(n15200), .ZN(
        P2_U2827) );
  INV_X1 U18518 ( .A(n15202), .ZN(n15217) );
  OAI211_X1 U18519 ( .C1(n15511), .C2(n15204), .A(n19420), .B(n15203), .ZN(
        n15216) );
  OR2_X1 U18520 ( .A1(n15309), .A2(n15206), .ZN(n15207) );
  NAND2_X1 U18521 ( .A1(n15205), .A2(n15207), .ZN(n16596) );
  INV_X1 U18522 ( .A(n16596), .ZN(n15214) );
  OAI22_X1 U18523 ( .A1(n19429), .A2(n15208), .B1(n15510), .B2(n19425), .ZN(
        n15213) );
  OR2_X1 U18524 ( .A1(n15387), .A2(n15209), .ZN(n15210) );
  AND2_X1 U18525 ( .A1(n15380), .A2(n15210), .ZN(n15751) );
  INV_X1 U18526 ( .A(n15751), .ZN(n16611) );
  INV_X1 U18527 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15211) );
  OAI22_X1 U18528 ( .A1(n16611), .A2(n19442), .B1(n19390), .B2(n15211), .ZN(
        n15212) );
  AOI211_X1 U18529 ( .C1(n15214), .C2(n19437), .A(n15213), .B(n15212), .ZN(
        n15215) );
  OAI211_X1 U18530 ( .C1(n15217), .C2(n19427), .A(n15216), .B(n15215), .ZN(
        P2_U2835) );
  INV_X1 U18531 ( .A(n15218), .ZN(n15231) );
  OAI211_X1 U18532 ( .C1(n15220), .C2(n15536), .A(n19420), .B(n15219), .ZN(
        n15230) );
  NAND2_X1 U18533 ( .A1(n15222), .A2(n15221), .ZN(n15223) );
  AND2_X1 U18534 ( .A1(n9708), .A2(n15223), .ZN(n16618) );
  AOI22_X1 U18535 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19459), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19443), .ZN(n15224) );
  OAI211_X1 U18536 ( .C1(n19425), .C2(n15535), .A(n15224), .B(n19424), .ZN(
        n15228) );
  NAND2_X1 U18537 ( .A1(n15316), .A2(n15225), .ZN(n15226) );
  NAND2_X1 U18538 ( .A1(n15311), .A2(n15226), .ZN(n16602) );
  NOR2_X1 U18539 ( .A1(n16602), .A2(n19453), .ZN(n15227) );
  AOI211_X1 U18540 ( .C1(n19450), .C2(n16618), .A(n15228), .B(n15227), .ZN(
        n15229) );
  OAI211_X1 U18541 ( .C1(n19427), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        P2_U2837) );
  OR2_X1 U18542 ( .A1(n14017), .A2(n15232), .ZN(n15233) );
  NAND2_X1 U18543 ( .A1(n15317), .A2(n15233), .ZN(n19470) );
  INV_X1 U18544 ( .A(n19470), .ZN(n15558) );
  NOR2_X1 U18545 ( .A1(n19425), .A2(n15552), .ZN(n15243) );
  AND2_X1 U18546 ( .A1(n15810), .A2(n15234), .ZN(n15235) );
  NOR2_X1 U18547 ( .A1(n15236), .A2(n15235), .ZN(n19498) );
  NAND2_X1 U18548 ( .A1(n19498), .A2(n19450), .ZN(n15241) );
  AOI22_X1 U18549 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19459), .ZN(n15240) );
  OR2_X1 U18550 ( .A1(n19416), .A2(n15237), .ZN(n19347) );
  XOR2_X1 U18551 ( .A(n19347), .B(n15554), .Z(n15238) );
  NAND2_X1 U18552 ( .A1(n19420), .A2(n15238), .ZN(n15239) );
  NAND4_X1 U18553 ( .A1(n15241), .A2(n15240), .A3(n19424), .A4(n15239), .ZN(
        n15242) );
  AOI211_X1 U18554 ( .C1(n15558), .C2(n19437), .A(n15243), .B(n15242), .ZN(
        n15244) );
  OAI21_X1 U18555 ( .B1(n15245), .B2(n19427), .A(n15244), .ZN(P2_U2839) );
  XNOR2_X1 U18556 ( .A(n9706), .B(n15246), .ZN(n16517) );
  OR2_X1 U18557 ( .A1(n15248), .A2(n15247), .ZN(n15326) );
  NAND3_X1 U18558 ( .A1(n15326), .A2(n15249), .A3(n19487), .ZN(n15251) );
  NAND2_X1 U18559 ( .A1(n19484), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15250) );
  OAI211_X1 U18560 ( .C1(n16517), .C2(n19484), .A(n15251), .B(n15250), .ZN(
        P2_U2858) );
  NAND2_X1 U18561 ( .A1(n15253), .A2(n15252), .ZN(n15255) );
  XNOR2_X1 U18562 ( .A(n15255), .B(n15254), .ZN(n15338) );
  NOR2_X1 U18563 ( .A1(n15256), .A2(n19484), .ZN(n15257) );
  AOI21_X1 U18564 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19484), .A(n15257), .ZN(
        n15258) );
  OAI21_X1 U18565 ( .B1(n15338), .B2(n19481), .A(n15258), .ZN(P2_U2859) );
  OAI21_X1 U18566 ( .B1(n15261), .B2(n15260), .A(n15259), .ZN(n15345) );
  NOR2_X1 U18567 ( .A1(n15432), .A2(n19484), .ZN(n15262) );
  AOI21_X1 U18568 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19484), .A(n15262), .ZN(
        n15263) );
  OAI21_X1 U18569 ( .B1(n15345), .B2(n19481), .A(n15263), .ZN(P2_U2860) );
  OAI21_X1 U18570 ( .B1(n15266), .B2(n15265), .A(n15264), .ZN(n15352) );
  NOR2_X1 U18571 ( .A1(n15276), .A2(n15267), .ZN(n15268) );
  NOR2_X1 U18572 ( .A1(n16540), .A2(n19484), .ZN(n15270) );
  AOI21_X1 U18573 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19484), .A(n15270), .ZN(
        n15271) );
  OAI21_X1 U18574 ( .B1(n15352), .B2(n19481), .A(n15271), .ZN(P2_U2861) );
  OAI21_X1 U18575 ( .B1(n15274), .B2(n15273), .A(n15272), .ZN(n15361) );
  AND2_X1 U18576 ( .A1(n15285), .A2(n15275), .ZN(n15277) );
  OR2_X1 U18577 ( .A1(n15277), .A2(n15276), .ZN(n16550) );
  MUX2_X1 U18578 ( .A(n16550), .B(n15278), .S(n19484), .Z(n15279) );
  OAI21_X1 U18579 ( .B1(n15361), .B2(n19481), .A(n15279), .ZN(P2_U2862) );
  AOI21_X1 U18580 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15283) );
  XOR2_X1 U18581 ( .A(n15284), .B(n15283), .Z(n15370) );
  INV_X1 U18582 ( .A(n15285), .ZN(n15286) );
  AOI21_X1 U18583 ( .B1(n15287), .B2(n15293), .A(n15286), .ZN(n16565) );
  NOR2_X1 U18584 ( .A1(n19490), .A2(n15288), .ZN(n15289) );
  AOI21_X1 U18585 ( .B1(n16565), .B2(n19490), .A(n15289), .ZN(n15290) );
  OAI21_X1 U18586 ( .B1(n15370), .B2(n19481), .A(n15290), .ZN(P2_U2863) );
  OR2_X1 U18587 ( .A1(n15480), .A2(n15291), .ZN(n15292) );
  NAND2_X1 U18588 ( .A1(n15293), .A2(n15292), .ZN(n15709) );
  AOI21_X1 U18589 ( .B1(n15296), .B2(n15295), .A(n15294), .ZN(n15377) );
  NAND2_X1 U18590 ( .A1(n15377), .A2(n19487), .ZN(n15298) );
  NAND2_X1 U18591 ( .A1(n19484), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15297) );
  OAI211_X1 U18592 ( .C1(n15709), .C2(n19484), .A(n15298), .B(n15297), .ZN(
        P2_U2864) );
  OAI21_X1 U18593 ( .B1(n15299), .B2(n15301), .A(n15300), .ZN(n15385) );
  NAND2_X1 U18594 ( .A1(n15205), .A2(n15302), .ZN(n15303) );
  NAND2_X1 U18595 ( .A1(n15479), .A2(n15303), .ZN(n15736) );
  NOR2_X1 U18596 ( .A1(n15736), .A2(n19484), .ZN(n15304) );
  AOI21_X1 U18597 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19484), .A(n15304), .ZN(
        n15305) );
  OAI21_X1 U18598 ( .B1(n15385), .B2(n19481), .A(n15305), .ZN(P2_U2866) );
  AND2_X1 U18599 ( .A1(n15307), .A2(n15306), .ZN(n16598) );
  OAI21_X1 U18600 ( .B1(n16598), .B2(n15308), .A(n16592), .ZN(n15395) );
  INV_X1 U18601 ( .A(n15309), .ZN(n15313) );
  NAND2_X1 U18602 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  NAND2_X1 U18603 ( .A1(n15313), .A2(n15312), .ZN(n19327) );
  NOR2_X1 U18604 ( .A1(n19327), .A2(n19484), .ZN(n15314) );
  AOI21_X1 U18605 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19484), .A(n15314), .ZN(
        n15315) );
  OAI21_X1 U18606 ( .B1(n15395), .B2(n19481), .A(n15315), .ZN(P2_U2868) );
  AOI21_X1 U18607 ( .B1(n15318), .B2(n15317), .A(n10132), .ZN(n19342) );
  INV_X1 U18608 ( .A(n19342), .ZN(n15796) );
  NOR2_X1 U18609 ( .A1(n15796), .A2(n19484), .ZN(n15319) );
  AOI21_X1 U18610 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19484), .A(n15319), .ZN(
        n15320) );
  OAI21_X1 U18611 ( .B1(n15321), .B2(n19481), .A(n15320), .ZN(P2_U2870) );
  NAND2_X1 U18612 ( .A1(n15323), .A2(n15322), .ZN(n15324) );
  NAND3_X1 U18613 ( .A1(n15326), .A2(n15249), .A3(n16619), .ZN(n15331) );
  OAI22_X1 U18614 ( .A1(n15390), .A2(n19510), .B1(n19537), .B2(n15327), .ZN(
        n15329) );
  INV_X1 U18615 ( .A(n19496), .ZN(n15366) );
  NOR2_X1 U18616 ( .A1(n15366), .A2(n16812), .ZN(n15328) );
  AOI211_X1 U18617 ( .C1(n19497), .C2(BUF2_REG_29__SCAN_IN), .A(n15329), .B(
        n15328), .ZN(n15330) );
  OAI211_X1 U18618 ( .C1(n19538), .C2(n16516), .A(n15331), .B(n15330), .ZN(
        P2_U2890) );
  INV_X1 U18619 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U18620 ( .A1(n19495), .A2(n19512), .B1(n19546), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15332) );
  OAI21_X1 U18621 ( .B1(n15356), .B2(n15333), .A(n15332), .ZN(n15336) );
  NOR2_X1 U18622 ( .A1(n15334), .A2(n19538), .ZN(n15335) );
  AOI211_X1 U18623 ( .C1(n19496), .C2(BUF1_REG_28__SCAN_IN), .A(n15336), .B(
        n15335), .ZN(n15337) );
  OAI21_X1 U18624 ( .B1(n15338), .B2(n19551), .A(n15337), .ZN(P2_U2891) );
  INV_X1 U18625 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U18626 ( .A1(n19495), .A2(n15339), .B1(n19546), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15340) );
  OAI21_X1 U18627 ( .B1(n15356), .B2(n15341), .A(n15340), .ZN(n15343) );
  NOR2_X1 U18628 ( .A1(n16536), .A2(n19538), .ZN(n15342) );
  AOI211_X1 U18629 ( .C1(n19496), .C2(BUF1_REG_27__SCAN_IN), .A(n15343), .B(
        n15342), .ZN(n15344) );
  OAI21_X1 U18630 ( .B1(n15345), .B2(n19551), .A(n15344), .ZN(P2_U2892) );
  AOI22_X1 U18631 ( .A1(n19495), .A2(n19517), .B1(n19546), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15346) );
  OAI21_X1 U18632 ( .B1(n15356), .B2(n17653), .A(n15346), .ZN(n15350) );
  NAND2_X1 U18633 ( .A1(n9722), .A2(n15347), .ZN(n15348) );
  NAND2_X1 U18634 ( .A1(n9707), .A2(n15348), .ZN(n16539) );
  NOR2_X1 U18635 ( .A1(n16539), .A2(n19538), .ZN(n15349) );
  AOI211_X1 U18636 ( .C1(n19496), .C2(BUF1_REG_26__SCAN_IN), .A(n15350), .B(
        n15349), .ZN(n15351) );
  OAI21_X1 U18637 ( .B1(n15352), .B2(n19551), .A(n15351), .ZN(P2_U2893) );
  INV_X1 U18638 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U18639 ( .A1(n19495), .A2(n15353), .B1(n19546), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15354) );
  OAI21_X1 U18640 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15359) );
  OAI21_X1 U18641 ( .B1(n15365), .B2(n15357), .A(n9722), .ZN(n16551) );
  NOR2_X1 U18642 ( .A1(n16551), .A2(n19538), .ZN(n15358) );
  AOI211_X1 U18643 ( .C1(n19496), .C2(BUF1_REG_25__SCAN_IN), .A(n15359), .B(
        n15358), .ZN(n15360) );
  OAI21_X1 U18644 ( .B1(n15361), .B2(n19551), .A(n15360), .ZN(P2_U2894) );
  INV_X1 U18645 ( .A(n19523), .ZN(n15362) );
  OAI22_X1 U18646 ( .A1(n15390), .A2(n15362), .B1(n19537), .B2(n13043), .ZN(
        n15368) );
  NOR2_X1 U18647 ( .A1(n15372), .A2(n15363), .ZN(n15364) );
  OR2_X1 U18648 ( .A1(n15365), .A2(n15364), .ZN(n16563) );
  OAI22_X1 U18649 ( .A1(n16563), .A2(n19538), .B1(n15366), .B2(n16822), .ZN(
        n15367) );
  AOI211_X1 U18650 ( .C1(n19497), .C2(BUF2_REG_24__SCAN_IN), .A(n15368), .B(
        n15367), .ZN(n15369) );
  OAI21_X1 U18651 ( .B1(n15370), .B2(n19551), .A(n15369), .ZN(P2_U2895) );
  AND2_X1 U18652 ( .A1(n15724), .A2(n15371), .ZN(n15373) );
  OR2_X1 U18653 ( .A1(n15373), .A2(n15372), .ZN(n16585) );
  AOI22_X1 U18654 ( .A1(n19495), .A2(n19661), .B1(n19546), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U18655 ( .A1(n19496), .A2(BUF1_REG_23__SCAN_IN), .B1(n19497), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15374) );
  OAI211_X1 U18656 ( .C1(n16585), .C2(n19538), .A(n15375), .B(n15374), .ZN(
        n15376) );
  AOI21_X1 U18657 ( .B1(n15377), .B2(n16619), .A(n15376), .ZN(n15378) );
  INV_X1 U18658 ( .A(n15378), .ZN(P2_U2896) );
  XNOR2_X1 U18659 ( .A(n15380), .B(n15379), .ZN(n15738) );
  INV_X1 U18660 ( .A(n15738), .ZN(n19312) );
  OAI22_X1 U18661 ( .A1(n15390), .A2(n19651), .B1(n19537), .B2(n15381), .ZN(
        n15382) );
  AOI21_X1 U18662 ( .B1(n19312), .B2(n19547), .A(n15382), .ZN(n15384) );
  AOI22_X1 U18663 ( .A1(n19496), .A2(BUF1_REG_21__SCAN_IN), .B1(n19497), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15383) );
  OAI211_X1 U18664 ( .C1(n15385), .C2(n19551), .A(n15384), .B(n15383), .ZN(
        P2_U2898) );
  AND2_X1 U18665 ( .A1(n9708), .A2(n15386), .ZN(n15388) );
  OR2_X1 U18666 ( .A1(n15388), .A2(n15387), .ZN(n19326) );
  INV_X1 U18667 ( .A(n19326), .ZN(n15392) );
  OAI22_X1 U18668 ( .A1(n15390), .A2(n19643), .B1(n19537), .B2(n15389), .ZN(
        n15391) );
  AOI21_X1 U18669 ( .B1(n19547), .B2(n15392), .A(n15391), .ZN(n15394) );
  AOI22_X1 U18670 ( .A1(n19496), .A2(BUF1_REG_19__SCAN_IN), .B1(n19497), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15393) );
  OAI211_X1 U18671 ( .C1(n15395), .C2(n19551), .A(n15394), .B(n15393), .ZN(
        P2_U2900) );
  INV_X1 U18672 ( .A(n19522), .ZN(n19555) );
  AOI21_X1 U18673 ( .B1(n16002), .B2(n15397), .A(n15396), .ZN(n19542) );
  XNOR2_X1 U18674 ( .A(n20248), .B(n20240), .ZN(n19541) );
  NOR2_X1 U18675 ( .A1(n19542), .A2(n19541), .ZN(n19540) );
  AOI21_X1 U18676 ( .B1(n20248), .B2(n20240), .A(n19540), .ZN(n15401) );
  NAND2_X1 U18677 ( .A1(n15398), .A2(n15399), .ZN(n15400) );
  INV_X1 U18678 ( .A(n15398), .ZN(n19488) );
  INV_X1 U18679 ( .A(n15399), .ZN(n15402) );
  NAND2_X1 U18680 ( .A1(n19488), .A2(n15402), .ZN(n19532) );
  OAI211_X1 U18681 ( .C1(n15401), .C2(n15400), .A(n16619), .B(n19532), .ZN(
        n15404) );
  AOI22_X1 U18682 ( .A1(n19547), .A2(n15402), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19546), .ZN(n15403) );
  OAI211_X1 U18683 ( .C1(n19555), .C2(n19647), .A(n15404), .B(n15403), .ZN(
        P2_U2915) );
  NAND2_X1 U18684 ( .A1(n15405), .A2(n15415), .ZN(n15410) );
  INV_X1 U18685 ( .A(n15406), .ZN(n15407) );
  NOR2_X1 U18686 ( .A1(n15408), .A2(n15407), .ZN(n15409) );
  XNOR2_X1 U18687 ( .A(n15410), .B(n15409), .ZN(n15657) );
  XNOR2_X1 U18688 ( .A(n15420), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15655) );
  NOR2_X1 U18689 ( .A1(n15644), .A2(n15640), .ZN(n15413) );
  XNOR2_X1 U18690 ( .A(n15423), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16510) );
  NAND2_X1 U18691 ( .A1(n19592), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15646) );
  NAND2_X1 U18692 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15411) );
  OAI211_X1 U18693 ( .C1(n19603), .C2(n16510), .A(n15646), .B(n15411), .ZN(
        n15412) );
  OAI21_X1 U18694 ( .B1(n15657), .B2(n16665), .A(n15414), .ZN(P2_U2984) );
  NAND2_X1 U18695 ( .A1(n15416), .A2(n15415), .ZN(n15418) );
  XOR2_X1 U18696 ( .A(n15418), .B(n15417), .Z(n15673) );
  INV_X1 U18697 ( .A(n15419), .ZN(n15422) );
  INV_X1 U18698 ( .A(n15420), .ZN(n15421) );
  AOI21_X1 U18699 ( .B1(n15663), .B2(n15422), .A(n15421), .ZN(n15671) );
  INV_X1 U18700 ( .A(n14445), .ZN(n15424) );
  AOI21_X1 U18701 ( .B1(n10016), .B2(n15424), .A(n15423), .ZN(n16493) );
  NAND2_X1 U18702 ( .A1(n19592), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15658) );
  OAI21_X1 U18703 ( .B1(n16670), .B2(n10016), .A(n15658), .ZN(n15425) );
  AOI21_X1 U18704 ( .B1(n16661), .B2(n16493), .A(n15425), .ZN(n15426) );
  OAI21_X1 U18705 ( .B1(n16517), .B2(n15640), .A(n15426), .ZN(n15427) );
  AOI21_X1 U18706 ( .B1(n15671), .B2(n19595), .A(n15427), .ZN(n15428) );
  OAI21_X1 U18707 ( .B1(n15673), .B2(n16665), .A(n15428), .ZN(P2_U2985) );
  NAND2_X1 U18708 ( .A1(n15429), .A2(n19598), .ZN(n15437) );
  OAI21_X1 U18709 ( .B1(n16670), .B2(n15431), .A(n15430), .ZN(n15434) );
  NOR2_X1 U18710 ( .A1(n15432), .A2(n15640), .ZN(n15433) );
  AOI211_X1 U18711 ( .C1(n16661), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        n15436) );
  OAI211_X1 U18712 ( .C1(n16664), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        P2_U2987) );
  OAI21_X1 U18713 ( .B1(n15450), .B2(n15447), .A(n15446), .ZN(n15439) );
  XOR2_X1 U18714 ( .A(n15440), .B(n15439), .Z(n15684) );
  INV_X1 U18715 ( .A(n15462), .ZN(n15441) );
  NAND2_X1 U18716 ( .A1(n15441), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15693) );
  AOI21_X1 U18717 ( .B1(n15677), .B2(n15693), .A(n9717), .ZN(n15681) );
  NOR2_X1 U18718 ( .A1(n16540), .A2(n15640), .ZN(n15444) );
  NAND2_X1 U18719 ( .A1(n19592), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15674) );
  NAND2_X1 U18720 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15442) );
  OAI211_X1 U18721 ( .C1(n19603), .C2(n16544), .A(n15674), .B(n15442), .ZN(
        n15443) );
  AOI211_X1 U18722 ( .C1(n15681), .C2(n19595), .A(n15444), .B(n15443), .ZN(
        n15445) );
  OAI21_X1 U18723 ( .B1(n15684), .B2(n16665), .A(n15445), .ZN(P2_U2988) );
  INV_X1 U18724 ( .A(n15446), .ZN(n15448) );
  NOR2_X1 U18725 ( .A1(n15448), .A2(n15447), .ZN(n15449) );
  XNOR2_X1 U18726 ( .A(n15450), .B(n15449), .ZN(n15696) );
  NAND2_X1 U18727 ( .A1(n19592), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15685) );
  OAI21_X1 U18728 ( .B1(n16670), .B2(n15451), .A(n15685), .ZN(n15453) );
  NOR2_X1 U18729 ( .A1(n16550), .A2(n15640), .ZN(n15452) );
  AOI211_X1 U18730 ( .C1(n16661), .C2(n15454), .A(n15453), .B(n15452), .ZN(
        n15456) );
  NAND2_X1 U18731 ( .A1(n15462), .A2(n15690), .ZN(n15692) );
  NAND3_X1 U18732 ( .A1(n15693), .A2(n19595), .A3(n15692), .ZN(n15455) );
  OAI211_X1 U18733 ( .C1(n15696), .C2(n16665), .A(n15456), .B(n15455), .ZN(
        P2_U2989) );
  XNOR2_X1 U18734 ( .A(n15457), .B(n15698), .ZN(n15458) );
  XNOR2_X1 U18735 ( .A(n15459), .B(n15458), .ZN(n15704) );
  NAND2_X1 U18736 ( .A1(n19592), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15701) );
  NAND2_X1 U18737 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15460) );
  OAI211_X1 U18738 ( .C1(n19603), .C2(n16568), .A(n15701), .B(n15460), .ZN(
        n15463) );
  INV_X1 U18739 ( .A(n15461), .ZN(n15788) );
  INV_X1 U18740 ( .A(n15699), .ZN(n15714) );
  NOR2_X1 U18741 ( .A1(n15487), .A2(n15714), .ZN(n15466) );
  XNOR2_X1 U18742 ( .A(n15465), .B(n15464), .ZN(n15721) );
  INV_X1 U18743 ( .A(n15487), .ZN(n15474) );
  NAND2_X1 U18744 ( .A1(n15474), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15473) );
  AOI21_X1 U18745 ( .B1(n15713), .B2(n15473), .A(n15466), .ZN(n15708) );
  NAND2_X1 U18746 ( .A1(n15708), .A2(n19595), .ZN(n15472) );
  NAND2_X1 U18747 ( .A1(n19592), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15716) );
  OAI21_X1 U18748 ( .B1(n16670), .B2(n15467), .A(n15716), .ZN(n15469) );
  NOR2_X1 U18749 ( .A1(n15709), .A2(n15640), .ZN(n15468) );
  AOI211_X1 U18750 ( .C1(n16661), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15471) );
  OAI211_X1 U18751 ( .C1(n15721), .C2(n16665), .A(n15472), .B(n15471), .ZN(
        P2_U2991) );
  OAI21_X1 U18752 ( .B1(n15474), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15473), .ZN(n15734) );
  NAND2_X1 U18753 ( .A1(n9744), .A2(n15476), .ZN(n15477) );
  XNOR2_X1 U18754 ( .A(n15475), .B(n15477), .ZN(n15732) );
  AND2_X1 U18755 ( .A1(n15479), .A2(n15478), .ZN(n15481) );
  OR2_X1 U18756 ( .A1(n15481), .A2(n15480), .ZN(n16590) );
  NOR2_X1 U18757 ( .A1(n19424), .A2(n15482), .ZN(n15726) );
  NOR2_X1 U18758 ( .A1(n19603), .A2(n16225), .ZN(n15483) );
  AOI211_X1 U18759 ( .C1(n19593), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15726), .B(n15483), .ZN(n15484) );
  OAI21_X1 U18760 ( .B1(n16590), .B2(n15640), .A(n15484), .ZN(n15485) );
  AOI21_X1 U18761 ( .B1(n15732), .B2(n19598), .A(n15485), .ZN(n15486) );
  OAI21_X1 U18762 ( .B1(n15734), .B2(n16664), .A(n15486), .ZN(P2_U2992) );
  OAI21_X1 U18763 ( .B1(n9716), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15487), .ZN(n15746) );
  NAND3_X1 U18764 ( .A1(n15560), .A2(n15562), .A3(n15572), .ZN(n15489) );
  NAND2_X1 U18765 ( .A1(n15489), .A2(n15488), .ZN(n15551) );
  INV_X1 U18766 ( .A(n15490), .ZN(n15491) );
  AOI21_X1 U18767 ( .B1(n15551), .B2(n15550), .A(n15491), .ZN(n15542) );
  NAND2_X1 U18768 ( .A1(n15492), .A2(n15493), .ZN(n15541) );
  INV_X1 U18769 ( .A(n15494), .ZN(n15519) );
  INV_X1 U18770 ( .A(n15530), .ZN(n15517) );
  INV_X1 U18771 ( .A(n15506), .ZN(n15496) );
  OAI21_X1 U18772 ( .B1(n15509), .B2(n15496), .A(n15507), .ZN(n15500) );
  NAND2_X1 U18773 ( .A1(n15498), .A2(n15497), .ZN(n15499) );
  XNOR2_X1 U18774 ( .A(n15500), .B(n15499), .ZN(n15735) );
  NAND2_X1 U18775 ( .A1(n15735), .A2(n19598), .ZN(n15505) );
  NAND2_X1 U18776 ( .A1(n19592), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15737) );
  OAI21_X1 U18777 ( .B1(n16670), .B2(n12791), .A(n15737), .ZN(n15502) );
  NOR2_X1 U18778 ( .A1(n15736), .A2(n15640), .ZN(n15501) );
  AOI211_X1 U18779 ( .C1(n16661), .C2(n15503), .A(n15502), .B(n15501), .ZN(
        n15504) );
  OAI211_X1 U18780 ( .C1(n16664), .C2(n15746), .A(n15505), .B(n15504), .ZN(
        P2_U2993) );
  NAND2_X1 U18781 ( .A1(n15507), .A2(n15506), .ZN(n15508) );
  XNOR2_X1 U18782 ( .A(n15509), .B(n15508), .ZN(n15758) );
  AOI21_X1 U18783 ( .B1(n15748), .B2(n15522), .A(n9716), .ZN(n15756) );
  NOR2_X1 U18784 ( .A1(n19424), .A2(n15510), .ZN(n15750) );
  NOR2_X1 U18785 ( .A1(n19603), .A2(n15511), .ZN(n15512) );
  AOI211_X1 U18786 ( .C1(n19593), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15750), .B(n15512), .ZN(n15513) );
  OAI21_X1 U18787 ( .B1(n16596), .B2(n15640), .A(n15513), .ZN(n15514) );
  AOI21_X1 U18788 ( .B1(n15756), .B2(n19595), .A(n15514), .ZN(n15515) );
  OAI21_X1 U18789 ( .B1(n15758), .B2(n16665), .A(n15515), .ZN(P2_U2994) );
  INV_X1 U18790 ( .A(n15516), .ZN(n15531) );
  AOI21_X1 U18791 ( .B1(n15533), .B2(n15517), .A(n15531), .ZN(n15521) );
  NAND2_X1 U18792 ( .A1(n15519), .A2(n15518), .ZN(n15520) );
  XNOR2_X1 U18793 ( .A(n15521), .B(n15520), .ZN(n15769) );
  INV_X1 U18794 ( .A(n15522), .ZN(n15524) );
  AOI21_X1 U18795 ( .B1(n15545), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U18796 ( .A1(n15524), .A2(n15523), .ZN(n15767) );
  NAND2_X1 U18797 ( .A1(n19592), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15759) );
  OAI21_X1 U18798 ( .B1(n16670), .B2(n19322), .A(n15759), .ZN(n15525) );
  AOI21_X1 U18799 ( .B1(n15526), .B2(n16661), .A(n15525), .ZN(n15527) );
  OAI21_X1 U18800 ( .B1(n19327), .B2(n15640), .A(n15527), .ZN(n15528) );
  AOI21_X1 U18801 ( .B1(n15767), .B2(n19595), .A(n15528), .ZN(n15529) );
  OAI21_X1 U18802 ( .B1(n15769), .B2(n16665), .A(n15529), .ZN(P2_U2995) );
  NOR2_X1 U18803 ( .A1(n15531), .A2(n15530), .ZN(n15532) );
  XNOR2_X1 U18804 ( .A(n15533), .B(n15532), .ZN(n15779) );
  XNOR2_X1 U18805 ( .A(n15545), .B(n15534), .ZN(n15777) );
  NOR2_X1 U18806 ( .A1(n19424), .A2(n15535), .ZN(n15772) );
  NOR2_X1 U18807 ( .A1(n15536), .A2(n19603), .ZN(n15537) );
  AOI211_X1 U18808 ( .C1(n19593), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15772), .B(n15537), .ZN(n15538) );
  OAI21_X1 U18809 ( .B1(n16602), .B2(n15640), .A(n15538), .ZN(n15539) );
  AOI21_X1 U18810 ( .B1(n15777), .B2(n19595), .A(n15539), .ZN(n15540) );
  OAI21_X1 U18811 ( .B1(n15779), .B2(n16665), .A(n15540), .ZN(P2_U2996) );
  XNOR2_X1 U18812 ( .A(n15542), .B(n15541), .ZN(n15798) );
  INV_X1 U18813 ( .A(n15543), .ZN(n19341) );
  NOR2_X1 U18814 ( .A1(n19424), .A2(n20206), .ZN(n15792) );
  AOI21_X1 U18815 ( .B1(n19593), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15792), .ZN(n15544) );
  OAI21_X1 U18816 ( .B1(n19341), .B2(n19603), .A(n15544), .ZN(n15548) );
  INV_X1 U18817 ( .A(n15781), .ZN(n15546) );
  AOI211_X1 U18818 ( .C1(n15790), .C2(n15546), .A(n16664), .B(n15545), .ZN(
        n15547) );
  OAI21_X1 U18819 ( .B1(n15798), .B2(n16665), .A(n15549), .ZN(P2_U2997) );
  XNOR2_X1 U18820 ( .A(n15551), .B(n15550), .ZN(n15808) );
  NOR2_X1 U18821 ( .A1(n19424), .A2(n15552), .ZN(n15802) );
  AOI21_X1 U18822 ( .B1(n19593), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15802), .ZN(n15553) );
  OAI21_X1 U18823 ( .B1(n19603), .B2(n15554), .A(n15553), .ZN(n15557) );
  AOI21_X1 U18824 ( .B1(n15787), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15555) );
  NOR3_X1 U18825 ( .A1(n15781), .A2(n15555), .A3(n16664), .ZN(n15556) );
  AOI211_X1 U18826 ( .C1(n19597), .C2(n15558), .A(n15557), .B(n15556), .ZN(
        n15559) );
  OAI21_X1 U18827 ( .B1(n15808), .B2(n16665), .A(n15559), .ZN(P2_U2998) );
  INV_X1 U18828 ( .A(n15560), .ZN(n15573) );
  NAND4_X1 U18829 ( .A1(n15573), .A2(n15572), .A3(n15571), .A4(n15584), .ZN(
        n15570) );
  NAND2_X1 U18830 ( .A1(n15570), .A2(n15572), .ZN(n15564) );
  NAND2_X1 U18831 ( .A1(n15562), .A2(n15561), .ZN(n15563) );
  XNOR2_X1 U18832 ( .A(n15564), .B(n15563), .ZN(n15822) );
  XNOR2_X1 U18833 ( .A(n15787), .B(n15784), .ZN(n15820) );
  NOR2_X1 U18834 ( .A1(n15809), .A2(n15640), .ZN(n15568) );
  NAND2_X1 U18835 ( .A1(n19592), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15813) );
  NAND2_X1 U18836 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15565) );
  OAI211_X1 U18837 ( .C1(n19603), .C2(n15566), .A(n15813), .B(n15565), .ZN(
        n15567) );
  AOI211_X1 U18838 ( .C1(n15820), .C2(n19595), .A(n15568), .B(n15567), .ZN(
        n15569) );
  OAI21_X1 U18839 ( .B1(n15822), .B2(n16665), .A(n15569), .ZN(P2_U2999) );
  INV_X1 U18840 ( .A(n15570), .ZN(n15575) );
  AOI22_X1 U18841 ( .A1(n15573), .A2(n15584), .B1(n15572), .B2(n15571), .ZN(
        n15574) );
  NOR2_X1 U18842 ( .A1(n15575), .A2(n15574), .ZN(n15838) );
  NOR2_X1 U18843 ( .A1(n19424), .A2(n15576), .ZN(n15829) );
  AOI21_X1 U18844 ( .B1(n19593), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15829), .ZN(n15577) );
  OAI21_X1 U18845 ( .B1(n19603), .B2(n15578), .A(n15577), .ZN(n15579) );
  AOI21_X1 U18846 ( .B1(n15580), .B2(n19597), .A(n15579), .ZN(n15582) );
  NAND2_X1 U18847 ( .A1(n15622), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15602) );
  INV_X1 U18848 ( .A(n15602), .ZN(n15623) );
  INV_X1 U18849 ( .A(n15826), .ZN(n15828) );
  NAND2_X1 U18850 ( .A1(n15623), .A2(n15828), .ZN(n15583) );
  AOI21_X1 U18851 ( .B1(n15583), .B2(n15827), .A(n15787), .ZN(n15835) );
  NAND2_X1 U18852 ( .A1(n15835), .A2(n19595), .ZN(n15581) );
  OAI211_X1 U18853 ( .C1(n15838), .C2(n16665), .A(n15582), .B(n15581), .ZN(
        P2_U3000) );
  NOR2_X1 U18854 ( .A1(n15602), .A2(n15858), .ZN(n15601) );
  OAI21_X1 U18855 ( .B1(n15601), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15583), .ZN(n15848) );
  INV_X1 U18856 ( .A(n15584), .ZN(n15585) );
  NOR2_X1 U18857 ( .A1(n15586), .A2(n15585), .ZN(n15587) );
  XNOR2_X1 U18858 ( .A(n15588), .B(n15587), .ZN(n15846) );
  NOR2_X1 U18859 ( .A1(n19424), .A2(n15589), .ZN(n15840) );
  NOR2_X1 U18860 ( .A1(n16670), .A2(n15590), .ZN(n15591) );
  AOI211_X1 U18861 ( .C1(n16661), .C2(n15592), .A(n15840), .B(n15591), .ZN(
        n15593) );
  OAI21_X1 U18862 ( .B1(n15594), .B2(n15640), .A(n15593), .ZN(n15595) );
  AOI21_X1 U18863 ( .B1(n15846), .B2(n19598), .A(n15595), .ZN(n15596) );
  OAI21_X1 U18864 ( .B1(n15848), .B2(n16664), .A(n15596), .ZN(P2_U3001) );
  NAND2_X1 U18865 ( .A1(n15598), .A2(n15597), .ZN(n15600) );
  XOR2_X1 U18866 ( .A(n15600), .B(n15599), .Z(n15862) );
  INV_X1 U18867 ( .A(n15601), .ZN(n15850) );
  NAND2_X1 U18868 ( .A1(n15602), .A2(n15858), .ZN(n15849) );
  NAND3_X1 U18869 ( .A1(n15850), .A2(n19595), .A3(n15849), .ZN(n15612) );
  OR2_X1 U18870 ( .A1(n15604), .A2(n15603), .ZN(n15605) );
  NAND2_X1 U18871 ( .A1(n15606), .A2(n15605), .ZN(n19475) );
  INV_X1 U18872 ( .A(n19475), .ZN(n15610) );
  NOR2_X1 U18873 ( .A1(n19424), .A2(n15607), .ZN(n15854) );
  AOI21_X1 U18874 ( .B1(n19593), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15854), .ZN(n15608) );
  OAI21_X1 U18875 ( .B1(n19603), .B2(n19359), .A(n15608), .ZN(n15609) );
  AOI21_X1 U18876 ( .B1(n15610), .B2(n19597), .A(n15609), .ZN(n15611) );
  OAI211_X1 U18877 ( .C1(n15862), .C2(n16665), .A(n15612), .B(n15611), .ZN(
        P2_U3002) );
  INV_X1 U18878 ( .A(n15613), .ZN(n15614) );
  INV_X1 U18879 ( .A(n15616), .ZN(n15915) );
  AOI211_X1 U18880 ( .C1(n15913), .C2(n15882), .A(n15881), .B(n15917), .ZN(
        n15621) );
  INV_X1 U18881 ( .A(n15617), .ZN(n15619) );
  NAND2_X1 U18882 ( .A1(n15619), .A2(n15618), .ZN(n15620) );
  XNOR2_X1 U18883 ( .A(n15621), .B(n15620), .ZN(n15880) );
  INV_X1 U18884 ( .A(n15622), .ZN(n15888) );
  AOI21_X1 U18885 ( .B1(n15875), .B2(n15888), .A(n15623), .ZN(n15878) );
  NAND2_X1 U18886 ( .A1(n19592), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n15870) );
  OAI21_X1 U18887 ( .B1(n16670), .B2(n15624), .A(n15870), .ZN(n15625) );
  AOI21_X1 U18888 ( .B1(n16661), .B2(n19373), .A(n15625), .ZN(n15626) );
  OAI21_X1 U18889 ( .B1(n15627), .B2(n15640), .A(n15626), .ZN(n15628) );
  AOI21_X1 U18890 ( .B1(n15878), .B2(n19595), .A(n15628), .ZN(n15629) );
  OAI21_X1 U18891 ( .B1(n15880), .B2(n16665), .A(n15629), .ZN(P2_U3003) );
  XNOR2_X1 U18892 ( .A(n15630), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15631) );
  XNOR2_X1 U18893 ( .A(n15632), .B(n15631), .ZN(n15935) );
  INV_X1 U18894 ( .A(n16641), .ZN(n15638) );
  NAND2_X1 U18895 ( .A1(n15633), .A2(n15634), .ZN(n15635) );
  OAI21_X1 U18896 ( .B1(n15636), .B2(n15638), .A(n15635), .ZN(n15637) );
  OAI21_X1 U18897 ( .B1(n16642), .B2(n15638), .A(n15637), .ZN(n15933) );
  OAI22_X1 U18898 ( .A1(n16670), .A2(n12692), .B1(n20194), .B2(n19424), .ZN(
        n15642) );
  INV_X1 U18899 ( .A(n19402), .ZN(n15639) );
  OAI22_X1 U18900 ( .A1(n15640), .A2(n19406), .B1(n19603), .B2(n15639), .ZN(
        n15641) );
  AOI211_X1 U18901 ( .C1(n15933), .C2(n19598), .A(n15642), .B(n15641), .ZN(
        n15643) );
  OAI21_X1 U18902 ( .B1(n15935), .B2(n16664), .A(n15643), .ZN(P2_U3007) );
  INV_X1 U18903 ( .A(n15644), .ZN(n15645) );
  OAI21_X1 U18904 ( .B1(n16506), .B2(n16677), .A(n15646), .ZN(n15651) );
  OAI21_X1 U18905 ( .B1(n15649), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10219), .ZN(n15650) );
  AOI21_X1 U18906 ( .B1(n15655), .B2(n19611), .A(n15654), .ZN(n15656) );
  OAI21_X1 U18907 ( .B1(n15657), .B2(n15974), .A(n15656), .ZN(P2_U3016) );
  OAI21_X1 U18908 ( .B1(n16516), .B2(n16677), .A(n15658), .ZN(n15666) );
  AOI21_X1 U18909 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15663), .A(
        n15662), .ZN(n15661) );
  AOI211_X1 U18910 ( .C1(n15663), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15664) );
  INV_X1 U18911 ( .A(n16517), .ZN(n15667) );
  AOI21_X1 U18912 ( .B1(n15671), .B2(n19611), .A(n15670), .ZN(n15672) );
  OAI21_X1 U18913 ( .B1(n15673), .B2(n15974), .A(n15672), .ZN(P2_U3017) );
  INV_X1 U18914 ( .A(n16540), .ZN(n15680) );
  OR2_X1 U18915 ( .A1(n15697), .A2(n15677), .ZN(n15675) );
  OAI211_X1 U18916 ( .C1(n16539), .C2(n16677), .A(n15675), .B(n15674), .ZN(
        n15679) );
  INV_X1 U18917 ( .A(n15691), .ZN(n15676) );
  AOI211_X1 U18918 ( .C1(n15677), .C2(n15690), .A(n9895), .B(n15676), .ZN(
        n15678) );
  AOI211_X1 U18919 ( .C1(n15680), .C2(n19613), .A(n15679), .B(n15678), .ZN(
        n15683) );
  NAND2_X1 U18920 ( .A1(n15681), .A2(n19611), .ZN(n15682) );
  OAI211_X1 U18921 ( .C1(n15684), .C2(n15974), .A(n15683), .B(n15682), .ZN(
        P2_U3020) );
  INV_X1 U18922 ( .A(n15697), .ZN(n15687) );
  OAI21_X1 U18923 ( .B1(n16551), .B2(n16677), .A(n15685), .ZN(n15686) );
  AOI21_X1 U18924 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15687), .A(
        n15686), .ZN(n15688) );
  OAI21_X1 U18925 ( .B1(n16550), .B2(n15927), .A(n15688), .ZN(n15689) );
  AOI21_X1 U18926 ( .B1(n15691), .B2(n15690), .A(n15689), .ZN(n15695) );
  NAND3_X1 U18927 ( .A1(n15693), .A2(n19611), .A3(n15692), .ZN(n15694) );
  OAI211_X1 U18928 ( .C1(n15696), .C2(n15974), .A(n15695), .B(n15694), .ZN(
        P2_U3021) );
  NOR2_X1 U18929 ( .A1(n15697), .A2(n15698), .ZN(n15703) );
  NOR2_X1 U18930 ( .A1(n15740), .A2(n15741), .ZN(n15727) );
  NAND3_X1 U18931 ( .A1(n15699), .A2(n15698), .A3(n15727), .ZN(n15700) );
  OAI211_X1 U18932 ( .C1(n16563), .C2(n16677), .A(n15701), .B(n15700), .ZN(
        n15702) );
  AOI211_X1 U18933 ( .C1(n16565), .C2(n19613), .A(n15703), .B(n15702), .ZN(
        n15706) );
  OR2_X1 U18934 ( .A1(n15704), .A2(n15974), .ZN(n15705) );
  OAI211_X1 U18935 ( .C1(n15707), .C2(n16684), .A(n15706), .B(n15705), .ZN(
        P2_U3022) );
  NAND2_X1 U18936 ( .A1(n15708), .A2(n19611), .ZN(n15720) );
  INV_X1 U18937 ( .A(n15709), .ZN(n16573) );
  OAI21_X1 U18938 ( .B1(n15780), .B2(n15710), .A(n15893), .ZN(n15764) );
  OAI21_X1 U18939 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15741), .A(
        n15764), .ZN(n15711) );
  AOI21_X1 U18940 ( .B1(n19617), .B2(n15712), .A(n15711), .ZN(n15739) );
  NOR2_X1 U18941 ( .A1(n15739), .A2(n15713), .ZN(n15718) );
  OAI211_X1 U18942 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15714), .B(n15727), .ZN(
        n15715) );
  OAI211_X1 U18943 ( .C1(n16585), .C2(n16677), .A(n15716), .B(n15715), .ZN(
        n15717) );
  AOI211_X1 U18944 ( .C1(n16573), .C2(n19613), .A(n15718), .B(n15717), .ZN(
        n15719) );
  OAI211_X1 U18945 ( .C1(n15721), .C2(n15974), .A(n15720), .B(n15719), .ZN(
        P2_U3023) );
  NOR2_X1 U18946 ( .A1(n16590), .A2(n15927), .ZN(n15731) );
  NAND2_X1 U18947 ( .A1(n10213), .A2(n15722), .ZN(n15723) );
  NAND2_X1 U18948 ( .A1(n15724), .A2(n15723), .ZN(n16604) );
  NOR2_X1 U18949 ( .A1(n16604), .A2(n16677), .ZN(n15725) );
  AOI211_X1 U18950 ( .C1(n15729), .C2(n15727), .A(n15726), .B(n15725), .ZN(
        n15728) );
  OAI21_X1 U18951 ( .B1(n15739), .B2(n15729), .A(n15728), .ZN(n15730) );
  AOI211_X1 U18952 ( .C1(n15732), .C2(n19606), .A(n15731), .B(n15730), .ZN(
        n15733) );
  OAI21_X1 U18953 ( .B1(n15734), .B2(n16684), .A(n15733), .ZN(P2_U3024) );
  NAND2_X1 U18954 ( .A1(n15735), .A2(n19606), .ZN(n15745) );
  INV_X1 U18955 ( .A(n15736), .ZN(n19313) );
  OAI21_X1 U18956 ( .B1(n15738), .B2(n16677), .A(n15737), .ZN(n15743) );
  AOI21_X1 U18957 ( .B1(n15741), .B2(n15740), .A(n15739), .ZN(n15742) );
  AOI211_X1 U18958 ( .C1(n19313), .C2(n19613), .A(n15743), .B(n15742), .ZN(
        n15744) );
  OAI211_X1 U18959 ( .C1(n15746), .C2(n16684), .A(n15745), .B(n15744), .ZN(
        P2_U3025) );
  OR2_X1 U18960 ( .A1(n15747), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15763) );
  AOI21_X1 U18961 ( .B1(n15763), .B2(n15764), .A(n15748), .ZN(n15755) );
  NAND4_X1 U18962 ( .A1(n15922), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15749), .A4(n15748), .ZN(n15753) );
  AOI21_X1 U18963 ( .B1(n15751), .B2(n19604), .A(n15750), .ZN(n15752) );
  OAI211_X1 U18964 ( .C1(n16596), .C2(n15927), .A(n15753), .B(n15752), .ZN(
        n15754) );
  AOI211_X1 U18965 ( .C1(n15756), .C2(n19611), .A(n15755), .B(n15754), .ZN(
        n15757) );
  OAI21_X1 U18966 ( .B1(n15758), .B2(n15974), .A(n15757), .ZN(P2_U3026) );
  INV_X1 U18967 ( .A(n19327), .ZN(n15761) );
  OAI21_X1 U18968 ( .B1(n19326), .B2(n16677), .A(n15759), .ZN(n15760) );
  AOI21_X1 U18969 ( .B1(n15761), .B2(n19613), .A(n15760), .ZN(n15762) );
  OAI211_X1 U18970 ( .C1(n15765), .C2(n15764), .A(n15763), .B(n15762), .ZN(
        n15766) );
  AOI21_X1 U18971 ( .B1(n15767), .B2(n19611), .A(n15766), .ZN(n15768) );
  OAI21_X1 U18972 ( .B1(n15769), .B2(n15974), .A(n15768), .ZN(P2_U3027) );
  INV_X1 U18973 ( .A(n15922), .ZN(n15863) );
  INV_X1 U18974 ( .A(n15770), .ZN(n15771) );
  NOR3_X1 U18975 ( .A1(n15863), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15771), .ZN(n15776) );
  OAI211_X1 U18976 ( .C1(n15780), .C2(n15771), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n15893), .ZN(n15774) );
  AOI21_X1 U18977 ( .B1(n19604), .B2(n16618), .A(n15772), .ZN(n15773) );
  OAI211_X1 U18978 ( .C1(n16602), .C2(n15927), .A(n15774), .B(n15773), .ZN(
        n15775) );
  AOI211_X1 U18979 ( .C1(n15777), .C2(n19611), .A(n15776), .B(n15775), .ZN(
        n15778) );
  OAI21_X1 U18980 ( .B1(n15779), .B2(n15974), .A(n15778), .ZN(P2_U3028) );
  INV_X1 U18981 ( .A(n15780), .ZN(n15912) );
  INV_X1 U18982 ( .A(n15893), .ZN(n15824) );
  AOI21_X1 U18983 ( .B1(n15912), .B2(n15788), .A(n15824), .ZN(n15815) );
  AOI21_X1 U18984 ( .B1(n16684), .B2(n15782), .A(n15781), .ZN(n15783) );
  INV_X1 U18985 ( .A(n15787), .ZN(n15789) );
  NAND2_X1 U18986 ( .A1(n15922), .A2(n15788), .ZN(n15818) );
  OAI21_X1 U18987 ( .B1(n15789), .B2(n16684), .A(n15818), .ZN(n15801) );
  NAND3_X1 U18988 ( .A1(n15801), .A2(n15791), .A3(n15790), .ZN(n15795) );
  INV_X1 U18989 ( .A(n19346), .ZN(n15793) );
  AOI21_X1 U18990 ( .B1(n19604), .B2(n15793), .A(n15792), .ZN(n15794) );
  OAI211_X1 U18991 ( .C1(n15796), .C2(n15927), .A(n15795), .B(n15794), .ZN(
        n15797) );
  INV_X1 U18992 ( .A(n15799), .ZN(n15806) );
  NAND3_X1 U18993 ( .A1(n15801), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15800), .ZN(n15804) );
  AOI21_X1 U18994 ( .B1(n19604), .B2(n19498), .A(n15802), .ZN(n15803) );
  OAI211_X1 U18995 ( .C1(n19470), .C2(n15927), .A(n15804), .B(n15803), .ZN(
        n15805) );
  AOI21_X1 U18996 ( .B1(n15806), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15805), .ZN(n15807) );
  OAI21_X1 U18997 ( .B1(n15808), .B2(n15974), .A(n15807), .ZN(P2_U3030) );
  INV_X1 U18998 ( .A(n15809), .ZN(n19355) );
  OAI21_X1 U18999 ( .B1(n15812), .B2(n15811), .A(n15810), .ZN(n19506) );
  OAI21_X1 U19000 ( .B1(n16677), .B2(n19506), .A(n15813), .ZN(n15814) );
  AOI21_X1 U19001 ( .B1(n19355), .B2(n19613), .A(n15814), .ZN(n15817) );
  NAND2_X1 U19002 ( .A1(n15815), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15816) );
  OAI211_X1 U19003 ( .C1(n15818), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15817), .B(n15816), .ZN(n15819) );
  AOI21_X1 U19004 ( .B1(n15820), .B2(n19611), .A(n15819), .ZN(n15821) );
  OAI21_X1 U19005 ( .B1(n15822), .B2(n15974), .A(n15821), .ZN(P2_U3031) );
  INV_X1 U19006 ( .A(n15825), .ZN(n15823) );
  NOR2_X1 U19007 ( .A1(n15863), .A2(n15823), .ZN(n15859) );
  AOI21_X1 U19008 ( .B1(n15912), .B2(n15825), .A(n15824), .ZN(n15851) );
  AOI21_X1 U19009 ( .B1(n15859), .B2(n15826), .A(n15851), .ZN(n15844) );
  INV_X1 U19010 ( .A(n15844), .ZN(n15834) );
  NAND3_X1 U19011 ( .A1(n15859), .A2(n15828), .A3(n15827), .ZN(n15831) );
  AOI21_X1 U19012 ( .B1(n19604), .B2(n19508), .A(n15829), .ZN(n15830) );
  OAI211_X1 U19013 ( .C1(n15832), .C2(n15927), .A(n15831), .B(n15830), .ZN(
        n15833) );
  AOI21_X1 U19014 ( .B1(n15834), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15833), .ZN(n15837) );
  NAND2_X1 U19015 ( .A1(n15835), .A2(n19611), .ZN(n15836) );
  OAI211_X1 U19016 ( .C1(n15838), .C2(n15974), .A(n15837), .B(n15836), .ZN(
        P2_U3032) );
  AOI21_X1 U19017 ( .B1(n15859), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15843) );
  NOR2_X1 U19018 ( .A1(n16677), .A2(n19511), .ZN(n15839) );
  AOI211_X1 U19019 ( .C1(n15841), .C2(n19613), .A(n15840), .B(n15839), .ZN(
        n15842) );
  OAI21_X1 U19020 ( .B1(n15844), .B2(n15843), .A(n15842), .ZN(n15845) );
  AOI21_X1 U19021 ( .B1(n15846), .B2(n19606), .A(n15845), .ZN(n15847) );
  OAI21_X1 U19022 ( .B1(n15848), .B2(n16684), .A(n15847), .ZN(P2_U3033) );
  NAND3_X1 U19023 ( .A1(n15850), .A2(n19611), .A3(n15849), .ZN(n15861) );
  NAND2_X1 U19024 ( .A1(n15851), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15856) );
  NOR2_X1 U19025 ( .A1(n15864), .A2(n15852), .ZN(n15853) );
  NOR2_X1 U19026 ( .A1(n12821), .A2(n15853), .ZN(n19513) );
  AOI21_X1 U19027 ( .B1(n19604), .B2(n19513), .A(n15854), .ZN(n15855) );
  OAI211_X1 U19028 ( .C1(n19475), .C2(n15927), .A(n15856), .B(n15855), .ZN(
        n15857) );
  AOI21_X1 U19029 ( .B1(n15859), .B2(n15858), .A(n15857), .ZN(n15860) );
  OAI211_X1 U19030 ( .C1(n15862), .C2(n15974), .A(n15861), .B(n15860), .ZN(
        P2_U3034) );
  NAND2_X1 U19031 ( .A1(n15912), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15894) );
  NOR3_X1 U19032 ( .A1(n15863), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15921), .ZN(n15901) );
  AOI21_X1 U19033 ( .B1(n15893), .B2(n15894), .A(n15901), .ZN(n15876) );
  INV_X1 U19034 ( .A(n15864), .ZN(n15869) );
  INV_X1 U19035 ( .A(n15865), .ZN(n15867) );
  NAND2_X1 U19036 ( .A1(n15895), .A2(n15906), .ZN(n15866) );
  NAND2_X1 U19037 ( .A1(n15867), .A2(n15866), .ZN(n15868) );
  NAND2_X1 U19038 ( .A1(n15869), .A2(n15868), .ZN(n19516) );
  OAI21_X1 U19039 ( .B1(n16677), .B2(n19516), .A(n15870), .ZN(n15871) );
  AOI21_X1 U19040 ( .B1(n19613), .B2(n19375), .A(n15871), .ZN(n15874) );
  NAND3_X1 U19041 ( .A1(n15922), .A2(n15872), .A3(n15875), .ZN(n15873) );
  OAI211_X1 U19042 ( .C1(n15876), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        n15877) );
  AOI21_X1 U19043 ( .B1(n15878), .B2(n19611), .A(n15877), .ZN(n15879) );
  OAI21_X1 U19044 ( .B1(n15880), .B2(n15974), .A(n15879), .ZN(P2_U3035) );
  OR2_X1 U19045 ( .A1(n15913), .A2(n15917), .ZN(n15884) );
  NAND2_X1 U19046 ( .A1(n10207), .A2(n15882), .ZN(n15883) );
  XNOR2_X1 U19047 ( .A(n15884), .B(n15883), .ZN(n16624) );
  INV_X1 U19048 ( .A(n16624), .ZN(n15904) );
  NAND2_X1 U19049 ( .A1(n15905), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15886) );
  NAND2_X1 U19050 ( .A1(n15886), .A2(n15885), .ZN(n15887) );
  NAND2_X1 U19051 ( .A1(n15888), .A2(n15887), .ZN(n16628) );
  INV_X1 U19052 ( .A(n16628), .ZN(n15902) );
  NAND2_X1 U19053 ( .A1(n15890), .A2(n15889), .ZN(n15891) );
  NAND2_X1 U19054 ( .A1(n15892), .A2(n15891), .ZN(n19478) );
  NAND3_X1 U19055 ( .A1(n15894), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15893), .ZN(n15899) );
  XNOR2_X1 U19056 ( .A(n15895), .B(n15906), .ZN(n19519) );
  INV_X1 U19057 ( .A(n19519), .ZN(n15897) );
  NOR2_X1 U19058 ( .A1(n12603), .A2(n19424), .ZN(n15896) );
  AOI21_X1 U19059 ( .B1(n19604), .B2(n15897), .A(n15896), .ZN(n15898) );
  OAI211_X1 U19060 ( .C1(n19478), .C2(n15927), .A(n15899), .B(n15898), .ZN(
        n15900) );
  AOI211_X1 U19061 ( .C1(n15902), .C2(n19611), .A(n15901), .B(n15900), .ZN(
        n15903) );
  OAI21_X1 U19062 ( .B1(n15904), .B2(n15974), .A(n15903), .ZN(P2_U3036) );
  XNOR2_X1 U19063 ( .A(n15905), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16632) );
  NOR2_X1 U19064 ( .A1(n12600), .A2(n19424), .ZN(n15910) );
  INV_X1 U19065 ( .A(n15906), .ZN(n15907) );
  OAI21_X1 U19066 ( .B1(n15908), .B2(n9745), .A(n15907), .ZN(n19521) );
  NOR2_X1 U19067 ( .A1(n16677), .A2(n19521), .ZN(n15909) );
  AOI211_X1 U19068 ( .C1(n19397), .C2(n19613), .A(n15910), .B(n15909), .ZN(
        n15911) );
  OAI21_X1 U19069 ( .B1(n15912), .B2(n15921), .A(n15911), .ZN(n15920) );
  INV_X1 U19070 ( .A(n15913), .ZN(n15918) );
  OAI21_X1 U19071 ( .B1(n15915), .B2(n15917), .A(n15914), .ZN(n15916) );
  OAI21_X1 U19072 ( .B1(n15918), .B2(n15917), .A(n15916), .ZN(n16633) );
  NOR2_X1 U19073 ( .A1(n16633), .A2(n15974), .ZN(n15919) );
  AOI211_X1 U19074 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        n15923) );
  OAI21_X1 U19075 ( .B1(n16632), .B2(n16684), .A(n15923), .ZN(P2_U3037) );
  NOR2_X1 U19076 ( .A1(n16673), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15932) );
  OAI21_X1 U19077 ( .B1(n15926), .B2(n15925), .A(n15924), .ZN(n19527) );
  NOR2_X1 U19078 ( .A1(n20194), .A2(n19424), .ZN(n15929) );
  NOR2_X1 U19079 ( .A1(n15927), .A2(n19406), .ZN(n15928) );
  AOI211_X1 U19080 ( .C1(n16671), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15929), .B(n15928), .ZN(n15930) );
  OAI21_X1 U19081 ( .B1(n19527), .B2(n16677), .A(n15930), .ZN(n15931) );
  AOI211_X1 U19082 ( .C1(n15933), .C2(n19606), .A(n15932), .B(n15931), .ZN(
        n15934) );
  OAI21_X1 U19083 ( .B1(n15935), .B2(n16684), .A(n15934), .ZN(P2_U3039) );
  XNOR2_X1 U19084 ( .A(n15937), .B(n15936), .ZN(n16654) );
  XNOR2_X1 U19085 ( .A(n15939), .B(n15938), .ZN(n19530) );
  INV_X1 U19086 ( .A(n19530), .ZN(n15949) );
  NAND4_X1 U19087 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15963), .A3(
        n15941), .A4(n15940), .ZN(n15944) );
  AOI22_X1 U19088 ( .A1(n19613), .A2(n19419), .B1(n19592), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U19089 ( .A1(n16671), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15942) );
  NAND3_X1 U19090 ( .A1(n15944), .A2(n15943), .A3(n15942), .ZN(n15948) );
  OAI21_X1 U19091 ( .B1(n15946), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15945), .ZN(n16657) );
  NOR2_X1 U19092 ( .A1(n16657), .A2(n16684), .ZN(n15947) );
  AOI211_X1 U19093 ( .C1(n19604), .C2(n15949), .A(n15948), .B(n15947), .ZN(
        n15950) );
  OAI21_X1 U19094 ( .B1(n15974), .B2(n16654), .A(n15950), .ZN(P2_U3040) );
  XNOR2_X1 U19095 ( .A(n15952), .B(n15951), .ZN(n16666) );
  INV_X1 U19096 ( .A(n15954), .ZN(n15957) );
  AND2_X1 U19097 ( .A1(n15954), .A2(n15953), .ZN(n15955) );
  OAI22_X1 U19098 ( .A1(n15958), .A2(n15957), .B1(n15956), .B2(n15955), .ZN(
        n16663) );
  INV_X1 U19099 ( .A(n16663), .ZN(n15972) );
  OAI21_X1 U19100 ( .B1(n15961), .B2(n15960), .A(n15959), .ZN(n19531) );
  AOI211_X1 U19101 ( .C1(n15965), .C2(n15964), .A(n15963), .B(n15962), .ZN(
        n15967) );
  INV_X1 U19102 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20190) );
  NOR2_X1 U19103 ( .A1(n20190), .A2(n19424), .ZN(n15966) );
  AOI211_X1 U19104 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15968), .A(
        n15967), .B(n15966), .ZN(n15970) );
  NAND2_X1 U19105 ( .A1(n19613), .A2(n19436), .ZN(n15969) );
  OAI211_X1 U19106 ( .C1(n19531), .C2(n16677), .A(n15970), .B(n15969), .ZN(
        n15971) );
  AOI21_X1 U19107 ( .B1(n15972), .B2(n19611), .A(n15971), .ZN(n15973) );
  OAI21_X1 U19108 ( .B1(n15974), .B2(n16666), .A(n15973), .ZN(P2_U3041) );
  AOI21_X1 U19109 ( .B1(n19416), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15975), .ZN(n15989) );
  NAND2_X1 U19110 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15976), .ZN(n15988) );
  INV_X1 U19111 ( .A(n15988), .ZN(n15983) );
  INV_X1 U19112 ( .A(n15977), .ZN(n15981) );
  INV_X1 U19113 ( .A(n15993), .ZN(n16710) );
  OAI22_X1 U19114 ( .A1(n16710), .A2(n15984), .B1(n15979), .B2(n15978), .ZN(
        n15980) );
  AOI22_X1 U19115 ( .A1(n19612), .A2(n16006), .B1(n15981), .B2(n15980), .ZN(
        n16714) );
  OAI22_X1 U19116 ( .A1(n20265), .A2(n16021), .B1(n19283), .B2(n16714), .ZN(
        n15982) );
  AOI21_X1 U19117 ( .B1(n15989), .B2(n15983), .A(n15982), .ZN(n15987) );
  NAND2_X1 U19118 ( .A1(n15986), .A2(n15984), .ZN(n15985) );
  OAI21_X1 U19119 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(P2_U3600) );
  NOR2_X1 U19120 ( .A1(n15989), .A2(n15988), .ZN(n16004) );
  INV_X1 U19121 ( .A(n15990), .ZN(n16699) );
  NOR2_X1 U19122 ( .A1(n15991), .A2(n16699), .ZN(n16011) );
  NOR2_X1 U19123 ( .A1(n15977), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16007) );
  NOR2_X1 U19124 ( .A1(n16007), .A2(n16013), .ZN(n15997) );
  NOR2_X1 U19125 ( .A1(n16011), .A2(n15997), .ZN(n16000) );
  INV_X1 U19126 ( .A(n15992), .ZN(n16012) );
  NAND2_X1 U19127 ( .A1(n15993), .A2(n16012), .ZN(n16008) );
  AND2_X1 U19128 ( .A1(n15996), .A2(n15995), .ZN(n16009) );
  INV_X1 U19129 ( .A(n15997), .ZN(n15998) );
  OAI22_X1 U19130 ( .A1(n16008), .A2(n15994), .B1(n16009), .B2(n15998), .ZN(
        n15999) );
  AOI211_X1 U19131 ( .C1(n16001), .C2(n16006), .A(n16000), .B(n15999), .ZN(
        n16692) );
  OAI22_X1 U19132 ( .A1(n16002), .A2(n16021), .B1(n19283), .B2(n16692), .ZN(
        n16003) );
  OAI21_X1 U19133 ( .B1(n16004), .B2(n16003), .A(n16022), .ZN(n16005) );
  OAI21_X1 U19134 ( .B1(n16022), .B2(n12397), .A(n16005), .ZN(P2_U3599) );
  NAND2_X1 U19135 ( .A1(n9675), .A2(n16006), .ZN(n16019) );
  INV_X1 U19136 ( .A(n16007), .ZN(n16014) );
  OAI211_X1 U19137 ( .C1(n16009), .C2(n16013), .A(n16008), .B(n16014), .ZN(
        n16010) );
  INV_X1 U19138 ( .A(n16010), .ZN(n16017) );
  OAI21_X1 U19139 ( .B1(n16710), .B2(n16012), .A(n16011), .ZN(n16015) );
  AOI21_X1 U19140 ( .B1(n16015), .B2(n16014), .A(n16013), .ZN(n16016) );
  MUX2_X1 U19141 ( .A(n16017), .B(n16016), .S(n12026), .Z(n16018) );
  NAND2_X1 U19142 ( .A1(n16019), .A2(n16018), .ZN(n16693) );
  INV_X1 U19143 ( .A(n16693), .ZN(n16020) );
  OAI22_X1 U19144 ( .A1(n20248), .A2(n16021), .B1(n19283), .B2(n16020), .ZN(
        n16023) );
  MUX2_X1 U19145 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16023), .S(
        n16022), .Z(P2_U3596) );
  NOR3_X1 U19146 ( .A1(n20262), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19786) );
  INV_X1 U19147 ( .A(n19786), .ZN(n19788) );
  NOR2_X1 U19148 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19788), .ZN(
        n19775) );
  INV_X1 U19149 ( .A(n19775), .ZN(n16044) );
  NAND2_X1 U19150 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16044), .ZN(n16024) );
  AND2_X1 U19151 ( .A1(n16026), .A2(n16025), .ZN(n16027) );
  OAI21_X1 U19152 ( .B1(n19760), .B2(n19800), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16031) );
  INV_X1 U19153 ( .A(n16029), .ZN(n19985) );
  AND2_X1 U19154 ( .A1(n19985), .A2(n16030), .ZN(n19995) );
  NAND2_X1 U19155 ( .A1(n19995), .A2(n20254), .ZN(n16034) );
  AOI22_X1 U19156 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n16044), .B1(n16031), 
        .B2(n16034), .ZN(n16032) );
  AND2_X1 U19157 ( .A1(n20098), .A2(n16032), .ZN(n16033) );
  INV_X1 U19158 ( .A(n19777), .ZN(n19764) );
  INV_X1 U19159 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16047) );
  OAI21_X1 U19160 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16034), .A(n19955), 
        .ZN(n16035) );
  AND2_X1 U19161 ( .A1(n16036), .A2(n16035), .ZN(n19776) );
  AND2_X1 U19162 ( .A1(n16039), .A2(n19658), .ZN(n20092) );
  INV_X1 U19163 ( .A(n20092), .ZN(n19832) );
  INV_X1 U19164 ( .A(n19657), .ZN(n16108) );
  INV_X1 U19165 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18604) );
  INV_X1 U19166 ( .A(n19656), .ZN(n16107) );
  OAI22_X2 U19167 ( .A1(n16822), .A2(n16108), .B1(n18604), .B2(n16107), .ZN(
        n20100) );
  AOI22_X1 U19168 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19656), .ZN(n20103) );
  INV_X1 U19169 ( .A(n20103), .ZN(n20019) );
  AOI22_X1 U19170 ( .A1(n19760), .A2(n20100), .B1(n19800), .B2(n20019), .ZN(
        n16043) );
  OAI21_X1 U19171 ( .B1(n19832), .B2(n16044), .A(n16043), .ZN(n16045) );
  AOI21_X1 U19172 ( .B1(n19776), .B2(n16038), .A(n16045), .ZN(n16046) );
  OAI21_X1 U19173 ( .B1(n19764), .B2(n16047), .A(n16046), .ZN(P2_U3080) );
  NOR2_X1 U19174 ( .A1(n20281), .A2(n19788), .ZN(n19805) );
  AOI21_X1 U19175 ( .B1(n19829), .B2(n19880), .A(n20049), .ZN(n16048) );
  NOR2_X1 U19176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19835), .ZN(
        n19824) );
  AOI221_X1 U19177 ( .B1(n19805), .B2(n20153), .C1(n16048), .C2(n20153), .A(
        n19824), .ZN(n16051) );
  INV_X1 U19178 ( .A(n16049), .ZN(n16050) );
  NOR3_X1 U19179 ( .A1(n16050), .A2(n19824), .A3(n19955), .ZN(n16053) );
  INV_X1 U19180 ( .A(n19826), .ZN(n16058) );
  AOI22_X1 U19181 ( .A1(n19817), .A2(n20100), .B1(n19868), .B2(n20019), .ZN(
        n16056) );
  NOR2_X1 U19182 ( .A1(n19805), .A2(n19824), .ZN(n16052) );
  OR2_X1 U19183 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n16052), .ZN(n16054) );
  AOI21_X1 U19184 ( .B1(n19955), .B2(n16054), .A(n16053), .ZN(n19825) );
  AOI22_X1 U19185 ( .A1(n19825), .A2(n16038), .B1(n20092), .B2(n19824), .ZN(
        n16055) );
  OAI211_X1 U19186 ( .C1(n16058), .C2(n16057), .A(n16056), .B(n16055), .ZN(
        P2_U3096) );
  NAND2_X1 U19187 ( .A1(n20046), .A2(n19667), .ZN(n19925) );
  NOR2_X1 U19188 ( .A1(n19914), .A2(n19896), .ZN(n16059) );
  OAI21_X1 U19189 ( .B1(n16059), .B2(n20049), .A(n20243), .ZN(n16066) );
  INV_X1 U19190 ( .A(n16066), .ZN(n16061) );
  NAND2_X1 U19191 ( .A1(n20262), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19947) );
  INV_X1 U19192 ( .A(n19947), .ZN(n19950) );
  NAND2_X1 U19193 ( .A1(n19950), .A2(n20272), .ZN(n16085) );
  NOR2_X1 U19194 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16085), .ZN(
        n19895) );
  NOR2_X1 U19195 ( .A1(n19839), .A2(n19895), .ZN(n16064) );
  AOI211_X1 U19196 ( .C1(n14292), .C2(n20153), .A(n19895), .B(n20243), .ZN(
        n16060) );
  INV_X1 U19197 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16069) );
  INV_X1 U19198 ( .A(n20100), .ZN(n16062) );
  INV_X1 U19199 ( .A(n19895), .ZN(n16072) );
  OAI22_X1 U19200 ( .A1(n16062), .A2(n19871), .B1(n19832), .B2(n16072), .ZN(
        n16063) );
  AOI21_X1 U19201 ( .B1(n19914), .B2(n20019), .A(n16063), .ZN(n16068) );
  OAI21_X1 U19202 ( .B1(n14292), .B2(n19895), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16065) );
  NAND2_X1 U19203 ( .A1(n19897), .A2(n16038), .ZN(n16067) );
  OAI211_X1 U19204 ( .C1(n19901), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        P2_U3112) );
  AOI22_X1 U19205 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19656), .ZN(n20066) );
  INV_X1 U19206 ( .A(n20066), .ZN(n20106) );
  NAND2_X1 U19207 ( .A1(n16070), .A2(n19658), .ZN(n20062) );
  AOI22_X1 U19208 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19656), .ZN(n20109) );
  NAND2_X1 U19209 ( .A1(n20023), .A2(n19896), .ZN(n16071) );
  OAI21_X1 U19210 ( .B1(n16072), .B2(n20062), .A(n16071), .ZN(n16073) );
  AOI21_X1 U19211 ( .B1(n19914), .B2(n20106), .A(n16073), .ZN(n16075) );
  NOR2_X2 U19212 ( .A1(n19556), .A2(n19782), .ZN(n20105) );
  NAND2_X1 U19213 ( .A1(n19897), .A2(n20105), .ZN(n16074) );
  OAI211_X1 U19214 ( .C1(n19901), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        P2_U3113) );
  OR2_X1 U19215 ( .A1(n20248), .A2(n20049), .ZN(n20094) );
  OAI21_X1 U19216 ( .B1(n19671), .B2(n20094), .A(n20243), .ZN(n16086) );
  INV_X1 U19217 ( .A(n16085), .ZN(n16077) );
  OR2_X1 U19218 ( .A1(n16086), .A2(n16077), .ZN(n16081) );
  NAND2_X1 U19219 ( .A1(n16083), .A2(n20153), .ZN(n16079) );
  NAND2_X1 U19220 ( .A1(n20272), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19668) );
  NOR2_X1 U19221 ( .A1(n19668), .A2(n19947), .ZN(n19920) );
  NOR2_X1 U19222 ( .A1(n19920), .A2(n20243), .ZN(n16078) );
  AOI21_X1 U19223 ( .B1(n16079), .B2(n16078), .A(n19782), .ZN(n16080) );
  NAND2_X1 U19224 ( .A1(n16081), .A2(n16080), .ZN(n19922) );
  INV_X1 U19225 ( .A(n19922), .ZN(n19907) );
  INV_X1 U19226 ( .A(n19920), .ZN(n19908) );
  OAI22_X1 U19227 ( .A1(n19925), .A2(n20109), .B1(n20062), .B2(n19908), .ZN(
        n16082) );
  AOI21_X1 U19228 ( .B1(n20106), .B2(n19942), .A(n16082), .ZN(n16088) );
  OAI21_X1 U19229 ( .B1(n16083), .B2(n19920), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16084) );
  OAI21_X1 U19230 ( .B1(n16086), .B2(n16085), .A(n16084), .ZN(n19921) );
  NAND2_X1 U19231 ( .A1(n19921), .A2(n20105), .ZN(n16087) );
  OAI211_X1 U19232 ( .C1(n19907), .C2(n16089), .A(n16088), .B(n16087), .ZN(
        P2_U3121) );
  AOI221_X1 U19233 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19975), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n19942), .A(n19920), .ZN(n16090) );
  MUX2_X1 U19234 ( .A(n14283), .B(n16090), .S(n19955), .Z(n16092) );
  NOR2_X1 U19235 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20272), .ZN(
        n19699) );
  AND2_X1 U19236 ( .A1(n19699), .A2(n19950), .ZN(n19940) );
  INV_X1 U19237 ( .A(n19940), .ZN(n16091) );
  OAI21_X1 U19238 ( .B1(n16092), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16091), 
        .ZN(n16093) );
  NAND2_X1 U19239 ( .A1(n16093), .A2(n20098), .ZN(n19943) );
  INV_X1 U19240 ( .A(n19943), .ZN(n19931) );
  AOI22_X1 U19241 ( .A1(n19942), .A2(n20100), .B1(n19975), .B2(n20019), .ZN(
        n16097) );
  INV_X1 U19242 ( .A(n14283), .ZN(n16094) );
  OAI21_X1 U19243 ( .B1(n16094), .B2(n19940), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16095) );
  OAI21_X1 U19244 ( .B1(n19947), .B2(n19700), .A(n16095), .ZN(n19941) );
  AOI22_X1 U19245 ( .A1(n19941), .A2(n16038), .B1(n20092), .B2(n19940), .ZN(
        n16096) );
  OAI211_X1 U19246 ( .C1(n19931), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P2_U3128) );
  NAND3_X1 U19247 ( .A1(n20272), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U19248 ( .B1(n20094), .B2(n19781), .A(n19984), .ZN(n16103) );
  NOR2_X1 U19249 ( .A1(n20281), .A2(n19984), .ZN(n20051) );
  INV_X1 U19250 ( .A(n20051), .ZN(n16099) );
  AND2_X1 U19251 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16099), .ZN(n16100) );
  NAND2_X1 U19252 ( .A1(n14296), .A2(n16100), .ZN(n16110) );
  OAI211_X1 U19253 ( .C1(n20051), .C2(n20153), .A(n16110), .B(n20098), .ZN(
        n16101) );
  INV_X1 U19254 ( .A(n16101), .ZN(n16102) );
  NAND2_X1 U19255 ( .A1(n16103), .A2(n16102), .ZN(n20041) );
  INV_X1 U19256 ( .A(n20041), .ZN(n20026) );
  AOI22_X1 U19257 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19656), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19657), .ZN(n20141) );
  INV_X1 U19258 ( .A(n20141), .ZN(n20009) );
  INV_X1 U19259 ( .A(n20090), .ZN(n20048) );
  INV_X1 U19260 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18634) );
  OAI22_X2 U19261 ( .A1(n16826), .A2(n16108), .B1(n18634), .B2(n16107), .ZN(
        n20138) );
  AOI22_X1 U19262 ( .A1(n20040), .A2(n20009), .B1(n20048), .B2(n20138), .ZN(
        n16112) );
  OAI21_X1 U19263 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19984), .A(n19955), 
        .ZN(n16109) );
  AND2_X1 U19264 ( .A1(n16110), .A2(n16109), .ZN(n20038) );
  NOR2_X2 U19265 ( .A1(n19528), .A2(n19782), .ZN(n20137) );
  NOR2_X2 U19266 ( .A1(n11844), .A2(n19637), .ZN(n20136) );
  AOI22_X1 U19267 ( .A1(n20038), .A2(n20137), .B1(n20136), .B2(n20051), .ZN(
        n16111) );
  OAI211_X1 U19268 ( .C1(n20026), .C2(n16113), .A(n16112), .B(n16111), .ZN(
        P2_U3158) );
  INV_X1 U19269 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17043) );
  INV_X1 U19270 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17383) );
  AND2_X1 U19271 ( .A1(n18642), .A2(n17437), .ZN(n17422) );
  NAND2_X1 U19272 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17409), .ZN(n17382) );
  NAND2_X1 U19273 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17381), .ZN(n17367) );
  INV_X1 U19274 ( .A(n16114), .ZN(n17363) );
  NOR2_X1 U19275 ( .A1(n17367), .A2(n17363), .ZN(n17357) );
  NAND2_X1 U19276 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17357), .ZN(n16190) );
  NOR2_X1 U19277 ( .A1(n17729), .A2(n17586), .ZN(n17617) );
  INV_X1 U19278 ( .A(n17617), .ZN(n17615) );
  NOR2_X1 U19279 ( .A1(n17618), .A2(n17357), .ZN(n17358) );
  INV_X1 U19280 ( .A(n17358), .ZN(n17365) );
  OAI21_X1 U19281 ( .B1(n17352), .B2(n17615), .A(n17365), .ZN(n17350) );
  AOI22_X1 U19282 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16118) );
  AOI22_X1 U19283 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U19284 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16116) );
  AOI22_X1 U19285 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16115) );
  NAND4_X1 U19286 ( .A1(n16118), .A2(n16117), .A3(n16116), .A4(n16115), .ZN(
        n16124) );
  AOI22_X1 U19287 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16122) );
  AOI22_X1 U19288 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16121) );
  AOI22_X1 U19289 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16120) );
  AOI22_X1 U19290 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16119) );
  NAND4_X1 U19291 ( .A1(n16122), .A2(n16121), .A3(n16120), .A4(n16119), .ZN(
        n16123) );
  NOR2_X1 U19292 ( .A1(n16124), .A2(n16123), .ZN(n16188) );
  AOI22_X1 U19293 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16128) );
  AOI22_X1 U19294 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U19295 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16126) );
  AOI22_X1 U19296 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16125) );
  NAND4_X1 U19297 ( .A1(n16128), .A2(n16127), .A3(n16126), .A4(n16125), .ZN(
        n16134) );
  AOI22_X1 U19298 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16132) );
  AOI22_X1 U19299 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U19300 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16130) );
  AOI22_X1 U19301 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16129) );
  NAND4_X1 U19302 ( .A1(n16132), .A2(n16131), .A3(n16130), .A4(n16129), .ZN(
        n16133) );
  NOR2_X1 U19303 ( .A1(n16134), .A2(n16133), .ZN(n17361) );
  AOI22_X1 U19304 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16138) );
  AOI22_X1 U19305 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17566), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17567), .ZN(n16137) );
  AOI22_X1 U19306 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16136) );
  AOI22_X1 U19307 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9651), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16135) );
  NAND4_X1 U19308 ( .A1(n16138), .A2(n16137), .A3(n16136), .A4(n16135), .ZN(
        n16144) );
  AOI22_X1 U19309 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16142) );
  AOI22_X1 U19310 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n11555), .ZN(n16141) );
  AOI22_X1 U19311 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17537), .ZN(n16140) );
  AOI22_X1 U19312 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17455), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11513), .ZN(n16139) );
  NAND4_X1 U19313 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        n16143) );
  NOR2_X1 U19314 ( .A1(n16144), .A2(n16143), .ZN(n17373) );
  AOI22_X1 U19315 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U19316 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16154) );
  AOI22_X1 U19317 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16145) );
  OAI21_X1 U19318 ( .B1(n17333), .B2(n16146), .A(n16145), .ZN(n16152) );
  AOI22_X1 U19319 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16150) );
  AOI22_X1 U19320 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16149) );
  AOI22_X1 U19321 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16148) );
  AOI22_X1 U19322 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16147) );
  NAND4_X1 U19323 ( .A1(n16150), .A2(n16149), .A3(n16148), .A4(n16147), .ZN(
        n16151) );
  AOI211_X1 U19324 ( .C1(n9653), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n16152), .B(n16151), .ZN(n16153) );
  NAND3_X1 U19325 ( .A1(n16155), .A2(n16154), .A3(n16153), .ZN(n17378) );
  AOI22_X1 U19326 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16165) );
  AOI22_X1 U19327 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16164) );
  AOI22_X1 U19328 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16163) );
  NOR2_X1 U19329 ( .A1(n10220), .A2(n17589), .ZN(n16161) );
  AOI22_X1 U19330 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16159) );
  AOI22_X1 U19331 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U19332 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16157) );
  AOI22_X1 U19333 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16156) );
  NAND4_X1 U19334 ( .A1(n16159), .A2(n16158), .A3(n16157), .A4(n16156), .ZN(
        n16160) );
  AOI211_X1 U19335 ( .C1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n17573), .A(
        n16161), .B(n16160), .ZN(n16162) );
  NAND4_X1 U19336 ( .A1(n16165), .A2(n16164), .A3(n16163), .A4(n16162), .ZN(
        n17379) );
  NAND2_X1 U19337 ( .A1(n17378), .A2(n17379), .ZN(n17377) );
  NOR2_X1 U19338 ( .A1(n17373), .A2(n17377), .ZN(n17372) );
  AOI22_X1 U19339 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16175) );
  AOI22_X1 U19340 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16174) );
  AOI22_X1 U19341 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16166) );
  OAI21_X1 U19342 ( .B1(n17333), .B2(n17612), .A(n16166), .ZN(n16172) );
  AOI22_X1 U19343 ( .A1(n11553), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16170) );
  AOI22_X1 U19344 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16169) );
  AOI22_X1 U19345 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U19346 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16167) );
  NAND4_X1 U19347 ( .A1(n16170), .A2(n16169), .A3(n16168), .A4(n16167), .ZN(
        n16171) );
  AOI211_X1 U19348 ( .C1(n17466), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n16172), .B(n16171), .ZN(n16173) );
  NAND3_X1 U19349 ( .A1(n16175), .A2(n16174), .A3(n16173), .ZN(n17369) );
  NAND2_X1 U19350 ( .A1(n17372), .A2(n17369), .ZN(n17368) );
  NOR2_X1 U19351 ( .A1(n17361), .A2(n17368), .ZN(n17360) );
  AOI22_X1 U19352 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16187) );
  INV_X1 U19353 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16178) );
  AOI22_X1 U19354 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16177) );
  AOI22_X1 U19355 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16176) );
  OAI211_X1 U19356 ( .C1(n16179), .C2(n16178), .A(n16177), .B(n16176), .ZN(
        n16185) );
  AOI22_X1 U19357 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U19358 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16182) );
  AOI22_X1 U19359 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U19360 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16180) );
  NAND4_X1 U19361 ( .A1(n16183), .A2(n16182), .A3(n16181), .A4(n16180), .ZN(
        n16184) );
  AOI211_X1 U19362 ( .C1(n17455), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n16185), .B(n16184), .ZN(n16186) );
  NAND2_X1 U19363 ( .A1(n16187), .A2(n16186), .ZN(n17355) );
  NAND2_X1 U19364 ( .A1(n17360), .A2(n17355), .ZN(n17354) );
  NOR2_X1 U19365 ( .A1(n16188), .A2(n17354), .ZN(n17349) );
  AOI21_X1 U19366 ( .B1(n16188), .B2(n17354), .A(n17349), .ZN(n17640) );
  AOI22_X1 U19367 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17350), .B1(n17640), 
        .B2(n17618), .ZN(n16189) );
  OAI21_X1 U19368 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16190), .A(n16189), .ZN(
        P3_U2675) );
  AOI22_X1 U19369 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16195) );
  AOI22_X1 U19370 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16194) );
  AOI22_X1 U19371 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U19372 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16192) );
  NAND4_X1 U19373 ( .A1(n16195), .A2(n16194), .A3(n16193), .A4(n16192), .ZN(
        n16202) );
  AOI22_X1 U19374 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U19375 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16196), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16199) );
  AOI22_X1 U19376 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16198) );
  AOI22_X1 U19377 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16197) );
  NAND4_X1 U19378 ( .A1(n16200), .A2(n16199), .A3(n16198), .A4(n16197), .ZN(
        n16201) );
  NOR2_X1 U19379 ( .A1(n16202), .A2(n16201), .ZN(n17719) );
  INV_X1 U19380 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17550) );
  AND3_X1 U19381 ( .A1(n17621), .A2(n17585), .A3(n16203), .ZN(n17591) );
  NAND2_X1 U19382 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17591), .ZN(n17583) );
  NOR2_X1 U19383 ( .A1(n17550), .A2(n17583), .ZN(n17565) );
  NAND2_X1 U19384 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17565), .ZN(n17548) );
  NOR2_X1 U19385 ( .A1(n16204), .A2(n17548), .ZN(n16205) );
  INV_X1 U19386 ( .A(n16205), .ZN(n17519) );
  INV_X1 U19387 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U19388 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17519), .B1(n16205), 
        .B2(n17504), .ZN(n16206) );
  AOI22_X1 U19389 ( .A1(n17618), .A2(n17719), .B1(n16206), .B2(n17596), .ZN(
        P3_U2690) );
  NAND2_X1 U19390 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18822) );
  AOI221_X1 U19391 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18822), .C1(n16208), 
        .C2(n18822), .A(n16207), .ZN(n18602) );
  NOR2_X1 U19392 ( .A1(n16209), .A2(n19076), .ZN(n16210) );
  OAI21_X1 U19393 ( .B1(n16210), .B2(n18897), .A(n18603), .ZN(n18600) );
  AOI22_X1 U19394 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18602), .B1(
        n18600), .B2(n19081), .ZN(P3_U2865) );
  INV_X1 U19395 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16796) );
  NAND2_X1 U19396 ( .A1(n17906), .A2(n16211), .ZN(n16284) );
  AOI21_X1 U19397 ( .B1(n16284), .B2(n16285), .A(n16212), .ZN(n16213) );
  XOR2_X1 U19398 ( .A(n16796), .B(n16213), .Z(n16791) );
  NOR2_X1 U19399 ( .A1(n18592), .A2(n18312), .ZN(n18538) );
  INV_X1 U19400 ( .A(n18538), .ZN(n18577) );
  NOR2_X1 U19401 ( .A1(n16796), .A2(n16216), .ZN(n16786) );
  NAND2_X1 U19402 ( .A1(n17746), .A2(n18590), .ZN(n18429) );
  NOR2_X1 U19403 ( .A1(n16774), .A2(n16796), .ZN(n16773) );
  NOR2_X1 U19404 ( .A1(n18304), .A2(n18592), .ZN(n18588) );
  INV_X1 U19405 ( .A(n18588), .ZN(n18435) );
  OAI22_X1 U19406 ( .A1(n16786), .A2(n18429), .B1(n16773), .B2(n18435), .ZN(
        n16291) );
  AOI211_X1 U19407 ( .C1(n18575), .C2(n16214), .A(n18569), .B(n16291), .ZN(
        n16215) );
  OAI21_X1 U19408 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18577), .A(
        n16215), .ZN(n16218) );
  NAND3_X1 U19409 ( .A1(n18575), .A2(n16769), .A3(n18291), .ZN(n16794) );
  INV_X1 U19410 ( .A(n16216), .ZN(n16788) );
  INV_X1 U19411 ( .A(n18429), .ZN(n18505) );
  NAND2_X1 U19412 ( .A1(n16788), .A2(n18505), .ZN(n16217) );
  OAI211_X1 U19413 ( .C1(n18435), .C2(n16774), .A(n16794), .B(n16217), .ZN(
        n16287) );
  AOI22_X1 U19414 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16218), .B1(
        n16287), .B2(n16796), .ZN(n16219) );
  NAND2_X1 U19415 ( .A1(n18570), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16780) );
  OAI211_X1 U19416 ( .C1(n18509), .C2(n16791), .A(n16219), .B(n16780), .ZN(
        P3_U2833) );
  AOI22_X1 U19417 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19443), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19444), .ZN(n16229) );
  OAI22_X1 U19418 ( .A1(n16220), .A2(n19427), .B1(n19390), .B2(n10020), .ZN(
        n16221) );
  INV_X1 U19419 ( .A(n16221), .ZN(n16228) );
  OAI22_X1 U19420 ( .A1(n16590), .A2(n19453), .B1(n16604), .B2(n19442), .ZN(
        n16222) );
  INV_X1 U19421 ( .A(n16222), .ZN(n16227) );
  OAI211_X1 U19422 ( .C1(n16225), .C2(n16224), .A(n19420), .B(n16223), .ZN(
        n16226) );
  NAND4_X1 U19423 ( .A1(n16229), .A2(n16228), .A3(n16227), .A4(n16226), .ZN(
        P2_U2833) );
  NAND2_X1 U19424 ( .A1(n16231), .A2(n16230), .ZN(n16237) );
  AOI21_X1 U19425 ( .B1(n16232), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20690), .ZN(n16233) );
  OAI211_X1 U19426 ( .C1(n16237), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16234), .B(n16233), .ZN(n16235) );
  INV_X1 U19427 ( .A(n16235), .ZN(n16236) );
  AOI21_X1 U19428 ( .B1(n16237), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16236), .ZN(n16238) );
  AOI222_X1 U19429 ( .A1(n20722), .A2(n16239), .B1(n20722), .B2(n16238), .C1(
        n16239), .C2(n16238), .ZN(n16243) );
  INV_X1 U19430 ( .A(n16243), .ZN(n16241) );
  OAI21_X1 U19431 ( .B1(n16241), .B2(n20862), .A(n16240), .ZN(n16242) );
  OAI21_X1 U19432 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16243), .A(
        n16242), .ZN(n16270) );
  INV_X1 U19433 ( .A(n16244), .ZN(n16269) );
  INV_X1 U19434 ( .A(n16245), .ZN(n16252) );
  INV_X1 U19435 ( .A(n16246), .ZN(n16248) );
  NAND3_X1 U19436 ( .A1(n16248), .A2(n12928), .A3(n16247), .ZN(n16250) );
  MUX2_X1 U19437 ( .A(n16250), .B(n16249), .S(n16254), .Z(n16251) );
  AOI21_X1 U19438 ( .B1(n12846), .B2(n16252), .A(n16251), .ZN(n21057) );
  INV_X1 U19439 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n16263) );
  INV_X1 U19440 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n16262) );
  OR2_X1 U19441 ( .A1(n16254), .A2(n16253), .ZN(n16258) );
  INV_X1 U19442 ( .A(n16255), .ZN(n16256) );
  NAND2_X1 U19443 ( .A1(n16256), .A2(n12928), .ZN(n16257) );
  NAND2_X1 U19444 ( .A1(n16258), .A2(n16257), .ZN(n20295) );
  NAND2_X1 U19445 ( .A1(n16260), .A2(n16259), .ZN(n21063) );
  AOI21_X1 U19446 ( .B1(n21063), .B2(n21061), .A(n20965), .ZN(n16261) );
  OR2_X1 U19447 ( .A1(n20295), .A2(n16261), .ZN(n20301) );
  AOI21_X1 U19448 ( .B1(n16263), .B2(n16262), .A(n20301), .ZN(n16265) );
  NOR2_X1 U19449 ( .A1(n16265), .A2(n16264), .ZN(n16266) );
  NAND3_X1 U19450 ( .A1(n16267), .A2(n21057), .A3(n16266), .ZN(n16268) );
  AOI211_X1 U19451 ( .C1(n16270), .C2(n20451), .A(n16269), .B(n16268), .ZN(
        n16283) );
  INV_X1 U19452 ( .A(n16283), .ZN(n16277) );
  NAND2_X1 U19453 ( .A1(n16272), .A2(n16271), .ZN(n16275) );
  NOR3_X1 U19454 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20769), .A3(n21064), 
        .ZN(n16273) );
  OAI22_X1 U19455 ( .A1(n16276), .A2(n16275), .B1(n16274), .B2(n16273), .ZN(
        n16488) );
  AOI221_X1 U19456 ( .B1(n10532), .B2(n16490), .C1(n16277), .C2(n16490), .A(
        n16488), .ZN(n16279) );
  NOR2_X1 U19457 ( .A1(n16279), .A2(n10532), .ZN(n20962) );
  OAI211_X1 U19458 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21064), .A(n20962), 
        .B(n16278), .ZN(n16489) );
  AOI21_X1 U19459 ( .B1(n21068), .B2(n21038), .A(n16279), .ZN(n16280) );
  OAI22_X1 U19460 ( .A1(n16281), .A2(n16489), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16280), .ZN(n16282) );
  OAI21_X1 U19461 ( .B1(n16283), .B2(n20294), .A(n16282), .ZN(P1_U3161) );
  NAND3_X1 U19462 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16289) );
  NAND2_X1 U19463 ( .A1(n16752), .A2(n16754), .ZN(n16286) );
  XNOR2_X1 U19464 ( .A(n16286), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16772) );
  INV_X1 U19465 ( .A(n18591), .ZN(n18581) );
  NOR2_X1 U19466 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16796), .ZN(
        n16768) );
  AOI22_X1 U19467 ( .A1(n18581), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16768), 
        .B2(n16287), .ZN(n16293) );
  AOI211_X1 U19468 ( .C1(n18499), .C2(n16289), .A(n18592), .B(n16288), .ZN(
        n16290) );
  NOR2_X1 U19469 ( .A1(n18570), .A2(n16290), .ZN(n16792) );
  OAI21_X1 U19470 ( .B1(n16792), .B2(n16291), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16292) );
  OAI211_X1 U19471 ( .C1(n16772), .C2(n18509), .A(n16293), .B(n16292), .ZN(
        P3_U2832) );
  INV_X1 U19472 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20979) );
  OAI221_X1 U19473 ( .B1(n20965), .B2(HOLD), .C1(n20965), .C2(n20979), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n16295) );
  INV_X1 U19474 ( .A(HOLD), .ZN(n20966) );
  OAI211_X1 U19475 ( .C1(n20979), .C2(n20966), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n16294) );
  NAND3_X1 U19476 ( .A1(n16295), .A2(n21061), .A3(n16294), .ZN(P1_U3195) );
  AND2_X1 U19477 ( .A1(n20391), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19478 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16735), .A3(n20155), 
        .ZN(n16725) );
  NOR3_X1 U19479 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATE2_REG_0__SCAN_IN), .ZN(n16296) );
  NOR4_X1 U19480 ( .A1(n16733), .A2(n16740), .A3(n16725), .A4(n16296), .ZN(
        P2_U3178) );
  INV_X1 U19481 ( .A(n20284), .ZN(n16297) );
  INV_X1 U19482 ( .A(n20279), .ZN(n20280) );
  NOR2_X1 U19483 ( .A1(n16298), .A2(n20280), .ZN(P2_U3047) );
  OAI221_X1 U19484 ( .B1(n16302), .B2(n16301), .C1(n16302), .C2(n16300), .A(
        n19251), .ZN(n17624) );
  INV_X1 U19485 ( .A(n17624), .ZN(n16303) );
  INV_X1 U19486 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17836) );
  NAND2_X1 U19487 ( .A1(n18642), .A2(n16303), .ZN(n17742) );
  NOR2_X1 U19488 ( .A1(n17836), .A2(n17742), .ZN(n17764) );
  NAND2_X1 U19489 ( .A1(n17763), .A2(n17775), .ZN(n17774) );
  AOI22_X1 U19490 ( .A1(n17772), .A2(BUF2_REG_0__SCAN_IN), .B1(n17771), .B2(
        n16304), .ZN(n16305) );
  OAI221_X1 U19491 ( .B1(n17774), .B2(n17836), .C1(n17774), .C2(n17742), .A(
        n16305), .ZN(P3_U2735) );
  INV_X1 U19492 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21009) );
  NAND2_X1 U19493 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16306) );
  OAI211_X1 U19494 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n16317), .B(n16306), .ZN(n16310) );
  OAI22_X1 U19495 ( .A1(n16307), .A2(n20363), .B1(n16419), .B2(n20377), .ZN(
        n16308) );
  AOI211_X1 U19496 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20334), .B(n16308), .ZN(n16309) );
  OAI211_X1 U19497 ( .C1(n16339), .C2(n20361), .A(n16310), .B(n16309), .ZN(
        n16311) );
  AOI21_X1 U19498 ( .B1(n16336), .B2(n20327), .A(n16311), .ZN(n16312) );
  OAI21_X1 U19499 ( .B1(n21009), .B2(n16321), .A(n16312), .ZN(P1_U2824) );
  INV_X1 U19500 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21007) );
  INV_X1 U19501 ( .A(n16313), .ZN(n16314) );
  AOI22_X1 U19502 ( .A1(n20346), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n20319), 
        .B2(n16314), .ZN(n16315) );
  OAI21_X1 U19503 ( .B1(n20377), .B2(n16426), .A(n16315), .ZN(n16316) );
  AOI211_X1 U19504 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20334), .B(n16316), .ZN(n16320) );
  AOI22_X1 U19505 ( .A1(n16318), .A2(n20327), .B1(n21007), .B2(n16317), .ZN(
        n16319) );
  OAI211_X1 U19506 ( .C1(n21007), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        P1_U2825) );
  NOR2_X1 U19507 ( .A1(n20361), .A2(n16359), .ZN(n16323) );
  OAI21_X1 U19508 ( .B1(n20321), .B2(n10929), .A(n20347), .ZN(n16322) );
  AOI211_X1 U19509 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n20346), .A(n16323), .B(
        n16322), .ZN(n16325) );
  NAND2_X1 U19510 ( .A1(n16438), .A2(n20345), .ZN(n16324) );
  OAI211_X1 U19511 ( .C1(n16326), .C2(n20999), .A(n16325), .B(n16324), .ZN(
        n16327) );
  AOI21_X1 U19512 ( .B1(n16356), .B2(n20327), .A(n16327), .ZN(n16328) );
  OAI21_X1 U19513 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16329), .A(n16328), 
        .ZN(P1_U2829) );
  AOI22_X1 U19514 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16338) );
  INV_X1 U19515 ( .A(n16330), .ZN(n16332) );
  OAI21_X1 U19516 ( .B1(n16333), .B2(n16332), .A(n16331), .ZN(n16335) );
  XNOR2_X1 U19517 ( .A(n16335), .B(n16334), .ZN(n16422) );
  AOI22_X1 U19518 ( .A1(n16336), .A2(n16364), .B1(n20302), .B2(n16422), .ZN(
        n16337) );
  OAI211_X1 U19519 ( .C1(n16370), .C2(n16339), .A(n16338), .B(n16337), .ZN(
        P1_U2983) );
  AOI22_X1 U19520 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U19521 ( .A1(n16341), .A2(n16364), .B1(n16361), .B2(n16340), .ZN(
        n16342) );
  OAI211_X1 U19522 ( .C1(n16344), .C2(n16349), .A(n16343), .B(n16342), .ZN(
        P1_U2985) );
  AOI22_X1 U19523 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16348) );
  AOI22_X1 U19524 ( .A1(n16346), .A2(n16364), .B1(n16361), .B2(n16345), .ZN(
        n16347) );
  OAI211_X1 U19525 ( .C1(n16350), .C2(n16349), .A(n16348), .B(n16347), .ZN(
        P1_U2987) );
  AOI22_X1 U19526 ( .A1(n16351), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20334), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16358) );
  NOR3_X1 U19527 ( .A1(n12829), .A2(n16352), .A3(n12917), .ZN(n16354) );
  NOR2_X1 U19528 ( .A1(n16354), .A2(n16353), .ZN(n16355) );
  XNOR2_X1 U19529 ( .A(n16355), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16440) );
  AOI22_X1 U19530 ( .A1(n16440), .A2(n20302), .B1(n16364), .B2(n16356), .ZN(
        n16357) );
  OAI211_X1 U19531 ( .C1(n16370), .C2(n16359), .A(n16358), .B(n16357), .ZN(
        P1_U2988) );
  INV_X1 U19532 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16368) );
  INV_X1 U19533 ( .A(n16360), .ZN(n16362) );
  AOI222_X1 U19534 ( .A1(n16365), .A2(n20302), .B1(n16364), .B2(n16363), .C1(
        n16362), .C2(n16361), .ZN(n16367) );
  OAI211_X1 U19535 ( .C1(n16368), .C2(n16375), .A(n16367), .B(n16366), .ZN(
        P1_U2992) );
  OAI22_X1 U19536 ( .A1(n20332), .A2(n16371), .B1(n20336), .B2(n16370), .ZN(
        n16372) );
  AOI21_X1 U19537 ( .B1(n16478), .B2(n20302), .A(n16372), .ZN(n16374) );
  INV_X1 U19538 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20987) );
  NOR2_X1 U19539 ( .A1(n20347), .A2(n20987), .ZN(n16474) );
  INV_X1 U19540 ( .A(n16474), .ZN(n16373) );
  OAI211_X1 U19541 ( .C1(n16376), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        P1_U2994) );
  INV_X1 U19542 ( .A(n16377), .ZN(n16382) );
  INV_X1 U19543 ( .A(n16378), .ZN(n16381) );
  INV_X1 U19544 ( .A(n16379), .ZN(n16380) );
  AOI222_X1 U19545 ( .A1(n16382), .A2(n20439), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16381), .C1(n20438), .C2(
        n16380), .ZN(n16386) );
  OAI211_X1 U19546 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16384), .B(n16383), .ZN(
        n16385) );
  OAI211_X1 U19547 ( .C1(n21168), .C2(n20347), .A(n16386), .B(n16385), .ZN(
        P1_U3009) );
  INV_X1 U19548 ( .A(n16387), .ZN(n16389) );
  AOI22_X1 U19549 ( .A1(n16389), .A2(n20439), .B1(n20438), .B2(n16388), .ZN(
        n16396) );
  INV_X1 U19550 ( .A(n16390), .ZN(n16392) );
  NOR2_X1 U19551 ( .A1(n20347), .A2(n21014), .ZN(n16391) );
  AOI221_X1 U19552 ( .B1(n16394), .B2(n16393), .C1(n16392), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16391), .ZN(n16395) );
  NAND2_X1 U19553 ( .A1(n16396), .A2(n16395), .ZN(P1_U3012) );
  NAND2_X1 U19554 ( .A1(n16398), .A2(n16418), .ZN(n16405) );
  AND2_X1 U19555 ( .A1(n16416), .A2(n16406), .ZN(n16397) );
  NOR2_X1 U19556 ( .A1(n16433), .A2(n16397), .ZN(n16415) );
  NOR2_X1 U19557 ( .A1(n16415), .A2(n16398), .ZN(n16401) );
  AND3_X1 U19558 ( .A1(n16399), .A2(n20439), .A3(n14948), .ZN(n16400) );
  AOI211_X1 U19559 ( .C1(n20438), .C2(n16402), .A(n16401), .B(n16400), .ZN(
        n16404) );
  NAND2_X1 U19560 ( .A1(n20334), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16403) );
  OAI211_X1 U19561 ( .C1(n16406), .C2(n16405), .A(n16404), .B(n16403), .ZN(
        P1_U3013) );
  NOR3_X1 U19562 ( .A1(n16417), .A2(n10739), .A3(n16424), .ZN(n16407) );
  AOI21_X1 U19563 ( .B1(n16407), .B2(n16418), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16414) );
  INV_X1 U19564 ( .A(n16408), .ZN(n16411) );
  INV_X1 U19565 ( .A(n16409), .ZN(n16410) );
  AOI22_X1 U19566 ( .A1(n16411), .A2(n20439), .B1(n20438), .B2(n16410), .ZN(
        n16413) );
  NAND2_X1 U19567 ( .A1(n20334), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16412) );
  OAI211_X1 U19568 ( .C1(n16415), .C2(n16414), .A(n16413), .B(n16412), .ZN(
        P1_U3014) );
  AOI21_X1 U19569 ( .B1(n16417), .B2(n16416), .A(n16433), .ZN(n16429) );
  NAND2_X1 U19570 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16418), .ZN(
        n16430) );
  AOI221_X1 U19571 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n10739), .C2(n16424), .A(
        n16430), .ZN(n16421) );
  OAI22_X1 U19572 ( .A1(n16419), .A2(n16466), .B1(n21009), .B2(n20347), .ZN(
        n16420) );
  AOI211_X1 U19573 ( .C1(n16422), .C2(n20439), .A(n16421), .B(n16420), .ZN(
        n16423) );
  OAI21_X1 U19574 ( .B1(n16429), .B2(n16424), .A(n16423), .ZN(P1_U3015) );
  OAI222_X1 U19575 ( .A1(n16426), .A2(n16466), .B1(n20347), .B2(n21007), .C1(
        n20431), .C2(n16425), .ZN(n16427) );
  INV_X1 U19576 ( .A(n16427), .ZN(n16428) );
  OAI221_X1 U19577 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16430), 
        .C1(n10739), .C2(n16429), .A(n16428), .ZN(P1_U3016) );
  AOI21_X1 U19578 ( .B1(n16432), .B2(n20438), .A(n16431), .ZN(n16436) );
  AOI22_X1 U19579 ( .A1(n16434), .A2(n20439), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16433), .ZN(n16435) );
  OAI211_X1 U19580 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16437), .A(
        n16436), .B(n16435), .ZN(P1_U3018) );
  AOI22_X1 U19581 ( .A1(n16438), .A2(n20438), .B1(n20334), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19582 ( .A1(n16440), .A2(n20439), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16439), .ZN(n16441) );
  OAI211_X1 U19583 ( .C1(n16444), .C2(n16443), .A(n16442), .B(n16441), .ZN(
        P1_U3020) );
  OAI211_X1 U19584 ( .C1(n16448), .C2(n16447), .A(n16446), .B(n16445), .ZN(
        n16450) );
  OAI21_X1 U19585 ( .B1(n16451), .B2(n16450), .A(n16449), .ZN(n16464) );
  INV_X1 U19586 ( .A(n16452), .ZN(n16457) );
  NAND3_X1 U19587 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16469), .ZN(n16459) );
  AOI221_X1 U19588 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12917), .C2(n14059), .A(
        n16459), .ZN(n16453) );
  AOI21_X1 U19589 ( .B1(n20334), .B2(P1_REIP_REG_10__SCAN_IN), .A(n16453), 
        .ZN(n16454) );
  OAI21_X1 U19590 ( .B1(n16455), .B2(n16466), .A(n16454), .ZN(n16456) );
  AOI21_X1 U19591 ( .B1(n16457), .B2(n20439), .A(n16456), .ZN(n16458) );
  OAI21_X1 U19592 ( .B1(n12917), .B2(n16464), .A(n16458), .ZN(P1_U3021) );
  INV_X1 U19593 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20995) );
  OAI22_X1 U19594 ( .A1(n20347), .A2(n20995), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16459), .ZN(n16462) );
  NOR2_X1 U19595 ( .A1(n16460), .A2(n20431), .ZN(n16461) );
  AOI211_X1 U19596 ( .C1(n20438), .C2(n20325), .A(n16462), .B(n16461), .ZN(
        n16463) );
  OAI21_X1 U19597 ( .B1(n14059), .B2(n16464), .A(n16463), .ZN(P1_U3022) );
  INV_X1 U19598 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20992) );
  OAI22_X1 U19599 ( .A1(n16466), .A2(n16465), .B1(n20992), .B2(n20347), .ZN(
        n16467) );
  AOI21_X1 U19600 ( .B1(n16468), .B2(n20439), .A(n16467), .ZN(n16471) );
  OAI221_X1 U19601 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16472), .C2(n10717), .A(
        n16469), .ZN(n16470) );
  OAI211_X1 U19602 ( .C1(n16473), .C2(n16472), .A(n16471), .B(n16470), .ZN(
        P1_U3023) );
  AOI21_X1 U19603 ( .B1(n20438), .B2(n20333), .A(n16474), .ZN(n16475) );
  OAI21_X1 U19604 ( .B1(n16476), .B2(n10669), .A(n16475), .ZN(n16477) );
  AOI21_X1 U19605 ( .B1(n16478), .B2(n20439), .A(n16477), .ZN(n16479) );
  OAI21_X1 U19606 ( .B1(n16481), .B2(n16480), .A(n16479), .ZN(P1_U3026) );
  INV_X1 U19607 ( .A(n16482), .ZN(n16483) );
  NAND3_X1 U19608 ( .A1(n16484), .A2(n21040), .A3(n16483), .ZN(n16485) );
  OAI21_X1 U19609 ( .B1(n21045), .B2(n16486), .A(n16485), .ZN(P1_U3468) );
  OAI221_X1 U19610 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n10532), .C2(n21064), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20963) );
  NAND2_X1 U19611 ( .A1(n16491), .A2(n20963), .ZN(n16487) );
  AOI22_X1 U19612 ( .A1(n16490), .A2(n16489), .B1(n16488), .B2(n16487), .ZN(
        P1_U3162) );
  OAI22_X1 U19613 ( .A1(n20962), .A2(n20811), .B1(n10532), .B2(n16491), .ZN(
        P1_U3466) );
  NAND2_X1 U19614 ( .A1(n16492), .A2(n9647), .ZN(n16520) );
  INV_X1 U19615 ( .A(n16493), .ZN(n16521) );
  NAND2_X1 U19616 ( .A1(n9647), .A2(n16519), .ZN(n16509) );
  NOR3_X1 U19617 ( .A1(n16495), .A2(n16586), .A3(n16494), .ZN(n16496) );
  AOI21_X1 U19618 ( .B1(n19444), .B2(P2_REIP_REG_31__SCAN_IN), .A(n16496), 
        .ZN(n16497) );
  OAI21_X1 U19619 ( .B1(n16498), .B2(n19427), .A(n16497), .ZN(n16499) );
  AOI21_X1 U19620 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19459), .A(
        n16499), .ZN(n16503) );
  INV_X1 U19621 ( .A(n16500), .ZN(n19491) );
  AOI22_X1 U19622 ( .A1(n16501), .A2(n19437), .B1(n19450), .B2(n19491), .ZN(
        n16502) );
  OAI211_X1 U19623 ( .C1(n16504), .C2(n16508), .A(n16503), .B(n16502), .ZN(
        P2_U2824) );
  AOI22_X1 U19624 ( .A1(n16505), .A2(n19448), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19443), .ZN(n16514) );
  AOI22_X1 U19625 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19459), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19444), .ZN(n16513) );
  OAI22_X1 U19626 ( .A1(n15644), .A2(n19453), .B1(n16506), .B2(n19442), .ZN(
        n16507) );
  INV_X1 U19627 ( .A(n16507), .ZN(n16512) );
  OAI211_X1 U19628 ( .C1(n16510), .C2(n16509), .A(n19438), .B(n16508), .ZN(
        n16511) );
  NAND4_X1 U19629 ( .A1(n16514), .A2(n16513), .A3(n16512), .A4(n16511), .ZN(
        P2_U2825) );
  AOI22_X1 U19630 ( .A1(n16515), .A2(n19448), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n19444), .ZN(n16525) );
  AOI22_X1 U19631 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19459), .ZN(n16524) );
  OAI22_X1 U19632 ( .A1(n16517), .A2(n19453), .B1(n19442), .B2(n16516), .ZN(
        n16518) );
  INV_X1 U19633 ( .A(n16518), .ZN(n16523) );
  OAI211_X1 U19634 ( .C1(n16521), .C2(n16520), .A(n19420), .B(n16519), .ZN(
        n16522) );
  NAND4_X1 U19635 ( .A1(n16525), .A2(n16524), .A3(n16523), .A4(n16522), .ZN(
        P2_U2826) );
  NOR2_X1 U19636 ( .A1(n16526), .A2(n19427), .ZN(n16529) );
  AOI22_X1 U19637 ( .A1(n19443), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19459), .ZN(n16527) );
  OAI21_X1 U19638 ( .B1(n19425), .B2(n20224), .A(n16527), .ZN(n16528) );
  AOI211_X1 U19639 ( .C1(n16530), .C2(n19437), .A(n16529), .B(n16528), .ZN(
        n16535) );
  OAI211_X1 U19640 ( .C1(n16533), .C2(n16532), .A(n19420), .B(n16531), .ZN(
        n16534) );
  OAI211_X1 U19641 ( .C1(n19442), .C2(n16536), .A(n16535), .B(n16534), .ZN(
        P2_U2828) );
  OAI22_X1 U19642 ( .A1(n16537), .A2(n19427), .B1(n20221), .B2(n19425), .ZN(
        n16538) );
  INV_X1 U19643 ( .A(n16538), .ZN(n16548) );
  AOI22_X1 U19644 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19459), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19443), .ZN(n16547) );
  OAI22_X1 U19645 ( .A1(n16540), .A2(n19453), .B1(n16539), .B2(n19442), .ZN(
        n16541) );
  INV_X1 U19646 ( .A(n16541), .ZN(n16546) );
  OAI211_X1 U19647 ( .C1(n16544), .C2(n16543), .A(n19420), .B(n16542), .ZN(
        n16545) );
  NAND4_X1 U19648 ( .A1(n16548), .A2(n16547), .A3(n16546), .A4(n16545), .ZN(
        P2_U2829) );
  AOI22_X1 U19649 ( .A1(n16549), .A2(n19448), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n19444), .ZN(n16560) );
  AOI22_X1 U19650 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19459), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19443), .ZN(n16559) );
  INV_X1 U19651 ( .A(n16550), .ZN(n16553) );
  INV_X1 U19652 ( .A(n16551), .ZN(n16552) );
  AOI22_X1 U19653 ( .A1(n16553), .A2(n19437), .B1(n16552), .B2(n19450), .ZN(
        n16558) );
  OAI211_X1 U19654 ( .C1(n16556), .C2(n16555), .A(n19420), .B(n16554), .ZN(
        n16557) );
  NAND4_X1 U19655 ( .A1(n16560), .A2(n16559), .A3(n16558), .A4(n16557), .ZN(
        P2_U2830) );
  INV_X1 U19656 ( .A(n16561), .ZN(n16562) );
  AOI22_X1 U19657 ( .A1(n16562), .A2(n19448), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n19444), .ZN(n16572) );
  AOI22_X1 U19658 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19459), .ZN(n16571) );
  INV_X1 U19659 ( .A(n16563), .ZN(n16564) );
  AOI22_X1 U19660 ( .A1(n16565), .A2(n19437), .B1(n16564), .B2(n19450), .ZN(
        n16570) );
  OAI211_X1 U19661 ( .C1(n16568), .C2(n16567), .A(n19420), .B(n16566), .ZN(
        n16569) );
  NAND4_X1 U19662 ( .A1(n16572), .A2(n16571), .A3(n16570), .A4(n16569), .ZN(
        P2_U2831) );
  NAND2_X1 U19663 ( .A1(n16573), .A2(n19437), .ZN(n16577) );
  OAI22_X1 U19664 ( .A1(n19429), .A2(n16574), .B1(n20215), .B2(n19425), .ZN(
        n16575) );
  AOI21_X1 U19665 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19459), .A(
        n16575), .ZN(n16576) );
  OAI211_X1 U19666 ( .C1(n16578), .C2(n19427), .A(n16577), .B(n16576), .ZN(
        n16579) );
  INV_X1 U19667 ( .A(n16579), .ZN(n16584) );
  OAI211_X1 U19668 ( .C1(n16582), .C2(n16581), .A(n19420), .B(n16580), .ZN(
        n16583) );
  OAI211_X1 U19669 ( .C1(n19442), .C2(n16585), .A(n16584), .B(n16583), .ZN(
        P2_U2832) );
  AOI22_X1 U19670 ( .A1(n19490), .A2(n16587), .B1(n16586), .B2(n19484), .ZN(
        P2_U2856) );
  AOI21_X1 U19671 ( .B1(n16588), .B2(n15300), .A(n9714), .ZN(n16606) );
  AOI22_X1 U19672 ( .A1(n16606), .A2(n19487), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19484), .ZN(n16589) );
  OAI21_X1 U19673 ( .B1(n19484), .B2(n16590), .A(n16589), .ZN(P2_U2865) );
  AND2_X1 U19674 ( .A1(n16592), .A2(n16591), .ZN(n16593) );
  OR2_X1 U19675 ( .A1(n16593), .A2(n15299), .ZN(n16612) );
  OAI22_X1 U19676 ( .A1(n16612), .A2(n19481), .B1(n19490), .B2(n15208), .ZN(
        n16594) );
  INV_X1 U19677 ( .A(n16594), .ZN(n16595) );
  OAI21_X1 U19678 ( .B1(n19484), .B2(n16596), .A(n16595), .ZN(P2_U2867) );
  INV_X1 U19679 ( .A(n16597), .ZN(n16600) );
  AOI21_X1 U19680 ( .B1(n16600), .B2(n16599), .A(n16598), .ZN(n16620) );
  AOI22_X1 U19681 ( .A1(n16620), .A2(n19487), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19484), .ZN(n16601) );
  OAI21_X1 U19682 ( .B1(n19484), .B2(n16602), .A(n16601), .ZN(P2_U2869) );
  AOI22_X1 U19683 ( .A1(n19495), .A2(n16603), .B1(n19546), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16609) );
  AOI22_X1 U19684 ( .A1(n19497), .A2(BUF2_REG_22__SCAN_IN), .B1(n19496), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16608) );
  INV_X1 U19685 ( .A(n16604), .ZN(n16605) );
  AOI22_X1 U19686 ( .A1(n16606), .A2(n16619), .B1(n19547), .B2(n16605), .ZN(
        n16607) );
  NAND3_X1 U19687 ( .A1(n16609), .A2(n16608), .A3(n16607), .ZN(P2_U2897) );
  AOI22_X1 U19688 ( .A1(n19495), .A2(n16610), .B1(n19546), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U19689 ( .A1(n19497), .A2(BUF2_REG_20__SCAN_IN), .B1(n19496), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16615) );
  OAI22_X1 U19690 ( .A1(n16612), .A2(n19551), .B1(n19538), .B2(n16611), .ZN(
        n16613) );
  INV_X1 U19691 ( .A(n16613), .ZN(n16614) );
  NAND3_X1 U19692 ( .A1(n16616), .A2(n16615), .A3(n16614), .ZN(P2_U2899) );
  AOI22_X1 U19693 ( .A1(n19495), .A2(n16617), .B1(n19546), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U19694 ( .A1(n19497), .A2(BUF2_REG_18__SCAN_IN), .B1(n19496), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16622) );
  AOI22_X1 U19695 ( .A1(n16620), .A2(n16619), .B1(n19547), .B2(n16618), .ZN(
        n16621) );
  NAND3_X1 U19696 ( .A1(n16623), .A2(n16622), .A3(n16621), .ZN(P2_U2901) );
  AOI22_X1 U19697 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19592), .ZN(n16631) );
  NAND2_X1 U19698 ( .A1(n16624), .A2(n19598), .ZN(n16627) );
  INV_X1 U19699 ( .A(n19478), .ZN(n16625) );
  NAND2_X1 U19700 ( .A1(n16625), .A2(n19597), .ZN(n16626) );
  OAI211_X1 U19701 ( .C1(n16628), .C2(n16664), .A(n16627), .B(n16626), .ZN(
        n16629) );
  INV_X1 U19702 ( .A(n16629), .ZN(n16630) );
  OAI211_X1 U19703 ( .C1(n19603), .C2(n19381), .A(n16631), .B(n16630), .ZN(
        P2_U3004) );
  AOI22_X1 U19704 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19592), .B1(n16661), 
        .B2(n19396), .ZN(n16636) );
  OAI22_X1 U19705 ( .A1(n16633), .A2(n16665), .B1(n16632), .B2(n16664), .ZN(
        n16634) );
  AOI21_X1 U19706 ( .B1(n19597), .B2(n19397), .A(n16634), .ZN(n16635) );
  OAI211_X1 U19707 ( .C1(n16670), .C2(n19389), .A(n16636), .B(n16635), .ZN(
        P2_U3005) );
  AOI22_X1 U19708 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19592), .ZN(n16652) );
  NAND2_X1 U19709 ( .A1(n16638), .A2(n16637), .ZN(n16639) );
  NAND2_X1 U19710 ( .A1(n16640), .A2(n16639), .ZN(n16685) );
  NAND2_X1 U19711 ( .A1(n16642), .A2(n16641), .ZN(n16647) );
  INV_X1 U19712 ( .A(n16643), .ZN(n16644) );
  NOR2_X1 U19713 ( .A1(n16645), .A2(n16644), .ZN(n16646) );
  XNOR2_X1 U19714 ( .A(n16647), .B(n16646), .ZN(n16680) );
  NAND2_X1 U19715 ( .A1(n16680), .A2(n19598), .ZN(n16649) );
  INV_X1 U19716 ( .A(n19486), .ZN(n16681) );
  NAND2_X1 U19717 ( .A1(n19597), .A2(n16681), .ZN(n16648) );
  OAI211_X1 U19718 ( .C1(n16685), .C2(n16664), .A(n16649), .B(n16648), .ZN(
        n16650) );
  INV_X1 U19719 ( .A(n16650), .ZN(n16651) );
  OAI211_X1 U19720 ( .C1(n19603), .C2(n16653), .A(n16652), .B(n16651), .ZN(
        P2_U3006) );
  AOI22_X1 U19721 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19592), .ZN(n16660) );
  OR2_X1 U19722 ( .A1(n16654), .A2(n16665), .ZN(n16656) );
  NAND2_X1 U19723 ( .A1(n19597), .A2(n19419), .ZN(n16655) );
  OAI211_X1 U19724 ( .C1(n16657), .C2(n16664), .A(n16656), .B(n16655), .ZN(
        n16658) );
  INV_X1 U19725 ( .A(n16658), .ZN(n16659) );
  OAI211_X1 U19726 ( .C1(n19603), .C2(n19417), .A(n16660), .B(n16659), .ZN(
        P2_U3008) );
  AOI22_X1 U19727 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n16662), .B1(n16661), 
        .B2(n19435), .ZN(n16669) );
  OAI22_X1 U19728 ( .A1(n16666), .A2(n16665), .B1(n16664), .B2(n16663), .ZN(
        n16667) );
  AOI21_X1 U19729 ( .B1(n19597), .B2(n19436), .A(n16667), .ZN(n16668) );
  OAI211_X1 U19730 ( .C1(n16670), .C2(n12686), .A(n16669), .B(n16668), .ZN(
        P2_U3009) );
  INV_X1 U19731 ( .A(n16671), .ZN(n16690) );
  INV_X1 U19732 ( .A(n16672), .ZN(n16674) );
  AOI211_X1 U19733 ( .C1(n16675), .C2(n16689), .A(n16674), .B(n16673), .ZN(
        n16679) );
  OAI22_X1 U19734 ( .A1(n16677), .A2(n16676), .B1(n13870), .B2(n19424), .ZN(
        n16678) );
  NOR2_X1 U19735 ( .A1(n16679), .A2(n16678), .ZN(n16688) );
  NAND2_X1 U19736 ( .A1(n16680), .A2(n19606), .ZN(n16683) );
  NAND2_X1 U19737 ( .A1(n19613), .A2(n16681), .ZN(n16682) );
  OAI211_X1 U19738 ( .C1(n16685), .C2(n16684), .A(n16683), .B(n16682), .ZN(
        n16686) );
  INV_X1 U19739 ( .A(n16686), .ZN(n16687) );
  OAI211_X1 U19740 ( .C1(n16690), .C2(n16689), .A(n16688), .B(n16687), .ZN(
        P2_U3038) );
  NOR2_X1 U19741 ( .A1(n16715), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16691) );
  AOI21_X1 U19742 ( .B1(n16692), .B2(n16715), .A(n16691), .ZN(n16723) );
  MUX2_X1 U19743 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16693), .S(
        n16715), .Z(n16722) );
  NOR4_X1 U19744 ( .A1(n16698), .A2(n9811), .A3(n16695), .A4(n16694), .ZN(
        n19287) );
  OR2_X1 U19745 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16704) );
  OAI22_X1 U19746 ( .A1(n13029), .A2(n16697), .B1(n9670), .B2(n16696), .ZN(
        n16703) );
  AOI22_X1 U19747 ( .A1(n16702), .A2(n16699), .B1(n12466), .B2(n16698), .ZN(
        n16700) );
  OAI21_X1 U19748 ( .B1(n16702), .B2(n16701), .A(n16700), .ZN(n20286) );
  AOI211_X1 U19749 ( .C1(n19287), .C2(n16704), .A(n16703), .B(n20286), .ZN(
        n16705) );
  OAI21_X1 U19750 ( .B1(n12444), .B2(n16715), .A(n16705), .ZN(n16721) );
  NAND2_X1 U19751 ( .A1(n20254), .A2(n20262), .ZN(n19730) );
  INV_X1 U19752 ( .A(n19730), .ZN(n19731) );
  INV_X1 U19753 ( .A(n16723), .ZN(n16707) );
  INV_X1 U19754 ( .A(n16722), .ZN(n16706) );
  OAI22_X1 U19755 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16707), .B1(
        n16706), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16717) );
  INV_X1 U19756 ( .A(n16714), .ZN(n16712) );
  OAI211_X1 U19757 ( .C1(n16710), .C2(n16709), .A(n16708), .B(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16711) );
  OAI21_X1 U19758 ( .B1(n16712), .B2(n20272), .A(n16711), .ZN(n16713) );
  OAI21_X1 U19759 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16714), .A(
        n16713), .ZN(n16716) );
  OAI211_X1 U19760 ( .C1(n19731), .C2(n16717), .A(n16716), .B(n16715), .ZN(
        n16719) );
  AOI22_X1 U19761 ( .A1(n16723), .A2(n19731), .B1(n16722), .B2(n20254), .ZN(
        n16718) );
  AOI21_X1 U19762 ( .B1(n16719), .B2(n16718), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16720) );
  AOI211_X1 U19763 ( .C1(n16723), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        n16739) );
  AOI211_X1 U19764 ( .C1(n16740), .C2(n20284), .A(n16725), .B(n16724), .ZN(
        n16738) );
  INV_X1 U19765 ( .A(n16726), .ZN(n16728) );
  NOR3_X1 U19766 ( .A1(n11925), .A2(n16728), .A3(n16727), .ZN(n16731) );
  INV_X1 U19767 ( .A(n16729), .ZN(n16730) );
  NOR3_X1 U19768 ( .A1(n16731), .A2(n16730), .A3(n19955), .ZN(n16734) );
  AOI22_X1 U19769 ( .A1(n20175), .A2(n16734), .B1(n16733), .B2(n16732), .ZN(
        n16736) );
  OAI221_X1 U19770 ( .B1(n16735), .B2(n16739), .C1(n16735), .C2(n20154), .A(
        n16734), .ZN(n20157) );
  NAND2_X1 U19771 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20157), .ZN(n16741) );
  OAI21_X1 U19772 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16736), .A(n16741), 
        .ZN(n16737) );
  OAI211_X1 U19773 ( .C1(n16739), .C2(n19286), .A(n16738), .B(n16737), .ZN(
        P2_U3176) );
  AOI21_X1 U19774 ( .B1(n16741), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16740), 
        .ZN(n16742) );
  INV_X1 U19775 ( .A(n16742), .ZN(P2_U3593) );
  INV_X1 U19776 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U19777 ( .A1(n16773), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16746) );
  XNOR2_X1 U19778 ( .A(n19218), .B(n16746), .ZN(n16804) );
  INV_X1 U19779 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16951) );
  INV_X1 U19780 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18249) );
  INV_X1 U19781 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17892) );
  INV_X1 U19782 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17992) );
  INV_X1 U19783 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18072) );
  NAND2_X1 U19784 ( .A1(n18213), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18202) );
  NAND4_X1 U19785 ( .A1(n18157), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17134) );
  NAND2_X1 U19786 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17135) );
  INV_X1 U19787 ( .A(n17135), .ZN(n18095) );
  INV_X1 U19788 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18032) );
  INV_X1 U19789 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17932) );
  NAND3_X1 U19790 ( .A1(n17930), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16748) );
  INV_X1 U19791 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16777) );
  INV_X1 U19792 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19192) );
  NOR2_X1 U19793 ( .A1(n19192), .A2(n18491), .ZN(n16798) );
  NAND2_X1 U19794 ( .A1(n19102), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19113) );
  AOI21_X1 U19795 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17969), .A(
        n18981), .ZN(n18009) );
  NAND2_X1 U19796 ( .A1(n16747), .A2(n18105), .ZN(n16764) );
  XNOR2_X1 U19797 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16750) );
  INV_X1 U19798 ( .A(n17969), .ZN(n17918) );
  NOR2_X1 U19799 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17918), .ZN(
        n16778) );
  INV_X1 U19800 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17014) );
  NOR2_X1 U19801 ( .A1(n18249), .A2(n16748), .ZN(n16937) );
  INV_X1 U19802 ( .A(n16937), .ZN(n17896) );
  NOR2_X1 U19803 ( .A1(n17014), .A2(n17896), .ZN(n16936) );
  NAND2_X1 U19804 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16936), .ZN(
        n16935) );
  NOR2_X1 U19805 ( .A1(n17892), .A2(n16935), .ZN(n16934) );
  NAND2_X1 U19806 ( .A1(n18981), .A2(n16749), .ZN(n16782) );
  OAI211_X1 U19807 ( .C1(n16934), .C2(n19113), .A(n18255), .B(n16782), .ZN(
        n16785) );
  NOR2_X1 U19808 ( .A1(n16778), .A2(n16785), .ZN(n16763) );
  OAI22_X1 U19809 ( .A1(n16764), .A2(n16750), .B1(n16763), .B2(n16951), .ZN(
        n16751) );
  AOI211_X1 U19810 ( .C1(n18115), .C2(n17271), .A(n16798), .B(n16751), .ZN(
        n16761) );
  NAND2_X1 U19811 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16753) );
  AOI22_X1 U19812 ( .A1(n18142), .A2(n16753), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n18155), .ZN(n16755) );
  NAND2_X1 U19813 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19218), .ZN(
        n16795) );
  NAND2_X1 U19814 ( .A1(n16786), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16757) );
  XOR2_X1 U19815 ( .A(n16757), .B(n19218), .Z(n16801) );
  INV_X1 U19816 ( .A(n16801), .ZN(n16758) );
  OAI211_X1 U19817 ( .C1(n18259), .C2(n16804), .A(n16761), .B(n16760), .ZN(
        P3_U2799) );
  OAI22_X1 U19818 ( .A1(n16773), .A2(n18259), .B1(n16786), .B2(n18084), .ZN(
        n16767) );
  INV_X1 U19819 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16964) );
  OAI21_X1 U19820 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16775), .A(
        n16762), .ZN(n16962) );
  OAI22_X1 U19821 ( .A1(n16763), .A2(n16964), .B1(n18044), .B2(n16962), .ZN(
        n16766) );
  INV_X1 U19822 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19194) );
  OAI22_X1 U19823 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16764), .B1(
        n18591), .B2(n19194), .ZN(n16765) );
  AOI211_X1 U19824 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16767), .A(
        n16766), .B(n16765), .ZN(n16771) );
  NAND3_X1 U19825 ( .A1(n16769), .A2(n16768), .A3(n18051), .ZN(n16770) );
  OAI211_X1 U19826 ( .C1(n16772), .C2(n18168), .A(n16771), .B(n16770), .ZN(
        P3_U2800) );
  AOI211_X1 U19827 ( .C1(n16774), .C2(n16796), .A(n16773), .B(n18259), .ZN(
        n16784) );
  INV_X1 U19828 ( .A(n16934), .ZN(n16776) );
  AOI21_X1 U19829 ( .B1(n16777), .B2(n16776), .A(n16775), .ZN(n16976) );
  OAI21_X1 U19830 ( .B1(n16778), .B2(n18115), .A(n16976), .ZN(n16779) );
  OAI211_X1 U19831 ( .C1(n16782), .C2(n16781), .A(n16780), .B(n16779), .ZN(
        n16783) );
  AOI211_X1 U19832 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16785), .A(
        n16784), .B(n16783), .ZN(n16790) );
  NOR2_X1 U19833 ( .A1(n16786), .A2(n18084), .ZN(n16787) );
  OAI21_X1 U19834 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16788), .A(
        n16787), .ZN(n16789) );
  OAI211_X1 U19835 ( .C1(n16791), .C2(n18168), .A(n16790), .B(n16789), .ZN(
        P3_U2801) );
  INV_X1 U19836 ( .A(n16792), .ZN(n16793) );
  OAI21_X1 U19837 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18577), .A(
        n16793), .ZN(n16799) );
  NOR3_X1 U19838 ( .A1(n16796), .A2(n16795), .A3(n16794), .ZN(n16797) );
  AOI211_X1 U19839 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16799), .A(
        n16798), .B(n16797), .ZN(n16803) );
  AOI22_X1 U19840 ( .A1(n16801), .A2(n18505), .B1(n16800), .B2(n18489), .ZN(
        n16802) );
  NOR3_X1 U19841 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16806) );
  NOR4_X1 U19842 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16805) );
  INV_X2 U19843 ( .A(n16902), .ZN(U215) );
  NAND4_X1 U19844 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16806), .A3(n16805), .A4(
        U215), .ZN(U213) );
  INV_X1 U19845 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16904) );
  INV_X2 U19846 ( .A(U214), .ZN(n16865) );
  INV_X1 U19847 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16905) );
  OAI222_X1 U19848 ( .A1(U212), .A2(n16904), .B1(n16867), .B2(n16808), .C1(
        U214), .C2(n16905), .ZN(U216) );
  AOI22_X1 U19849 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16864), .ZN(n16809) );
  OAI21_X1 U19850 ( .B1(n16810), .B2(n16867), .A(n16809), .ZN(U217) );
  AOI22_X1 U19851 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16864), .ZN(n16811) );
  OAI21_X1 U19852 ( .B1(n16812), .B2(n16867), .A(n16811), .ZN(U218) );
  AOI22_X1 U19853 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16864), .ZN(n16813) );
  OAI21_X1 U19854 ( .B1(n16814), .B2(n16867), .A(n16813), .ZN(U219) );
  AOI22_X1 U19855 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16864), .ZN(n16815) );
  OAI21_X1 U19856 ( .B1(n16816), .B2(n16867), .A(n16815), .ZN(U220) );
  AOI22_X1 U19857 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16864), .ZN(n16817) );
  OAI21_X1 U19858 ( .B1(n16818), .B2(n16867), .A(n16817), .ZN(U221) );
  AOI22_X1 U19859 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16864), .ZN(n16819) );
  OAI21_X1 U19860 ( .B1(n16820), .B2(n16867), .A(n16819), .ZN(U222) );
  AOI22_X1 U19861 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16864), .ZN(n16821) );
  OAI21_X1 U19862 ( .B1(n16822), .B2(n16867), .A(n16821), .ZN(U223) );
  AOI22_X1 U19863 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16864), .ZN(n16823) );
  OAI21_X1 U19864 ( .B1(n16824), .B2(n16867), .A(n16823), .ZN(U224) );
  AOI22_X1 U19865 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16864), .ZN(n16825) );
  OAI21_X1 U19866 ( .B1(n16826), .B2(n16867), .A(n16825), .ZN(U225) );
  AOI22_X1 U19867 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16864), .ZN(n16827) );
  OAI21_X1 U19868 ( .B1(n16828), .B2(n16867), .A(n16827), .ZN(U226) );
  AOI22_X1 U19869 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16864), .ZN(n16829) );
  OAI21_X1 U19870 ( .B1(n16830), .B2(n16867), .A(n16829), .ZN(U227) );
  AOI22_X1 U19871 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16864), .ZN(n16831) );
  OAI21_X1 U19872 ( .B1(n16832), .B2(n16867), .A(n16831), .ZN(U228) );
  AOI22_X1 U19873 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16864), .ZN(n16833) );
  OAI21_X1 U19874 ( .B1(n16834), .B2(n16867), .A(n16833), .ZN(U229) );
  AOI22_X1 U19875 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16864), .ZN(n16835) );
  OAI21_X1 U19876 ( .B1(n16836), .B2(n16867), .A(n16835), .ZN(U230) );
  AOI22_X1 U19877 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16864), .ZN(n16837) );
  OAI21_X1 U19878 ( .B1(n16838), .B2(n16867), .A(n16837), .ZN(U231) );
  AOI22_X1 U19879 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16864), .ZN(n16839) );
  OAI21_X1 U19880 ( .B1(n13624), .B2(n16867), .A(n16839), .ZN(U232) );
  AOI22_X1 U19881 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16864), .ZN(n16840) );
  OAI21_X1 U19882 ( .B1(n16841), .B2(n16867), .A(n16840), .ZN(U233) );
  AOI22_X1 U19883 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16864), .ZN(n16842) );
  OAI21_X1 U19884 ( .B1(n16843), .B2(n16867), .A(n16842), .ZN(U234) );
  AOI22_X1 U19885 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16864), .ZN(n16844) );
  OAI21_X1 U19886 ( .B1(n16845), .B2(n16867), .A(n16844), .ZN(U235) );
  AOI22_X1 U19887 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16864), .ZN(n16846) );
  OAI21_X1 U19888 ( .B1(n16847), .B2(n16867), .A(n16846), .ZN(U236) );
  AOI22_X1 U19889 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16864), .ZN(n16848) );
  OAI21_X1 U19890 ( .B1(n16849), .B2(n16867), .A(n16848), .ZN(U237) );
  AOI22_X1 U19891 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16864), .ZN(n16850) );
  OAI21_X1 U19892 ( .B1(n12974), .B2(n16867), .A(n16850), .ZN(U238) );
  AOI22_X1 U19893 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16864), .ZN(n16851) );
  OAI21_X1 U19894 ( .B1(n16852), .B2(n16867), .A(n16851), .ZN(U239) );
  AOI22_X1 U19895 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16864), .ZN(n16853) );
  OAI21_X1 U19896 ( .B1(n12982), .B2(n16867), .A(n16853), .ZN(U240) );
  INV_X1 U19897 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U19898 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16864), .ZN(n16854) );
  OAI21_X1 U19899 ( .B1(n16855), .B2(n16867), .A(n16854), .ZN(U241) );
  AOI22_X1 U19900 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16864), .ZN(n16856) );
  OAI21_X1 U19901 ( .B1(n13423), .B2(n16867), .A(n16856), .ZN(U242) );
  AOI22_X1 U19902 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16864), .ZN(n16857) );
  OAI21_X1 U19903 ( .B1(n13410), .B2(n16867), .A(n16857), .ZN(U243) );
  INV_X1 U19904 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U19905 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16864), .ZN(n16858) );
  OAI21_X1 U19906 ( .B1(n16859), .B2(n16867), .A(n16858), .ZN(U244) );
  INV_X1 U19907 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U19908 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16864), .ZN(n16860) );
  OAI21_X1 U19909 ( .B1(n16861), .B2(n16867), .A(n16860), .ZN(U245) );
  INV_X1 U19910 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U19911 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16864), .ZN(n16862) );
  OAI21_X1 U19912 ( .B1(n16863), .B2(n16867), .A(n16862), .ZN(U246) );
  INV_X1 U19913 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U19914 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16865), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16864), .ZN(n16866) );
  OAI21_X1 U19915 ( .B1(n16868), .B2(n16867), .A(n16866), .ZN(U247) );
  OAI22_X1 U19916 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16902), .ZN(n16869) );
  INV_X1 U19917 ( .A(n16869), .ZN(U251) );
  OAI22_X1 U19918 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16902), .ZN(n16870) );
  INV_X1 U19919 ( .A(n16870), .ZN(U252) );
  OAI22_X1 U19920 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16902), .ZN(n16871) );
  INV_X1 U19921 ( .A(n16871), .ZN(U253) );
  OAI22_X1 U19922 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16902), .ZN(n16872) );
  INV_X1 U19923 ( .A(n16872), .ZN(U254) );
  OAI22_X1 U19924 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16902), .ZN(n16873) );
  INV_X1 U19925 ( .A(n16873), .ZN(U255) );
  OAI22_X1 U19926 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16902), .ZN(n16874) );
  INV_X1 U19927 ( .A(n16874), .ZN(U256) );
  OAI22_X1 U19928 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16902), .ZN(n16875) );
  INV_X1 U19929 ( .A(n16875), .ZN(U257) );
  OAI22_X1 U19930 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16902), .ZN(n16876) );
  INV_X1 U19931 ( .A(n16876), .ZN(U258) );
  OAI22_X1 U19932 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16902), .ZN(n16877) );
  INV_X1 U19933 ( .A(n16877), .ZN(U259) );
  OAI22_X1 U19934 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16896), .ZN(n16878) );
  INV_X1 U19935 ( .A(n16878), .ZN(U260) );
  OAI22_X1 U19936 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16896), .ZN(n16879) );
  INV_X1 U19937 ( .A(n16879), .ZN(U261) );
  OAI22_X1 U19938 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16902), .ZN(n16880) );
  INV_X1 U19939 ( .A(n16880), .ZN(U262) );
  OAI22_X1 U19940 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16902), .ZN(n16881) );
  INV_X1 U19941 ( .A(n16881), .ZN(U263) );
  OAI22_X1 U19942 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16902), .ZN(n16882) );
  INV_X1 U19943 ( .A(n16882), .ZN(U264) );
  OAI22_X1 U19944 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16902), .ZN(n16883) );
  INV_X1 U19945 ( .A(n16883), .ZN(U265) );
  OAI22_X1 U19946 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16896), .ZN(n16884) );
  INV_X1 U19947 ( .A(n16884), .ZN(U266) );
  OAI22_X1 U19948 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16896), .ZN(n16885) );
  INV_X1 U19949 ( .A(n16885), .ZN(U267) );
  OAI22_X1 U19950 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16896), .ZN(n16886) );
  INV_X1 U19951 ( .A(n16886), .ZN(U268) );
  OAI22_X1 U19952 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16896), .ZN(n16887) );
  INV_X1 U19953 ( .A(n16887), .ZN(U269) );
  OAI22_X1 U19954 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16896), .ZN(n16888) );
  INV_X1 U19955 ( .A(n16888), .ZN(U270) );
  OAI22_X1 U19956 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16896), .ZN(n16889) );
  INV_X1 U19957 ( .A(n16889), .ZN(U271) );
  OAI22_X1 U19958 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16902), .ZN(n16890) );
  INV_X1 U19959 ( .A(n16890), .ZN(U272) );
  OAI22_X1 U19960 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16902), .ZN(n16891) );
  INV_X1 U19961 ( .A(n16891), .ZN(U273) );
  OAI22_X1 U19962 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16896), .ZN(n16892) );
  INV_X1 U19963 ( .A(n16892), .ZN(U274) );
  OAI22_X1 U19964 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16902), .ZN(n16893) );
  INV_X1 U19965 ( .A(n16893), .ZN(U275) );
  OAI22_X1 U19966 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16902), .ZN(n16894) );
  INV_X1 U19967 ( .A(n16894), .ZN(U276) );
  OAI22_X1 U19968 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16902), .ZN(n16895) );
  INV_X1 U19969 ( .A(n16895), .ZN(U277) );
  OAI22_X1 U19970 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16896), .ZN(n16897) );
  INV_X1 U19971 ( .A(n16897), .ZN(U278) );
  OAI22_X1 U19972 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16902), .ZN(n16898) );
  INV_X1 U19973 ( .A(n16898), .ZN(U279) );
  OAI22_X1 U19974 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16902), .ZN(n16899) );
  INV_X1 U19975 ( .A(n16899), .ZN(U280) );
  OAI22_X1 U19976 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16902), .ZN(n16901) );
  INV_X1 U19977 ( .A(n16901), .ZN(U281) );
  INV_X1 U19978 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U19979 ( .A1(n16902), .A2(n16904), .B1(n17630), .B2(U215), .ZN(U282) );
  INV_X1 U19980 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16903) );
  AOI222_X1 U19981 ( .A1(n16905), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16904), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16903), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16906) );
  INV_X2 U19982 ( .A(n16908), .ZN(n16907) );
  INV_X1 U19983 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19151) );
  INV_X1 U19984 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20198) );
  AOI22_X1 U19985 ( .A1(n16907), .A2(n19151), .B1(n20198), .B2(n16908), .ZN(
        U347) );
  INV_X1 U19986 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19149) );
  INV_X1 U19987 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20197) );
  AOI22_X1 U19988 ( .A1(n16907), .A2(n19149), .B1(n20197), .B2(n16908), .ZN(
        U348) );
  INV_X1 U19989 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19146) );
  INV_X1 U19990 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U19991 ( .A1(n16907), .A2(n19146), .B1(n20196), .B2(n16908), .ZN(
        U349) );
  INV_X1 U19992 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19145) );
  INV_X1 U19993 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20195) );
  AOI22_X1 U19994 ( .A1(n16907), .A2(n19145), .B1(n20195), .B2(n16908), .ZN(
        U350) );
  INV_X1 U19995 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19143) );
  INV_X1 U19996 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20193) );
  AOI22_X1 U19997 ( .A1(n16907), .A2(n19143), .B1(n20193), .B2(n16908), .ZN(
        U351) );
  INV_X1 U19998 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19140) );
  INV_X1 U19999 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U20000 ( .A1(n16907), .A2(n19140), .B1(n20191), .B2(n16908), .ZN(
        U352) );
  INV_X1 U20001 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19139) );
  INV_X1 U20002 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20189) );
  AOI22_X1 U20003 ( .A1(n16907), .A2(n19139), .B1(n20189), .B2(n16908), .ZN(
        U353) );
  INV_X1 U20004 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19137) );
  AOI22_X1 U20005 ( .A1(n16907), .A2(n19137), .B1(n20188), .B2(n16908), .ZN(
        U354) );
  INV_X1 U20006 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19191) );
  INV_X1 U20007 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20227) );
  AOI22_X1 U20008 ( .A1(n16907), .A2(n19191), .B1(n20227), .B2(n16908), .ZN(
        U356) );
  INV_X1 U20009 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19187) );
  INV_X1 U20010 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U20011 ( .A1(n16907), .A2(n19187), .B1(n20225), .B2(n16908), .ZN(
        U357) );
  INV_X1 U20012 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19186) );
  INV_X1 U20013 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20223) );
  AOI22_X1 U20014 ( .A1(n16907), .A2(n19186), .B1(n20223), .B2(n16908), .ZN(
        U358) );
  INV_X1 U20015 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19184) );
  INV_X1 U20016 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20222) );
  AOI22_X1 U20017 ( .A1(n16907), .A2(n19184), .B1(n20222), .B2(n16908), .ZN(
        U359) );
  INV_X1 U20018 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19182) );
  INV_X1 U20019 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20220) );
  AOI22_X1 U20020 ( .A1(n16907), .A2(n19182), .B1(n20220), .B2(n16908), .ZN(
        U360) );
  INV_X1 U20021 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19179) );
  INV_X1 U20022 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U20023 ( .A1(n16907), .A2(n19179), .B1(n20218), .B2(n16908), .ZN(
        U361) );
  INV_X1 U20024 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19177) );
  INV_X1 U20025 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U20026 ( .A1(n16907), .A2(n19177), .B1(n20216), .B2(n16908), .ZN(
        U362) );
  INV_X1 U20027 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19175) );
  INV_X1 U20028 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U20029 ( .A1(n16907), .A2(n19175), .B1(n20214), .B2(n16908), .ZN(
        U363) );
  INV_X1 U20030 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19173) );
  INV_X1 U20031 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20213) );
  AOI22_X1 U20032 ( .A1(n16907), .A2(n19173), .B1(n20213), .B2(n16908), .ZN(
        U364) );
  INV_X1 U20033 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19135) );
  INV_X1 U20034 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20186) );
  AOI22_X1 U20035 ( .A1(n16907), .A2(n19135), .B1(n20186), .B2(n16908), .ZN(
        U365) );
  INV_X1 U20036 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19170) );
  INV_X1 U20037 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20211) );
  AOI22_X1 U20038 ( .A1(n16907), .A2(n19170), .B1(n20211), .B2(n16908), .ZN(
        U366) );
  INV_X1 U20039 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19169) );
  INV_X1 U20040 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U20041 ( .A1(n16907), .A2(n19169), .B1(n20210), .B2(n16908), .ZN(
        U367) );
  INV_X1 U20042 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19167) );
  INV_X1 U20043 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U20044 ( .A1(n16907), .A2(n19167), .B1(n20208), .B2(n16908), .ZN(
        U368) );
  INV_X1 U20045 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19165) );
  INV_X1 U20046 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20207) );
  AOI22_X1 U20047 ( .A1(n16907), .A2(n19165), .B1(n20207), .B2(n16908), .ZN(
        U369) );
  INV_X1 U20048 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19163) );
  INV_X1 U20049 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20205) );
  AOI22_X1 U20050 ( .A1(n16907), .A2(n19163), .B1(n20205), .B2(n16908), .ZN(
        U370) );
  INV_X1 U20051 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19161) );
  INV_X1 U20052 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20204) );
  AOI22_X1 U20053 ( .A1(n16907), .A2(n19161), .B1(n20204), .B2(n16908), .ZN(
        U371) );
  INV_X1 U20054 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19158) );
  INV_X1 U20055 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20202) );
  AOI22_X1 U20056 ( .A1(n16907), .A2(n19158), .B1(n20202), .B2(n16908), .ZN(
        U372) );
  INV_X1 U20057 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19157) );
  INV_X1 U20058 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20201) );
  AOI22_X1 U20059 ( .A1(n16907), .A2(n19157), .B1(n20201), .B2(n16908), .ZN(
        U373) );
  INV_X1 U20060 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19155) );
  INV_X1 U20061 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20200) );
  AOI22_X1 U20062 ( .A1(n16907), .A2(n19155), .B1(n20200), .B2(n16908), .ZN(
        U374) );
  INV_X1 U20063 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19153) );
  INV_X1 U20064 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20199) );
  AOI22_X1 U20065 ( .A1(n16907), .A2(n19153), .B1(n20199), .B2(n16908), .ZN(
        U375) );
  INV_X1 U20066 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19133) );
  INV_X1 U20067 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20185) );
  AOI22_X1 U20068 ( .A1(n16907), .A2(n19133), .B1(n20185), .B2(n16908), .ZN(
        U376) );
  INV_X1 U20069 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19132) );
  NAND2_X1 U20070 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19132), .ZN(n19118) );
  AOI22_X1 U20071 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19118), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19130), .ZN(n19203) );
  AOI21_X1 U20072 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19203), .ZN(n16909) );
  INV_X1 U20073 ( .A(n16909), .ZN(P3_U2633) );
  NAND2_X1 U20074 ( .A1(n19251), .A2(n19039), .ZN(n17839) );
  OAI21_X1 U20075 ( .B1(n16917), .B2(n17839), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16910) );
  OAI21_X1 U20076 ( .B1(n16911), .B2(n19105), .A(n16910), .ZN(P3_U2634) );
  AOI21_X1 U20077 ( .B1(n19130), .B2(n19132), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16912) );
  AOI22_X1 U20078 ( .A1(n19265), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16912), 
        .B2(n19266), .ZN(P3_U2635) );
  NOR2_X1 U20079 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16913) );
  OAI21_X1 U20080 ( .B1(n16913), .B2(BS16), .A(n19203), .ZN(n19201) );
  OAI21_X1 U20081 ( .B1(n19203), .B2(n19255), .A(n19201), .ZN(P3_U2636) );
  INV_X1 U20082 ( .A(n16914), .ZN(n16916) );
  NOR3_X1 U20083 ( .A1(n16917), .A2(n16916), .A3(n16915), .ZN(n19042) );
  NOR2_X1 U20084 ( .A1(n19042), .A2(n19100), .ZN(n19247) );
  OAI21_X1 U20085 ( .B1(n19247), .B2(n18598), .A(n16918), .ZN(P3_U2637) );
  NOR4_X1 U20086 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16922) );
  NOR4_X1 U20087 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16921) );
  NOR4_X1 U20088 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16920) );
  NOR4_X1 U20089 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16919) );
  NAND4_X1 U20090 ( .A1(n16922), .A2(n16921), .A3(n16920), .A4(n16919), .ZN(
        n16928) );
  NOR4_X1 U20091 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16926) );
  AOI211_X1 U20092 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16925) );
  NOR4_X1 U20093 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16924) );
  NOR4_X1 U20094 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16923) );
  NAND4_X1 U20095 ( .A1(n16926), .A2(n16925), .A3(n16924), .A4(n16923), .ZN(
        n16927) );
  NOR2_X1 U20096 ( .A1(n16928), .A2(n16927), .ZN(n19241) );
  INV_X1 U20097 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16930) );
  NOR3_X1 U20098 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16931) );
  OAI21_X1 U20099 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16931), .A(n19241), .ZN(
        n16929) );
  OAI21_X1 U20100 ( .B1(n19241), .B2(n16930), .A(n16929), .ZN(P3_U2638) );
  INV_X1 U20101 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19237) );
  INV_X1 U20102 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19202) );
  AOI21_X1 U20103 ( .B1(n19237), .B2(n19202), .A(n16931), .ZN(n16933) );
  INV_X1 U20104 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16932) );
  INV_X1 U20105 ( .A(n19241), .ZN(n19244) );
  AOI22_X1 U20106 ( .A1(n19241), .A2(n16933), .B1(n16932), .B2(n19244), .ZN(
        P3_U2639) );
  AOI21_X1 U20107 ( .B1(n17892), .B2(n16935), .A(n16934), .ZN(n17902) );
  OAI21_X1 U20108 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16936), .A(
        n16935), .ZN(n17909) );
  INV_X1 U20109 ( .A(n17909), .ZN(n16995) );
  AOI21_X1 U20110 ( .B1(n17014), .B2(n17896), .A(n16936), .ZN(n17927) );
  INV_X1 U20111 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17933) );
  INV_X1 U20112 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17944) );
  NOR2_X1 U20113 ( .A1(n18249), .A2(n17960), .ZN(n17931) );
  NAND2_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17931), .ZN(
        n16939) );
  OR2_X1 U20115 ( .A1(n17944), .A2(n16939), .ZN(n16938) );
  AOI21_X1 U20116 ( .B1(n17933), .B2(n16938), .A(n16937), .ZN(n17936) );
  XOR2_X1 U20117 ( .A(n17944), .B(n16939), .Z(n17947) );
  OAI21_X1 U20118 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17931), .A(
        n16939), .ZN(n16940) );
  INV_X1 U20119 ( .A(n16940), .ZN(n17957) );
  INV_X1 U20120 ( .A(n16941), .ZN(n18008) );
  NOR2_X1 U20121 ( .A1(n18249), .A2(n18008), .ZN(n18007) );
  NAND3_X1 U20122 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n18007), .ZN(n17967) );
  NOR2_X1 U20123 ( .A1(n17992), .A2(n17967), .ZN(n16943) );
  NAND2_X1 U20124 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16943), .ZN(
        n16942) );
  AOI21_X1 U20125 ( .B1(n10083), .B2(n16942), .A(n17931), .ZN(n17972) );
  XOR2_X1 U20126 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16943), .Z(
        n17989) );
  AOI21_X1 U20127 ( .B1(n17992), .B2(n17967), .A(n16943), .ZN(n17996) );
  INV_X1 U20128 ( .A(n17967), .ZN(n16944) );
  INV_X1 U20129 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18057) );
  NAND2_X1 U20130 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18041), .ZN(
        n18042) );
  NOR2_X1 U20131 ( .A1(n18057), .A2(n18042), .ZN(n17121) );
  INV_X1 U20132 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17307) );
  NAND2_X1 U20133 ( .A1(n17121), .A2(n17307), .ZN(n17087) );
  NAND2_X1 U20134 ( .A1(n17271), .A2(n17087), .ZN(n17122) );
  OAI21_X1 U20135 ( .B1(n16944), .B2(n9731), .A(n17122), .ZN(n17068) );
  NOR2_X1 U20136 ( .A1(n17996), .A2(n17068), .ZN(n17067) );
  NOR2_X1 U20137 ( .A1(n17067), .A2(n9731), .ZN(n17057) );
  NOR2_X1 U20138 ( .A1(n17989), .A2(n17057), .ZN(n17056) );
  NOR2_X1 U20139 ( .A1(n17035), .A2(n9731), .ZN(n17029) );
  NOR2_X1 U20140 ( .A1(n17947), .A2(n17029), .ZN(n17028) );
  NOR2_X1 U20141 ( .A1(n17028), .A2(n9731), .ZN(n17017) );
  NOR2_X1 U20142 ( .A1(n17936), .A2(n17017), .ZN(n17016) );
  NOR2_X1 U20143 ( .A1(n17016), .A2(n9731), .ZN(n17008) );
  NOR2_X1 U20144 ( .A1(n17927), .A2(n17008), .ZN(n17007) );
  NOR2_X1 U20145 ( .A1(n17007), .A2(n9731), .ZN(n16994) );
  NOR2_X1 U20146 ( .A1(n16995), .A2(n16994), .ZN(n16993) );
  NOR2_X1 U20147 ( .A1(n16993), .A2(n9731), .ZN(n16986) );
  NAND2_X1 U20148 ( .A1(n16962), .A2(n16963), .ZN(n16960) );
  NAND4_X1 U20149 ( .A1(n19268), .A2(n19102), .A3(n19255), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17223) );
  INV_X1 U20150 ( .A(n17223), .ZN(n17278) );
  NAND2_X1 U20151 ( .A1(n17271), .A2(n17278), .ZN(n17306) );
  INV_X1 U20152 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16950) );
  NOR2_X1 U20153 ( .A1(n16950), .A2(n19256), .ZN(n16947) );
  OAI211_X2 U20154 ( .C1(P3_STATEBS16_REG_SCAN_IN), .C2(n19122), .A(n16949), 
        .B(n16947), .ZN(n17314) );
  NOR3_X1 U20155 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17291) );
  NAND2_X1 U20156 ( .A1(n17291), .A2(n17281), .ZN(n17279) );
  NOR2_X1 U20157 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17279), .ZN(n17256) );
  NAND2_X1 U20158 ( .A1(n17256), .A2(n17252), .ZN(n17251) );
  NAND2_X1 U20159 ( .A1(n17236), .A2(n17216), .ZN(n17218) );
  NAND2_X1 U20160 ( .A1(n17210), .A2(n17550), .ZN(n17198) );
  INV_X1 U20161 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17533) );
  NAND2_X1 U20162 ( .A1(n17180), .A2(n17533), .ZN(n17176) );
  NAND2_X1 U20163 ( .A1(n17160), .A2(n17504), .ZN(n17152) );
  INV_X1 U20164 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17478) );
  NAND2_X1 U20165 ( .A1(n17132), .A2(n17478), .ZN(n17128) );
  INV_X1 U20166 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17104) );
  NAND2_X1 U20167 ( .A1(n17113), .A2(n17104), .ZN(n17102) );
  NAND2_X1 U20168 ( .A1(n17093), .A2(n17424), .ZN(n17081) );
  INV_X1 U20169 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17408) );
  NAND2_X1 U20170 ( .A1(n17064), .A2(n17408), .ZN(n17060) );
  NAND2_X1 U20171 ( .A1(n17049), .A2(n17043), .ZN(n17042) );
  NOR2_X1 U20172 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17042), .ZN(n17015) );
  NAND2_X1 U20173 ( .A1(n17015), .A2(n17362), .ZN(n17006) );
  NOR2_X1 U20174 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17006), .ZN(n17005) );
  INV_X1 U20175 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17356) );
  NAND2_X1 U20176 ( .A1(n17005), .A2(n17356), .ZN(n16999) );
  NOR2_X1 U20177 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16999), .ZN(n16984) );
  NAND2_X1 U20178 ( .A1(n16984), .A2(n17351), .ZN(n16961) );
  NOR2_X1 U20179 ( .A1(n17314), .A2(n16961), .ZN(n16969) );
  INV_X1 U20180 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16954) );
  AOI211_X1 U20181 ( .C1(n19256), .C2(n19254), .A(n19122), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16948) );
  INV_X1 U20182 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19181) );
  INV_X1 U20183 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19176) );
  INV_X1 U20184 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19171) );
  INV_X1 U20185 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19156) );
  INV_X1 U20186 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19138) );
  NAND3_X1 U20187 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17263) );
  NOR2_X1 U20188 ( .A1(n19138), .A2(n17263), .ZN(n17245) );
  NAND2_X1 U20189 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17245), .ZN(n17169) );
  INV_X1 U20190 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19147) );
  NAND2_X1 U20191 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17205) );
  NOR2_X1 U20192 ( .A1(n19147), .A2(n17205), .ZN(n17168) );
  NAND4_X1 U20193 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17168), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17148) );
  NOR2_X1 U20194 ( .A1(n17169), .A2(n17148), .ZN(n17162) );
  NAND2_X1 U20195 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17162), .ZN(n17143) );
  NOR2_X1 U20196 ( .A1(n19156), .A2(n17143), .ZN(n17133) );
  NAND2_X1 U20197 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17133), .ZN(n17106) );
  INV_X1 U20198 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19166) );
  NAND3_X1 U20199 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17085) );
  NOR2_X1 U20200 ( .A1(n19166), .A2(n17085), .ZN(n17074) );
  NAND2_X1 U20201 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17074), .ZN(n17066) );
  NOR3_X1 U20202 ( .A1(n19171), .A2(n17106), .A3(n17066), .ZN(n17048) );
  NAND3_X1 U20203 ( .A1(n17048), .A2(P3_REIP_REG_22__SCAN_IN), .A3(
        P3_REIP_REG_21__SCAN_IN), .ZN(n17039) );
  NOR2_X1 U20204 ( .A1(n19176), .A2(n17039), .ZN(n17037) );
  NAND2_X1 U20205 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17037), .ZN(n17018) );
  NOR2_X1 U20206 ( .A1(n19181), .A2(n17018), .ZN(n17004) );
  NAND2_X1 U20207 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17004), .ZN(n16956) );
  NOR2_X1 U20208 ( .A1(n17308), .A2(n16956), .ZN(n16983) );
  NAND4_X1 U20209 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16983), .ZN(n16955) );
  NOR3_X1 U20210 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19194), .A3(n16955), 
        .ZN(n16953) );
  INV_X1 U20211 ( .A(n17278), .ZN(n19109) );
  NAND2_X1 U20212 ( .A1(n19268), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18975) );
  OR2_X1 U20213 ( .A1(n19105), .A2(n18975), .ZN(n19098) );
  INV_X1 U20214 ( .A(n16948), .ZN(n19093) );
  OAI211_X2 U20215 ( .C1(n16950), .C2(n19256), .A(n19093), .B(n16949), .ZN(
        n17315) );
  OAI22_X1 U20216 ( .A1(n16951), .A2(n17305), .B1(n16950), .B2(n17315), .ZN(
        n16952) );
  AOI211_X1 U20217 ( .C1(n16969), .C2(n16954), .A(n16953), .B(n16952), .ZN(
        n16959) );
  NOR2_X1 U20218 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16955), .ZN(n16967) );
  NAND3_X1 U20219 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16957) );
  AND2_X1 U20220 ( .A1(n17294), .A2(n16956), .ZN(n17003) );
  NOR2_X1 U20221 ( .A1(n17255), .A2(n17003), .ZN(n17002) );
  INV_X1 U20222 ( .A(n17002), .ZN(n17011) );
  AOI21_X1 U20223 ( .B1(n17294), .B2(n16957), .A(n17011), .ZN(n16965) );
  INV_X1 U20224 ( .A(n16965), .ZN(n16979) );
  OAI21_X1 U20225 ( .B1(n16967), .B2(n16979), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16958) );
  OAI211_X1 U20226 ( .C1(n16960), .C2(n17306), .A(n16959), .B(n16958), .ZN(
        P3_U2640) );
  NAND2_X1 U20227 ( .A1(n17280), .A2(n16961), .ZN(n16972) );
  XOR2_X1 U20228 ( .A(n16963), .B(n16962), .Z(n16968) );
  OAI22_X1 U20229 ( .A1(n16965), .A2(n19194), .B1(n16964), .B2(n17305), .ZN(
        n16966) );
  OAI21_X1 U20230 ( .B1(n17285), .B2(n16969), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16970) );
  NAND3_X1 U20231 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16983), .ZN(n16982) );
  AOI22_X1 U20232 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17286), .B1(
        n17285), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16981) );
  INV_X1 U20233 ( .A(n16984), .ZN(n16973) );
  AOI21_X1 U20234 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16973), .A(n16972), .ZN(
        n16978) );
  AOI211_X1 U20235 ( .C1(n16976), .C2(n16975), .A(n16974), .B(n19109), .ZN(
        n16977) );
  AOI211_X1 U20236 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16979), .A(n16978), 
        .B(n16977), .ZN(n16980) );
  OAI211_X1 U20237 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16982), .A(n16981), 
        .B(n16980), .ZN(P3_U2642) );
  NAND2_X1 U20238 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16983), .ZN(n16992) );
  AOI22_X1 U20239 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17286), .B1(
        n17285), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16991) );
  INV_X1 U20240 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19185) );
  NAND2_X1 U20241 ( .A1(n16983), .A2(n19185), .ZN(n16996) );
  NAND2_X1 U20242 ( .A1(n17002), .A2(n16996), .ZN(n16989) );
  AOI211_X1 U20243 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16999), .A(n16984), .B(
        n17314), .ZN(n16988) );
  AOI211_X1 U20244 ( .C1(n17902), .C2(n16986), .A(n16985), .B(n19109), .ZN(
        n16987) );
  AOI211_X1 U20245 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16989), .A(n16988), 
        .B(n16987), .ZN(n16990) );
  OAI211_X1 U20246 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16992), .A(n16991), 
        .B(n16990), .ZN(P3_U2643) );
  AOI211_X1 U20247 ( .C1(n16995), .C2(n16994), .A(n16993), .B(n19109), .ZN(
        n16998) );
  OAI21_X1 U20248 ( .B1(n17356), .B2(n17315), .A(n16996), .ZN(n16997) );
  AOI211_X1 U20249 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16998), .B(n16997), .ZN(n17001) );
  OAI211_X1 U20250 ( .C1(n17005), .C2(n17356), .A(n17280), .B(n16999), .ZN(
        n17000) );
  OAI211_X1 U20251 ( .C1(n17002), .C2(n19185), .A(n17001), .B(n17000), .ZN(
        P3_U2644) );
  AOI22_X1 U20252 ( .A1(n17285), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n17004), 
        .B2(n17003), .ZN(n17013) );
  AOI211_X1 U20253 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17006), .A(n17005), .B(
        n17314), .ZN(n17010) );
  AOI211_X1 U20254 ( .C1(n17927), .C2(n17008), .A(n17007), .B(n19109), .ZN(
        n17009) );
  AOI211_X1 U20255 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17011), .A(n17010), 
        .B(n17009), .ZN(n17012) );
  OAI211_X1 U20256 ( .C1(n17014), .C2(n17305), .A(n17013), .B(n17012), .ZN(
        P3_U2645) );
  OR2_X1 U20257 ( .A1(n17314), .A2(n17015), .ZN(n17027) );
  AOI21_X1 U20258 ( .B1(n17280), .B2(n17015), .A(n17285), .ZN(n17025) );
  AOI211_X1 U20259 ( .C1(n17936), .C2(n17017), .A(n17016), .B(n17223), .ZN(
        n17023) );
  NOR2_X1 U20260 ( .A1(n17308), .A2(n17018), .ZN(n17021) );
  INV_X1 U20261 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19178) );
  OAI21_X1 U20262 ( .B1(n17037), .B2(n17308), .A(n17318), .ZN(n17034) );
  AOI21_X1 U20263 ( .B1(n17294), .B2(n19178), .A(n17034), .ZN(n17019) );
  INV_X1 U20264 ( .A(n17019), .ZN(n17020) );
  MUX2_X1 U20265 ( .A(n17021), .B(n17020), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n17022) );
  AOI211_X1 U20266 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17023), .B(n17022), .ZN(n17024) );
  OAI221_X1 U20267 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17027), .C1(n17362), 
        .C2(n17025), .A(n17024), .ZN(P3_U2646) );
  NOR2_X1 U20268 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17308), .ZN(n17026) );
  AOI22_X1 U20269 ( .A1(n17285), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17037), 
        .B2(n17026), .ZN(n17033) );
  AOI21_X1 U20270 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17042), .A(n17027), .ZN(
        n17031) );
  AOI211_X1 U20271 ( .C1(n17947), .C2(n17029), .A(n17028), .B(n17223), .ZN(
        n17030) );
  AOI211_X1 U20272 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17034), .A(n17031), 
        .B(n17030), .ZN(n17032) );
  OAI211_X1 U20273 ( .C1(n17944), .C2(n17305), .A(n17033), .B(n17032), .ZN(
        P3_U2647) );
  INV_X1 U20274 ( .A(n17034), .ZN(n17046) );
  AOI211_X1 U20275 ( .C1(n17957), .C2(n17036), .A(n17035), .B(n17223), .ZN(
        n17041) );
  OR2_X1 U20276 ( .A1(n17308), .A2(n17037), .ZN(n17038) );
  OAI22_X1 U20277 ( .A1(n17315), .A2(n17043), .B1(n17039), .B2(n17038), .ZN(
        n17040) );
  AOI211_X1 U20278 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17041), .B(n17040), .ZN(n17045) );
  OAI211_X1 U20279 ( .C1(n17049), .C2(n17043), .A(n17280), .B(n17042), .ZN(
        n17044) );
  OAI211_X1 U20280 ( .C1(n17046), .C2(n19176), .A(n17045), .B(n17044), .ZN(
        P3_U2648) );
  INV_X1 U20281 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19174) );
  INV_X1 U20282 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19172) );
  NAND2_X1 U20283 ( .A1(n17294), .A2(n17048), .ZN(n17063) );
  AOI221_X1 U20284 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n19174), .C2(n19172), .A(n17063), .ZN(n17047) );
  AOI21_X1 U20285 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17285), .A(n17047), .ZN(
        n17055) );
  OAI21_X1 U20286 ( .B1(n17048), .B2(n17308), .A(n17318), .ZN(n17071) );
  AOI211_X1 U20287 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17060), .A(n17049), .B(
        n17314), .ZN(n17053) );
  AOI211_X1 U20288 ( .C1(n17972), .C2(n17051), .A(n17050), .B(n17223), .ZN(
        n17052) );
  AOI211_X1 U20289 ( .C1(n17071), .C2(P3_REIP_REG_22__SCAN_IN), .A(n17053), 
        .B(n17052), .ZN(n17054) );
  OAI211_X1 U20290 ( .C1(n10083), .C2(n17305), .A(n17055), .B(n17054), .ZN(
        P3_U2649) );
  AOI211_X1 U20291 ( .C1(n17989), .C2(n17057), .A(n17056), .B(n17223), .ZN(
        n17059) );
  OAI22_X1 U20292 ( .A1(n10082), .A2(n17305), .B1(n17315), .B2(n17408), .ZN(
        n17058) );
  AOI211_X1 U20293 ( .C1(n17071), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17059), 
        .B(n17058), .ZN(n17062) );
  OAI211_X1 U20294 ( .C1(n17064), .C2(n17408), .A(n17280), .B(n17060), .ZN(
        n17061) );
  OAI211_X1 U20295 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17063), .A(n17062), 
        .B(n17061), .ZN(P3_U2650) );
  AOI211_X1 U20296 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17081), .A(n17064), .B(
        n17314), .ZN(n17065) );
  AOI21_X1 U20297 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17285), .A(n17065), .ZN(
        n17073) );
  NAND3_X1 U20298 ( .A1(n17294), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n17133), 
        .ZN(n17123) );
  NOR2_X1 U20299 ( .A1(n17066), .A2(n17123), .ZN(n17070) );
  AOI211_X1 U20300 ( .C1(n17996), .C2(n17068), .A(n17067), .B(n19109), .ZN(
        n17069) );
  AOI221_X1 U20301 ( .B1(n17071), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n17070), 
        .C2(n19171), .A(n17069), .ZN(n17072) );
  OAI211_X1 U20302 ( .C1(n17992), .C2(n17305), .A(n17073), .B(n17072), .ZN(
        P3_U2651) );
  AOI22_X1 U20303 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17286), .B1(
        n17285), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17084) );
  INV_X1 U20304 ( .A(n17074), .ZN(n17076) );
  NAND2_X1 U20305 ( .A1(n17318), .A2(n17308), .ZN(n17316) );
  AOI21_X1 U20306 ( .B1(n17294), .B2(n17106), .A(n17255), .ZN(n17138) );
  INV_X1 U20307 ( .A(n17138), .ZN(n17127) );
  AOI21_X1 U20308 ( .B1(n17076), .B2(n17316), .A(n17127), .ZN(n17075) );
  INV_X1 U20309 ( .A(n17075), .ZN(n17097) );
  NOR3_X1 U20310 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17076), .A3(n17123), 
        .ZN(n17080) );
  NAND2_X1 U20311 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18007), .ZN(
        n17086) );
  OAI21_X1 U20312 ( .B1(n17087), .B2(n17086), .A(n17271), .ZN(n17090) );
  INV_X1 U20313 ( .A(n17086), .ZN(n17077) );
  OAI21_X1 U20314 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17077), .A(
        n17967), .ZN(n18013) );
  OAI21_X1 U20315 ( .B1(n17090), .B2(n18013), .A(n17278), .ZN(n17078) );
  AOI21_X1 U20316 ( .B1(n17090), .B2(n18013), .A(n17078), .ZN(n17079) );
  AOI211_X1 U20317 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17097), .A(n17080), 
        .B(n17079), .ZN(n17083) );
  OAI211_X1 U20318 ( .C1(n17093), .C2(n17424), .A(n17280), .B(n17081), .ZN(
        n17082) );
  NAND4_X1 U20319 ( .A1(n17084), .A2(n17083), .A3(n18491), .A4(n17082), .ZN(
        P3_U2652) );
  INV_X1 U20320 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17099) );
  OAI21_X1 U20321 ( .B1(n17085), .B2(n17123), .A(n19166), .ZN(n17096) );
  OAI21_X1 U20322 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18007), .A(
        n17086), .ZN(n18019) );
  NOR2_X1 U20323 ( .A1(n19109), .A2(n17271), .ZN(n17225) );
  INV_X1 U20324 ( .A(n17225), .ZN(n17301) );
  NOR2_X1 U20325 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17087), .ZN(
        n17088) );
  OAI21_X1 U20326 ( .B1(n17088), .B2(n18019), .A(n17278), .ZN(n17089) );
  AOI22_X1 U20327 ( .A1(n17090), .A2(n18019), .B1(n17301), .B2(n17089), .ZN(
        n17095) );
  AOI21_X1 U20328 ( .B1(n17102), .B2(P3_EBX_REG_18__SCAN_IN), .A(n17314), .ZN(
        n17091) );
  INV_X1 U20329 ( .A(n17091), .ZN(n17092) );
  INV_X1 U20330 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18022) );
  OAI22_X1 U20331 ( .A1(n17093), .A2(n17092), .B1(n18022), .B2(n17305), .ZN(
        n17094) );
  AOI211_X1 U20332 ( .C1(n17097), .C2(n17096), .A(n17095), .B(n17094), .ZN(
        n17098) );
  OAI211_X1 U20333 ( .C1(n17315), .C2(n17099), .A(n17098), .B(n18591), .ZN(
        P3_U2653) );
  OR2_X1 U20334 ( .A1(n18249), .A2(n18031), .ZN(n17100) );
  OAI21_X1 U20335 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17121), .A(
        n17100), .ZN(n18043) );
  AOI21_X1 U20336 ( .B1(n17122), .B2(n18043), .A(n9731), .ZN(n17101) );
  AOI21_X1 U20337 ( .B1(n18032), .B2(n17100), .A(n18007), .ZN(n18034) );
  XNOR2_X1 U20338 ( .A(n17101), .B(n18034), .ZN(n17112) );
  OAI211_X1 U20339 ( .C1(n17113), .C2(n17104), .A(n17280), .B(n17102), .ZN(
        n17103) );
  OAI211_X1 U20340 ( .C1(n17315), .C2(n17104), .A(n18491), .B(n17103), .ZN(
        n17110) );
  NAND2_X1 U20341 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17105) );
  NOR2_X1 U20342 ( .A1(n17105), .A2(n17123), .ZN(n17108) );
  AOI221_X1 U20343 ( .B1(n17106), .B2(n17294), .C1(n17105), .C2(n17294), .A(
        n17255), .ZN(n17120) );
  INV_X1 U20344 ( .A(n17120), .ZN(n17107) );
  MUX2_X1 U20345 ( .A(n17108), .B(n17107), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n17109) );
  AOI211_X1 U20346 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n17286), .A(
        n17110), .B(n17109), .ZN(n17111) );
  OAI21_X1 U20347 ( .B1(n19109), .B2(n17112), .A(n17111), .ZN(P3_U2654) );
  INV_X1 U20348 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19162) );
  INV_X1 U20349 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19160) );
  NOR3_X1 U20350 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19160), .A3(n17123), 
        .ZN(n17116) );
  AOI211_X1 U20351 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17128), .A(n17113), .B(
        n17314), .ZN(n17115) );
  INV_X1 U20352 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18045) );
  OAI22_X1 U20353 ( .A1(n18045), .A2(n17305), .B1(n17315), .B2(n17479), .ZN(
        n17114) );
  NOR4_X1 U20354 ( .A1(n18570), .A2(n17116), .A3(n17115), .A4(n17114), .ZN(
        n17119) );
  NAND2_X1 U20355 ( .A1(n17122), .A2(n18043), .ZN(n17117) );
  OAI211_X1 U20356 ( .C1(n17122), .C2(n18043), .A(n17278), .B(n17117), .ZN(
        n17118) );
  OAI211_X1 U20357 ( .C1(n17120), .C2(n19162), .A(n17119), .B(n17118), .ZN(
        P3_U2655) );
  AOI22_X1 U20358 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17286), .B1(
        n17285), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17131) );
  AOI21_X1 U20359 ( .B1(n18057), .B2(n18042), .A(n17121), .ZN(n18060) );
  NOR3_X1 U20360 ( .A1(n18060), .A2(n17122), .A3(n17223), .ZN(n17126) );
  AOI21_X1 U20361 ( .B1(n17271), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17223), .ZN(n17310) );
  INV_X1 U20362 ( .A(n17310), .ZN(n17149) );
  OAI21_X1 U20363 ( .B1(n18057), .B2(n9731), .A(n18060), .ZN(n17124) );
  OAI22_X1 U20364 ( .A1(n17149), .A2(n17124), .B1(P3_REIP_REG_15__SCAN_IN), 
        .B2(n17123), .ZN(n17125) );
  AOI211_X1 U20365 ( .C1(n17127), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17126), 
        .B(n17125), .ZN(n17130) );
  OAI211_X1 U20366 ( .C1(n17132), .C2(n17478), .A(n17280), .B(n17128), .ZN(
        n17129) );
  NAND4_X1 U20367 ( .A1(n17131), .A2(n17130), .A3(n18491), .A4(n17129), .ZN(
        P3_U2656) );
  INV_X1 U20368 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17477) );
  AOI211_X1 U20369 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17152), .A(n17132), .B(
        n17314), .ZN(n17141) );
  AOI21_X1 U20370 ( .B1(n17294), .B2(n17133), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n17139) );
  NOR2_X1 U20371 ( .A1(n18249), .A2(n18171), .ZN(n17208) );
  INV_X1 U20372 ( .A(n17208), .ZN(n17233) );
  NOR2_X1 U20373 ( .A1(n17134), .A2(n17233), .ZN(n17170) );
  INV_X1 U20374 ( .A(n17170), .ZN(n18091) );
  NOR3_X1 U20375 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17135), .A3(
        n18091), .ZN(n17146) );
  NOR2_X1 U20376 ( .A1(n17146), .A2(n9731), .ZN(n17136) );
  NOR2_X1 U20377 ( .A1(n17135), .A2(n18091), .ZN(n17145) );
  OAI21_X1 U20378 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17145), .A(
        n18042), .ZN(n18088) );
  XOR2_X1 U20379 ( .A(n17136), .B(n18088), .Z(n17137) );
  OAI22_X1 U20380 ( .A1(n17139), .A2(n17138), .B1(n19109), .B2(n17137), .ZN(
        n17140) );
  AOI211_X1 U20381 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17141), .B(n17140), .ZN(n17142) );
  OAI211_X1 U20382 ( .C1(n17315), .C2(n17477), .A(n17142), .B(n18591), .ZN(
        P3_U2657) );
  NOR3_X1 U20383 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17308), .A3(n17143), 
        .ZN(n17144) );
  AOI211_X1 U20384 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17286), .A(
        n18570), .B(n17144), .ZN(n17156) );
  INV_X1 U20385 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18093) );
  NAND2_X1 U20386 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17170), .ZN(
        n17157) );
  AOI21_X1 U20387 ( .B1(n18093), .B2(n17157), .A(n17145), .ZN(n18098) );
  NOR3_X1 U20388 ( .A1(n18098), .A2(n17146), .A3(n17306), .ZN(n17147) );
  AOI21_X1 U20389 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17285), .A(n17147), .ZN(
        n17155) );
  OR2_X1 U20390 ( .A1(n17169), .A2(n17255), .ZN(n17227) );
  OAI21_X1 U20391 ( .B1(n17148), .B2(n17227), .A(n17316), .ZN(n17173) );
  OAI21_X1 U20392 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17308), .A(n17173), 
        .ZN(n17151) );
  AOI21_X1 U20393 ( .B1(n17157), .B2(n17301), .A(n17149), .ZN(n17150) );
  AOI22_X1 U20394 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17151), .B1(n18098), 
        .B2(n17150), .ZN(n17154) );
  OAI211_X1 U20395 ( .C1(n17160), .C2(n17504), .A(n17280), .B(n17152), .ZN(
        n17153) );
  NAND4_X1 U20396 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        P3_U2658) );
  OAI21_X1 U20397 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18091), .A(
        n17271), .ZN(n17159) );
  OAI21_X1 U20398 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17170), .A(
        n17157), .ZN(n17158) );
  INV_X1 U20399 ( .A(n17158), .ZN(n18114) );
  XOR2_X1 U20400 ( .A(n17159), .B(n18114), .Z(n17167) );
  AOI211_X1 U20401 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17176), .A(n17160), .B(
        n17314), .ZN(n17165) );
  INV_X1 U20402 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19154) );
  NOR2_X1 U20403 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17308), .ZN(n17161) );
  AOI22_X1 U20404 ( .A1(n17285), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n17162), 
        .B2(n17161), .ZN(n17163) );
  OAI211_X1 U20405 ( .C1(n19154), .C2(n17173), .A(n17163), .B(n18591), .ZN(
        n17164) );
  AOI211_X1 U20406 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17165), .B(n17164), .ZN(n17166) );
  OAI21_X1 U20407 ( .B1(n17167), .B2(n17223), .A(n17166), .ZN(P3_U2659) );
  INV_X1 U20408 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17179) );
  INV_X1 U20409 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19150) );
  INV_X1 U20410 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19148) );
  NOR2_X1 U20411 ( .A1(n19150), .A2(n19148), .ZN(n17184) );
  INV_X1 U20412 ( .A(n17168), .ZN(n17182) );
  OR2_X1 U20413 ( .A1(n17308), .A2(n17169), .ZN(n17228) );
  NOR2_X1 U20414 ( .A1(n17182), .A2(n17228), .ZN(n17203) );
  AOI21_X1 U20415 ( .B1(n17184), .B2(n17203), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17174) );
  INV_X1 U20416 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18145) );
  NAND2_X1 U20417 ( .A1(n18157), .A2(n17208), .ZN(n17207) );
  NOR2_X1 U20418 ( .A1(n18145), .A2(n17207), .ZN(n17194) );
  NAND2_X1 U20419 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17194), .ZN(
        n17185) );
  AOI21_X1 U20420 ( .B1(n17179), .B2(n17185), .A(n17170), .ZN(n18123) );
  OAI21_X1 U20421 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17185), .A(
        n17271), .ZN(n17171) );
  XOR2_X1 U20422 ( .A(n18123), .B(n17171), .Z(n17172) );
  OAI22_X1 U20423 ( .A1(n17174), .A2(n17173), .B1(n19109), .B2(n17172), .ZN(
        n17175) );
  AOI211_X1 U20424 ( .C1(n17285), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18581), .B(
        n17175), .ZN(n17178) );
  OAI211_X1 U20425 ( .C1(n17180), .C2(n17533), .A(n17280), .B(n17176), .ZN(
        n17177) );
  OAI211_X1 U20426 ( .C1(n17305), .C2(n17179), .A(n17178), .B(n17177), .ZN(
        P3_U2660) );
  INV_X1 U20427 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17193) );
  AOI211_X1 U20428 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17198), .A(n17180), .B(
        n17314), .ZN(n17181) );
  AOI211_X1 U20429 ( .C1(n17285), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18570), .B(
        n17181), .ZN(n17192) );
  OAI21_X1 U20430 ( .B1(n17182), .B2(n17227), .A(n17316), .ZN(n17215) );
  INV_X1 U20431 ( .A(n17215), .ZN(n17190) );
  INV_X1 U20432 ( .A(n17203), .ZN(n17183) );
  AOI211_X1 U20433 ( .C1(n19150), .C2(n19148), .A(n17184), .B(n17183), .ZN(
        n17189) );
  OAI21_X1 U20434 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17194), .A(
        n17185), .ZN(n18131) );
  INV_X1 U20435 ( .A(n17194), .ZN(n17186) );
  OAI21_X1 U20436 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17186), .A(
        n17271), .ZN(n17195) );
  OAI21_X1 U20437 ( .B1(n18131), .B2(n17195), .A(n17278), .ZN(n17187) );
  AOI21_X1 U20438 ( .B1(n18131), .B2(n17195), .A(n17187), .ZN(n17188) );
  AOI211_X1 U20439 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n17190), .A(n17189), 
        .B(n17188), .ZN(n17191) );
  OAI211_X1 U20440 ( .C1(n17193), .C2(n17305), .A(n17192), .B(n17191), .ZN(
        P3_U2661) );
  AOI21_X1 U20441 ( .B1(n18145), .B2(n17207), .A(n17194), .ZN(n17196) );
  INV_X1 U20442 ( .A(n17196), .ZN(n18147) );
  AOI221_X1 U20443 ( .B1(n17196), .B2(n17271), .C1(n18147), .C2(n17195), .A(
        n17223), .ZN(n17202) );
  NOR3_X1 U20444 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19109), .A3(
        n17207), .ZN(n17197) );
  AOI221_X1 U20445 ( .B1(n17286), .B2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C1(
        n17197), .C2(n18145), .A(n18581), .ZN(n17200) );
  OAI211_X1 U20446 ( .C1(n17210), .C2(n17550), .A(n17280), .B(n17198), .ZN(
        n17199) );
  OAI211_X1 U20447 ( .C1(n17550), .C2(n17315), .A(n17200), .B(n17199), .ZN(
        n17201) );
  AOI211_X1 U20448 ( .C1(n17203), .C2(n19148), .A(n17202), .B(n17201), .ZN(
        n17204) );
  OAI21_X1 U20449 ( .B1(n19148), .B2(n17215), .A(n17204), .ZN(P3_U2662) );
  NOR3_X1 U20450 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17205), .A3(n17228), .ZN(
        n17206) );
  AOI211_X1 U20451 ( .C1(n17285), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18570), .B(
        n17206), .ZN(n17214) );
  INV_X1 U20452 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18174) );
  NOR2_X1 U20453 ( .A1(n18174), .A2(n17233), .ZN(n17221) );
  OAI21_X1 U20454 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17221), .A(
        n17207), .ZN(n18158) );
  NAND2_X1 U20455 ( .A1(n17208), .A2(n17307), .ZN(n17237) );
  OAI21_X1 U20456 ( .B1(n18174), .B2(n17237), .A(n17271), .ZN(n17222) );
  OAI21_X1 U20457 ( .B1(n18158), .B2(n17222), .A(n17278), .ZN(n17209) );
  AOI21_X1 U20458 ( .B1(n18158), .B2(n17222), .A(n17209), .ZN(n17212) );
  AOI211_X1 U20459 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17218), .A(n17210), .B(
        n17314), .ZN(n17211) );
  AOI211_X1 U20460 ( .C1(n17286), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17212), .B(n17211), .ZN(n17213) );
  OAI211_X1 U20461 ( .C1(n19147), .C2(n17215), .A(n17214), .B(n17213), .ZN(
        P3_U2663) );
  OAI21_X1 U20462 ( .B1(n17216), .B2(n17236), .A(n17280), .ZN(n17217) );
  INV_X1 U20463 ( .A(n17217), .ZN(n17219) );
  AOI22_X1 U20464 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17286), .B1(
        n17219), .B2(n17218), .ZN(n17232) );
  INV_X1 U20465 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19142) );
  NOR3_X1 U20466 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n19142), .A3(n17228), .ZN(
        n17220) );
  AOI211_X1 U20467 ( .C1(n17285), .C2(P3_EBX_REG_7__SCAN_IN), .A(n18570), .B(
        n17220), .ZN(n17231) );
  AOI21_X1 U20468 ( .B1(n18174), .B2(n17233), .A(n17221), .ZN(n18179) );
  INV_X1 U20469 ( .A(n17222), .ZN(n17226) );
  AOI21_X1 U20470 ( .B1(n18179), .B2(n17237), .A(n17223), .ZN(n17224) );
  OAI22_X1 U20471 ( .A1(n18179), .A2(n17226), .B1(n17225), .B2(n17224), .ZN(
        n17230) );
  NAND2_X1 U20472 ( .A1(n17316), .A2(n17227), .ZN(n17248) );
  INV_X1 U20473 ( .A(n17248), .ZN(n17241) );
  NOR2_X1 U20474 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17228), .ZN(n17235) );
  OAI21_X1 U20475 ( .B1(n17241), .B2(n17235), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n17229) );
  NAND4_X1 U20476 ( .A1(n17232), .A2(n17231), .A3(n17230), .A4(n17229), .ZN(
        P3_U2664) );
  AND2_X1 U20477 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18190), .ZN(
        n17246) );
  OAI21_X1 U20478 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17246), .A(
        n17233), .ZN(n18193) );
  OAI21_X1 U20479 ( .B1(n17246), .B2(n9731), .A(n17310), .ZN(n17244) );
  AOI211_X1 U20480 ( .C1(n17285), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18570), .B(
        n17235), .ZN(n17243) );
  AOI211_X1 U20481 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17251), .A(n17236), .B(
        n17314), .ZN(n17240) );
  NAND2_X1 U20482 ( .A1(n18193), .A2(n17237), .ZN(n17238) );
  OAI22_X1 U20483 ( .A1(n10091), .A2(n17305), .B1(n17306), .B2(n17238), .ZN(
        n17239) );
  AOI211_X1 U20484 ( .C1(n17241), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17240), .B(
        n17239), .ZN(n17242) );
  OAI211_X1 U20485 ( .C1(n18193), .C2(n17244), .A(n17243), .B(n17242), .ZN(
        P3_U2665) );
  AOI21_X1 U20486 ( .B1(n17294), .B2(n17245), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n17249) );
  OR2_X1 U20487 ( .A1(n18249), .A2(n18202), .ZN(n17260) );
  AOI21_X1 U20488 ( .B1(n18201), .B2(n17260), .A(n17246), .ZN(n18203) );
  OAI21_X1 U20489 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17260), .A(
        n17271), .ZN(n17261) );
  XOR2_X1 U20490 ( .A(n18203), .B(n17261), .Z(n17247) );
  OAI22_X1 U20491 ( .A1(n17249), .A2(n17248), .B1(n19109), .B2(n17247), .ZN(
        n17250) );
  AOI211_X1 U20492 ( .C1(n17285), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18581), .B(
        n17250), .ZN(n17254) );
  OAI211_X1 U20493 ( .C1(n17256), .C2(n17252), .A(n17280), .B(n17251), .ZN(
        n17253) );
  OAI211_X1 U20494 ( .C1(n17305), .C2(n18201), .A(n17254), .B(n17253), .ZN(
        P3_U2666) );
  AOI21_X1 U20495 ( .B1(n17294), .B2(n17263), .A(n17255), .ZN(n17273) );
  AOI211_X1 U20496 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17279), .A(n17256), .B(
        n17314), .ZN(n17259) );
  NOR2_X1 U20497 ( .A1(n18610), .A2(n19249), .ZN(n19273) );
  INV_X1 U20498 ( .A(n19273), .ZN(n17321) );
  INV_X1 U20499 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19045) );
  OAI221_X1 U20500 ( .B1(n17321), .B2(n17257), .C1(n17321), .C2(n19045), .A(
        n18591), .ZN(n17258) );
  AOI211_X1 U20501 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17285), .A(n17259), .B(
        n17258), .ZN(n17269) );
  AND2_X1 U20502 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18213), .ZN(
        n17270) );
  OAI21_X1 U20503 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17270), .A(
        n17260), .ZN(n18217) );
  INV_X1 U20504 ( .A(n18217), .ZN(n17262) );
  NAND2_X1 U20505 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17307), .ZN(
        n17289) );
  INV_X1 U20506 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17264) );
  NAND2_X1 U20507 ( .A1(n18213), .A2(n17264), .ZN(n18221) );
  OAI22_X1 U20508 ( .A1(n17262), .A2(n17261), .B1(n17289), .B2(n18221), .ZN(
        n17267) );
  NOR3_X1 U20509 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17308), .A3(n17263), .ZN(
        n17266) );
  OAI22_X1 U20510 ( .A1(n17264), .A2(n17305), .B1(n18217), .B2(n17301), .ZN(
        n17265) );
  AOI211_X1 U20511 ( .C1(n17278), .C2(n17267), .A(n17266), .B(n17265), .ZN(
        n17268) );
  OAI211_X1 U20512 ( .C1(n19138), .C2(n17273), .A(n17269), .B(n17268), .ZN(
        P3_U2667) );
  NAND2_X1 U20513 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19056), .ZN(
        n17287) );
  AOI21_X1 U20514 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17287), .A(
        n17466), .ZN(n19208) );
  NAND2_X1 U20515 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17284) );
  AOI21_X1 U20516 ( .B1(n17274), .B2(n17284), .A(n17270), .ZN(n18225) );
  OAI21_X1 U20517 ( .B1(n18236), .B2(n17289), .A(n17271), .ZN(n17272) );
  XNOR2_X1 U20518 ( .A(n18225), .B(n17272), .ZN(n17277) );
  INV_X1 U20519 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19136) );
  NAND2_X1 U20520 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17293) );
  AOI221_X1 U20521 ( .B1(n17308), .B2(n19136), .C1(n17293), .C2(n19136), .A(
        n17273), .ZN(n17276) );
  OAI22_X1 U20522 ( .A1(n17274), .A2(n17305), .B1(n17315), .B2(n17281), .ZN(
        n17275) );
  AOI211_X1 U20523 ( .C1(n17278), .C2(n17277), .A(n17276), .B(n17275), .ZN(
        n17283) );
  OAI211_X1 U20524 ( .C1(n17291), .C2(n17281), .A(n17280), .B(n17279), .ZN(
        n17282) );
  OAI211_X1 U20525 ( .C1(n19208), .C2(n17321), .A(n17283), .B(n17282), .ZN(
        P3_U2668) );
  OAI21_X1 U20526 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17284), .ZN(n18243) );
  AOI22_X1 U20527 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17286), .B1(
        n17285), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17300) );
  INV_X1 U20528 ( .A(n17287), .ZN(n19055) );
  AOI21_X1 U20529 ( .B1(n9868), .B2(n19065), .A(n19055), .ZN(n19219) );
  INV_X1 U20530 ( .A(n18243), .ZN(n17290) );
  NOR2_X1 U20531 ( .A1(n18236), .A2(n17289), .ZN(n17288) );
  AOI211_X1 U20532 ( .C1(n17290), .C2(n17289), .A(n17288), .B(n17306), .ZN(
        n17298) );
  INV_X1 U20533 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19134) );
  INV_X1 U20534 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17620) );
  INV_X1 U20535 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17614) );
  NAND2_X1 U20536 ( .A1(n17620), .A2(n17614), .ZN(n17303) );
  AOI211_X1 U20537 ( .C1(n17303), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17314), .B(
        n17291), .ZN(n17292) );
  INV_X1 U20538 ( .A(n17292), .ZN(n17296) );
  OAI211_X1 U20539 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17294), .B(n17293), .ZN(n17295) );
  OAI211_X1 U20540 ( .C1(n19134), .C2(n17318), .A(n17296), .B(n17295), .ZN(
        n17297) );
  AOI211_X1 U20541 ( .C1(n19273), .C2(n19219), .A(n17298), .B(n17297), .ZN(
        n17299) );
  OAI211_X1 U20542 ( .C1(n18243), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        P3_U2669) );
  NAND2_X1 U20543 ( .A1(n19065), .A2(n17302), .ZN(n19222) );
  OAI21_X1 U20544 ( .B1(n17614), .B2(n17620), .A(n17303), .ZN(n17616) );
  OAI22_X1 U20545 ( .A1(n17314), .A2(n17616), .B1(n17318), .B2(n19237), .ZN(
        n17304) );
  INV_X1 U20546 ( .A(n17304), .ZN(n17313) );
  OAI21_X1 U20547 ( .B1(n17307), .B2(n17306), .A(n17305), .ZN(n17311) );
  OAI22_X1 U20548 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17308), .B1(n17315), 
        .B2(n17614), .ZN(n17309) );
  AOI221_X1 U20549 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17311), .C1(
        n18249), .C2(n17310), .A(n17309), .ZN(n17312) );
  OAI211_X1 U20550 ( .C1(n19222), .C2(n17321), .A(n17313), .B(n17312), .ZN(
        P3_U2670) );
  NAND2_X1 U20551 ( .A1(n17315), .A2(n17314), .ZN(n17317) );
  AOI22_X1 U20552 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17317), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17316), .ZN(n17320) );
  NAND3_X1 U20553 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19212), .A3(
        n17318), .ZN(n17319) );
  OAI211_X1 U20554 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17321), .A(
        n17320), .B(n17319), .ZN(P3_U2671) );
  AOI22_X1 U20555 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20556 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20557 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20558 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17322) );
  NAND4_X1 U20559 ( .A1(n17325), .A2(n17324), .A3(n17323), .A4(n17322), .ZN(
        n17331) );
  AOI22_X1 U20560 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20561 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20562 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20563 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17326) );
  NAND4_X1 U20564 ( .A1(n17329), .A2(n17328), .A3(n17327), .A4(n17326), .ZN(
        n17330) );
  NOR2_X1 U20565 ( .A1(n17331), .A2(n17330), .ZN(n17343) );
  AOI22_X1 U20566 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20567 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17341) );
  AOI22_X1 U20568 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17332) );
  OAI21_X1 U20569 ( .B1(n17333), .B2(n17593), .A(n17332), .ZN(n17339) );
  AOI22_X1 U20570 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20571 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20572 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17335) );
  AOI22_X1 U20573 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17334) );
  NAND4_X1 U20574 ( .A1(n17337), .A2(n17336), .A3(n17335), .A4(n17334), .ZN(
        n17338) );
  AOI211_X1 U20575 ( .C1(n17567), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17339), .B(n17338), .ZN(n17340) );
  NAND3_X1 U20576 ( .A1(n17342), .A2(n17341), .A3(n17340), .ZN(n17348) );
  NAND2_X1 U20577 ( .A1(n17349), .A2(n17348), .ZN(n17347) );
  XNOR2_X1 U20578 ( .A(n17343), .B(n17347), .ZN(n17631) );
  NOR2_X1 U20579 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17344), .ZN(n17346) );
  OAI22_X1 U20580 ( .A1(n17631), .A2(n17596), .B1(n17346), .B2(n17345), .ZN(
        P3_U2673) );
  OAI21_X1 U20581 ( .B1(n17349), .B2(n17348), .A(n17347), .ZN(n17639) );
  OAI222_X1 U20582 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17357), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n17352), .C1(n17351), .C2(n17350), .ZN(
        n17353) );
  OAI21_X1 U20583 ( .B1(n17639), .B2(n17596), .A(n17353), .ZN(P3_U2674) );
  OAI21_X1 U20584 ( .B1(n17360), .B2(n17355), .A(n17354), .ZN(n17648) );
  AOI22_X1 U20585 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17358), .B1(n17357), 
        .B2(n17356), .ZN(n17359) );
  OAI21_X1 U20586 ( .B1(n17648), .B2(n17596), .A(n17359), .ZN(P3_U2676) );
  AOI21_X1 U20587 ( .B1(n17361), .B2(n17368), .A(n17360), .ZN(n17649) );
  NOR2_X1 U20588 ( .A1(n17362), .A2(n17367), .ZN(n17371) );
  AOI22_X1 U20589 ( .A1(n17649), .A2(n17618), .B1(n17371), .B2(n17363), .ZN(
        n17364) );
  OAI21_X1 U20590 ( .B1(n17366), .B2(n17365), .A(n17364), .ZN(P3_U2677) );
  INV_X1 U20591 ( .A(n17367), .ZN(n17376) );
  AOI21_X1 U20592 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17596), .A(n17376), .ZN(
        n17370) );
  OAI21_X1 U20593 ( .B1(n17372), .B2(n17369), .A(n17368), .ZN(n17658) );
  OAI22_X1 U20594 ( .A1(n17371), .A2(n17370), .B1(n17658), .B2(n17596), .ZN(
        P3_U2678) );
  AOI21_X1 U20595 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17596), .A(n17381), .ZN(
        n17375) );
  AOI21_X1 U20596 ( .B1(n17373), .B2(n17377), .A(n17372), .ZN(n17659) );
  INV_X1 U20597 ( .A(n17659), .ZN(n17374) );
  OAI22_X1 U20598 ( .A1(n17376), .A2(n17375), .B1(n17374), .B2(n17596), .ZN(
        P3_U2679) );
  NOR2_X1 U20599 ( .A1(n17383), .A2(n17382), .ZN(n17396) );
  AOI21_X1 U20600 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17596), .A(n17396), .ZN(
        n17380) );
  OAI21_X1 U20601 ( .B1(n17379), .B2(n17378), .A(n17377), .ZN(n17670) );
  OAI22_X1 U20602 ( .A1(n17381), .A2(n17380), .B1(n17670), .B2(n17596), .ZN(
        P3_U2680) );
  OAI21_X1 U20603 ( .B1(n17383), .B2(n17618), .A(n17382), .ZN(n17384) );
  INV_X1 U20604 ( .A(n17384), .ZN(n17395) );
  AOI22_X1 U20605 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20606 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20607 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20608 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17385) );
  NAND4_X1 U20609 ( .A1(n17388), .A2(n17387), .A3(n17386), .A4(n17385), .ZN(
        n17394) );
  AOI22_X1 U20610 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20611 ( .A1(n17552), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20612 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20613 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17389) );
  NAND4_X1 U20614 ( .A1(n17392), .A2(n17391), .A3(n17390), .A4(n17389), .ZN(
        n17393) );
  NOR2_X1 U20615 ( .A1(n17394), .A2(n17393), .ZN(n17672) );
  OAI22_X1 U20616 ( .A1(n17396), .A2(n17395), .B1(n17672), .B2(n17596), .ZN(
        P3_U2681) );
  AOI22_X1 U20617 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20618 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20619 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11489), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20620 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17397) );
  NAND4_X1 U20621 ( .A1(n17400), .A2(n17399), .A3(n17398), .A4(n17397), .ZN(
        n17406) );
  AOI22_X1 U20622 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20623 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11551), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U20624 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20625 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17401) );
  NAND4_X1 U20626 ( .A1(n17404), .A2(n17403), .A3(n17402), .A4(n17401), .ZN(
        n17405) );
  NOR2_X1 U20627 ( .A1(n17406), .A2(n17405), .ZN(n17680) );
  AND2_X1 U20628 ( .A1(n17596), .A2(n17407), .ZN(n17421) );
  AOI22_X1 U20629 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17421), .B1(n17409), 
        .B2(n17408), .ZN(n17410) );
  OAI21_X1 U20630 ( .B1(n17680), .B2(n17596), .A(n17410), .ZN(P3_U2682) );
  AOI22_X1 U20631 ( .A1(n11489), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11551), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20632 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20633 ( .A1(n17552), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20634 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17411) );
  NAND4_X1 U20635 ( .A1(n17414), .A2(n17413), .A3(n17412), .A4(n17411), .ZN(
        n17420) );
  AOI22_X1 U20636 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20637 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U20638 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17416) );
  AOI22_X1 U20639 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17415) );
  NAND4_X1 U20640 ( .A1(n17418), .A2(n17417), .A3(n17416), .A4(n17415), .ZN(
        n17419) );
  NOR2_X1 U20641 ( .A1(n17420), .A2(n17419), .ZN(n17684) );
  OAI21_X1 U20642 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17422), .A(n17421), .ZN(
        n17423) );
  OAI21_X1 U20643 ( .B1(n17684), .B2(n17596), .A(n17423), .ZN(P3_U2683) );
  AOI21_X1 U20644 ( .B1(n17424), .B2(n17448), .A(n17618), .ZN(n17425) );
  INV_X1 U20645 ( .A(n17425), .ZN(n17436) );
  AOI22_X1 U20646 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U20647 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20648 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20649 ( .A1(n11489), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11551), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17426) );
  NAND4_X1 U20650 ( .A1(n17429), .A2(n17428), .A3(n17427), .A4(n17426), .ZN(
        n17435) );
  AOI22_X1 U20651 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20652 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20653 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20654 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17430) );
  NAND4_X1 U20655 ( .A1(n17433), .A2(n17432), .A3(n17431), .A4(n17430), .ZN(
        n17434) );
  NOR2_X1 U20656 ( .A1(n17435), .A2(n17434), .ZN(n17689) );
  OAI22_X1 U20657 ( .A1(n17437), .A2(n17436), .B1(n17689), .B2(n17596), .ZN(
        P3_U2684) );
  AOI22_X1 U20658 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U20659 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20660 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20661 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9666), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17438) );
  NAND4_X1 U20662 ( .A1(n17441), .A2(n17440), .A3(n17439), .A4(n17438), .ZN(
        n17447) );
  AOI22_X1 U20663 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20664 ( .A1(n11489), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20665 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20666 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17442) );
  NAND4_X1 U20667 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17446) );
  NOR2_X1 U20668 ( .A1(n17447), .A2(n17446), .ZN(n17694) );
  OAI21_X1 U20669 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17449), .A(n17448), .ZN(
        n17450) );
  AOI22_X1 U20670 ( .A1(n17618), .A2(n17694), .B1(n17450), .B2(n17596), .ZN(
        P3_U2685) );
  AOI22_X1 U20671 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9666), .ZN(n17454) );
  AOI22_X1 U20672 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17552), .ZN(n17453) );
  AOI22_X1 U20673 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17574), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17553), .ZN(n17452) );
  AOI22_X1 U20674 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17451) );
  NAND4_X1 U20675 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17461) );
  AOI22_X1 U20676 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20677 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11489), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17537), .ZN(n17458) );
  AOI22_X1 U20678 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9651), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9653), .ZN(n17457) );
  AOI22_X1 U20679 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17455), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n11513), .ZN(n17456) );
  NAND4_X1 U20680 ( .A1(n17459), .A2(n17458), .A3(n17457), .A4(n17456), .ZN(
        n17460) );
  NOR2_X1 U20681 ( .A1(n17461), .A2(n17460), .ZN(n17700) );
  OAI211_X1 U20682 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17463), .A(n17617), .B(
        n17462), .ZN(n17465) );
  NAND2_X1 U20683 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17586), .ZN(n17464) );
  OAI211_X1 U20684 ( .C1(n17700), .C2(n17596), .A(n17465), .B(n17464), .ZN(
        P3_U2686) );
  AOI22_X1 U20685 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9666), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20686 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U20687 ( .A1(n11512), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20688 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11551), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17467) );
  NAND4_X1 U20689 ( .A1(n17470), .A2(n17469), .A3(n17468), .A4(n17467), .ZN(
        n17476) );
  AOI22_X1 U20690 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20691 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U20692 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20693 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17471) );
  NAND4_X1 U20694 ( .A1(n17474), .A2(n17473), .A3(n17472), .A4(n17471), .ZN(
        n17475) );
  NOR2_X1 U20695 ( .A1(n17476), .A2(n17475), .ZN(n17707) );
  NOR3_X1 U20696 ( .A1(n17477), .A2(n17504), .A3(n17519), .ZN(n17481) );
  INV_X1 U20697 ( .A(n17481), .ZN(n17505) );
  NOR2_X1 U20698 ( .A1(n17478), .A2(n17505), .ZN(n17493) );
  XOR2_X1 U20699 ( .A(n17479), .B(n17493), .Z(n17480) );
  AOI22_X1 U20700 ( .A1(n17618), .A2(n17707), .B1(n17480), .B2(n17596), .ZN(
        P3_U2687) );
  OAI21_X1 U20701 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17481), .A(n17596), .ZN(
        n17492) );
  AOI22_X1 U20702 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9651), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U20703 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20704 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20705 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17482) );
  NAND4_X1 U20706 ( .A1(n17485), .A2(n17484), .A3(n17483), .A4(n17482), .ZN(
        n17491) );
  AOI22_X1 U20707 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17489) );
  AOI22_X1 U20708 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20709 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U20710 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17486) );
  NAND4_X1 U20711 ( .A1(n17489), .A2(n17488), .A3(n17487), .A4(n17486), .ZN(
        n17490) );
  NOR2_X1 U20712 ( .A1(n17491), .A2(n17490), .ZN(n17711) );
  OAI22_X1 U20713 ( .A1(n17493), .A2(n17492), .B1(n17711), .B2(n17596), .ZN(
        P3_U2688) );
  AOI22_X1 U20714 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20715 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17502) );
  AOI22_X1 U20716 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20717 ( .B1(n17522), .B2(n17593), .A(n17494), .ZN(n17500) );
  AOI22_X1 U20718 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20719 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20720 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U20721 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17495) );
  NAND4_X1 U20722 ( .A1(n17498), .A2(n17497), .A3(n17496), .A4(n17495), .ZN(
        n17499) );
  AOI211_X1 U20723 ( .C1(n11487), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17500), .B(n17499), .ZN(n17501) );
  NAND3_X1 U20724 ( .A1(n17503), .A2(n17502), .A3(n17501), .ZN(n17713) );
  INV_X1 U20725 ( .A(n17713), .ZN(n17508) );
  NOR2_X1 U20726 ( .A1(n17504), .A2(n17519), .ZN(n17506) );
  OAI21_X1 U20727 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17506), .A(n17505), .ZN(
        n17507) );
  AOI22_X1 U20728 ( .A1(n17618), .A2(n17508), .B1(n17507), .B2(n17596), .ZN(
        P3_U2689) );
  AOI22_X1 U20729 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20730 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U20731 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17510) );
  AOI22_X1 U20732 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17509) );
  NAND4_X1 U20733 ( .A1(n17512), .A2(n17511), .A3(n17510), .A4(n17509), .ZN(
        n17518) );
  AOI22_X1 U20734 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U20735 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17515) );
  AOI22_X1 U20736 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20737 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17513) );
  NAND4_X1 U20738 ( .A1(n17516), .A2(n17515), .A3(n17514), .A4(n17513), .ZN(
        n17517) );
  NOR2_X1 U20739 ( .A1(n17518), .A2(n17517), .ZN(n17723) );
  NOR2_X1 U20740 ( .A1(n17533), .A2(n17548), .ZN(n17532) );
  OAI21_X1 U20741 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17532), .A(n17519), .ZN(
        n17520) );
  AOI22_X1 U20742 ( .A1(n17618), .A2(n17723), .B1(n17520), .B2(n17596), .ZN(
        P3_U2691) );
  AOI22_X1 U20743 ( .A1(n9666), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20744 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20745 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16191), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20746 ( .B1(n17522), .B2(n17608), .A(n17521), .ZN(n17528) );
  AOI22_X1 U20747 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U20748 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20749 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U20750 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17523) );
  NAND4_X1 U20751 ( .A1(n17526), .A2(n17525), .A3(n17524), .A4(n17523), .ZN(
        n17527) );
  AOI211_X1 U20752 ( .C1(n17566), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17528), .B(n17527), .ZN(n17529) );
  NAND3_X1 U20753 ( .A1(n17531), .A2(n17530), .A3(n17529), .ZN(n17726) );
  INV_X1 U20754 ( .A(n17532), .ZN(n17535) );
  AOI21_X1 U20755 ( .B1(n17533), .B2(n17548), .A(n17618), .ZN(n17534) );
  AOI22_X1 U20756 ( .A1(n17726), .A2(n17618), .B1(n17535), .B2(n17534), .ZN(
        n17536) );
  INV_X1 U20757 ( .A(n17536), .ZN(P3_U2692) );
  AOI22_X1 U20758 ( .A1(n17537), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20759 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17566), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17540) );
  AOI22_X1 U20760 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17574), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20761 ( .A1(n11555), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17538) );
  NAND4_X1 U20762 ( .A1(n17541), .A2(n17540), .A3(n17539), .A4(n17538), .ZN(
        n17547) );
  AOI22_X1 U20763 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17545) );
  AOI22_X1 U20764 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U20765 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20766 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17542) );
  NAND4_X1 U20767 ( .A1(n17545), .A2(n17544), .A3(n17543), .A4(n17542), .ZN(
        n17546) );
  NOR2_X1 U20768 ( .A1(n17547), .A2(n17546), .ZN(n17730) );
  OAI21_X1 U20769 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17565), .A(n17548), .ZN(
        n17549) );
  AOI22_X1 U20770 ( .A1(n17618), .A2(n17730), .B1(n17549), .B2(n17596), .ZN(
        P3_U2693) );
  AOI21_X1 U20771 ( .B1(n17550), .B2(n17583), .A(n17618), .ZN(n17551) );
  INV_X1 U20772 ( .A(n17551), .ZN(n17564) );
  AOI22_X1 U20773 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9666), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U20774 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17574), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17552), .ZN(n17556) );
  AOI22_X1 U20775 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20776 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9651), .ZN(n17554) );
  NAND4_X1 U20777 ( .A1(n17557), .A2(n17556), .A3(n17555), .A4(n17554), .ZN(
        n17563) );
  AOI22_X1 U20778 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17561) );
  AOI22_X1 U20779 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11489), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17566), .ZN(n17560) );
  AOI22_X1 U20780 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9653), .ZN(n17559) );
  AOI22_X1 U20781 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11513), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17455), .ZN(n17558) );
  NAND4_X1 U20782 ( .A1(n17561), .A2(n17560), .A3(n17559), .A4(n17558), .ZN(
        n17562) );
  NOR2_X1 U20783 ( .A1(n17563), .A2(n17562), .ZN(n17734) );
  OAI22_X1 U20784 ( .A1(n17565), .A2(n17564), .B1(n17734), .B2(n17596), .ZN(
        P3_U2694) );
  AOI22_X1 U20785 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11555), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17571) );
  AOI22_X1 U20786 ( .A1(n17566), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U20787 ( .A1(n11509), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17567), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U20788 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17537), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17568) );
  NAND4_X1 U20789 ( .A1(n17571), .A2(n17570), .A3(n17569), .A4(n17568), .ZN(
        n17582) );
  AOI22_X1 U20790 ( .A1(n17573), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17572), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U20791 ( .A1(n17574), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17552), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17579) );
  AOI22_X1 U20792 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17575), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U20793 ( .A1(n17576), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11513), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17577) );
  NAND4_X1 U20794 ( .A1(n17580), .A2(n17579), .A3(n17578), .A4(n17577), .ZN(
        n17581) );
  NOR2_X1 U20795 ( .A1(n17582), .A2(n17581), .ZN(n17741) );
  OAI21_X1 U20796 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17591), .A(n17583), .ZN(
        n17584) );
  AOI22_X1 U20797 ( .A1(n17618), .A2(n17741), .B1(n17584), .B2(n17596), .ZN(
        P3_U2695) );
  INV_X1 U20798 ( .A(n17585), .ZN(n17603) );
  NOR2_X1 U20799 ( .A1(n17586), .A2(n17603), .ZN(n17595) );
  AND2_X1 U20800 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17595), .ZN(n17599) );
  NAND2_X1 U20801 ( .A1(n18642), .A2(n17599), .ZN(n17594) );
  NOR2_X1 U20802 ( .A1(n17587), .A2(n17594), .ZN(n17588) );
  OAI21_X1 U20803 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17588), .A(n17596), .ZN(
        n17590) );
  OAI22_X1 U20804 ( .A1(n17591), .A2(n17590), .B1(n17589), .B2(n17596), .ZN(
        P3_U2696) );
  NAND3_X1 U20805 ( .A1(n17594), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17596), .ZN(
        n17592) );
  OAI221_X1 U20806 ( .B1(n17594), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17596), 
        .C2(n17593), .A(n17592), .ZN(P3_U2697) );
  OAI21_X1 U20807 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17595), .A(n17596), .ZN(
        n17598) );
  INV_X1 U20808 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17597) );
  OAI22_X1 U20809 ( .A1(n17599), .A2(n17598), .B1(n17597), .B2(n17596), .ZN(
        P3_U2698) );
  INV_X1 U20810 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17605) );
  NOR2_X1 U20811 ( .A1(n17600), .A2(n17615), .ZN(n17610) );
  NAND2_X1 U20812 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17610), .ZN(n17606) );
  OAI21_X1 U20813 ( .B1(n17618), .B2(n17601), .A(n17606), .ZN(n17602) );
  OAI21_X1 U20814 ( .B1(n17615), .B2(n17603), .A(n17602), .ZN(n17604) );
  OAI21_X1 U20815 ( .B1(n17596), .B2(n17605), .A(n17604), .ZN(P3_U2699) );
  OAI211_X1 U20816 ( .C1(n17610), .C2(P3_EBX_REG_3__SCAN_IN), .A(n17596), .B(
        n17606), .ZN(n17607) );
  OAI21_X1 U20817 ( .B1(n17596), .B2(n17608), .A(n17607), .ZN(P3_U2700) );
  NOR2_X1 U20818 ( .A1(n17620), .A2(n17614), .ZN(n17609) );
  AOI221_X1 U20819 ( .B1(n17609), .B2(n17621), .C1(n17729), .C2(n17621), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17611) );
  AOI211_X1 U20820 ( .C1(n17618), .C2(n17612), .A(n17611), .B(n17610), .ZN(
        P3_U2701) );
  OAI222_X1 U20821 ( .A1(n17616), .A2(n17615), .B1(n17614), .B2(n17621), .C1(
        n17613), .C2(n17596), .ZN(P3_U2702) );
  AOI22_X1 U20822 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17618), .B1(
        n17617), .B2(n17620), .ZN(n17619) );
  OAI21_X1 U20823 ( .B1(n17621), .B2(n17620), .A(n17619), .ZN(P3_U2703) );
  INV_X1 U20824 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17853) );
  INV_X1 U20825 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17787) );
  INV_X1 U20826 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17789) );
  INV_X1 U20827 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17791) );
  INV_X1 U20828 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17806) );
  NAND3_X1 U20829 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .ZN(n17744) );
  NAND2_X1 U20830 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17745) );
  NOR2_X1 U20831 ( .A1(n17744), .A2(n17745), .ZN(n17623) );
  NAND4_X1 U20832 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17623), .ZN(n17743) );
  NOR2_X1 U20833 ( .A1(n17624), .A2(n17743), .ZN(n17738) );
  NAND2_X1 U20834 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17712) );
  NAND4_X1 U20835 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17625)
         );
  NAND2_X1 U20836 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17714), .ZN(n17708) );
  NOR2_X2 U20837 ( .A1(n17806), .A2(n17708), .ZN(n17703) );
  INV_X1 U20838 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17793) );
  INV_X1 U20839 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17795) );
  INV_X1 U20840 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17797) );
  INV_X1 U20841 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17842) );
  NOR4_X1 U20842 ( .A1(n17793), .A2(n17795), .A3(n17797), .A4(n17842), .ZN(
        n17626) );
  NAND4_X1 U20843 ( .A1(n17703), .A2(P3_EAX_REG_19__SCAN_IN), .A3(
        P3_EAX_REG_18__SCAN_IN), .A4(n17626), .ZN(n17666) );
  NAND2_X1 U20844 ( .A1(n18642), .A2(n17665), .ZN(n17660) );
  NOR2_X2 U20845 ( .A1(n17787), .A2(n17661), .ZN(n17654) );
  NOR2_X2 U20846 ( .A1(n17853), .A2(n17650), .ZN(n17644) );
  NAND2_X1 U20847 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17644), .ZN(n17641) );
  NAND2_X1 U20848 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17636), .ZN(n17635) );
  NOR2_X1 U20849 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17635), .ZN(n17628) );
  NAND2_X1 U20850 ( .A1(n17763), .A2(n17635), .ZN(n17634) );
  OAI21_X1 U20851 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17742), .A(n17634), .ZN(
        n17627) );
  AOI22_X1 U20852 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17628), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17627), .ZN(n17629) );
  OAI21_X1 U20853 ( .B1(n17630), .B2(n17671), .A(n17629), .ZN(P3_U2704) );
  INV_X1 U20854 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17857) );
  NOR2_X2 U20855 ( .A1(n18627), .A2(n17763), .ZN(n17702) );
  OAI22_X1 U20856 ( .A1(n17631), .A2(n17766), .B1(n12670), .B2(n17671), .ZN(
        n17632) );
  AOI21_X1 U20857 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17702), .A(n17632), .ZN(
        n17633) );
  OAI221_X1 U20858 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17635), .C1(n17857), 
        .C2(n17634), .A(n17633), .ZN(P3_U2705) );
  AOI22_X1 U20859 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17701), .ZN(n17638) );
  OAI211_X1 U20860 ( .C1(n17636), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17763), .B(
        n17635), .ZN(n17637) );
  OAI211_X1 U20861 ( .C1(n17639), .C2(n17766), .A(n17638), .B(n17637), .ZN(
        P3_U2706) );
  AOI22_X1 U20862 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17702), .B1(n17771), .B2(
        n17640), .ZN(n17643) );
  OAI211_X1 U20863 ( .C1(n17644), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17763), .B(
        n17641), .ZN(n17642) );
  OAI211_X1 U20864 ( .C1(n17671), .C2(n15333), .A(n17643), .B(n17642), .ZN(
        P3_U2707) );
  AOI22_X1 U20865 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17701), .ZN(n17647) );
  AOI211_X1 U20866 ( .C1(n17853), .C2(n17650), .A(n17644), .B(n17715), .ZN(
        n17645) );
  INV_X1 U20867 ( .A(n17645), .ZN(n17646) );
  OAI211_X1 U20868 ( .C1(n17648), .C2(n17766), .A(n17647), .B(n17646), .ZN(
        P3_U2708) );
  INV_X1 U20869 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17653) );
  AOI22_X1 U20870 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17702), .B1(n17771), .B2(
        n17649), .ZN(n17652) );
  OAI211_X1 U20871 ( .C1(n17654), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17763), .B(
        n17650), .ZN(n17651) );
  OAI211_X1 U20872 ( .C1(n17671), .C2(n17653), .A(n17652), .B(n17651), .ZN(
        P3_U2709) );
  AOI22_X1 U20873 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17701), .ZN(n17657) );
  AOI211_X1 U20874 ( .C1(n17787), .C2(n17661), .A(n17654), .B(n17715), .ZN(
        n17655) );
  INV_X1 U20875 ( .A(n17655), .ZN(n17656) );
  OAI211_X1 U20876 ( .C1(n17658), .C2(n17766), .A(n17657), .B(n17656), .ZN(
        P3_U2710) );
  AOI22_X1 U20877 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17702), .B1(n17771), .B2(
        n17659), .ZN(n17664) );
  OAI21_X1 U20878 ( .B1(n17789), .B2(n17715), .A(n17660), .ZN(n17662) );
  NAND2_X1 U20879 ( .A1(n17662), .A2(n17661), .ZN(n17663) );
  OAI211_X1 U20880 ( .C1(n17671), .C2(n18604), .A(n17664), .B(n17663), .ZN(
        P3_U2711) );
  AOI211_X1 U20881 ( .C1(n17791), .C2(n17666), .A(n17715), .B(n17665), .ZN(
        n17667) );
  AOI21_X1 U20882 ( .B1(n17701), .B2(BUF2_REG_23__SCAN_IN), .A(n17667), .ZN(
        n17669) );
  NAND2_X1 U20883 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17702), .ZN(n17668) );
  OAI211_X1 U20884 ( .C1(n17670), .C2(n17766), .A(n17669), .B(n17668), .ZN(
        P3_U2712) );
  INV_X1 U20885 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17800) );
  INV_X1 U20886 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17802) );
  NAND2_X1 U20887 ( .A1(n18642), .A2(n17703), .ZN(n17695) );
  NAND2_X1 U20888 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17685), .ZN(n17681) );
  NAND2_X1 U20889 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17677), .ZN(n17676) );
  NAND2_X1 U20890 ( .A1(n17676), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17675) );
  OAI22_X1 U20891 ( .A1(n17672), .A2(n17766), .B1(n18634), .B2(n17671), .ZN(
        n17673) );
  AOI21_X1 U20892 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17702), .A(n17673), .ZN(
        n17674) );
  OAI221_X1 U20893 ( .B1(n17676), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17675), 
        .C2(n17715), .A(n17674), .ZN(P3_U2713) );
  AOI22_X1 U20894 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17701), .ZN(n17679) );
  OAI211_X1 U20895 ( .C1(n17677), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17763), .B(
        n17676), .ZN(n17678) );
  OAI211_X1 U20896 ( .C1(n17680), .C2(n17766), .A(n17679), .B(n17678), .ZN(
        P3_U2714) );
  AOI22_X1 U20897 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17701), .ZN(n17683) );
  OAI211_X1 U20898 ( .C1(n17685), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17763), .B(
        n17681), .ZN(n17682) );
  OAI211_X1 U20899 ( .C1(n17684), .C2(n17766), .A(n17683), .B(n17682), .ZN(
        P3_U2715) );
  AOI22_X1 U20900 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17701), .ZN(n17688) );
  NAND2_X1 U20901 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17691), .ZN(n17690) );
  AOI211_X1 U20902 ( .C1(n17800), .C2(n17690), .A(n17685), .B(n17715), .ZN(
        n17686) );
  INV_X1 U20903 ( .A(n17686), .ZN(n17687) );
  OAI211_X1 U20904 ( .C1(n17689), .C2(n17766), .A(n17688), .B(n17687), .ZN(
        P3_U2716) );
  AOI22_X1 U20905 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17701), .ZN(n17693) );
  OAI211_X1 U20906 ( .C1(n17691), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17763), .B(
        n17690), .ZN(n17692) );
  OAI211_X1 U20907 ( .C1(n17694), .C2(n17766), .A(n17693), .B(n17692), .ZN(
        P3_U2717) );
  AOI22_X1 U20908 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17701), .ZN(n17699) );
  OAI21_X1 U20909 ( .B1(n17842), .B2(n17715), .A(n17695), .ZN(n17697) );
  NAND2_X1 U20910 ( .A1(n17697), .A2(n17696), .ZN(n17698) );
  OAI211_X1 U20911 ( .C1(n17700), .C2(n17766), .A(n17699), .B(n17698), .ZN(
        P3_U2718) );
  AOI22_X1 U20912 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17702), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17701), .ZN(n17706) );
  AOI211_X1 U20913 ( .C1(n17806), .C2(n17708), .A(n17715), .B(n17703), .ZN(
        n17704) );
  INV_X1 U20914 ( .A(n17704), .ZN(n17705) );
  OAI211_X1 U20915 ( .C1(n17707), .C2(n17766), .A(n17706), .B(n17705), .ZN(
        P3_U2719) );
  OAI211_X1 U20916 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17714), .A(n17763), .B(
        n17708), .ZN(n17710) );
  NAND2_X1 U20917 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17772), .ZN(n17709) );
  OAI211_X1 U20918 ( .C1(n17711), .C2(n17766), .A(n17710), .B(n17709), .ZN(
        P3_U2720) );
  INV_X1 U20919 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17874) );
  OR3_X1 U20920 ( .A1(n17729), .A2(n17737), .A3(n17712), .ZN(n17728) );
  NOR2_X1 U20921 ( .A1(n17874), .A2(n17728), .ZN(n17722) );
  NAND2_X1 U20922 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17725), .ZN(n17718) );
  AOI22_X1 U20923 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17772), .B1(n17771), .B2(
        n17713), .ZN(n17717) );
  INV_X1 U20924 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17883) );
  OR3_X1 U20925 ( .A1(n17883), .A2(n17715), .A3(n17714), .ZN(n17716) );
  OAI211_X1 U20926 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17718), .A(n17717), .B(
        n17716), .ZN(P3_U2721) );
  INV_X1 U20927 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17881) );
  INV_X1 U20928 ( .A(n17718), .ZN(n17721) );
  AOI21_X1 U20929 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17763), .A(n17725), .ZN(
        n17720) );
  OAI222_X1 U20930 ( .A1(n17769), .A2(n17881), .B1(n17721), .B2(n17720), .C1(
        n17766), .C2(n17719), .ZN(P3_U2722) );
  INV_X1 U20931 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17876) );
  AOI21_X1 U20932 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17763), .A(n17722), .ZN(
        n17724) );
  OAI222_X1 U20933 ( .A1(n17769), .A2(n17876), .B1(n17725), .B2(n17724), .C1(
        n17766), .C2(n17723), .ZN(P3_U2723) );
  NAND2_X1 U20934 ( .A1(n17763), .A2(n17728), .ZN(n17732) );
  AOI22_X1 U20935 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17772), .B1(n17771), .B2(
        n17726), .ZN(n17727) );
  OAI221_X1 U20936 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17728), .C1(n17874), 
        .C2(n17732), .A(n17727), .ZN(P3_U2724) );
  INV_X1 U20937 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17872) );
  NOR2_X1 U20938 ( .A1(n17729), .A2(n17737), .ZN(n17733) );
  AOI21_X1 U20939 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17733), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17731) );
  OAI222_X1 U20940 ( .A1(n17769), .A2(n17872), .B1(n17732), .B2(n17731), .C1(
        n17766), .C2(n17730), .ZN(P3_U2725) );
  INV_X1 U20941 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17870) );
  INV_X1 U20942 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17817) );
  NOR2_X1 U20943 ( .A1(n17737), .A2(n17817), .ZN(n17736) );
  AOI21_X1 U20944 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17763), .A(n17733), .ZN(
        n17735) );
  OAI222_X1 U20945 ( .A1(n17769), .A2(n17870), .B1(n17736), .B2(n17735), .C1(
        n17766), .C2(n17734), .ZN(P3_U2726) );
  OAI211_X1 U20946 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17738), .A(n17763), .B(
        n17737), .ZN(n17740) );
  NAND2_X1 U20947 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17772), .ZN(n17739) );
  OAI211_X1 U20948 ( .C1(n17741), .C2(n17766), .A(n17740), .B(n17739), .ZN(
        P3_U2727) );
  INV_X1 U20949 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18639) );
  NOR2_X1 U20950 ( .A1(n17743), .A2(n17742), .ZN(n17748) );
  NOR2_X1 U20951 ( .A1(n17744), .A2(n17775), .ZN(n17761) );
  INV_X1 U20952 ( .A(n17761), .ZN(n17755) );
  NOR2_X1 U20953 ( .A1(n17745), .A2(n17755), .ZN(n17753) );
  AOI22_X1 U20954 ( .A1(n17753), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17763), .ZN(n17747) );
  OAI222_X1 U20955 ( .A1(n17769), .A2(n18639), .B1(n17748), .B2(n17747), .C1(
        n17766), .C2(n17746), .ZN(P3_U2728) );
  INV_X1 U20956 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18635) );
  AOI21_X1 U20957 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17763), .A(n17753), .ZN(
        n17751) );
  AND2_X1 U20958 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17753), .ZN(n17750) );
  OAI222_X1 U20959 ( .A1(n17769), .A2(n18635), .B1(n17751), .B2(n17750), .C1(
        n17766), .C2(n17749), .ZN(P3_U2729) );
  INV_X1 U20960 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18628) );
  AOI22_X1 U20961 ( .A1(n17761), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17763), .ZN(n17754) );
  OAI222_X1 U20962 ( .A1(n17769), .A2(n18628), .B1(n17754), .B2(n17753), .C1(
        n17766), .C2(n17752), .ZN(P3_U2730) );
  INV_X1 U20963 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18624) );
  AOI21_X1 U20964 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17763), .A(n17761), .ZN(
        n17758) );
  INV_X1 U20965 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17827) );
  NOR2_X1 U20966 ( .A1(n17827), .A2(n17755), .ZN(n17757) );
  OAI222_X1 U20967 ( .A1(n17769), .A2(n18624), .B1(n17758), .B2(n17757), .C1(
        n17766), .C2(n17756), .ZN(P3_U2731) );
  INV_X1 U20968 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18620) );
  NAND2_X1 U20969 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n17759) );
  NOR2_X1 U20970 ( .A1(n17759), .A2(n17775), .ZN(n17768) );
  AOI21_X1 U20971 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17763), .A(n17768), .ZN(
        n17762) );
  OAI222_X1 U20972 ( .A1(n17769), .A2(n18620), .B1(n17762), .B2(n17761), .C1(
        n17766), .C2(n17760), .ZN(P3_U2732) );
  INV_X1 U20973 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18615) );
  AOI22_X1 U20974 ( .A1(n17764), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17763), .ZN(n17767) );
  OAI222_X1 U20975 ( .A1(n18615), .A2(n17769), .B1(n17768), .B2(n17767), .C1(
        n17766), .C2(n17765), .ZN(P3_U2733) );
  INV_X1 U20976 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U20977 ( .A1(n17772), .A2(BUF2_REG_1__SCAN_IN), .B1(n17771), .B2(
        n17770), .ZN(n17773) );
  OAI221_X1 U20978 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17775), .C1(n17860), 
        .C2(n17774), .A(n17773), .ZN(P3_U2734) );
  NOR2_X2 U20979 ( .A1(n19216), .A2(n19113), .ZN(n19253) );
  INV_X1 U20980 ( .A(n17839), .ZN(n17837) );
  NOR2_X4 U20981 ( .A1(n19253), .A2(n17777), .ZN(n17798) );
  AND2_X1 U20982 ( .A1(n17798), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20983 ( .A1(n17777), .A2(n18610), .ZN(n17805) );
  AOI22_X1 U20984 ( .A1(n19253), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17798), .ZN(n17778) );
  OAI21_X1 U20985 ( .B1(n17857), .B2(n17805), .A(n17778), .ZN(P3_U2737) );
  INV_X1 U20986 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U20987 ( .A1(n19253), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17779) );
  OAI21_X1 U20988 ( .B1(n17780), .B2(n17805), .A(n17779), .ZN(P3_U2738) );
  INV_X1 U20989 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17782) );
  AOI22_X1 U20990 ( .A1(n19253), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17781) );
  OAI21_X1 U20991 ( .B1(n17782), .B2(n17805), .A(n17781), .ZN(P3_U2739) );
  AOI22_X1 U20992 ( .A1(n19253), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17783) );
  OAI21_X1 U20993 ( .B1(n17853), .B2(n17805), .A(n17783), .ZN(P3_U2740) );
  INV_X1 U20994 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17785) );
  AOI22_X1 U20995 ( .A1(n19253), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17784) );
  OAI21_X1 U20996 ( .B1(n17785), .B2(n17805), .A(n17784), .ZN(P3_U2741) );
  AOI22_X1 U20997 ( .A1(n19253), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17786) );
  OAI21_X1 U20998 ( .B1(n17787), .B2(n17805), .A(n17786), .ZN(P3_U2742) );
  AOI22_X1 U20999 ( .A1(n19253), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17788) );
  OAI21_X1 U21000 ( .B1(n17789), .B2(n17805), .A(n17788), .ZN(P3_U2743) );
  CLKBUF_X1 U21001 ( .A(n19253), .Z(n17833) );
  AOI22_X1 U21002 ( .A1(n17833), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17790) );
  OAI21_X1 U21003 ( .B1(n17791), .B2(n17805), .A(n17790), .ZN(P3_U2744) );
  AOI22_X1 U21004 ( .A1(n17833), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17792) );
  OAI21_X1 U21005 ( .B1(n17793), .B2(n17805), .A(n17792), .ZN(P3_U2745) );
  AOI22_X1 U21006 ( .A1(n17833), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17794) );
  OAI21_X1 U21007 ( .B1(n17795), .B2(n17805), .A(n17794), .ZN(P3_U2746) );
  AOI22_X1 U21008 ( .A1(n17833), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17796) );
  OAI21_X1 U21009 ( .B1(n17797), .B2(n17805), .A(n17796), .ZN(P3_U2747) );
  AOI22_X1 U21010 ( .A1(n17833), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17799) );
  OAI21_X1 U21011 ( .B1(n17800), .B2(n17805), .A(n17799), .ZN(P3_U2748) );
  AOI22_X1 U21012 ( .A1(n17833), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17801) );
  OAI21_X1 U21013 ( .B1(n17802), .B2(n17805), .A(n17801), .ZN(P3_U2749) );
  AOI22_X1 U21014 ( .A1(n17833), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17803) );
  OAI21_X1 U21015 ( .B1(n17842), .B2(n17805), .A(n17803), .ZN(P3_U2750) );
  AOI22_X1 U21016 ( .A1(n17833), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17804) );
  OAI21_X1 U21017 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(P3_U2751) );
  INV_X1 U21018 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17888) );
  AOI22_X1 U21019 ( .A1(n17833), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17807) );
  OAI21_X1 U21020 ( .B1(n17888), .B2(n17835), .A(n17807), .ZN(P3_U2752) );
  AOI22_X1 U21021 ( .A1(n17833), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17808) );
  OAI21_X1 U21022 ( .B1(n17883), .B2(n17835), .A(n17808), .ZN(P3_U2753) );
  INV_X1 U21023 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17810) );
  AOI22_X1 U21024 ( .A1(n17833), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17809) );
  OAI21_X1 U21025 ( .B1(n17810), .B2(n17835), .A(n17809), .ZN(P3_U2754) );
  INV_X1 U21026 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U21027 ( .A1(n17833), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17811) );
  OAI21_X1 U21028 ( .B1(n17812), .B2(n17835), .A(n17811), .ZN(P3_U2755) );
  AOI22_X1 U21029 ( .A1(n17833), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17813) );
  OAI21_X1 U21030 ( .B1(n17874), .B2(n17835), .A(n17813), .ZN(P3_U2756) );
  INV_X1 U21031 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U21032 ( .A1(n17833), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17814) );
  OAI21_X1 U21033 ( .B1(n17815), .B2(n17835), .A(n17814), .ZN(P3_U2757) );
  AOI22_X1 U21034 ( .A1(n17833), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17816) );
  OAI21_X1 U21035 ( .B1(n17817), .B2(n17835), .A(n17816), .ZN(P3_U2758) );
  INV_X1 U21036 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U21037 ( .A1(n17833), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17818) );
  OAI21_X1 U21038 ( .B1(n17819), .B2(n17835), .A(n17818), .ZN(P3_U2759) );
  INV_X1 U21039 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U21040 ( .A1(n17833), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17820) );
  OAI21_X1 U21041 ( .B1(n17821), .B2(n17835), .A(n17820), .ZN(P3_U2760) );
  INV_X1 U21042 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17823) );
  AOI22_X1 U21043 ( .A1(n17833), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17822) );
  OAI21_X1 U21044 ( .B1(n17823), .B2(n17835), .A(n17822), .ZN(P3_U2761) );
  INV_X1 U21045 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U21046 ( .A1(n17833), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17824) );
  OAI21_X1 U21047 ( .B1(n17825), .B2(n17835), .A(n17824), .ZN(P3_U2762) );
  AOI22_X1 U21048 ( .A1(n17833), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17826) );
  OAI21_X1 U21049 ( .B1(n17827), .B2(n17835), .A(n17826), .ZN(P3_U2763) );
  INV_X1 U21050 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U21051 ( .A1(n17833), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U21052 ( .B1(n17829), .B2(n17835), .A(n17828), .ZN(P3_U2764) );
  INV_X1 U21053 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U21054 ( .A1(n17833), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U21055 ( .B1(n17831), .B2(n17835), .A(n17830), .ZN(P3_U2765) );
  AOI22_X1 U21056 ( .A1(n17833), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17832) );
  OAI21_X1 U21057 ( .B1(n17860), .B2(n17835), .A(n17832), .ZN(P3_U2766) );
  AOI22_X1 U21058 ( .A1(n17833), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17798), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17834) );
  OAI21_X1 U21059 ( .B1(n17836), .B2(n17835), .A(n17834), .ZN(P3_U2767) );
  INV_X1 U21060 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18605) );
  OAI211_X1 U21061 ( .C1(n19257), .C2(n19256), .A(n17838), .B(n17837), .ZN(
        n17884) );
  OR2_X1 U21062 ( .A1(n19094), .A2(n17839), .ZN(n17887) );
  AOI22_X1 U21063 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17877), .ZN(n17840) );
  OAI21_X1 U21064 ( .B1(n18605), .B2(n17880), .A(n17840), .ZN(P3_U2768) );
  AOI22_X1 U21065 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17885), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17877), .ZN(n17841) );
  OAI21_X1 U21066 ( .B1(n17842), .B2(n17887), .A(n17841), .ZN(P3_U2769) );
  AOI22_X1 U21067 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17877), .ZN(n17843) );
  OAI21_X1 U21068 ( .B1(n18615), .B2(n17880), .A(n17843), .ZN(P3_U2770) );
  AOI22_X1 U21069 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17877), .ZN(n17844) );
  OAI21_X1 U21070 ( .B1(n18620), .B2(n17880), .A(n17844), .ZN(P3_U2771) );
  AOI22_X1 U21071 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17877), .ZN(n17845) );
  OAI21_X1 U21072 ( .B1(n18624), .B2(n17880), .A(n17845), .ZN(P3_U2772) );
  AOI22_X1 U21073 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17877), .ZN(n17846) );
  OAI21_X1 U21074 ( .B1(n18628), .B2(n17880), .A(n17846), .ZN(P3_U2773) );
  AOI22_X1 U21075 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17877), .ZN(n17847) );
  OAI21_X1 U21076 ( .B1(n18635), .B2(n17880), .A(n17847), .ZN(P3_U2774) );
  AOI22_X1 U21077 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17877), .ZN(n17848) );
  OAI21_X1 U21078 ( .B1(n18639), .B2(n17880), .A(n17848), .ZN(P3_U2775) );
  INV_X1 U21079 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U21080 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17877), .ZN(n17849) );
  OAI21_X1 U21081 ( .B1(n17868), .B2(n17880), .A(n17849), .ZN(P3_U2776) );
  AOI22_X1 U21082 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17877), .ZN(n17850) );
  OAI21_X1 U21083 ( .B1(n17870), .B2(n17880), .A(n17850), .ZN(P3_U2777) );
  AOI22_X1 U21084 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17877), .ZN(n17851) );
  OAI21_X1 U21085 ( .B1(n17872), .B2(n17880), .A(n17851), .ZN(P3_U2778) );
  AOI22_X1 U21086 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17885), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17877), .ZN(n17852) );
  OAI21_X1 U21087 ( .B1(n17853), .B2(n17887), .A(n17852), .ZN(P3_U2779) );
  AOI22_X1 U21088 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17877), .ZN(n17854) );
  OAI21_X1 U21089 ( .B1(n17876), .B2(n17880), .A(n17854), .ZN(P3_U2780) );
  AOI22_X1 U21090 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17878), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17877), .ZN(n17855) );
  OAI21_X1 U21091 ( .B1(n17881), .B2(n17880), .A(n17855), .ZN(P3_U2781) );
  AOI22_X1 U21092 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17885), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17877), .ZN(n17856) );
  OAI21_X1 U21093 ( .B1(n17857), .B2(n17887), .A(n17856), .ZN(P3_U2782) );
  AOI22_X1 U21094 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17877), .ZN(n17858) );
  OAI21_X1 U21095 ( .B1(n18605), .B2(n17880), .A(n17858), .ZN(P3_U2783) );
  AOI22_X1 U21096 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17885), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17877), .ZN(n17859) );
  OAI21_X1 U21097 ( .B1(n17860), .B2(n17887), .A(n17859), .ZN(P3_U2784) );
  AOI22_X1 U21098 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17884), .ZN(n17861) );
  OAI21_X1 U21099 ( .B1(n18615), .B2(n17880), .A(n17861), .ZN(P3_U2785) );
  AOI22_X1 U21100 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17884), .ZN(n17862) );
  OAI21_X1 U21101 ( .B1(n18620), .B2(n17880), .A(n17862), .ZN(P3_U2786) );
  AOI22_X1 U21102 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17884), .ZN(n17863) );
  OAI21_X1 U21103 ( .B1(n18624), .B2(n17880), .A(n17863), .ZN(P3_U2787) );
  AOI22_X1 U21104 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17884), .ZN(n17864) );
  OAI21_X1 U21105 ( .B1(n18628), .B2(n17880), .A(n17864), .ZN(P3_U2788) );
  AOI22_X1 U21106 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17884), .ZN(n17865) );
  OAI21_X1 U21107 ( .B1(n18635), .B2(n17880), .A(n17865), .ZN(P3_U2789) );
  AOI22_X1 U21108 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17884), .ZN(n17866) );
  OAI21_X1 U21109 ( .B1(n18639), .B2(n17880), .A(n17866), .ZN(P3_U2790) );
  AOI22_X1 U21110 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17884), .ZN(n17867) );
  OAI21_X1 U21111 ( .B1(n17868), .B2(n17880), .A(n17867), .ZN(P3_U2791) );
  AOI22_X1 U21112 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17877), .ZN(n17869) );
  OAI21_X1 U21113 ( .B1(n17870), .B2(n17880), .A(n17869), .ZN(P3_U2792) );
  AOI22_X1 U21114 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17877), .ZN(n17871) );
  OAI21_X1 U21115 ( .B1(n17872), .B2(n17880), .A(n17871), .ZN(P3_U2793) );
  AOI22_X1 U21116 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17885), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17884), .ZN(n17873) );
  OAI21_X1 U21117 ( .B1(n17874), .B2(n17887), .A(n17873), .ZN(P3_U2794) );
  AOI22_X1 U21118 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17877), .ZN(n17875) );
  OAI21_X1 U21119 ( .B1(n17876), .B2(n17880), .A(n17875), .ZN(P3_U2795) );
  AOI22_X1 U21120 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17878), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17877), .ZN(n17879) );
  OAI21_X1 U21121 ( .B1(n17881), .B2(n17880), .A(n17879), .ZN(P3_U2796) );
  AOI22_X1 U21122 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17885), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17884), .ZN(n17882) );
  OAI21_X1 U21123 ( .B1(n17883), .B2(n17887), .A(n17882), .ZN(P3_U2797) );
  AOI22_X1 U21124 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17885), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17884), .ZN(n17886) );
  OAI21_X1 U21125 ( .B1(n17888), .B2(n17887), .A(n17886), .ZN(P3_U2798) );
  NAND2_X1 U21126 ( .A1(n18331), .A2(n18051), .ZN(n18017) );
  NAND2_X1 U21127 ( .A1(n18105), .A2(n17892), .ZN(n17899) );
  NOR3_X1 U21128 ( .A1(n18009), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17893), .ZN(n17911) );
  INV_X1 U21129 ( .A(n19113), .ZN(n18092) );
  INV_X1 U21130 ( .A(n18156), .ZN(n18212) );
  OAI21_X1 U21131 ( .B1(n17894), .B2(n18212), .A(n18255), .ZN(n17895) );
  AOI21_X1 U21132 ( .B1(n18092), .B2(n17896), .A(n17895), .ZN(n17921) );
  OAI21_X1 U21133 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17918), .A(
        n17921), .ZN(n17912) );
  OAI21_X1 U21134 ( .B1(n17911), .B2(n17912), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17898) );
  OAI211_X1 U21135 ( .C1(n17900), .C2(n17899), .A(n17898), .B(n17897), .ZN(
        n17901) );
  NAND2_X1 U21136 ( .A1(n18259), .A2(n18084), .ZN(n18001) );
  NAND2_X1 U21137 ( .A1(n17937), .A2(n17903), .ZN(n18268) );
  OR3_X1 U21138 ( .A1(n18290), .A2(n18272), .A3(n18324), .ZN(n18267) );
  AOI22_X1 U21139 ( .A1(n18248), .A2(n18268), .B1(n18165), .B2(n18267), .ZN(
        n17924) );
  NAND2_X1 U21140 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17924), .ZN(
        n17914) );
  NAND3_X1 U21141 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18001), .A3(
        n17914), .ZN(n17904) );
  NOR2_X1 U21142 ( .A1(n17907), .A2(n17906), .ZN(n17908) );
  XOR2_X1 U21143 ( .A(n17908), .B(n18142), .Z(n18278) );
  OAI22_X1 U21144 ( .A1(n18591), .A2(n19185), .B1(n18044), .B2(n17909), .ZN(
        n17910) );
  AOI211_X1 U21145 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17912), .A(
        n17911), .B(n17910), .ZN(n17917) );
  NOR2_X1 U21146 ( .A1(n17913), .A2(n18040), .ZN(n17965) );
  OAI221_X1 U21147 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17915), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17965), .A(n17914), .ZN(
        n17916) );
  OAI211_X1 U21148 ( .C1(n18278), .C2(n18168), .A(n17917), .B(n17916), .ZN(
        P3_U2803) );
  INV_X1 U21149 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18282) );
  NAND3_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18282), .ZN(n18288) );
  NAND2_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17965), .ZN(
        n17953) );
  NAND2_X1 U21152 ( .A1(n18044), .A2(n17918), .ZN(n18029) );
  AOI21_X1 U21153 ( .B1(n17919), .B2(n18981), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17920) );
  INV_X1 U21154 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19183) );
  OAI22_X1 U21155 ( .A1(n17921), .A2(n17920), .B1(n18591), .B2(n19183), .ZN(
        n17926) );
  AOI21_X1 U21156 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17923), .A(
        n17922), .ZN(n18281) );
  OAI22_X1 U21157 ( .A1(n17924), .A2(n18282), .B1(n18281), .B2(n18168), .ZN(
        n17925) );
  AOI211_X1 U21158 ( .C1(n17927), .C2(n18029), .A(n17926), .B(n17925), .ZN(
        n17928) );
  OAI21_X1 U21159 ( .B1(n18288), .B2(n17953), .A(n17928), .ZN(P3_U2804) );
  NAND2_X1 U21160 ( .A1(n18292), .A2(n18402), .ZN(n17929) );
  XOR2_X1 U21161 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17929), .Z(
        n18302) );
  NAND2_X1 U21162 ( .A1(n17930), .A2(n18105), .ZN(n17945) );
  AOI221_X1 U21163 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n17944), .C2(n17933), .A(
        n17945), .ZN(n17935) );
  OR2_X1 U21164 ( .A1(n18636), .A2(n17930), .ZN(n17961) );
  OAI211_X1 U21165 ( .C1(n17931), .C2(n19113), .A(n18255), .B(n17961), .ZN(
        n17958) );
  AOI21_X1 U21166 ( .B1(n17969), .B2(n17932), .A(n17958), .ZN(n17943) );
  OAI22_X1 U21167 ( .A1(n17943), .A2(n17933), .B1(n18591), .B2(n19181), .ZN(
        n17934) );
  AOI211_X1 U21168 ( .C1(n17936), .C2(n18115), .A(n17935), .B(n17934), .ZN(
        n17942) );
  NAND3_X1 U21169 ( .A1(n17937), .A2(n18280), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17938) );
  XOR2_X1 U21170 ( .A(n17938), .B(n18289), .Z(n18299) );
  AOI21_X1 U21171 ( .B1(n17949), .B2(n18155), .A(n17939), .ZN(n17940) );
  XOR2_X1 U21172 ( .A(n17940), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18298) );
  AOI22_X1 U21173 ( .A1(n18248), .A2(n18299), .B1(n18150), .B2(n18298), .ZN(
        n17941) );
  OAI211_X1 U21174 ( .C1(n18084), .C2(n18302), .A(n17942), .B(n17941), .ZN(
        P3_U2805) );
  NAND2_X1 U21175 ( .A1(n18570), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18315) );
  OAI221_X1 U21176 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17945), .C1(
        n17944), .C2(n17943), .A(n18315), .ZN(n17946) );
  AOI21_X1 U21177 ( .B1(n18115), .B2(n17947), .A(n17946), .ZN(n17952) );
  INV_X1 U21178 ( .A(n18280), .ZN(n17948) );
  NOR2_X1 U21179 ( .A1(n18410), .A2(n17948), .ZN(n18305) );
  NOR2_X1 U21180 ( .A1(n18324), .A2(n17948), .ZN(n18303) );
  OAI22_X1 U21181 ( .A1(n18305), .A2(n18259), .B1(n18303), .B2(n18084), .ZN(
        n17963) );
  OAI21_X1 U21182 ( .B1(n17950), .B2(n18310), .A(n17949), .ZN(n18314) );
  AOI22_X1 U21183 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17963), .B1(
        n18150), .B2(n18314), .ZN(n17951) );
  OAI211_X1 U21184 ( .C1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17953), .A(
        n17952), .B(n17951), .ZN(P3_U2806) );
  AOI22_X1 U21185 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18155), .B1(
        n17954), .B2(n17973), .ZN(n17955) );
  NAND2_X1 U21186 ( .A1(n17997), .A2(n17955), .ZN(n17956) );
  XOR2_X1 U21187 ( .A(n17956), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18323) );
  AOI22_X1 U21188 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17958), .B1(
        n17957), .B2(n18029), .ZN(n17959) );
  NAND2_X1 U21189 ( .A1(n18570), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18322) );
  OAI211_X1 U21190 ( .C1(n17961), .C2(n17960), .A(n17959), .B(n18322), .ZN(
        n17962) );
  AOI221_X1 U21191 ( .B1(n17965), .B2(n17964), .C1(n17963), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17962), .ZN(n17966) );
  OAI21_X1 U21192 ( .B1(n18168), .B2(n18323), .A(n17966), .ZN(P3_U2807) );
  NAND2_X1 U21193 ( .A1(n18092), .A2(n17967), .ZN(n17968) );
  OAI211_X1 U21194 ( .C1(n9767), .C2(n18212), .A(n18255), .B(n17968), .ZN(
        n17995) );
  AOI21_X1 U21195 ( .B1(n17969), .B2(n17992), .A(n17995), .ZN(n17981) );
  NAND2_X1 U21196 ( .A1(n18570), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18338) );
  INV_X1 U21197 ( .A(n18338), .ZN(n17971) );
  NAND2_X1 U21198 ( .A1(n9767), .A2(n18105), .ZN(n17982) );
  AOI221_X1 U21199 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n10082), .C2(n10083), .A(
        n17982), .ZN(n17970) );
  AOI211_X1 U21200 ( .C1(n17972), .C2(n18115), .A(n17971), .B(n17970), .ZN(
        n17980) );
  INV_X1 U21201 ( .A(n17973), .ZN(n17974) );
  OAI221_X1 U21202 ( .B1(n17974), .B2(n18334), .C1(n17974), .C2(n18049), .A(
        n17997), .ZN(n17975) );
  XOR2_X1 U21203 ( .A(n18262), .B(n17975), .Z(n18337) );
  INV_X1 U21204 ( .A(n18334), .ZN(n18264) );
  NOR2_X1 U21205 ( .A1(n18264), .A2(n18040), .ZN(n17977) );
  AOI22_X1 U21206 ( .A1(n18410), .A2(n18248), .B1(n18324), .B2(n18165), .ZN(
        n18054) );
  INV_X1 U21207 ( .A(n18054), .ZN(n18000) );
  AOI21_X1 U21208 ( .B1(n18264), .B2(n18001), .A(n18000), .ZN(n17991) );
  INV_X1 U21209 ( .A(n17991), .ZN(n17976) );
  MUX2_X1 U21210 ( .A(n17977), .B(n17976), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17978) );
  AOI21_X1 U21211 ( .B1(n18150), .B2(n18337), .A(n17978), .ZN(n17979) );
  OAI211_X1 U21212 ( .C1(n17981), .C2(n10083), .A(n17980), .B(n17979), .ZN(
        P3_U2808) );
  NAND2_X1 U21213 ( .A1(n18570), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18348) );
  OAI221_X1 U21214 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17982), .C1(
        n10082), .C2(n17981), .A(n18348), .ZN(n17988) );
  NOR3_X1 U21215 ( .A1(n18018), .A2(n18155), .A3(n17983), .ZN(n18005) );
  AOI22_X1 U21216 ( .A1(n17986), .A2(n18005), .B1(n18025), .B2(n17984), .ZN(
        n17985) );
  XOR2_X1 U21217 ( .A(n17985), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n18341) );
  NAND2_X1 U21218 ( .A1(n17986), .A2(n18344), .ZN(n18350) );
  OAI22_X1 U21219 ( .A1(n18341), .A2(n18168), .B1(n18017), .B2(n18350), .ZN(
        n17987) );
  AOI211_X1 U21220 ( .C1(n18115), .C2(n17989), .A(n17988), .B(n17987), .ZN(
        n17990) );
  OAI21_X1 U21221 ( .B1(n17991), .B2(n18344), .A(n17990), .ZN(P3_U2809) );
  OAI21_X1 U21222 ( .B1(n18636), .B2(n17993), .A(n17992), .ZN(n17994) );
  AOI22_X1 U21223 ( .A1(n17996), .A2(n18029), .B1(n17995), .B2(n17994), .ZN(
        n18004) );
  INV_X1 U21224 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18332) );
  OAI221_X1 U21225 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18024), 
        .C1(n18367), .C2(n18005), .A(n17997), .ZN(n17998) );
  XOR2_X1 U21226 ( .A(n18332), .B(n17998), .Z(n18359) );
  NOR2_X1 U21227 ( .A1(n17999), .A2(n18367), .ZN(n18352) );
  INV_X1 U21228 ( .A(n18352), .ZN(n18329) );
  AOI21_X1 U21229 ( .B1(n18001), .B2(n18329), .A(n18000), .ZN(n18016) );
  NAND2_X1 U21230 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18332), .ZN(
        n18363) );
  OAI22_X1 U21231 ( .A1(n18016), .A2(n18332), .B1(n18017), .B2(n18363), .ZN(
        n18002) );
  AOI21_X1 U21232 ( .B1(n18150), .B2(n18359), .A(n18002), .ZN(n18003) );
  OAI211_X1 U21233 ( .C1(n18591), .C2(n19171), .A(n18004), .B(n18003), .ZN(
        P3_U2810) );
  AOI21_X1 U21234 ( .B1(n18024), .B2(n18025), .A(n18005), .ZN(n18006) );
  XOR2_X1 U21235 ( .A(n18367), .B(n18006), .Z(n18364) );
  INV_X1 U21236 ( .A(n18189), .ZN(n18250) );
  OAI21_X1 U21237 ( .B1(n18226), .B2(n18008), .A(n18250), .ZN(n18030) );
  OAI21_X1 U21238 ( .B1(n18007), .B2(n19113), .A(n18030), .ZN(n18021) );
  AOI22_X1 U21239 ( .A1(n18581), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18021), .ZN(n18012) );
  NOR2_X1 U21240 ( .A1(n18009), .A2(n18008), .ZN(n18023) );
  NAND2_X1 U21241 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18010) );
  OAI211_X1 U21242 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18023), .B(n18010), .ZN(n18011) );
  OAI211_X1 U21243 ( .C1(n18044), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        n18014) );
  AOI21_X1 U21244 ( .B1(n18150), .B2(n18364), .A(n18014), .ZN(n18015) );
  OAI221_X1 U21245 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18017), 
        .C1(n18367), .C2(n18016), .A(n18015), .ZN(P3_U2811) );
  NAND2_X1 U21246 ( .A1(n18375), .A2(n18018), .ZN(n18382) );
  OAI22_X1 U21247 ( .A1(n18591), .A2(n19166), .B1(n18044), .B2(n18019), .ZN(
        n18020) );
  AOI221_X1 U21248 ( .B1(n18023), .B2(n18022), .C1(n18021), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18020), .ZN(n18028) );
  OAI21_X1 U21249 ( .B1(n18375), .B2(n18040), .A(n18054), .ZN(n18037) );
  AOI21_X1 U21250 ( .B1(n18142), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n18024), .ZN(n18026) );
  XOR2_X1 U21251 ( .A(n18026), .B(n18025), .Z(n18378) );
  AOI22_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18037), .B1(
        n18150), .B2(n18378), .ZN(n18027) );
  OAI211_X1 U21253 ( .C1(n18040), .C2(n18382), .A(n18028), .B(n18027), .ZN(
        P3_U2812) );
  NAND2_X1 U21254 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18383), .ZN(
        n18389) );
  INV_X1 U21255 ( .A(n18029), .ZN(n18244) );
  INV_X1 U21256 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19164) );
  NOR2_X1 U21257 ( .A1(n18591), .A2(n19164), .ZN(n18386) );
  AOI221_X1 U21258 ( .B1(n18636), .B2(n18032), .C1(n18031), .C2(n18032), .A(
        n18030), .ZN(n18033) );
  AOI211_X1 U21259 ( .C1(n18034), .C2(n18029), .A(n18386), .B(n18033), .ZN(
        n18039) );
  OAI21_X1 U21260 ( .B1(n18036), .B2(n18383), .A(n18035), .ZN(n18387) );
  AOI22_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18037), .B1(
        n18150), .B2(n18387), .ZN(n18038) );
  OAI211_X1 U21262 ( .C1(n18040), .C2(n18389), .A(n18039), .B(n18038), .ZN(
        P3_U2813) );
  NAND2_X1 U21263 ( .A1(n18041), .A2(n18105), .ZN(n18058) );
  AOI221_X1 U21264 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n18057), .C2(n18045), .A(
        n18058), .ZN(n18047) );
  OAI21_X1 U21265 ( .B1(n18041), .B2(n18212), .A(n18255), .ZN(n18075) );
  AOI21_X1 U21266 ( .B1(n18092), .B2(n18042), .A(n18075), .ZN(n18056) );
  OAI22_X1 U21267 ( .A1(n18056), .A2(n18045), .B1(n18044), .B2(n18043), .ZN(
        n18046) );
  AOI211_X1 U21268 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n18570), .A(n18047), 
        .B(n18046), .ZN(n18053) );
  NOR2_X1 U21269 ( .A1(n18155), .A2(n18460), .ZN(n18133) );
  INV_X1 U21270 ( .A(n18133), .ZN(n18141) );
  OAI22_X1 U21271 ( .A1(n18142), .A2(n18049), .B1(n18048), .B2(n18141), .ZN(
        n18050) );
  XOR2_X1 U21272 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18050), .Z(
        n18395) );
  AOI22_X1 U21273 ( .A1(n18150), .A2(n18395), .B1(n18051), .B2(n18398), .ZN(
        n18052) );
  OAI211_X1 U21274 ( .C1(n18054), .C2(n18398), .A(n18053), .B(n18052), .ZN(
        P3_U2814) );
  INV_X1 U21275 ( .A(n18415), .ZN(n18417) );
  NAND4_X1 U21276 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18417), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n18079), .ZN(n18080) );
  NAND2_X1 U21277 ( .A1(n18401), .A2(n18080), .ZN(n18409) );
  INV_X1 U21278 ( .A(n18409), .ZN(n18071) );
  NAND2_X1 U21279 ( .A1(n18248), .A2(n18410), .ZN(n18070) );
  NAND2_X1 U21280 ( .A1(n18570), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18055) );
  OAI221_X1 U21281 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18058), .C1(
        n18057), .C2(n18056), .A(n18055), .ZN(n18059) );
  AOI21_X1 U21282 ( .B1(n18115), .B2(n18060), .A(n18059), .ZN(n18069) );
  INV_X1 U21283 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18449) );
  INV_X1 U21284 ( .A(n18103), .ZN(n18448) );
  NAND3_X1 U21285 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18061), .ZN(n18063) );
  NOR3_X1 U21286 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18142), .A3(
        n9987), .ZN(n18132) );
  INV_X1 U21287 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18135) );
  NAND2_X1 U21288 ( .A1(n18132), .A2(n18135), .ZN(n18117) );
  NOR2_X1 U21289 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18117), .ZN(
        n18102) );
  NAND2_X1 U21290 ( .A1(n18102), .A2(n18420), .ZN(n18077) );
  OAI21_X1 U21291 ( .B1(n18448), .B2(n18063), .A(n18077), .ZN(n18064) );
  OAI221_X1 U21292 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18426), 
        .C1(n18449), .C2(n18142), .A(n18064), .ZN(n18065) );
  XOR2_X1 U21293 ( .A(n18401), .B(n18065), .Z(n18405) );
  NOR2_X1 U21294 ( .A1(n18402), .A2(n18084), .ZN(n18067) );
  NAND4_X1 U21295 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18417), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n18066), .ZN(n18082) );
  NAND2_X1 U21296 ( .A1(n18401), .A2(n18082), .ZN(n18404) );
  AOI22_X1 U21297 ( .A1(n18150), .A2(n18405), .B1(n18067), .B2(n18404), .ZN(
        n18068) );
  OAI211_X1 U21298 ( .C1(n18071), .C2(n18070), .A(n18069), .B(n18068), .ZN(
        P3_U2815) );
  OAI21_X1 U21299 ( .B1(n18636), .B2(n18073), .A(n18072), .ZN(n18074) );
  AOI22_X1 U21300 ( .A1(n18581), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18075), 
        .B2(n18074), .ZN(n18087) );
  OAI22_X1 U21301 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18077), .B1(
        n18141), .B2(n18076), .ZN(n18078) );
  XOR2_X1 U21302 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18078), .Z(
        n18427) );
  NAND2_X1 U21303 ( .A1(n18417), .A2(n18079), .ZN(n18441) );
  NOR2_X1 U21304 ( .A1(n18420), .A2(n18441), .ZN(n18081) );
  OAI21_X1 U21305 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18081), .A(
        n18080), .ZN(n18434) );
  NOR2_X1 U21306 ( .A1(n18415), .A2(n18460), .ZN(n18439) );
  INV_X1 U21307 ( .A(n18439), .ZN(n18089) );
  NOR2_X1 U21308 ( .A1(n18420), .A2(n18089), .ZN(n18083) );
  OAI21_X1 U21309 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18083), .A(
        n18082), .ZN(n18428) );
  OAI22_X1 U21310 ( .A1(n18259), .A2(n18434), .B1(n18084), .B2(n18428), .ZN(
        n18085) );
  AOI21_X1 U21311 ( .B1(n18150), .B2(n18427), .A(n18085), .ZN(n18086) );
  OAI211_X1 U21312 ( .C1(n18244), .C2(n18088), .A(n18087), .B(n18086), .ZN(
        P3_U2816) );
  AOI22_X1 U21313 ( .A1(n18248), .A2(n18441), .B1(n18165), .B2(n18089), .ZN(
        n18109) );
  NOR2_X1 U21314 ( .A1(n18591), .A2(n19156), .ZN(n18097) );
  OAI211_X1 U21315 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18120), .B(n18105), .ZN(n18094) );
  OAI21_X1 U21316 ( .B1(n18120), .B2(n18212), .A(n18255), .ZN(n18090) );
  AOI21_X1 U21317 ( .B1(n18092), .B2(n18091), .A(n18090), .ZN(n18106) );
  OAI22_X1 U21318 ( .A1(n18095), .A2(n18094), .B1(n18106), .B2(n18093), .ZN(
        n18096) );
  AOI211_X1 U21319 ( .C1(n18115), .C2(n18098), .A(n18097), .B(n18096), .ZN(
        n18101) );
  AOI22_X1 U21320 ( .A1(n18133), .A2(n18417), .B1(n18102), .B2(n18449), .ZN(
        n18099) );
  XOR2_X1 U21321 ( .A(n18420), .B(n18099), .Z(n18445) );
  NOR2_X1 U21322 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18415), .ZN(
        n18444) );
  AOI22_X1 U21323 ( .A1(n18150), .A2(n18445), .B1(n18444), .B2(n18127), .ZN(
        n18100) );
  OAI211_X1 U21324 ( .C1(n18109), .C2(n18420), .A(n18101), .B(n18100), .ZN(
        P3_U2817) );
  AOI21_X1 U21325 ( .B1(n18133), .B2(n18103), .A(n18102), .ZN(n18104) );
  XOR2_X1 U21326 ( .A(n18104), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18458) );
  NAND2_X1 U21327 ( .A1(n18120), .A2(n18105), .ZN(n18108) );
  INV_X1 U21328 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18107) );
  NAND2_X1 U21329 ( .A1(n18570), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18456) );
  OAI221_X1 U21330 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18108), .C1(
        n18107), .C2(n18106), .A(n18456), .ZN(n18113) );
  INV_X1 U21331 ( .A(n18127), .ZN(n18153) );
  NOR2_X1 U21332 ( .A1(n18153), .A2(n18448), .ZN(n18111) );
  INV_X1 U21333 ( .A(n18109), .ZN(n18110) );
  MUX2_X1 U21334 ( .A(n18111), .B(n18110), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18112) );
  AOI211_X1 U21335 ( .C1(n18115), .C2(n18114), .A(n18113), .B(n18112), .ZN(
        n18116) );
  OAI21_X1 U21336 ( .B1(n18458), .B2(n18168), .A(n18116), .ZN(P3_U2818) );
  OAI21_X1 U21337 ( .B1(n18128), .B2(n18141), .A(n18117), .ZN(n18118) );
  XOR2_X1 U21338 ( .A(n18118), .B(n18436), .Z(n18472) );
  NOR3_X1 U21339 ( .A1(n18636), .A2(n18171), .A3(n18174), .ZN(n18160) );
  NAND2_X1 U21340 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18160), .ZN(
        n18146) );
  NOR2_X1 U21341 ( .A1(n18145), .A2(n18146), .ZN(n18144) );
  NAND2_X1 U21342 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18144), .ZN(
        n18129) );
  NAND2_X1 U21343 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18250), .ZN(
        n18119) );
  AOI22_X1 U21344 ( .A1(n18981), .A2(n18120), .B1(n18129), .B2(n18119), .ZN(
        n18122) );
  INV_X1 U21345 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19152) );
  NOR2_X1 U21346 ( .A1(n18491), .A2(n19152), .ZN(n18121) );
  AOI211_X1 U21347 ( .C1(n18123), .C2(n18029), .A(n18122), .B(n18121), .ZN(
        n18126) );
  INV_X1 U21348 ( .A(n18128), .ZN(n18465) );
  AOI22_X1 U21349 ( .A1(n18248), .A2(n18462), .B1(n18165), .B2(n18460), .ZN(
        n18152) );
  OAI21_X1 U21350 ( .B1(n18465), .B2(n18153), .A(n18152), .ZN(n18124) );
  NOR2_X1 U21351 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18128), .ZN(
        n18459) );
  AOI22_X1 U21352 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18124), .B1(
        n18459), .B2(n18127), .ZN(n18125) );
  OAI211_X1 U21353 ( .C1(n18472), .C2(n18168), .A(n18126), .B(n18125), .ZN(
        P3_U2819) );
  NAND2_X1 U21354 ( .A1(n18128), .A2(n18127), .ZN(n18139) );
  OAI211_X1 U21355 ( .C1(n18144), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18250), .B(n18129), .ZN(n18130) );
  OAI21_X1 U21356 ( .B1(n18244), .B2(n18131), .A(n18130), .ZN(n18137) );
  AOI21_X1 U21357 ( .B1(n18133), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18132), .ZN(n18134) );
  XOR2_X1 U21358 ( .A(n18134), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18480) );
  OAI22_X1 U21359 ( .A1(n18480), .A2(n18168), .B1(n18152), .B2(n18135), .ZN(
        n18136) );
  AOI211_X1 U21360 ( .C1(n18570), .C2(P3_REIP_REG_10__SCAN_IN), .A(n18137), 
        .B(n18136), .ZN(n18138) );
  OAI21_X1 U21361 ( .B1(n18140), .B2(n18139), .A(n18138), .ZN(P3_U2820) );
  INV_X1 U21362 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18486) );
  OAI21_X1 U21363 ( .B1(n9987), .B2(n18142), .A(n18141), .ZN(n18143) );
  XOR2_X1 U21364 ( .A(n18143), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18488) );
  AOI211_X1 U21365 ( .C1(n18146), .C2(n18145), .A(n18189), .B(n18144), .ZN(
        n18149) );
  OAI22_X1 U21366 ( .A1(n18244), .A2(n18147), .B1(n18591), .B2(n19148), .ZN(
        n18148) );
  AOI211_X1 U21367 ( .C1(n18150), .C2(n18488), .A(n18149), .B(n18148), .ZN(
        n18151) );
  OAI221_X1 U21368 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18153), .C1(
        n18486), .C2(n18152), .A(n18151), .ZN(P3_U2821) );
  AOI21_X1 U21369 ( .B1(n18155), .B2(n18164), .A(n18154), .ZN(n18510) );
  AOI21_X1 U21370 ( .B1(n18156), .B2(n18171), .A(n18226), .ZN(n18172) );
  OAI21_X1 U21371 ( .B1(n18157), .B2(n18636), .A(n18172), .ZN(n18161) );
  OAI22_X1 U21372 ( .A1(n18244), .A2(n18158), .B1(n18591), .B2(n19147), .ZN(
        n18159) );
  AOI221_X1 U21373 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18161), .C1(
        n18160), .C2(n18161), .A(n18159), .ZN(n18167) );
  AOI21_X1 U21374 ( .B1(n18163), .B2(n18502), .A(n18162), .ZN(n18504) );
  INV_X1 U21375 ( .A(n18164), .ZN(n18506) );
  AOI22_X1 U21376 ( .A1(n18248), .A2(n18504), .B1(n18165), .B2(n18506), .ZN(
        n18166) );
  OAI211_X1 U21377 ( .C1(n18510), .C2(n18168), .A(n18167), .B(n18166), .ZN(
        P3_U2822) );
  INV_X1 U21378 ( .A(n18228), .ZN(n18258) );
  OAI21_X1 U21379 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18170), .A(
        n18169), .ZN(n18518) );
  NOR2_X1 U21380 ( .A1(n18636), .A2(n18171), .ZN(n18175) );
  INV_X1 U21381 ( .A(n18172), .ZN(n18173) );
  INV_X1 U21382 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19144) );
  NOR2_X1 U21383 ( .A1(n18491), .A2(n19144), .ZN(n18511) );
  AOI221_X1 U21384 ( .B1(n18175), .B2(n18174), .C1(n18173), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18511), .ZN(n18181) );
  NAND2_X1 U21385 ( .A1(n18177), .A2(n18176), .ZN(n18178) );
  INV_X1 U21386 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18513) );
  XOR2_X1 U21387 ( .A(n18178), .B(n18513), .Z(n18514) );
  AOI22_X1 U21388 ( .A1(n18248), .A2(n18514), .B1(n18179), .B2(n18029), .ZN(
        n18180) );
  OAI211_X1 U21389 ( .C1(n18258), .C2(n18518), .A(n18181), .B(n18180), .ZN(
        P3_U2823) );
  NAND2_X1 U21390 ( .A1(n18981), .A2(n18190), .ZN(n18185) );
  OAI21_X1 U21391 ( .B1(n18184), .B2(n18183), .A(n18182), .ZN(n18527) );
  OAI22_X1 U21392 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18185), .B1(
        n18258), .B2(n18527), .ZN(n18186) );
  AOI21_X1 U21393 ( .B1(n18570), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18186), .ZN(
        n18192) );
  AOI21_X1 U21394 ( .B1(n18188), .B2(n18522), .A(n18187), .ZN(n18524) );
  AOI21_X1 U21395 ( .B1(n18190), .B2(n18981), .A(n18189), .ZN(n18205) );
  AOI22_X1 U21396 ( .A1(n18248), .A2(n18524), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18205), .ZN(n18191) );
  OAI211_X1 U21397 ( .C1(n18244), .C2(n18193), .A(n18192), .B(n18191), .ZN(
        P3_U2824) );
  OAI21_X1 U21398 ( .B1(n18196), .B2(n18195), .A(n18194), .ZN(n18197) );
  XOR2_X1 U21399 ( .A(n18197), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18534) );
  AOI21_X1 U21400 ( .B1(n18200), .B2(n18199), .A(n18198), .ZN(n18528) );
  AOI22_X1 U21401 ( .A1(n18248), .A2(n18528), .B1(n18570), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18207) );
  OAI21_X1 U21402 ( .B1(n18226), .B2(n18202), .A(n18201), .ZN(n18204) );
  AOI22_X1 U21403 ( .A1(n18205), .A2(n18204), .B1(n18203), .B2(n18029), .ZN(
        n18206) );
  OAI211_X1 U21404 ( .C1(n18258), .C2(n18534), .A(n18207), .B(n18206), .ZN(
        P3_U2825) );
  OAI21_X1 U21405 ( .B1(n18210), .B2(n18209), .A(n18208), .ZN(n18211) );
  XOR2_X1 U21406 ( .A(n18211), .B(n18544), .Z(n18541) );
  AOI22_X1 U21407 ( .A1(n18248), .A2(n18541), .B1(n18570), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18220) );
  OAI21_X1 U21408 ( .B1(n18213), .B2(n18212), .A(n18255), .ZN(n18227) );
  OAI21_X1 U21409 ( .B1(n18216), .B2(n18215), .A(n18214), .ZN(n18539) );
  OAI22_X1 U21410 ( .A1(n18244), .A2(n18217), .B1(n18258), .B2(n18539), .ZN(
        n18218) );
  AOI21_X1 U21411 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18227), .A(
        n18218), .ZN(n18219) );
  OAI211_X1 U21412 ( .C1(n18636), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2826) );
  AOI21_X1 U21413 ( .B1(n18224), .B2(n18223), .A(n18222), .ZN(n18554) );
  AOI22_X1 U21414 ( .A1(n18248), .A2(n18554), .B1(n18225), .B2(n18029), .ZN(
        n18231) );
  NOR2_X1 U21415 ( .A1(n18226), .A2(n18236), .ZN(n18235) );
  OAI21_X1 U21416 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18235), .A(
        n18227), .ZN(n18230) );
  NAND2_X1 U21417 ( .A1(n18570), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18551) );
  OAI211_X1 U21418 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18547), .A(
        n18228), .B(n18546), .ZN(n18229) );
  NAND4_X1 U21419 ( .A1(n18231), .A2(n18230), .A3(n18551), .A4(n18229), .ZN(
        P3_U2827) );
  AOI21_X1 U21420 ( .B1(n18234), .B2(n18233), .A(n18232), .ZN(n18563) );
  AOI21_X1 U21421 ( .B1(n18636), .B2(n18236), .A(n18235), .ZN(n18241) );
  OAI21_X1 U21422 ( .B1(n18239), .B2(n18238), .A(n18237), .ZN(n18573) );
  OAI22_X1 U21423 ( .A1(n18258), .A2(n18573), .B1(n18591), .B2(n19134), .ZN(
        n18240) );
  AOI211_X1 U21424 ( .C1(n18563), .C2(n18248), .A(n18241), .B(n18240), .ZN(
        n18242) );
  OAI21_X1 U21425 ( .B1(n18244), .B2(n18243), .A(n18242), .ZN(P3_U2828) );
  OAI21_X1 U21426 ( .B1(n18246), .B2(n18253), .A(n18245), .ZN(n18585) );
  NAND2_X1 U21427 ( .A1(n19232), .A2(n18254), .ZN(n18247) );
  XNOR2_X1 U21428 ( .A(n18247), .B(n18246), .ZN(n18580) );
  AOI22_X1 U21429 ( .A1(n18248), .A2(n18580), .B1(n18581), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U21430 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18250), .B1(
        n18029), .B2(n18249), .ZN(n18251) );
  OAI211_X1 U21431 ( .C1(n18258), .C2(n18585), .A(n18252), .B(n18251), .ZN(
        P3_U2829) );
  AOI21_X1 U21432 ( .B1(n18254), .B2(n19232), .A(n18253), .ZN(n18589) );
  INV_X1 U21433 ( .A(n18589), .ZN(n18587) );
  NAND3_X1 U21434 ( .A1(n19216), .A2(n19113), .A3(n18255), .ZN(n18256) );
  AOI22_X1 U21435 ( .A1(n18581), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18256), .ZN(n18257) );
  OAI221_X1 U21436 ( .B1(n18589), .B2(n18259), .C1(n18587), .C2(n18258), .A(
        n18257), .ZN(P3_U2830) );
  NOR2_X1 U21437 ( .A1(n18260), .A2(n18264), .ZN(n18336) );
  NAND2_X1 U21438 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18336), .ZN(
        n18318) );
  NOR2_X1 U21439 ( .A1(n18261), .A2(n18318), .ZN(n18274) );
  NOR2_X1 U21440 ( .A1(n18593), .A2(n19070), .ZN(n18497) );
  INV_X1 U21441 ( .A(n18497), .ZN(n18557) );
  AOI221_X1 U21442 ( .B1(n18325), .B2(n19070), .C1(n18263), .C2(n19070), .A(
        n18262), .ZN(n18327) );
  NOR2_X1 U21443 ( .A1(n18264), .A2(n18391), .ZN(n18265) );
  AOI21_X1 U21444 ( .B1(n18327), .B2(n18265), .A(n18497), .ZN(n18307) );
  AOI21_X1 U21445 ( .B1(n18266), .B2(n18557), .A(n18307), .ZN(n18295) );
  AOI22_X1 U21446 ( .A1(n19035), .A2(n18268), .B1(n18461), .B2(n18267), .ZN(
        n18269) );
  NAND2_X1 U21447 ( .A1(n18295), .A2(n18269), .ZN(n18270) );
  AOI211_X1 U21448 ( .C1(n18272), .C2(n18557), .A(n18271), .B(n18270), .ZN(
        n18283) );
  INV_X1 U21449 ( .A(n18283), .ZN(n18273) );
  MUX2_X1 U21450 ( .A(n18274), .B(n18273), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18275) );
  AOI22_X1 U21451 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18569), .B1(
        n18575), .B2(n18275), .ZN(n18277) );
  NAND2_X1 U21452 ( .A1(n18581), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18276) );
  OAI211_X1 U21453 ( .C1(n18278), .C2(n18509), .A(n18277), .B(n18276), .ZN(
        P3_U2835) );
  NAND2_X1 U21454 ( .A1(n18280), .A2(n18279), .ZN(n18317) );
  INV_X1 U21455 ( .A(n18281), .ZN(n18285) );
  AOI211_X1 U21456 ( .C1(n18575), .C2(n18283), .A(n18581), .B(n18282), .ZN(
        n18284) );
  AOI21_X1 U21457 ( .B1(n18489), .B2(n18285), .A(n18284), .ZN(n18287) );
  NAND2_X1 U21458 ( .A1(n18581), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18286) );
  OAI211_X1 U21459 ( .C1(n18288), .C2(n18317), .A(n18287), .B(n18286), .ZN(
        P3_U2836) );
  NOR2_X1 U21460 ( .A1(n18591), .A2(n19181), .ZN(n18297) );
  AOI221_X1 U21461 ( .B1(n18290), .B2(n19051), .C1(n18328), .C2(n19051), .A(
        n18289), .ZN(n18294) );
  AOI21_X1 U21462 ( .B1(n18292), .B2(n18291), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18293) );
  AOI211_X1 U21463 ( .C1(n18295), .C2(n18294), .A(n18293), .B(n18592), .ZN(
        n18296) );
  AOI211_X1 U21464 ( .C1(n18569), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18297), .B(n18296), .ZN(n18301) );
  AOI22_X1 U21465 ( .A1(n18588), .A2(n18299), .B1(n18489), .B2(n18298), .ZN(
        n18300) );
  OAI211_X1 U21466 ( .C1(n18429), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2837) );
  OAI22_X1 U21467 ( .A1(n18305), .A2(n18304), .B1(n18303), .B2(n18438), .ZN(
        n18306) );
  NOR3_X1 U21468 ( .A1(n18569), .A2(n18307), .A3(n18306), .ZN(n18311) );
  OAI211_X1 U21469 ( .C1(n18308), .C2(n19068), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18311), .ZN(n18309) );
  AND2_X1 U21470 ( .A1(n18491), .A2(n18309), .ZN(n18319) );
  AOI21_X1 U21471 ( .B1(n18312), .B2(n18311), .A(n18310), .ZN(n18313) );
  AOI22_X1 U21472 ( .A1(n18489), .A2(n18314), .B1(n18319), .B2(n18313), .ZN(
        n18316) );
  OAI211_X1 U21473 ( .C1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n18317), .A(
        n18316), .B(n18315), .ZN(P3_U2838) );
  NOR2_X1 U21474 ( .A1(n18569), .A2(n18318), .ZN(n18320) );
  OAI21_X1 U21475 ( .B1(n18320), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18319), .ZN(n18321) );
  OAI211_X1 U21476 ( .C1(n18323), .C2(n18509), .A(n18322), .B(n18321), .ZN(
        P3_U2839) );
  AOI22_X1 U21477 ( .A1(n19035), .A2(n18410), .B1(n18461), .B2(n18324), .ZN(
        n18351) );
  AOI22_X1 U21478 ( .A1(n19051), .A2(n18325), .B1(n18593), .B2(n18344), .ZN(
        n18326) );
  NAND3_X1 U21479 ( .A1(n18327), .A2(n18351), .A3(n18326), .ZN(n18335) );
  NOR2_X1 U21480 ( .A1(n19035), .A2(n18461), .ZN(n18464) );
  NAND2_X1 U21481 ( .A1(n19051), .A2(n18328), .ZN(n18374) );
  OAI21_X1 U21482 ( .B1(n18391), .B2(n18329), .A(n18593), .ZN(n18330) );
  OAI211_X1 U21483 ( .C1(n18331), .C2(n19068), .A(n18374), .B(n18330), .ZN(
        n18354) );
  AOI21_X1 U21484 ( .B1(n18593), .B2(n18332), .A(n18354), .ZN(n18333) );
  OAI21_X1 U21485 ( .B1(n18334), .B2(n18464), .A(n18333), .ZN(n18342) );
  OAI22_X1 U21486 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18336), .B1(
        n18335), .B2(n18342), .ZN(n18340) );
  AOI22_X1 U21487 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18569), .B1(
        n18489), .B2(n18337), .ZN(n18339) );
  OAI211_X1 U21488 ( .C1(n18592), .C2(n18340), .A(n18339), .B(n18338), .ZN(
        P3_U2840) );
  INV_X1 U21489 ( .A(n18341), .ZN(n18347) );
  NAND2_X1 U21490 ( .A1(n19047), .A2(n19068), .ZN(n18574) );
  NAND2_X1 U21491 ( .A1(n18575), .A2(n18351), .ZN(n18394) );
  AOI211_X1 U21492 ( .C1(n18343), .C2(n18574), .A(n18394), .B(n18342), .ZN(
        n18345) );
  AOI211_X1 U21493 ( .C1(n18345), .C2(n18355), .A(n18581), .B(n18344), .ZN(
        n18346) );
  AOI21_X1 U21494 ( .B1(n18489), .B2(n18347), .A(n18346), .ZN(n18349) );
  OAI211_X1 U21495 ( .C1(n18350), .C2(n18366), .A(n18349), .B(n18348), .ZN(
        P3_U2841) );
  OAI211_X1 U21496 ( .C1(n18352), .C2(n18464), .A(n18351), .B(n18576), .ZN(
        n18353) );
  NOR2_X1 U21497 ( .A1(n18354), .A2(n18353), .ZN(n18356) );
  AOI21_X1 U21498 ( .B1(n18356), .B2(n18355), .A(n18570), .ZN(n18357) );
  NOR2_X1 U21499 ( .A1(n18357), .A2(n18367), .ZN(n18368) );
  AOI21_X1 U21500 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18574), .A(n18357), 
        .ZN(n18358) );
  NOR2_X1 U21501 ( .A1(n18368), .A2(n18358), .ZN(n18360) );
  AOI22_X1 U21502 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18360), .B1(
        n18489), .B2(n18359), .ZN(n18362) );
  NAND2_X1 U21503 ( .A1(n18581), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18361) );
  OAI211_X1 U21504 ( .C1(n18363), .C2(n18366), .A(n18362), .B(n18361), .ZN(
        P3_U2842) );
  AOI22_X1 U21505 ( .A1(n18581), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18489), 
        .B2(n18364), .ZN(n18365) );
  OAI221_X1 U21506 ( .B1(n18368), .B2(n18367), .C1(n18368), .C2(n18366), .A(
        n18365), .ZN(P3_U2843) );
  NAND2_X1 U21507 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18535) );
  OAI22_X1 U21508 ( .A1(n18536), .A2(n19068), .B1(n18535), .B2(n18560), .ZN(
        n18549) );
  NAND2_X1 U21509 ( .A1(n18369), .A2(n18549), .ZN(n18521) );
  NOR2_X1 U21510 ( .A1(n18370), .A2(n18521), .ZN(n18400) );
  NOR2_X1 U21511 ( .A1(n18400), .A2(n18371), .ZN(n18450) );
  NAND2_X1 U21512 ( .A1(n18372), .A2(n18487), .ZN(n18399) );
  NAND2_X1 U21513 ( .A1(n19070), .A2(n19232), .ZN(n18565) );
  NAND3_X1 U21514 ( .A1(n18373), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18565), .ZN(n18377) );
  AOI22_X1 U21515 ( .A1(n18375), .A2(n18374), .B1(n18464), .B2(n19068), .ZN(
        n18376) );
  AOI211_X1 U21516 ( .C1(n18557), .C2(n18377), .A(n18376), .B(n18394), .ZN(
        n18384) );
  AOI221_X1 U21517 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18384), 
        .C1(n18497), .C2(n18384), .A(n18581), .ZN(n18379) );
  AOI22_X1 U21518 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18379), .B1(
        n18489), .B2(n18378), .ZN(n18381) );
  NAND2_X1 U21519 ( .A1(n18581), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18380) );
  OAI211_X1 U21520 ( .C1(n18382), .C2(n18399), .A(n18381), .B(n18380), .ZN(
        P3_U2844) );
  NOR3_X1 U21521 ( .A1(n18581), .A2(n18384), .A3(n18383), .ZN(n18385) );
  AOI211_X1 U21522 ( .C1(n18489), .C2(n18387), .A(n18386), .B(n18385), .ZN(
        n18388) );
  OAI21_X1 U21523 ( .B1(n18399), .B2(n18389), .A(n18388), .ZN(P3_U2845) );
  OAI21_X1 U21524 ( .B1(n18493), .B2(n18498), .A(n18593), .ZN(n18418) );
  INV_X1 U21525 ( .A(n18418), .ZN(n18390) );
  NOR2_X1 U21526 ( .A1(n18416), .A2(n19068), .ZN(n18467) );
  NOR2_X1 U21527 ( .A1(n18390), .A2(n18467), .ZN(n18482) );
  INV_X1 U21528 ( .A(n18593), .ZN(n19072) );
  OAI21_X1 U21529 ( .B1(n19072), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n19047), .ZN(n18484) );
  OAI22_X1 U21530 ( .A1(n19232), .A2(n18391), .B1(n18401), .B2(n18484), .ZN(
        n18392) );
  OAI211_X1 U21531 ( .C1(n18475), .C2(n18393), .A(n18482), .B(n18392), .ZN(
        n18407) );
  OAI221_X1 U21532 ( .B1(n18394), .B2(n18499), .C1(n18394), .C2(n18407), .A(
        n18491), .ZN(n18397) );
  AOI22_X1 U21533 ( .A1(n18581), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18489), 
        .B2(n18395), .ZN(n18396) );
  OAI221_X1 U21534 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18399), 
        .C1(n18398), .C2(n18397), .A(n18396), .ZN(P3_U2846) );
  NAND2_X1 U21535 ( .A1(n18422), .A2(n18400), .ZN(n18424) );
  OAI21_X1 U21536 ( .B1(n18426), .B2(n18424), .A(n18401), .ZN(n18408) );
  NOR2_X1 U21537 ( .A1(n18402), .A2(n18438), .ZN(n18403) );
  AOI222_X1 U21538 ( .A1(n18408), .A2(n18407), .B1(n18406), .B2(n18405), .C1(
        n18404), .C2(n18403), .ZN(n18413) );
  AOI22_X1 U21539 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18569), .B1(
        n18581), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18412) );
  NAND3_X1 U21540 ( .A1(n18588), .A2(n18410), .A3(n18409), .ZN(n18411) );
  OAI211_X1 U21541 ( .C1(n18413), .C2(n18592), .A(n18412), .B(n18411), .ZN(
        P3_U2847) );
  NAND2_X1 U21542 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18414), .ZN(
        n18483) );
  NOR2_X1 U21543 ( .A1(n18415), .A2(n18483), .ZN(n18453) );
  NOR2_X1 U21544 ( .A1(n19047), .A2(n18453), .ZN(n18443) );
  AOI21_X1 U21545 ( .B1(n18417), .B2(n18416), .A(n19068), .ZN(n18419) );
  OAI21_X1 U21546 ( .B1(n19072), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n18418), .ZN(n18477) );
  AOI211_X1 U21547 ( .C1(n18420), .C2(n18574), .A(n18419), .B(n18477), .ZN(
        n18421) );
  OAI211_X1 U21548 ( .C1(n19072), .C2(n18422), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18421), .ZN(n18423) );
  OAI21_X1 U21549 ( .B1(n18443), .B2(n18423), .A(n18575), .ZN(n18425) );
  AOI222_X1 U21550 ( .A1(n18426), .A2(n18425), .B1(n18426), .B2(n18424), .C1(
        n18425), .C2(n18576), .ZN(n18432) );
  INV_X1 U21551 ( .A(n18427), .ZN(n18430) );
  OAI22_X1 U21552 ( .A1(n18430), .A2(n18509), .B1(n18429), .B2(n18428), .ZN(
        n18431) );
  AOI211_X1 U21553 ( .C1(n18570), .C2(P3_REIP_REG_14__SCAN_IN), .A(n18432), 
        .B(n18431), .ZN(n18433) );
  OAI21_X1 U21554 ( .B1(n18435), .B2(n18434), .A(n18433), .ZN(P3_U2848) );
  AOI21_X1 U21555 ( .B1(n18593), .B2(n18436), .A(n18449), .ZN(n18452) );
  NOR2_X1 U21556 ( .A1(n19072), .A2(n18465), .ZN(n18437) );
  AOI211_X1 U21557 ( .C1(n19051), .C2(n18448), .A(n18437), .B(n18477), .ZN(
        n18468) );
  OAI21_X1 U21558 ( .B1(n18439), .B2(n18438), .A(n18468), .ZN(n18440) );
  AOI211_X1 U21559 ( .C1(n19035), .C2(n18441), .A(n18467), .B(n18440), .ZN(
        n18451) );
  OAI211_X1 U21560 ( .C1(n18475), .C2(n18452), .A(n18575), .B(n18451), .ZN(
        n18442) );
  OAI21_X1 U21561 ( .B1(n18443), .B2(n18442), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18447) );
  AOI22_X1 U21562 ( .A1(n18489), .A2(n18445), .B1(n18487), .B2(n18444), .ZN(
        n18446) );
  OAI221_X1 U21563 ( .B1(n18570), .B2(n18447), .C1(n18491), .C2(n19156), .A(
        n18446), .ZN(P3_U2849) );
  AOI221_X1 U21564 ( .B1(n18450), .B2(n18449), .C1(n18448), .C2(n18449), .A(
        n18592), .ZN(n18455) );
  OAI211_X1 U21565 ( .C1(n18453), .C2(n19047), .A(n18452), .B(n18451), .ZN(
        n18454) );
  AOI22_X1 U21566 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18569), .B1(
        n18455), .B2(n18454), .ZN(n18457) );
  OAI211_X1 U21567 ( .C1(n18458), .C2(n18509), .A(n18457), .B(n18456), .ZN(
        P3_U2850) );
  AOI22_X1 U21568 ( .A1(n18581), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18487), 
        .B2(n18459), .ZN(n18471) );
  AOI22_X1 U21569 ( .A1(n19035), .A2(n18462), .B1(n18461), .B2(n18460), .ZN(
        n18481) );
  OAI21_X1 U21570 ( .B1(n18486), .B2(n18483), .A(n19070), .ZN(n18463) );
  OAI211_X1 U21571 ( .C1(n18465), .C2(n18464), .A(n18481), .B(n18463), .ZN(
        n18466) );
  NOR3_X1 U21572 ( .A1(n18467), .A2(n18592), .A3(n18466), .ZN(n18474) );
  OAI211_X1 U21573 ( .C1(n19047), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18468), .B(n18474), .ZN(n18469) );
  NAND3_X1 U21574 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18491), .A3(
        n18469), .ZN(n18470) );
  OAI211_X1 U21575 ( .C1(n18472), .C2(n18509), .A(n18471), .B(n18470), .ZN(
        P3_U2851) );
  NOR2_X1 U21576 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18486), .ZN(
        n18473) );
  AOI22_X1 U21577 ( .A1(n18581), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18487), 
        .B2(n18473), .ZN(n18479) );
  OAI21_X1 U21578 ( .B1(n18475), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18474), .ZN(n18476) );
  OAI211_X1 U21579 ( .C1(n18477), .C2(n18476), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18591), .ZN(n18478) );
  OAI211_X1 U21580 ( .C1(n18480), .C2(n18509), .A(n18479), .B(n18478), .ZN(
        P3_U2852) );
  NAND3_X1 U21581 ( .A1(n18482), .A2(n18481), .A3(n18576), .ZN(n18485) );
  OAI221_X1 U21582 ( .B1(n18485), .B2(n18484), .C1(n18485), .C2(n18483), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18492) );
  AOI22_X1 U21583 ( .A1(n18489), .A2(n18488), .B1(n18487), .B2(n18486), .ZN(
        n18490) );
  OAI221_X1 U21584 ( .B1(n18570), .B2(n18492), .C1(n18491), .C2(n19148), .A(
        n18490), .ZN(P3_U2853) );
  NOR3_X1 U21585 ( .A1(n18592), .A2(n18498), .A3(n18521), .ZN(n18503) );
  INV_X1 U21586 ( .A(n18493), .ZN(n18496) );
  NAND2_X1 U21587 ( .A1(n19051), .A2(n18494), .ZN(n18495) );
  OAI211_X1 U21588 ( .C1(n18497), .C2(n18496), .A(n18565), .B(n18495), .ZN(
        n18519) );
  AOI21_X1 U21589 ( .B1(n18499), .B2(n18498), .A(n18519), .ZN(n18512) );
  OAI21_X1 U21590 ( .B1(n18512), .B2(n18577), .A(n18576), .ZN(n18501) );
  NOR2_X1 U21591 ( .A1(n18591), .A2(n19147), .ZN(n18500) );
  AOI221_X1 U21592 ( .B1(n18503), .B2(n18502), .C1(n18501), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18500), .ZN(n18508) );
  AOI22_X1 U21593 ( .A1(n18506), .A2(n18505), .B1(n18588), .B2(n18504), .ZN(
        n18507) );
  OAI211_X1 U21594 ( .C1(n18510), .C2(n18509), .A(n18508), .B(n18507), .ZN(
        P3_U2854) );
  INV_X1 U21595 ( .A(n18590), .ZN(n18584) );
  AOI21_X1 U21596 ( .B1(n18569), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18511), .ZN(n18517) );
  AOI221_X1 U21597 ( .B1(n18522), .B2(n18513), .C1(n18521), .C2(n18513), .A(
        n18512), .ZN(n18515) );
  AOI22_X1 U21598 ( .A1(n18575), .A2(n18515), .B1(n18588), .B2(n18514), .ZN(
        n18516) );
  OAI211_X1 U21599 ( .C1(n18584), .C2(n18518), .A(n18517), .B(n18516), .ZN(
        P3_U2855) );
  AOI21_X1 U21600 ( .B1(n18519), .B2(n18575), .A(n18569), .ZN(n18520) );
  INV_X1 U21601 ( .A(n18520), .ZN(n18531) );
  AOI22_X1 U21602 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18531), .B1(
        n18570), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18526) );
  NOR2_X1 U21603 ( .A1(n18592), .A2(n18521), .ZN(n18523) );
  AOI22_X1 U21604 ( .A1(n18524), .A2(n18588), .B1(n18523), .B2(n18522), .ZN(
        n18525) );
  OAI211_X1 U21605 ( .C1(n18584), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        P3_U2856) );
  AOI22_X1 U21606 ( .A1(n18581), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18588), 
        .B2(n18528), .ZN(n18533) );
  NAND3_X1 U21607 ( .A1(n18575), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18549), .ZN(n18545) );
  NOR2_X1 U21608 ( .A1(n18544), .A2(n18545), .ZN(n18530) );
  AOI22_X1 U21609 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18531), .B1(
        n18530), .B2(n18529), .ZN(n18532) );
  OAI211_X1 U21610 ( .C1(n18584), .C2(n18534), .A(n18533), .B(n18532), .ZN(
        P3_U2857) );
  AOI22_X1 U21611 ( .A1(n19051), .A2(n18536), .B1(n18535), .B2(n18557), .ZN(
        n18537) );
  NAND3_X1 U21612 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18537), .A3(
        n18565), .ZN(n18548) );
  AOI21_X1 U21613 ( .B1(n18538), .B2(n18548), .A(n18569), .ZN(n18543) );
  OAI22_X1 U21614 ( .A1(n18591), .A2(n19138), .B1(n18584), .B2(n18539), .ZN(
        n18540) );
  AOI21_X1 U21615 ( .B1(n18588), .B2(n18541), .A(n18540), .ZN(n18542) );
  OAI221_X1 U21616 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18545), .C1(
        n18544), .C2(n18543), .A(n18542), .ZN(P3_U2858) );
  OAI21_X1 U21617 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18547), .A(
        n18546), .ZN(n18552) );
  OAI211_X1 U21618 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18549), .A(
        n18575), .B(n18548), .ZN(n18550) );
  OAI211_X1 U21619 ( .C1(n18584), .C2(n18552), .A(n18551), .B(n18550), .ZN(
        n18553) );
  AOI21_X1 U21620 ( .B1(n18588), .B2(n18554), .A(n18553), .ZN(n18555) );
  OAI21_X1 U21621 ( .B1(n18556), .B2(n18576), .A(n18555), .ZN(P3_U2859) );
  INV_X1 U21622 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19217) );
  NOR2_X1 U21623 ( .A1(n19232), .A2(n19217), .ZN(n18558) );
  AOI22_X1 U21624 ( .A1(n19051), .A2(n18558), .B1(n19217), .B2(n18557), .ZN(
        n18566) );
  NOR2_X1 U21625 ( .A1(n19068), .A2(n18559), .ZN(n18562) );
  NOR3_X1 U21626 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19217), .A3(
        n18560), .ZN(n18561) );
  AOI211_X1 U21627 ( .C1(n18563), .C2(n19035), .A(n18562), .B(n18561), .ZN(
        n18564) );
  OAI221_X1 U21628 ( .B1(n18567), .B2(n18566), .C1(n18567), .C2(n18565), .A(
        n18564), .ZN(n18568) );
  AOI22_X1 U21629 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18569), .B1(
        n18575), .B2(n18568), .ZN(n18572) );
  NAND2_X1 U21630 ( .A1(n18570), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18571) );
  OAI211_X1 U21631 ( .C1(n18584), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2860) );
  NAND3_X1 U21632 ( .A1(n18575), .A2(n19232), .A3(n18574), .ZN(n18595) );
  AOI21_X1 U21633 ( .B1(n18576), .B2(n18595), .A(n19217), .ZN(n18579) );
  AOI211_X1 U21634 ( .C1(n19072), .C2(n19232), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18577), .ZN(n18578) );
  AOI211_X1 U21635 ( .C1(n18588), .C2(n18580), .A(n18579), .B(n18578), .ZN(
        n18583) );
  NAND2_X1 U21636 ( .A1(n18581), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18582) );
  OAI211_X1 U21637 ( .C1(n18585), .C2(n18584), .A(n18583), .B(n18582), .ZN(
        P3_U2861) );
  INV_X1 U21638 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19243) );
  NOR2_X1 U21639 ( .A1(n18591), .A2(n19243), .ZN(n18586) );
  AOI221_X1 U21640 ( .B1(n18590), .B2(n18589), .C1(n18588), .C2(n18587), .A(
        n18586), .ZN(n18596) );
  OAI211_X1 U21641 ( .C1(n18593), .C2(n18592), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18591), .ZN(n18594) );
  NAND3_X1 U21642 ( .A1(n18596), .A2(n18595), .A3(n18594), .ZN(P3_U2862) );
  INV_X1 U21643 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18895) );
  AOI211_X1 U21644 ( .C1(n18598), .C2(n18597), .A(n19268), .B(n19216), .ZN(
        n19095) );
  OAI21_X1 U21645 ( .B1(n19095), .B2(n18646), .A(n18603), .ZN(n18599) );
  OAI221_X1 U21646 ( .B1(n18895), .B2(n19250), .C1(n18895), .C2(n18603), .A(
        n18599), .ZN(P3_U2863) );
  INV_X1 U21647 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19084) );
  NAND2_X1 U21648 ( .A1(n19081), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18872) );
  INV_X1 U21649 ( .A(n18872), .ZN(n18896) );
  NAND2_X1 U21650 ( .A1(n19084), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18778) );
  INV_X1 U21651 ( .A(n18778), .ZN(n18777) );
  NOR2_X1 U21652 ( .A1(n18896), .A2(n18777), .ZN(n18601) );
  OAI22_X1 U21653 ( .A1(n18602), .A2(n19084), .B1(n18601), .B2(n18600), .ZN(
        P3_U2866) );
  NOR2_X1 U21654 ( .A1(n19085), .A2(n18603), .ZN(P3_U2867) );
  NAND2_X1 U21655 ( .A1(n18981), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18985) );
  NAND2_X1 U21656 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18606) );
  NAND2_X1 U21657 ( .A1(n18895), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18846) );
  NOR2_X2 U21658 ( .A1(n18606), .A2(n18846), .ZN(n18969) );
  INV_X1 U21659 ( .A(n18969), .ZN(n18966) );
  NOR2_X1 U21660 ( .A1(n18606), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18980) );
  NAND2_X1 U21661 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18980), .ZN(
        n19034) );
  INV_X1 U21662 ( .A(n19034), .ZN(n19018) );
  NOR2_X2 U21663 ( .A1(n18604), .A2(n18636), .ZN(n18977) );
  NOR2_X2 U21664 ( .A1(n18947), .A2(n18605), .ZN(n18976) );
  NAND2_X1 U21665 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19075) );
  NOR2_X2 U21666 ( .A1(n19075), .A2(n18606), .ZN(n19029) );
  INV_X1 U21667 ( .A(n19029), .ZN(n19023) );
  NAND2_X1 U21668 ( .A1(n19076), .A2(n18895), .ZN(n19077) );
  NAND2_X1 U21669 ( .A1(n19081), .A2(n19084), .ZN(n18731) );
  NOR2_X2 U21670 ( .A1(n19077), .A2(n18731), .ZN(n18704) );
  INV_X1 U21671 ( .A(n18704), .ZN(n18686) );
  INV_X1 U21672 ( .A(n18975), .ZN(n19103) );
  AOI21_X1 U21673 ( .B1(n19023), .B2(n18686), .A(n19103), .ZN(n18640) );
  AOI22_X1 U21674 ( .A1(n19018), .A2(n18977), .B1(n18976), .B2(n18640), .ZN(
        n18612) );
  NAND2_X1 U21675 ( .A1(n19076), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18730) );
  AND2_X1 U21676 ( .A1(n18846), .A2(n18730), .ZN(n18899) );
  NOR2_X1 U21677 ( .A1(n18899), .A2(n18606), .ZN(n18945) );
  AOI21_X1 U21678 ( .B1(n19023), .B2(n18686), .A(n18947), .ZN(n18666) );
  NAND2_X1 U21679 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18607) );
  AOI22_X1 U21680 ( .A1(n18981), .A2(n18945), .B1(n18666), .B2(n18607), .ZN(
        n18643) );
  NAND2_X1 U21681 ( .A1(n18609), .A2(n18608), .ZN(n18641) );
  INV_X1 U21682 ( .A(n18641), .ZN(n18633) );
  NAND2_X1 U21683 ( .A1(n18610), .A2(n18633), .ZN(n18853) );
  INV_X1 U21684 ( .A(n18853), .ZN(n18982) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18643), .B1(
        n18704), .B2(n18982), .ZN(n18611) );
  OAI211_X1 U21686 ( .C1(n18985), .C2(n18966), .A(n18612), .B(n18611), .ZN(
        P3_U2868) );
  NAND2_X1 U21687 ( .A1(n18981), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18991) );
  NAND2_X1 U21688 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18981), .ZN(n18878) );
  INV_X1 U21689 ( .A(n18878), .ZN(n18987) );
  INV_X1 U21690 ( .A(n18947), .ZN(n18901) );
  AND2_X1 U21691 ( .A1(n18901), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18986) );
  AOI22_X1 U21692 ( .A1(n19018), .A2(n18987), .B1(n18640), .B2(n18986), .ZN(
        n18614) );
  NOR2_X2 U21693 ( .A1(n19256), .A2(n18641), .ZN(n18988) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18643), .B1(
        n18704), .B2(n18988), .ZN(n18613) );
  OAI211_X1 U21695 ( .C1(n18966), .C2(n18991), .A(n18614), .B(n18613), .ZN(
        P3_U2869) );
  NAND2_X1 U21696 ( .A1(n18981), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18997) );
  NAND2_X1 U21697 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18981), .ZN(n18931) );
  INV_X1 U21698 ( .A(n18931), .ZN(n18992) );
  NOR2_X2 U21699 ( .A1(n18947), .A2(n18615), .ZN(n18993) );
  AOI22_X1 U21700 ( .A1(n19018), .A2(n18992), .B1(n18640), .B2(n18993), .ZN(
        n18618) );
  NOR2_X2 U21701 ( .A1(n18616), .A2(n18641), .ZN(n18994) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18643), .B1(
        n18704), .B2(n18994), .ZN(n18617) );
  OAI211_X1 U21703 ( .C1(n18966), .C2(n18997), .A(n18618), .B(n18617), .ZN(
        P3_U2870) );
  NAND2_X1 U21704 ( .A1(n18633), .A2(n18619), .ZN(n19003) );
  AND2_X1 U21705 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n18981), .ZN(n18999) );
  NOR2_X2 U21706 ( .A1(n18620), .A2(n18947), .ZN(n18998) );
  AOI22_X1 U21707 ( .A1(n18969), .A2(n18999), .B1(n18640), .B2(n18998), .ZN(
        n18622) );
  NOR2_X2 U21708 ( .A1(n15341), .A2(n18636), .ZN(n19000) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18643), .B1(
        n19018), .B2(n19000), .ZN(n18621) );
  OAI211_X1 U21710 ( .C1(n18686), .C2(n19003), .A(n18622), .B(n18621), .ZN(
        P3_U2871) );
  NAND2_X1 U21711 ( .A1(n18633), .A2(n18623), .ZN(n19009) );
  AND2_X1 U21712 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18981), .ZN(n19005) );
  NOR2_X2 U21713 ( .A1(n18624), .A2(n18947), .ZN(n19004) );
  AOI22_X1 U21714 ( .A1(n18969), .A2(n19005), .B1(n18640), .B2(n19004), .ZN(
        n18626) );
  NOR2_X2 U21715 ( .A1(n15333), .A2(n18636), .ZN(n19006) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18643), .B1(
        n19018), .B2(n19006), .ZN(n18625) );
  OAI211_X1 U21717 ( .C1(n18686), .C2(n19009), .A(n18626), .B(n18625), .ZN(
        P3_U2872) );
  NAND2_X1 U21718 ( .A1(n18633), .A2(n18627), .ZN(n19015) );
  AND2_X1 U21719 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18981), .ZN(n19012) );
  NOR2_X2 U21720 ( .A1(n18628), .A2(n18947), .ZN(n19010) );
  AOI22_X1 U21721 ( .A1(n18969), .A2(n19012), .B1(n18640), .B2(n19010), .ZN(
        n18631) );
  INV_X1 U21722 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18629) );
  NOR2_X2 U21723 ( .A1(n18629), .A2(n18636), .ZN(n19011) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18643), .B1(
        n19018), .B2(n19011), .ZN(n18630) );
  OAI211_X1 U21725 ( .C1(n18686), .C2(n19015), .A(n18631), .B(n18630), .ZN(
        P3_U2873) );
  NAND2_X1 U21726 ( .A1(n18633), .A2(n18632), .ZN(n19022) );
  NOR2_X2 U21727 ( .A1(n18634), .A2(n18636), .ZN(n19017) );
  NOR2_X2 U21728 ( .A1(n18635), .A2(n18947), .ZN(n19016) );
  AOI22_X1 U21729 ( .A1(n18969), .A2(n19017), .B1(n18640), .B2(n19016), .ZN(
        n18638) );
  NOR2_X2 U21730 ( .A1(n12670), .A2(n18636), .ZN(n19019) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18643), .B1(
        n19018), .B2(n19019), .ZN(n18637) );
  OAI211_X1 U21732 ( .C1(n18686), .C2(n19022), .A(n18638), .B(n18637), .ZN(
        P3_U2874) );
  NAND2_X1 U21733 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18981), .ZN(n19033) );
  NAND2_X1 U21734 ( .A1(n18981), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18974) );
  INV_X1 U21735 ( .A(n18974), .ZN(n19027) );
  NOR2_X2 U21736 ( .A1(n18639), .A2(n18947), .ZN(n19025) );
  AOI22_X1 U21737 ( .A1(n19018), .A2(n19027), .B1(n18640), .B2(n19025), .ZN(
        n18645) );
  NOR2_X2 U21738 ( .A1(n18642), .A2(n18641), .ZN(n19028) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18643), .B1(
        n18704), .B2(n19028), .ZN(n18644) );
  OAI211_X1 U21740 ( .C1(n18966), .C2(n19033), .A(n18645), .B(n18644), .ZN(
        P3_U2875) );
  NAND2_X1 U21741 ( .A1(n19076), .A2(n18975), .ZN(n18821) );
  NOR2_X1 U21742 ( .A1(n18731), .A2(n18821), .ZN(n18661) );
  AOI22_X1 U21743 ( .A1(n18969), .A2(n18977), .B1(n18976), .B2(n18661), .ZN(
        n18648) );
  NOR2_X1 U21744 ( .A1(n19084), .A2(n18822), .ZN(n18978) );
  INV_X1 U21745 ( .A(n18731), .ZN(n18688) );
  NOR2_X1 U21746 ( .A1(n18947), .A2(n18646), .ZN(n18979) );
  INV_X1 U21747 ( .A(n18979), .ZN(n18687) );
  NOR2_X1 U21748 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18687), .ZN(
        n18732) );
  AOI22_X1 U21749 ( .A1(n18981), .A2(n18978), .B1(n18688), .B2(n18732), .ZN(
        n18662) );
  INV_X1 U21750 ( .A(n18730), .ZN(n18825) );
  NAND2_X1 U21751 ( .A1(n18688), .A2(n18825), .ZN(n18729) );
  INV_X1 U21752 ( .A(n18729), .ZN(n18722) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18662), .B1(
        n18982), .B2(n18722), .ZN(n18647) );
  OAI211_X1 U21754 ( .C1(n18985), .C2(n19023), .A(n18648), .B(n18647), .ZN(
        P3_U2876) );
  INV_X1 U21755 ( .A(n18991), .ZN(n18875) );
  AOI22_X1 U21756 ( .A1(n19029), .A2(n18875), .B1(n18986), .B2(n18661), .ZN(
        n18650) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18662), .B1(
        n18988), .B2(n18722), .ZN(n18649) );
  OAI211_X1 U21758 ( .C1(n18966), .C2(n18878), .A(n18650), .B(n18649), .ZN(
        P3_U2877) );
  INV_X1 U21759 ( .A(n18997), .ZN(n18927) );
  AOI22_X1 U21760 ( .A1(n19029), .A2(n18927), .B1(n18993), .B2(n18661), .ZN(
        n18652) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18662), .B1(
        n18994), .B2(n18722), .ZN(n18651) );
  OAI211_X1 U21762 ( .C1(n18966), .C2(n18931), .A(n18652), .B(n18651), .ZN(
        P3_U2878) );
  AOI22_X1 U21763 ( .A1(n18969), .A2(n19000), .B1(n18998), .B2(n18661), .ZN(
        n18654) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18662), .B1(
        n19029), .B2(n18999), .ZN(n18653) );
  OAI211_X1 U21765 ( .C1(n19003), .C2(n18729), .A(n18654), .B(n18653), .ZN(
        P3_U2879) );
  AOI22_X1 U21766 ( .A1(n18969), .A2(n19006), .B1(n19004), .B2(n18661), .ZN(
        n18656) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18662), .B1(
        n19029), .B2(n19005), .ZN(n18655) );
  OAI211_X1 U21768 ( .C1(n19009), .C2(n18729), .A(n18656), .B(n18655), .ZN(
        P3_U2880) );
  AOI22_X1 U21769 ( .A1(n19029), .A2(n19012), .B1(n19010), .B2(n18661), .ZN(
        n18658) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18662), .B1(
        n18969), .B2(n19011), .ZN(n18657) );
  OAI211_X1 U21771 ( .C1(n19015), .C2(n18729), .A(n18658), .B(n18657), .ZN(
        P3_U2881) );
  AOI22_X1 U21772 ( .A1(n18969), .A2(n19019), .B1(n19016), .B2(n18661), .ZN(
        n18660) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18662), .B1(
        n19029), .B2(n19017), .ZN(n18659) );
  OAI211_X1 U21774 ( .C1(n19022), .C2(n18729), .A(n18660), .B(n18659), .ZN(
        P3_U2882) );
  INV_X1 U21775 ( .A(n19033), .ZN(n18968) );
  AOI22_X1 U21776 ( .A1(n19029), .A2(n18968), .B1(n19025), .B2(n18661), .ZN(
        n18664) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18662), .B1(
        n19028), .B2(n18722), .ZN(n18663) );
  OAI211_X1 U21778 ( .C1(n18966), .C2(n18974), .A(n18664), .B(n18663), .ZN(
        P3_U2883) );
  NOR2_X2 U21779 ( .A1(n18846), .A2(n18731), .ZN(n18746) );
  INV_X1 U21780 ( .A(n18746), .ZN(n18753) );
  INV_X1 U21781 ( .A(n18985), .ZN(n18850) );
  AOI21_X1 U21782 ( .B1(n18729), .B2(n18753), .A(n19103), .ZN(n18682) );
  AOI22_X1 U21783 ( .A1(n18850), .A2(n18704), .B1(n18976), .B2(n18682), .ZN(
        n18669) );
  OAI21_X1 U21784 ( .B1(n18722), .B2(n18746), .A(n18901), .ZN(n18708) );
  INV_X1 U21785 ( .A(n18708), .ZN(n18667) );
  NAND2_X1 U21786 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18753), .ZN(n18665) );
  OAI221_X1 U21787 ( .B1(n18667), .B2(n18666), .C1(n18667), .C2(n18897), .A(
        n18665), .ZN(n18683) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18683), .B1(
        n19029), .B2(n18977), .ZN(n18668) );
  OAI211_X1 U21789 ( .C1(n18853), .C2(n18753), .A(n18669), .B(n18668), .ZN(
        P3_U2884) );
  AOI22_X1 U21790 ( .A1(n19029), .A2(n18987), .B1(n18986), .B2(n18682), .ZN(
        n18671) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18683), .B1(
        n18988), .B2(n18746), .ZN(n18670) );
  OAI211_X1 U21792 ( .C1(n18686), .C2(n18991), .A(n18671), .B(n18670), .ZN(
        P3_U2885) );
  AOI22_X1 U21793 ( .A1(n19029), .A2(n18992), .B1(n18993), .B2(n18682), .ZN(
        n18673) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18683), .B1(
        n18994), .B2(n18746), .ZN(n18672) );
  OAI211_X1 U21795 ( .C1(n18686), .C2(n18997), .A(n18673), .B(n18672), .ZN(
        P3_U2886) );
  AOI22_X1 U21796 ( .A1(n18704), .A2(n18999), .B1(n18998), .B2(n18682), .ZN(
        n18675) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18683), .B1(
        n19029), .B2(n19000), .ZN(n18674) );
  OAI211_X1 U21798 ( .C1(n19003), .C2(n18753), .A(n18675), .B(n18674), .ZN(
        P3_U2887) );
  AOI22_X1 U21799 ( .A1(n19029), .A2(n19006), .B1(n19004), .B2(n18682), .ZN(
        n18677) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18683), .B1(
        n18704), .B2(n19005), .ZN(n18676) );
  OAI211_X1 U21801 ( .C1(n19009), .C2(n18753), .A(n18677), .B(n18676), .ZN(
        P3_U2888) );
  AOI22_X1 U21802 ( .A1(n19029), .A2(n19011), .B1(n19010), .B2(n18682), .ZN(
        n18679) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18683), .B1(
        n18704), .B2(n19012), .ZN(n18678) );
  OAI211_X1 U21804 ( .C1(n19015), .C2(n18753), .A(n18679), .B(n18678), .ZN(
        P3_U2889) );
  AOI22_X1 U21805 ( .A1(n19029), .A2(n19019), .B1(n19016), .B2(n18682), .ZN(
        n18681) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18683), .B1(
        n18704), .B2(n19017), .ZN(n18680) );
  OAI211_X1 U21807 ( .C1(n19022), .C2(n18753), .A(n18681), .B(n18680), .ZN(
        P3_U2890) );
  AOI22_X1 U21808 ( .A1(n19029), .A2(n19027), .B1(n19025), .B2(n18682), .ZN(
        n18685) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18683), .B1(
        n19028), .B2(n18746), .ZN(n18684) );
  OAI211_X1 U21810 ( .C1(n18686), .C2(n19033), .A(n18685), .B(n18684), .ZN(
        P3_U2891) );
  AOI22_X1 U21811 ( .A1(n18704), .A2(n18977), .B1(n18976), .B2(n18703), .ZN(
        n18690) );
  AOI21_X1 U21812 ( .B1(n19076), .B2(n18847), .A(n18687), .ZN(n18776) );
  NAND2_X1 U21813 ( .A1(n18688), .A2(n18776), .ZN(n18705) );
  NOR2_X2 U21814 ( .A1(n19075), .A2(n18731), .ZN(n18768) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18705), .B1(
        n18982), .B2(n18768), .ZN(n18689) );
  OAI211_X1 U21816 ( .C1(n18985), .C2(n18729), .A(n18690), .B(n18689), .ZN(
        P3_U2892) );
  AOI22_X1 U21817 ( .A1(n18704), .A2(n18987), .B1(n18986), .B2(n18703), .ZN(
        n18692) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18705), .B1(
        n18988), .B2(n18768), .ZN(n18691) );
  OAI211_X1 U21819 ( .C1(n18991), .C2(n18729), .A(n18692), .B(n18691), .ZN(
        P3_U2893) );
  AOI22_X1 U21820 ( .A1(n18704), .A2(n18992), .B1(n18993), .B2(n18703), .ZN(
        n18694) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18705), .B1(
        n18994), .B2(n18768), .ZN(n18693) );
  OAI211_X1 U21822 ( .C1(n18997), .C2(n18729), .A(n18694), .B(n18693), .ZN(
        P3_U2894) );
  INV_X1 U21823 ( .A(n18768), .ZN(n18775) );
  AOI22_X1 U21824 ( .A1(n18999), .A2(n18722), .B1(n18998), .B2(n18703), .ZN(
        n18696) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n19000), .ZN(n18695) );
  OAI211_X1 U21826 ( .C1(n19003), .C2(n18775), .A(n18696), .B(n18695), .ZN(
        P3_U2895) );
  AOI22_X1 U21827 ( .A1(n19005), .A2(n18722), .B1(n19004), .B2(n18703), .ZN(
        n18698) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n19006), .ZN(n18697) );
  OAI211_X1 U21829 ( .C1(n19009), .C2(n18775), .A(n18698), .B(n18697), .ZN(
        P3_U2896) );
  AOI22_X1 U21830 ( .A1(n19012), .A2(n18722), .B1(n19010), .B2(n18703), .ZN(
        n18700) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18705), .B1(
        n18704), .B2(n19011), .ZN(n18699) );
  OAI211_X1 U21832 ( .C1(n19015), .C2(n18775), .A(n18700), .B(n18699), .ZN(
        P3_U2897) );
  AOI22_X1 U21833 ( .A1(n18704), .A2(n19019), .B1(n19016), .B2(n18703), .ZN(
        n18702) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18705), .B1(
        n19017), .B2(n18722), .ZN(n18701) );
  OAI211_X1 U21835 ( .C1(n19022), .C2(n18775), .A(n18702), .B(n18701), .ZN(
        P3_U2898) );
  AOI22_X1 U21836 ( .A1(n18704), .A2(n19027), .B1(n19025), .B2(n18703), .ZN(
        n18707) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18705), .B1(
        n19028), .B2(n18768), .ZN(n18706) );
  OAI211_X1 U21838 ( .C1(n19033), .C2(n18729), .A(n18707), .B(n18706), .ZN(
        P3_U2899) );
  NOR2_X2 U21839 ( .A1(n19077), .A2(n18778), .ZN(n18791) );
  INV_X1 U21840 ( .A(n18791), .ZN(n18798) );
  NOR2_X1 U21841 ( .A1(n18768), .A2(n18791), .ZN(n18754) );
  NOR2_X1 U21842 ( .A1(n19103), .A2(n18754), .ZN(n18725) );
  AOI22_X1 U21843 ( .A1(n18977), .A2(n18722), .B1(n18976), .B2(n18725), .ZN(
        n18711) );
  OAI22_X1 U21844 ( .A1(n18754), .A2(n18947), .B1(n18847), .B2(n18708), .ZN(
        n18709) );
  OAI21_X1 U21845 ( .B1(n18791), .B2(n19206), .A(n18709), .ZN(n18726) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18726), .B1(
        n18850), .B2(n18746), .ZN(n18710) );
  OAI211_X1 U21847 ( .C1(n18853), .C2(n18798), .A(n18711), .B(n18710), .ZN(
        P3_U2900) );
  AOI22_X1 U21848 ( .A1(n18987), .A2(n18722), .B1(n18986), .B2(n18725), .ZN(
        n18713) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18726), .B1(
        n18988), .B2(n18791), .ZN(n18712) );
  OAI211_X1 U21850 ( .C1(n18991), .C2(n18753), .A(n18713), .B(n18712), .ZN(
        P3_U2901) );
  AOI22_X1 U21851 ( .A1(n18927), .A2(n18746), .B1(n18993), .B2(n18725), .ZN(
        n18715) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18726), .B1(
        n18994), .B2(n18791), .ZN(n18714) );
  OAI211_X1 U21853 ( .C1(n18931), .C2(n18729), .A(n18715), .B(n18714), .ZN(
        P3_U2902) );
  AOI22_X1 U21854 ( .A1(n18999), .A2(n18746), .B1(n18998), .B2(n18725), .ZN(
        n18717) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18726), .B1(
        n19000), .B2(n18722), .ZN(n18716) );
  OAI211_X1 U21856 ( .C1(n19003), .C2(n18798), .A(n18717), .B(n18716), .ZN(
        P3_U2903) );
  AOI22_X1 U21857 ( .A1(n19006), .A2(n18722), .B1(n19004), .B2(n18725), .ZN(
        n18719) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18726), .B1(
        n19005), .B2(n18746), .ZN(n18718) );
  OAI211_X1 U21859 ( .C1(n19009), .C2(n18798), .A(n18719), .B(n18718), .ZN(
        P3_U2904) );
  AOI22_X1 U21860 ( .A1(n19012), .A2(n18746), .B1(n19010), .B2(n18725), .ZN(
        n18721) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18726), .B1(
        n19011), .B2(n18722), .ZN(n18720) );
  OAI211_X1 U21862 ( .C1(n19015), .C2(n18798), .A(n18721), .B(n18720), .ZN(
        P3_U2905) );
  AOI22_X1 U21863 ( .A1(n19017), .A2(n18746), .B1(n19016), .B2(n18725), .ZN(
        n18724) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18726), .B1(
        n19019), .B2(n18722), .ZN(n18723) );
  OAI211_X1 U21865 ( .C1(n19022), .C2(n18798), .A(n18724), .B(n18723), .ZN(
        P3_U2906) );
  AOI22_X1 U21866 ( .A1(n18968), .A2(n18746), .B1(n19025), .B2(n18725), .ZN(
        n18728) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18726), .B1(
        n19028), .B2(n18791), .ZN(n18727) );
  OAI211_X1 U21868 ( .C1(n18974), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        P3_U2907) );
  NOR2_X2 U21869 ( .A1(n18778), .A2(n18730), .ZN(n18817) );
  INV_X1 U21870 ( .A(n18817), .ZN(n18807) );
  NOR2_X1 U21871 ( .A1(n18778), .A2(n18821), .ZN(n18749) );
  AOI22_X1 U21872 ( .A1(n18850), .A2(n18768), .B1(n18976), .B2(n18749), .ZN(
        n18735) );
  NOR2_X1 U21873 ( .A1(n19076), .A2(n18731), .ZN(n18733) );
  AOI22_X1 U21874 ( .A1(n18981), .A2(n18733), .B1(n18777), .B2(n18732), .ZN(
        n18750) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18750), .B1(
        n18977), .B2(n18746), .ZN(n18734) );
  OAI211_X1 U21876 ( .C1(n18853), .C2(n18807), .A(n18735), .B(n18734), .ZN(
        P3_U2908) );
  AOI22_X1 U21877 ( .A1(n18875), .A2(n18768), .B1(n18986), .B2(n18749), .ZN(
        n18737) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18750), .B1(
        n18988), .B2(n18817), .ZN(n18736) );
  OAI211_X1 U21879 ( .C1(n18878), .C2(n18753), .A(n18737), .B(n18736), .ZN(
        P3_U2909) );
  AOI22_X1 U21880 ( .A1(n18993), .A2(n18749), .B1(n18992), .B2(n18746), .ZN(
        n18739) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18750), .B1(
        n18994), .B2(n18817), .ZN(n18738) );
  OAI211_X1 U21882 ( .C1(n18997), .C2(n18775), .A(n18739), .B(n18738), .ZN(
        P3_U2910) );
  AOI22_X1 U21883 ( .A1(n19000), .A2(n18746), .B1(n18998), .B2(n18749), .ZN(
        n18741) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18750), .B1(
        n18999), .B2(n18768), .ZN(n18740) );
  OAI211_X1 U21885 ( .C1(n19003), .C2(n18807), .A(n18741), .B(n18740), .ZN(
        P3_U2911) );
  AOI22_X1 U21886 ( .A1(n19005), .A2(n18768), .B1(n19004), .B2(n18749), .ZN(
        n18743) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18750), .B1(
        n19006), .B2(n18746), .ZN(n18742) );
  OAI211_X1 U21888 ( .C1(n19009), .C2(n18807), .A(n18743), .B(n18742), .ZN(
        P3_U2912) );
  AOI22_X1 U21889 ( .A1(n19012), .A2(n18768), .B1(n19010), .B2(n18749), .ZN(
        n18745) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18750), .B1(
        n19011), .B2(n18746), .ZN(n18744) );
  OAI211_X1 U21891 ( .C1(n19015), .C2(n18807), .A(n18745), .B(n18744), .ZN(
        P3_U2913) );
  AOI22_X1 U21892 ( .A1(n19019), .A2(n18746), .B1(n19016), .B2(n18749), .ZN(
        n18748) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18750), .B1(
        n19017), .B2(n18768), .ZN(n18747) );
  OAI211_X1 U21894 ( .C1(n19022), .C2(n18807), .A(n18748), .B(n18747), .ZN(
        P3_U2914) );
  AOI22_X1 U21895 ( .A1(n18968), .A2(n18768), .B1(n19025), .B2(n18749), .ZN(
        n18752) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18750), .B1(
        n19028), .B2(n18817), .ZN(n18751) );
  OAI211_X1 U21897 ( .C1(n18974), .C2(n18753), .A(n18752), .B(n18751), .ZN(
        P3_U2915) );
  NOR2_X2 U21898 ( .A1(n18778), .A2(n18846), .ZN(n18842) );
  INV_X1 U21899 ( .A(n18842), .ZN(n18832) );
  AOI21_X1 U21900 ( .B1(n18807), .B2(n18832), .A(n19103), .ZN(n18771) );
  AOI22_X1 U21901 ( .A1(n18850), .A2(n18791), .B1(n18976), .B2(n18771), .ZN(
        n18757) );
  AOI221_X1 U21902 ( .B1(n18754), .B2(n18807), .C1(n18847), .C2(n18807), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18755) );
  OAI21_X1 U21903 ( .B1(n18842), .B2(n18755), .A(n18901), .ZN(n18772) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18772), .B1(
        n18977), .B2(n18768), .ZN(n18756) );
  OAI211_X1 U21905 ( .C1(n18853), .C2(n18832), .A(n18757), .B(n18756), .ZN(
        P3_U2916) );
  AOI22_X1 U21906 ( .A1(n18987), .A2(n18768), .B1(n18986), .B2(n18771), .ZN(
        n18759) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18772), .B1(
        n18988), .B2(n18842), .ZN(n18758) );
  OAI211_X1 U21908 ( .C1(n18991), .C2(n18798), .A(n18759), .B(n18758), .ZN(
        P3_U2917) );
  AOI22_X1 U21909 ( .A1(n18993), .A2(n18771), .B1(n18992), .B2(n18768), .ZN(
        n18761) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18772), .B1(
        n18994), .B2(n18842), .ZN(n18760) );
  OAI211_X1 U21911 ( .C1(n18997), .C2(n18798), .A(n18761), .B(n18760), .ZN(
        P3_U2918) );
  AOI22_X1 U21912 ( .A1(n18999), .A2(n18791), .B1(n18998), .B2(n18771), .ZN(
        n18763) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18772), .B1(
        n19000), .B2(n18768), .ZN(n18762) );
  OAI211_X1 U21914 ( .C1(n19003), .C2(n18832), .A(n18763), .B(n18762), .ZN(
        P3_U2919) );
  AOI22_X1 U21915 ( .A1(n19006), .A2(n18768), .B1(n19004), .B2(n18771), .ZN(
        n18765) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18772), .B1(
        n19005), .B2(n18791), .ZN(n18764) );
  OAI211_X1 U21917 ( .C1(n19009), .C2(n18832), .A(n18765), .B(n18764), .ZN(
        P3_U2920) );
  AOI22_X1 U21918 ( .A1(n19011), .A2(n18768), .B1(n19010), .B2(n18771), .ZN(
        n18767) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18772), .B1(
        n19012), .B2(n18791), .ZN(n18766) );
  OAI211_X1 U21920 ( .C1(n19015), .C2(n18832), .A(n18767), .B(n18766), .ZN(
        P3_U2921) );
  AOI22_X1 U21921 ( .A1(n19019), .A2(n18768), .B1(n19016), .B2(n18771), .ZN(
        n18770) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18772), .B1(
        n19017), .B2(n18791), .ZN(n18769) );
  OAI211_X1 U21923 ( .C1(n19022), .C2(n18832), .A(n18770), .B(n18769), .ZN(
        P3_U2922) );
  AOI22_X1 U21924 ( .A1(n18968), .A2(n18791), .B1(n19025), .B2(n18771), .ZN(
        n18774) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18772), .B1(
        n19028), .B2(n18842), .ZN(n18773) );
  OAI211_X1 U21926 ( .C1(n18974), .C2(n18775), .A(n18774), .B(n18773), .ZN(
        P3_U2923) );
  AOI22_X1 U21927 ( .A1(n18977), .A2(n18791), .B1(n18976), .B2(n18794), .ZN(
        n18780) );
  NAND2_X1 U21928 ( .A1(n18777), .A2(n18776), .ZN(n18795) );
  NOR2_X2 U21929 ( .A1(n19075), .A2(n18778), .ZN(n18868) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18795), .B1(
        n18982), .B2(n18868), .ZN(n18779) );
  OAI211_X1 U21931 ( .C1(n18985), .C2(n18807), .A(n18780), .B(n18779), .ZN(
        P3_U2924) );
  AOI22_X1 U21932 ( .A1(n18987), .A2(n18791), .B1(n18986), .B2(n18794), .ZN(
        n18782) );
  AOI22_X1 U21933 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18795), .B1(
        n18988), .B2(n18868), .ZN(n18781) );
  OAI211_X1 U21934 ( .C1(n18991), .C2(n18807), .A(n18782), .B(n18781), .ZN(
        P3_U2925) );
  AOI22_X1 U21935 ( .A1(n18927), .A2(n18817), .B1(n18993), .B2(n18794), .ZN(
        n18784) );
  AOI22_X1 U21936 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18795), .B1(
        n18994), .B2(n18868), .ZN(n18783) );
  OAI211_X1 U21937 ( .C1(n18931), .C2(n18798), .A(n18784), .B(n18783), .ZN(
        P3_U2926) );
  INV_X1 U21938 ( .A(n18868), .ZN(n18856) );
  AOI22_X1 U21939 ( .A1(n18999), .A2(n18817), .B1(n18998), .B2(n18794), .ZN(
        n18786) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18795), .B1(
        n19000), .B2(n18791), .ZN(n18785) );
  OAI211_X1 U21941 ( .C1(n19003), .C2(n18856), .A(n18786), .B(n18785), .ZN(
        P3_U2927) );
  AOI22_X1 U21942 ( .A1(n19006), .A2(n18791), .B1(n19004), .B2(n18794), .ZN(
        n18788) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18795), .B1(
        n19005), .B2(n18817), .ZN(n18787) );
  OAI211_X1 U21944 ( .C1(n19009), .C2(n18856), .A(n18788), .B(n18787), .ZN(
        P3_U2928) );
  AOI22_X1 U21945 ( .A1(n19011), .A2(n18791), .B1(n19010), .B2(n18794), .ZN(
        n18790) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18795), .B1(
        n19012), .B2(n18817), .ZN(n18789) );
  OAI211_X1 U21947 ( .C1(n19015), .C2(n18856), .A(n18790), .B(n18789), .ZN(
        P3_U2929) );
  AOI22_X1 U21948 ( .A1(n19017), .A2(n18817), .B1(n19016), .B2(n18794), .ZN(
        n18793) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18795), .B1(
        n19019), .B2(n18791), .ZN(n18792) );
  OAI211_X1 U21950 ( .C1(n19022), .C2(n18856), .A(n18793), .B(n18792), .ZN(
        P3_U2930) );
  AOI22_X1 U21951 ( .A1(n18968), .A2(n18817), .B1(n19025), .B2(n18794), .ZN(
        n18797) );
  AOI22_X1 U21952 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18795), .B1(
        n19028), .B2(n18868), .ZN(n18796) );
  OAI211_X1 U21953 ( .C1(n18974), .C2(n18798), .A(n18797), .B(n18796), .ZN(
        P3_U2931) );
  NOR2_X2 U21954 ( .A1(n19077), .A2(n18872), .ZN(n18887) );
  INV_X1 U21955 ( .A(n18887), .ZN(n18894) );
  NOR2_X1 U21956 ( .A1(n18817), .A2(n18842), .ZN(n18799) );
  NOR2_X1 U21957 ( .A1(n18868), .A2(n18887), .ZN(n18848) );
  OAI21_X1 U21958 ( .B1(n18799), .B2(n18847), .A(n18848), .ZN(n18800) );
  OAI211_X1 U21959 ( .C1(n18887), .C2(n19206), .A(n18901), .B(n18800), .ZN(
        n18818) );
  NOR2_X1 U21960 ( .A1(n19103), .A2(n18848), .ZN(n18816) );
  AOI22_X1 U21961 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18818), .B1(
        n18976), .B2(n18816), .ZN(n18802) );
  AOI22_X1 U21962 ( .A1(n18850), .A2(n18842), .B1(n18977), .B2(n18817), .ZN(
        n18801) );
  OAI211_X1 U21963 ( .C1(n18853), .C2(n18894), .A(n18802), .B(n18801), .ZN(
        P3_U2932) );
  AOI22_X1 U21964 ( .A1(n18875), .A2(n18842), .B1(n18986), .B2(n18816), .ZN(
        n18804) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18818), .B1(
        n18988), .B2(n18887), .ZN(n18803) );
  OAI211_X1 U21966 ( .C1(n18878), .C2(n18807), .A(n18804), .B(n18803), .ZN(
        P3_U2933) );
  AOI22_X1 U21967 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18818), .B1(
        n18993), .B2(n18816), .ZN(n18806) );
  AOI22_X1 U21968 ( .A1(n18927), .A2(n18842), .B1(n18994), .B2(n18887), .ZN(
        n18805) );
  OAI211_X1 U21969 ( .C1(n18931), .C2(n18807), .A(n18806), .B(n18805), .ZN(
        P3_U2934) );
  AOI22_X1 U21970 ( .A1(n18999), .A2(n18842), .B1(n18998), .B2(n18816), .ZN(
        n18809) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18818), .B1(
        n19000), .B2(n18817), .ZN(n18808) );
  OAI211_X1 U21972 ( .C1(n19003), .C2(n18894), .A(n18809), .B(n18808), .ZN(
        P3_U2935) );
  AOI22_X1 U21973 ( .A1(n19005), .A2(n18842), .B1(n19004), .B2(n18816), .ZN(
        n18811) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18818), .B1(
        n19006), .B2(n18817), .ZN(n18810) );
  OAI211_X1 U21975 ( .C1(n19009), .C2(n18894), .A(n18811), .B(n18810), .ZN(
        P3_U2936) );
  AOI22_X1 U21976 ( .A1(n19011), .A2(n18817), .B1(n19010), .B2(n18816), .ZN(
        n18813) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18818), .B1(
        n19012), .B2(n18842), .ZN(n18812) );
  OAI211_X1 U21978 ( .C1(n19015), .C2(n18894), .A(n18813), .B(n18812), .ZN(
        P3_U2937) );
  AOI22_X1 U21979 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18818), .B1(
        n19016), .B2(n18816), .ZN(n18815) );
  AOI22_X1 U21980 ( .A1(n19019), .A2(n18817), .B1(n19017), .B2(n18842), .ZN(
        n18814) );
  OAI211_X1 U21981 ( .C1(n19022), .C2(n18894), .A(n18815), .B(n18814), .ZN(
        P3_U2938) );
  AOI22_X1 U21982 ( .A1(n19027), .A2(n18817), .B1(n19025), .B2(n18816), .ZN(
        n18820) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18818), .B1(
        n19028), .B2(n18887), .ZN(n18819) );
  OAI211_X1 U21984 ( .C1(n19033), .C2(n18832), .A(n18820), .B(n18819), .ZN(
        P3_U2939) );
  NOR2_X1 U21985 ( .A1(n18872), .A2(n18821), .ZN(n18841) );
  AOI22_X1 U21986 ( .A1(n18977), .A2(n18842), .B1(n18976), .B2(n18841), .ZN(
        n18827) );
  NOR2_X1 U21987 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18822), .ZN(
        n18824) );
  NOR2_X1 U21988 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18872), .ZN(
        n18823) );
  AOI22_X1 U21989 ( .A1(n18981), .A2(n18824), .B1(n18979), .B2(n18823), .ZN(
        n18843) );
  NAND2_X1 U21990 ( .A1(n18896), .A2(n18825), .ZN(n18908) );
  INV_X1 U21991 ( .A(n18908), .ZN(n18918) );
  AOI22_X1 U21992 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18843), .B1(
        n18982), .B2(n18918), .ZN(n18826) );
  OAI211_X1 U21993 ( .C1(n18985), .C2(n18856), .A(n18827), .B(n18826), .ZN(
        P3_U2940) );
  AOI22_X1 U21994 ( .A1(n18875), .A2(n18868), .B1(n18986), .B2(n18841), .ZN(
        n18829) );
  AOI22_X1 U21995 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18843), .B1(
        n18988), .B2(n18918), .ZN(n18828) );
  OAI211_X1 U21996 ( .C1(n18878), .C2(n18832), .A(n18829), .B(n18828), .ZN(
        P3_U2941) );
  AOI22_X1 U21997 ( .A1(n18927), .A2(n18868), .B1(n18993), .B2(n18841), .ZN(
        n18831) );
  AOI22_X1 U21998 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18843), .B1(
        n18994), .B2(n18918), .ZN(n18830) );
  OAI211_X1 U21999 ( .C1(n18931), .C2(n18832), .A(n18831), .B(n18830), .ZN(
        P3_U2942) );
  AOI22_X1 U22000 ( .A1(n18999), .A2(n18868), .B1(n18998), .B2(n18841), .ZN(
        n18834) );
  AOI22_X1 U22001 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18843), .B1(
        n19000), .B2(n18842), .ZN(n18833) );
  OAI211_X1 U22002 ( .C1(n19003), .C2(n18908), .A(n18834), .B(n18833), .ZN(
        P3_U2943) );
  AOI22_X1 U22003 ( .A1(n19005), .A2(n18868), .B1(n19004), .B2(n18841), .ZN(
        n18836) );
  AOI22_X1 U22004 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18843), .B1(
        n19006), .B2(n18842), .ZN(n18835) );
  OAI211_X1 U22005 ( .C1(n19009), .C2(n18908), .A(n18836), .B(n18835), .ZN(
        P3_U2944) );
  AOI22_X1 U22006 ( .A1(n19012), .A2(n18868), .B1(n19010), .B2(n18841), .ZN(
        n18838) );
  AOI22_X1 U22007 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18843), .B1(
        n19011), .B2(n18842), .ZN(n18837) );
  OAI211_X1 U22008 ( .C1(n19015), .C2(n18908), .A(n18838), .B(n18837), .ZN(
        P3_U2945) );
  AOI22_X1 U22009 ( .A1(n19019), .A2(n18842), .B1(n19016), .B2(n18841), .ZN(
        n18840) );
  AOI22_X1 U22010 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18843), .B1(
        n19017), .B2(n18868), .ZN(n18839) );
  OAI211_X1 U22011 ( .C1(n19022), .C2(n18908), .A(n18840), .B(n18839), .ZN(
        P3_U2946) );
  AOI22_X1 U22012 ( .A1(n19027), .A2(n18842), .B1(n19025), .B2(n18841), .ZN(
        n18845) );
  AOI22_X1 U22013 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18843), .B1(
        n19028), .B2(n18918), .ZN(n18844) );
  OAI211_X1 U22014 ( .C1(n19033), .C2(n18856), .A(n18845), .B(n18844), .ZN(
        P3_U2947) );
  NOR2_X2 U22015 ( .A1(n18872), .A2(n18846), .ZN(n18941) );
  INV_X1 U22016 ( .A(n18941), .ZN(n18930) );
  AOI21_X1 U22017 ( .B1(n18908), .B2(n18930), .A(n19103), .ZN(n18867) );
  AOI22_X1 U22018 ( .A1(n18977), .A2(n18868), .B1(n18976), .B2(n18867), .ZN(
        n18852) );
  OAI211_X1 U22019 ( .C1(n18848), .C2(n18847), .A(n18908), .B(n18930), .ZN(
        n18849) );
  OAI211_X1 U22020 ( .C1(n18941), .C2(n19206), .A(n18901), .B(n18849), .ZN(
        n18869) );
  AOI22_X1 U22021 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18869), .B1(
        n18850), .B2(n18887), .ZN(n18851) );
  OAI211_X1 U22022 ( .C1(n18853), .C2(n18930), .A(n18852), .B(n18851), .ZN(
        P3_U2948) );
  AOI22_X1 U22023 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18869), .B1(
        n18986), .B2(n18867), .ZN(n18855) );
  AOI22_X1 U22024 ( .A1(n18875), .A2(n18887), .B1(n18988), .B2(n18941), .ZN(
        n18854) );
  OAI211_X1 U22025 ( .C1(n18878), .C2(n18856), .A(n18855), .B(n18854), .ZN(
        P3_U2949) );
  AOI22_X1 U22026 ( .A1(n18993), .A2(n18867), .B1(n18992), .B2(n18868), .ZN(
        n18858) );
  AOI22_X1 U22027 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18869), .B1(
        n18994), .B2(n18941), .ZN(n18857) );
  OAI211_X1 U22028 ( .C1(n18997), .C2(n18894), .A(n18858), .B(n18857), .ZN(
        P3_U2950) );
  AOI22_X1 U22029 ( .A1(n18999), .A2(n18887), .B1(n18998), .B2(n18867), .ZN(
        n18860) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18869), .B1(
        n19000), .B2(n18868), .ZN(n18859) );
  OAI211_X1 U22031 ( .C1(n19003), .C2(n18930), .A(n18860), .B(n18859), .ZN(
        P3_U2951) );
  AOI22_X1 U22032 ( .A1(n19005), .A2(n18887), .B1(n19004), .B2(n18867), .ZN(
        n18862) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18869), .B1(
        n19006), .B2(n18868), .ZN(n18861) );
  OAI211_X1 U22034 ( .C1(n19009), .C2(n18930), .A(n18862), .B(n18861), .ZN(
        P3_U2952) );
  AOI22_X1 U22035 ( .A1(n19012), .A2(n18887), .B1(n19010), .B2(n18867), .ZN(
        n18864) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18869), .B1(
        n19011), .B2(n18868), .ZN(n18863) );
  OAI211_X1 U22037 ( .C1(n19015), .C2(n18930), .A(n18864), .B(n18863), .ZN(
        P3_U2953) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18869), .B1(
        n19016), .B2(n18867), .ZN(n18866) );
  AOI22_X1 U22039 ( .A1(n19019), .A2(n18868), .B1(n19017), .B2(n18887), .ZN(
        n18865) );
  OAI211_X1 U22040 ( .C1(n19022), .C2(n18930), .A(n18866), .B(n18865), .ZN(
        P3_U2954) );
  AOI22_X1 U22041 ( .A1(n19027), .A2(n18868), .B1(n19025), .B2(n18867), .ZN(
        n18871) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18869), .B1(
        n19028), .B2(n18941), .ZN(n18870) );
  OAI211_X1 U22043 ( .C1(n19033), .C2(n18894), .A(n18871), .B(n18870), .ZN(
        P3_U2955) );
  NOR2_X1 U22044 ( .A1(n19076), .A2(n18872), .ZN(n18922) );
  AND2_X1 U22045 ( .A1(n18975), .A2(n18922), .ZN(n18890) );
  AOI22_X1 U22046 ( .A1(n18977), .A2(n18887), .B1(n18976), .B2(n18890), .ZN(
        n18874) );
  OAI211_X1 U22047 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18981), .A(
        n18979), .B(n18896), .ZN(n18891) );
  NOR2_X2 U22048 ( .A1(n19075), .A2(n18872), .ZN(n18963) );
  AOI22_X1 U22049 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18891), .B1(
        n18982), .B2(n18963), .ZN(n18873) );
  OAI211_X1 U22050 ( .C1(n18985), .C2(n18908), .A(n18874), .B(n18873), .ZN(
        P3_U2956) );
  AOI22_X1 U22051 ( .A1(n18875), .A2(n18918), .B1(n18986), .B2(n18890), .ZN(
        n18877) );
  AOI22_X1 U22052 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18891), .B1(
        n18988), .B2(n18963), .ZN(n18876) );
  OAI211_X1 U22053 ( .C1(n18878), .C2(n18894), .A(n18877), .B(n18876), .ZN(
        P3_U2957) );
  AOI22_X1 U22054 ( .A1(n18993), .A2(n18890), .B1(n18992), .B2(n18887), .ZN(
        n18880) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18891), .B1(
        n18994), .B2(n18963), .ZN(n18879) );
  OAI211_X1 U22056 ( .C1(n18997), .C2(n18908), .A(n18880), .B(n18879), .ZN(
        P3_U2958) );
  INV_X1 U22057 ( .A(n18963), .ZN(n18973) );
  AOI22_X1 U22058 ( .A1(n19000), .A2(n18887), .B1(n18998), .B2(n18890), .ZN(
        n18882) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18891), .B1(
        n18999), .B2(n18918), .ZN(n18881) );
  OAI211_X1 U22060 ( .C1(n19003), .C2(n18973), .A(n18882), .B(n18881), .ZN(
        P3_U2959) );
  AOI22_X1 U22061 ( .A1(n19005), .A2(n18918), .B1(n19004), .B2(n18890), .ZN(
        n18884) );
  AOI22_X1 U22062 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18891), .B1(
        n19006), .B2(n18887), .ZN(n18883) );
  OAI211_X1 U22063 ( .C1(n19009), .C2(n18973), .A(n18884), .B(n18883), .ZN(
        P3_U2960) );
  AOI22_X1 U22064 ( .A1(n19011), .A2(n18887), .B1(n19010), .B2(n18890), .ZN(
        n18886) );
  AOI22_X1 U22065 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18891), .B1(
        n19012), .B2(n18918), .ZN(n18885) );
  OAI211_X1 U22066 ( .C1(n19015), .C2(n18973), .A(n18886), .B(n18885), .ZN(
        P3_U2961) );
  AOI22_X1 U22067 ( .A1(n19017), .A2(n18918), .B1(n19016), .B2(n18890), .ZN(
        n18889) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18891), .B1(
        n19019), .B2(n18887), .ZN(n18888) );
  OAI211_X1 U22069 ( .C1(n19022), .C2(n18973), .A(n18889), .B(n18888), .ZN(
        P3_U2962) );
  AOI22_X1 U22070 ( .A1(n18968), .A2(n18918), .B1(n19025), .B2(n18890), .ZN(
        n18893) );
  AOI22_X1 U22071 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18891), .B1(
        n19028), .B2(n18963), .ZN(n18892) );
  OAI211_X1 U22072 ( .C1(n18974), .C2(n18894), .A(n18893), .B(n18892), .ZN(
        P3_U2963) );
  NAND2_X1 U22073 ( .A1(n18895), .A2(n18980), .ZN(n18956) );
  INV_X1 U22074 ( .A(n18956), .ZN(n19026) );
  NAND2_X1 U22075 ( .A1(n18897), .A2(n18896), .ZN(n18898) );
  NOR2_X1 U22076 ( .A1(n18963), .A2(n19026), .ZN(n18948) );
  OAI21_X1 U22077 ( .B1(n18899), .B2(n18898), .A(n18948), .ZN(n18900) );
  OAI211_X1 U22078 ( .C1(n19026), .C2(n19206), .A(n18901), .B(n18900), .ZN(
        n18919) );
  NOR2_X1 U22079 ( .A1(n19103), .A2(n18948), .ZN(n18917) );
  AOI22_X1 U22080 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18919), .B1(
        n18976), .B2(n18917), .ZN(n18903) );
  AOI22_X1 U22081 ( .A1(n18982), .A2(n19026), .B1(n18977), .B2(n18918), .ZN(
        n18902) );
  OAI211_X1 U22082 ( .C1(n18985), .C2(n18930), .A(n18903), .B(n18902), .ZN(
        P3_U2964) );
  AOI22_X1 U22083 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18919), .B1(
        n18986), .B2(n18917), .ZN(n18905) );
  AOI22_X1 U22084 ( .A1(n18988), .A2(n19026), .B1(n18987), .B2(n18918), .ZN(
        n18904) );
  OAI211_X1 U22085 ( .C1(n18991), .C2(n18930), .A(n18905), .B(n18904), .ZN(
        P3_U2965) );
  AOI22_X1 U22086 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18919), .B1(
        n18993), .B2(n18917), .ZN(n18907) );
  AOI22_X1 U22087 ( .A1(n18927), .A2(n18941), .B1(n18994), .B2(n19026), .ZN(
        n18906) );
  OAI211_X1 U22088 ( .C1(n18931), .C2(n18908), .A(n18907), .B(n18906), .ZN(
        P3_U2966) );
  AOI22_X1 U22089 ( .A1(n19000), .A2(n18918), .B1(n18998), .B2(n18917), .ZN(
        n18910) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18919), .B1(
        n18999), .B2(n18941), .ZN(n18909) );
  OAI211_X1 U22091 ( .C1(n19003), .C2(n18956), .A(n18910), .B(n18909), .ZN(
        P3_U2967) );
  AOI22_X1 U22092 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18919), .B1(
        n19004), .B2(n18917), .ZN(n18912) );
  AOI22_X1 U22093 ( .A1(n19006), .A2(n18918), .B1(n19005), .B2(n18941), .ZN(
        n18911) );
  OAI211_X1 U22094 ( .C1(n19009), .C2(n18956), .A(n18912), .B(n18911), .ZN(
        P3_U2968) );
  AOI22_X1 U22095 ( .A1(n19011), .A2(n18918), .B1(n19010), .B2(n18917), .ZN(
        n18914) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18919), .B1(
        n19012), .B2(n18941), .ZN(n18913) );
  OAI211_X1 U22097 ( .C1(n19015), .C2(n18956), .A(n18914), .B(n18913), .ZN(
        P3_U2969) );
  AOI22_X1 U22098 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18919), .B1(
        n19016), .B2(n18917), .ZN(n18916) );
  AOI22_X1 U22099 ( .A1(n19019), .A2(n18918), .B1(n19017), .B2(n18941), .ZN(
        n18915) );
  OAI211_X1 U22100 ( .C1(n19022), .C2(n18956), .A(n18916), .B(n18915), .ZN(
        P3_U2970) );
  AOI22_X1 U22101 ( .A1(n19027), .A2(n18918), .B1(n19025), .B2(n18917), .ZN(
        n18921) );
  AOI22_X1 U22102 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18919), .B1(
        n19028), .B2(n19026), .ZN(n18920) );
  OAI211_X1 U22103 ( .C1(n19033), .C2(n18930), .A(n18921), .B(n18920), .ZN(
        P3_U2971) );
  AND2_X1 U22104 ( .A1(n18975), .A2(n18980), .ZN(n18940) );
  AOI22_X1 U22105 ( .A1(n18977), .A2(n18941), .B1(n18976), .B2(n18940), .ZN(
        n18924) );
  AOI22_X1 U22106 ( .A1(n18981), .A2(n18922), .B1(n18980), .B2(n18979), .ZN(
        n18942) );
  AOI22_X1 U22107 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18942), .B1(
        n18982), .B2(n19018), .ZN(n18923) );
  OAI211_X1 U22108 ( .C1(n18985), .C2(n18973), .A(n18924), .B(n18923), .ZN(
        P3_U2972) );
  AOI22_X1 U22109 ( .A1(n18987), .A2(n18941), .B1(n18986), .B2(n18940), .ZN(
        n18926) );
  AOI22_X1 U22110 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18942), .B1(
        n19018), .B2(n18988), .ZN(n18925) );
  OAI211_X1 U22111 ( .C1(n18991), .C2(n18973), .A(n18926), .B(n18925), .ZN(
        P3_U2973) );
  AOI22_X1 U22112 ( .A1(n18927), .A2(n18963), .B1(n18993), .B2(n18940), .ZN(
        n18929) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18942), .B1(
        n19018), .B2(n18994), .ZN(n18928) );
  OAI211_X1 U22114 ( .C1(n18931), .C2(n18930), .A(n18929), .B(n18928), .ZN(
        P3_U2974) );
  AOI22_X1 U22115 ( .A1(n18999), .A2(n18963), .B1(n18998), .B2(n18940), .ZN(
        n18933) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18942), .B1(
        n19000), .B2(n18941), .ZN(n18932) );
  OAI211_X1 U22117 ( .C1(n19034), .C2(n19003), .A(n18933), .B(n18932), .ZN(
        P3_U2975) );
  AOI22_X1 U22118 ( .A1(n19006), .A2(n18941), .B1(n19004), .B2(n18940), .ZN(
        n18935) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18942), .B1(
        n19005), .B2(n18963), .ZN(n18934) );
  OAI211_X1 U22120 ( .C1(n19034), .C2(n19009), .A(n18935), .B(n18934), .ZN(
        P3_U2976) );
  AOI22_X1 U22121 ( .A1(n19011), .A2(n18941), .B1(n19010), .B2(n18940), .ZN(
        n18937) );
  AOI22_X1 U22122 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18942), .B1(
        n19012), .B2(n18963), .ZN(n18936) );
  OAI211_X1 U22123 ( .C1(n19034), .C2(n19015), .A(n18937), .B(n18936), .ZN(
        P3_U2977) );
  AOI22_X1 U22124 ( .A1(n19019), .A2(n18941), .B1(n19016), .B2(n18940), .ZN(
        n18939) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18942), .B1(
        n19017), .B2(n18963), .ZN(n18938) );
  OAI211_X1 U22126 ( .C1(n19034), .C2(n19022), .A(n18939), .B(n18938), .ZN(
        P3_U2978) );
  AOI22_X1 U22127 ( .A1(n19027), .A2(n18941), .B1(n19025), .B2(n18940), .ZN(
        n18944) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18942), .B1(
        n19018), .B2(n19028), .ZN(n18943) );
  OAI211_X1 U22129 ( .C1(n19033), .C2(n18973), .A(n18944), .B(n18943), .ZN(
        P3_U2979) );
  INV_X1 U22130 ( .A(n18945), .ZN(n18946) );
  NOR2_X1 U22131 ( .A1(n19103), .A2(n18946), .ZN(n18967) );
  AOI22_X1 U22132 ( .A1(n18977), .A2(n18963), .B1(n18976), .B2(n18967), .ZN(
        n18951) );
  OAI22_X1 U22133 ( .A1(n18948), .A2(n18636), .B1(n18947), .B2(n18946), .ZN(
        n18949) );
  OAI21_X1 U22134 ( .B1(n18969), .B2(n19206), .A(n18949), .ZN(n18970) );
  AOI22_X1 U22135 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18970), .B1(
        n18969), .B2(n18982), .ZN(n18950) );
  OAI211_X1 U22136 ( .C1(n18985), .C2(n18956), .A(n18951), .B(n18950), .ZN(
        P3_U2980) );
  AOI22_X1 U22137 ( .A1(n18987), .A2(n18963), .B1(n18986), .B2(n18967), .ZN(
        n18953) );
  AOI22_X1 U22138 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18970), .B1(
        n18969), .B2(n18988), .ZN(n18952) );
  OAI211_X1 U22139 ( .C1(n18991), .C2(n18956), .A(n18953), .B(n18952), .ZN(
        P3_U2981) );
  AOI22_X1 U22140 ( .A1(n18993), .A2(n18967), .B1(n18992), .B2(n18963), .ZN(
        n18955) );
  AOI22_X1 U22141 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18970), .B1(
        n18969), .B2(n18994), .ZN(n18954) );
  OAI211_X1 U22142 ( .C1(n18997), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        P3_U2982) );
  AOI22_X1 U22143 ( .A1(n19000), .A2(n18963), .B1(n18998), .B2(n18967), .ZN(
        n18958) );
  AOI22_X1 U22144 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18970), .B1(
        n18999), .B2(n19026), .ZN(n18957) );
  OAI211_X1 U22145 ( .C1(n18966), .C2(n19003), .A(n18958), .B(n18957), .ZN(
        P3_U2983) );
  AOI22_X1 U22146 ( .A1(n19006), .A2(n18963), .B1(n19004), .B2(n18967), .ZN(
        n18960) );
  AOI22_X1 U22147 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18970), .B1(
        n19005), .B2(n19026), .ZN(n18959) );
  OAI211_X1 U22148 ( .C1(n18966), .C2(n19009), .A(n18960), .B(n18959), .ZN(
        P3_U2984) );
  AOI22_X1 U22149 ( .A1(n19011), .A2(n18963), .B1(n19010), .B2(n18967), .ZN(
        n18962) );
  AOI22_X1 U22150 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18970), .B1(
        n19012), .B2(n19026), .ZN(n18961) );
  OAI211_X1 U22151 ( .C1(n18966), .C2(n19015), .A(n18962), .B(n18961), .ZN(
        P3_U2985) );
  AOI22_X1 U22152 ( .A1(n19017), .A2(n19026), .B1(n19016), .B2(n18967), .ZN(
        n18965) );
  AOI22_X1 U22153 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18970), .B1(
        n19019), .B2(n18963), .ZN(n18964) );
  OAI211_X1 U22154 ( .C1(n18966), .C2(n19022), .A(n18965), .B(n18964), .ZN(
        P3_U2986) );
  AOI22_X1 U22155 ( .A1(n18968), .A2(n19026), .B1(n19025), .B2(n18967), .ZN(
        n18972) );
  AOI22_X1 U22156 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18970), .B1(
        n18969), .B2(n19028), .ZN(n18971) );
  OAI211_X1 U22157 ( .C1(n18974), .C2(n18973), .A(n18972), .B(n18971), .ZN(
        P3_U2987) );
  AND2_X1 U22158 ( .A1(n18975), .A2(n18978), .ZN(n19024) );
  AOI22_X1 U22159 ( .A1(n18977), .A2(n19026), .B1(n18976), .B2(n19024), .ZN(
        n18984) );
  AOI22_X1 U22160 ( .A1(n18981), .A2(n18980), .B1(n18979), .B2(n18978), .ZN(
        n19030) );
  AOI22_X1 U22161 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18982), .ZN(n18983) );
  OAI211_X1 U22162 ( .C1(n18985), .C2(n19034), .A(n18984), .B(n18983), .ZN(
        P3_U2988) );
  AOI22_X1 U22163 ( .A1(n18987), .A2(n19026), .B1(n18986), .B2(n19024), .ZN(
        n18990) );
  AOI22_X1 U22164 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18988), .ZN(n18989) );
  OAI211_X1 U22165 ( .C1(n19034), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P3_U2989) );
  AOI22_X1 U22166 ( .A1(n18993), .A2(n19024), .B1(n18992), .B2(n19026), .ZN(
        n18996) );
  AOI22_X1 U22167 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n18994), .ZN(n18995) );
  OAI211_X1 U22168 ( .C1(n19034), .C2(n18997), .A(n18996), .B(n18995), .ZN(
        P3_U2990) );
  AOI22_X1 U22169 ( .A1(n19018), .A2(n18999), .B1(n18998), .B2(n19024), .ZN(
        n19002) );
  AOI22_X1 U22170 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19030), .B1(
        n19000), .B2(n19026), .ZN(n19001) );
  OAI211_X1 U22171 ( .C1(n19023), .C2(n19003), .A(n19002), .B(n19001), .ZN(
        P3_U2991) );
  AOI22_X1 U22172 ( .A1(n19018), .A2(n19005), .B1(n19004), .B2(n19024), .ZN(
        n19008) );
  AOI22_X1 U22173 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19030), .B1(
        n19006), .B2(n19026), .ZN(n19007) );
  OAI211_X1 U22174 ( .C1(n19023), .C2(n19009), .A(n19008), .B(n19007), .ZN(
        P3_U2992) );
  AOI22_X1 U22175 ( .A1(n19011), .A2(n19026), .B1(n19010), .B2(n19024), .ZN(
        n19014) );
  AOI22_X1 U22176 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19030), .B1(
        n19018), .B2(n19012), .ZN(n19013) );
  OAI211_X1 U22177 ( .C1(n19023), .C2(n19015), .A(n19014), .B(n19013), .ZN(
        P3_U2993) );
  AOI22_X1 U22178 ( .A1(n19018), .A2(n19017), .B1(n19016), .B2(n19024), .ZN(
        n19021) );
  AOI22_X1 U22179 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19030), .B1(
        n19019), .B2(n19026), .ZN(n19020) );
  OAI211_X1 U22180 ( .C1(n19023), .C2(n19022), .A(n19021), .B(n19020), .ZN(
        P3_U2994) );
  AOI22_X1 U22181 ( .A1(n19027), .A2(n19026), .B1(n19025), .B2(n19024), .ZN(
        n19032) );
  AOI22_X1 U22182 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19030), .B1(
        n19029), .B2(n19028), .ZN(n19031) );
  OAI211_X1 U22183 ( .C1(n19034), .C2(n19033), .A(n19032), .B(n19031), .ZN(
        P3_U2995) );
  NOR2_X1 U22184 ( .A1(n19051), .A2(n19035), .ZN(n19037) );
  OAI222_X1 U22185 ( .A1(n19041), .A2(n19040), .B1(n19039), .B2(n19038), .C1(
        n19037), .C2(n19036), .ZN(n19248) );
  OAI21_X1 U22186 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19042), .ZN(n19044) );
  OAI211_X1 U22187 ( .C1(n19069), .C2(n19045), .A(n19044), .B(n19043), .ZN(
        n19090) );
  INV_X1 U22188 ( .A(n19069), .ZN(n19079) );
  NAND2_X1 U22189 ( .A1(n9868), .A2(n19065), .ZN(n19050) );
  OAI21_X1 U22190 ( .B1(n19235), .B2(n19047), .A(n19046), .ZN(n19061) );
  NOR2_X1 U22191 ( .A1(n19061), .A2(n19048), .ZN(n19073) );
  INV_X1 U22192 ( .A(n19073), .ZN(n19049) );
  AOI22_X1 U22193 ( .A1(n19051), .A2(n19050), .B1(n19056), .B2(n19049), .ZN(
        n19207) );
  NOR2_X1 U22194 ( .A1(n19079), .A2(n19207), .ZN(n19059) );
  AOI21_X1 U22195 ( .B1(n19054), .B2(n19053), .A(n19052), .ZN(n19063) );
  OAI22_X1 U22196 ( .A1(n19072), .A2(n19056), .B1(n19055), .B2(n19063), .ZN(
        n19057) );
  AOI21_X1 U22197 ( .B1(n9868), .B2(n19065), .A(n19057), .ZN(n19211) );
  NAND2_X1 U22198 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19211), .ZN(
        n19058) );
  OAI22_X1 U22199 ( .A1(n19059), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19079), .B2(n19058), .ZN(n19088) );
  NAND2_X1 U22200 ( .A1(n19229), .A2(n9868), .ZN(n19060) );
  OAI221_X1 U22201 ( .B1(n19229), .B2(n9868), .C1(n19062), .C2(n19061), .A(
        n19060), .ZN(n19067) );
  INV_X1 U22202 ( .A(n19063), .ZN(n19064) );
  NAND3_X1 U22203 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19065), .A3(
        n19064), .ZN(n19066) );
  OAI211_X1 U22204 ( .C1(n19219), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        n19220) );
  MUX2_X1 U22205 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19220), .S(
        n19069), .Z(n19083) );
  NOR2_X1 U22206 ( .A1(n19071), .A2(n19070), .ZN(n19074) );
  AOI22_X1 U22207 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19072), .B1(
        n19074), .B2(n19235), .ZN(n19231) );
  OAI22_X1 U22208 ( .A1(n19074), .A2(n19222), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19073), .ZN(n19227) );
  AOI222_X1 U22209 ( .A1(n19231), .A2(n19227), .B1(n19231), .B2(n19076), .C1(
        n19227), .C2(n19075), .ZN(n19078) );
  OAI21_X1 U22210 ( .B1(n19079), .B2(n19078), .A(n19077), .ZN(n19082) );
  AND2_X1 U22211 ( .A1(n19083), .A2(n19082), .ZN(n19080) );
  OAI221_X1 U22212 ( .B1(n19083), .B2(n19082), .C1(n19081), .C2(n19080), .A(
        n19085), .ZN(n19087) );
  AOI21_X1 U22213 ( .B1(n19085), .B2(n19084), .A(n19083), .ZN(n19086) );
  AOI222_X1 U22214 ( .A1(n19088), .A2(n19087), .B1(n19088), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19087), .C2(n19086), .ZN(
        n19089) );
  NOR4_X1 U22215 ( .A1(n19091), .A2(n19248), .A3(n19090), .A4(n19089), .ZN(
        n19101) );
  AOI22_X1 U22216 ( .A1(n19230), .A2(n19260), .B1(n19122), .B2(n19253), .ZN(
        n19092) );
  INV_X1 U22217 ( .A(n19092), .ZN(n19097) );
  OAI211_X1 U22218 ( .C1(n19094), .C2(n19093), .A(n19251), .B(n19101), .ZN(
        n19205) );
  OAI21_X1 U22219 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19257), .A(n19205), 
        .ZN(n19104) );
  NOR2_X1 U22220 ( .A1(n19095), .A2(n19104), .ZN(n19096) );
  OAI211_X1 U22221 ( .C1(n19101), .C2(n19100), .A(n19099), .B(n19098), .ZN(
        P3_U2996) );
  NAND2_X1 U22222 ( .A1(n19122), .A2(n19253), .ZN(n19108) );
  NOR4_X1 U22223 ( .A1(n19102), .A2(n19216), .A3(n19257), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19111) );
  INV_X1 U22224 ( .A(n19111), .ZN(n19107) );
  OR3_X1 U22225 ( .A1(n19105), .A2(n19104), .A3(n19103), .ZN(n19106) );
  NAND4_X1 U22226 ( .A1(n19109), .A2(n19108), .A3(n19107), .A4(n19106), .ZN(
        P3_U2997) );
  OAI21_X1 U22227 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19110), .ZN(n19112) );
  AOI21_X1 U22228 ( .B1(n19113), .B2(n19112), .A(n19111), .ZN(P3_U2998) );
  INV_X1 U22229 ( .A(n19203), .ZN(n19114) );
  AND2_X1 U22230 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19114), .ZN(
        P3_U2999) );
  AND2_X1 U22231 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19114), .ZN(
        P3_U3000) );
  AND2_X1 U22232 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19114), .ZN(
        P3_U3001) );
  AND2_X1 U22233 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19114), .ZN(
        P3_U3002) );
  AND2_X1 U22234 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19114), .ZN(
        P3_U3003) );
  AND2_X1 U22235 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19114), .ZN(
        P3_U3004) );
  AND2_X1 U22236 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19114), .ZN(
        P3_U3005) );
  AND2_X1 U22237 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19114), .ZN(
        P3_U3006) );
  AND2_X1 U22238 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19114), .ZN(
        P3_U3007) );
  AND2_X1 U22239 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19114), .ZN(
        P3_U3008) );
  AND2_X1 U22240 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19114), .ZN(
        P3_U3009) );
  AND2_X1 U22241 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19114), .ZN(
        P3_U3010) );
  AND2_X1 U22242 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19114), .ZN(
        P3_U3011) );
  AND2_X1 U22243 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19114), .ZN(
        P3_U3012) );
  AND2_X1 U22244 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19114), .ZN(
        P3_U3013) );
  AND2_X1 U22245 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19114), .ZN(
        P3_U3014) );
  AND2_X1 U22246 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19114), .ZN(
        P3_U3015) );
  AND2_X1 U22247 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19114), .ZN(
        P3_U3016) );
  AND2_X1 U22248 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19114), .ZN(
        P3_U3017) );
  AND2_X1 U22249 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19114), .ZN(
        P3_U3018) );
  AND2_X1 U22250 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19114), .ZN(
        P3_U3019) );
  AND2_X1 U22251 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19114), .ZN(
        P3_U3020) );
  AND2_X1 U22252 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19114), .ZN(P3_U3021) );
  AND2_X1 U22253 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19114), .ZN(P3_U3022) );
  AND2_X1 U22254 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19114), .ZN(P3_U3023) );
  AND2_X1 U22255 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19114), .ZN(P3_U3024) );
  AND2_X1 U22256 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19114), .ZN(P3_U3025) );
  AND2_X1 U22257 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19114), .ZN(P3_U3026) );
  AND2_X1 U22258 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19114), .ZN(P3_U3027) );
  AND2_X1 U22259 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19114), .ZN(P3_U3028) );
  INV_X1 U22260 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19119) );
  NOR2_X1 U22261 ( .A1(n19132), .A2(n20966), .ZN(n19128) );
  INV_X1 U22262 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19115) );
  NOR2_X1 U22263 ( .A1(n19128), .A2(n19115), .ZN(n19121) );
  OAI21_X1 U22264 ( .B1(n19119), .B2(n20966), .A(n19121), .ZN(n19116) );
  AOI22_X1 U22265 ( .A1(n19130), .A2(n19132), .B1(n19266), .B2(n19116), .ZN(
        n19117) );
  NAND3_X1 U22266 ( .A1(NA), .A2(n19130), .A3(n19119), .ZN(n19125) );
  OAI211_X1 U22267 ( .C1(n19257), .C2(n19118), .A(n19117), .B(n19125), .ZN(
        P3_U3029) );
  NOR2_X1 U22268 ( .A1(n19119), .A2(n20966), .ZN(n19120) );
  AOI22_X1 U22269 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19121), .B1(n19120), 
        .B2(n19132), .ZN(n19123) );
  NAND2_X1 U22270 ( .A1(n19122), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19126) );
  NAND3_X1 U22271 ( .A1(n19123), .A2(n19254), .A3(n19126), .ZN(P3_U3030) );
  INV_X1 U22272 ( .A(n19126), .ZN(n19124) );
  AOI21_X1 U22273 ( .B1(n19130), .B2(n19125), .A(n19124), .ZN(n19131) );
  OAI22_X1 U22274 ( .A1(NA), .A2(n19126), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19127) );
  OAI22_X1 U22275 ( .A1(n19128), .A2(n19127), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19129) );
  OAI22_X1 U22276 ( .A1(n19131), .A2(n19132), .B1(n19130), .B2(n19129), .ZN(
        P3_U3031) );
  OAI222_X1 U22277 ( .A1(n19237), .A2(n19189), .B1(n19133), .B2(n19265), .C1(
        n19134), .C2(n19180), .ZN(P3_U3032) );
  OAI222_X1 U22278 ( .A1(n19180), .A2(n19136), .B1(n19135), .B2(n19265), .C1(
        n19134), .C2(n19189), .ZN(P3_U3033) );
  OAI222_X1 U22279 ( .A1(n19180), .A2(n19138), .B1(n19137), .B2(n19265), .C1(
        n19136), .C2(n19189), .ZN(P3_U3034) );
  INV_X1 U22280 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19141) );
  OAI222_X1 U22281 ( .A1(n19180), .A2(n19141), .B1(n19139), .B2(n19265), .C1(
        n19138), .C2(n19189), .ZN(P3_U3035) );
  OAI222_X1 U22282 ( .A1(n19141), .A2(n19189), .B1(n19140), .B2(n19265), .C1(
        n19142), .C2(n19180), .ZN(P3_U3036) );
  OAI222_X1 U22283 ( .A1(n19180), .A2(n19144), .B1(n19143), .B2(n19265), .C1(
        n19142), .C2(n19189), .ZN(P3_U3037) );
  OAI222_X1 U22284 ( .A1(n19180), .A2(n19147), .B1(n19145), .B2(n19265), .C1(
        n19144), .C2(n19189), .ZN(P3_U3038) );
  OAI222_X1 U22285 ( .A1(n19147), .A2(n19189), .B1(n19146), .B2(n19265), .C1(
        n19148), .C2(n19180), .ZN(P3_U3039) );
  OAI222_X1 U22286 ( .A1(n19180), .A2(n19150), .B1(n19149), .B2(n19265), .C1(
        n19148), .C2(n19189), .ZN(P3_U3040) );
  OAI222_X1 U22287 ( .A1(n19180), .A2(n19152), .B1(n19151), .B2(n19265), .C1(
        n19150), .C2(n19189), .ZN(P3_U3041) );
  OAI222_X1 U22288 ( .A1(n19180), .A2(n19154), .B1(n19153), .B2(n19265), .C1(
        n19152), .C2(n19189), .ZN(P3_U3042) );
  OAI222_X1 U22289 ( .A1(n19180), .A2(n19156), .B1(n19155), .B2(n19265), .C1(
        n19154), .C2(n19189), .ZN(P3_U3043) );
  INV_X1 U22290 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19159) );
  OAI222_X1 U22291 ( .A1(n19180), .A2(n19159), .B1(n19157), .B2(n19265), .C1(
        n19156), .C2(n19189), .ZN(P3_U3044) );
  OAI222_X1 U22292 ( .A1(n19159), .A2(n19189), .B1(n19158), .B2(n19265), .C1(
        n19160), .C2(n19180), .ZN(P3_U3045) );
  OAI222_X1 U22293 ( .A1(n19180), .A2(n19162), .B1(n19161), .B2(n19265), .C1(
        n19160), .C2(n19195), .ZN(P3_U3046) );
  OAI222_X1 U22294 ( .A1(n19180), .A2(n19164), .B1(n19163), .B2(n19265), .C1(
        n19162), .C2(n19195), .ZN(P3_U3047) );
  OAI222_X1 U22295 ( .A1(n19180), .A2(n19166), .B1(n19165), .B2(n19265), .C1(
        n19164), .C2(n19195), .ZN(P3_U3048) );
  INV_X1 U22296 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19168) );
  OAI222_X1 U22297 ( .A1(n19180), .A2(n19168), .B1(n19167), .B2(n19265), .C1(
        n19166), .C2(n19195), .ZN(P3_U3049) );
  OAI222_X1 U22298 ( .A1(n19180), .A2(n19171), .B1(n19169), .B2(n19265), .C1(
        n19168), .C2(n19195), .ZN(P3_U3050) );
  OAI222_X1 U22299 ( .A1(n19171), .A2(n19189), .B1(n19170), .B2(n19265), .C1(
        n19172), .C2(n19180), .ZN(P3_U3051) );
  OAI222_X1 U22300 ( .A1(n19180), .A2(n19174), .B1(n19173), .B2(n19265), .C1(
        n19172), .C2(n19195), .ZN(P3_U3052) );
  OAI222_X1 U22301 ( .A1(n19180), .A2(n19176), .B1(n19175), .B2(n19265), .C1(
        n19174), .C2(n19195), .ZN(P3_U3053) );
  OAI222_X1 U22302 ( .A1(n19180), .A2(n19178), .B1(n19177), .B2(n19265), .C1(
        n19176), .C2(n19195), .ZN(P3_U3054) );
  OAI222_X1 U22303 ( .A1(n19180), .A2(n19181), .B1(n19179), .B2(n19265), .C1(
        n19178), .C2(n19195), .ZN(P3_U3055) );
  OAI222_X1 U22304 ( .A1(n19180), .A2(n19183), .B1(n19182), .B2(n19265), .C1(
        n19181), .C2(n19189), .ZN(P3_U3056) );
  OAI222_X1 U22305 ( .A1(n19180), .A2(n19185), .B1(n19184), .B2(n19265), .C1(
        n19183), .C2(n19189), .ZN(P3_U3057) );
  INV_X1 U22306 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19188) );
  OAI222_X1 U22307 ( .A1(n19180), .A2(n19188), .B1(n19186), .B2(n19265), .C1(
        n19185), .C2(n19189), .ZN(P3_U3058) );
  INV_X1 U22308 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19190) );
  OAI222_X1 U22309 ( .A1(n19188), .A2(n19189), .B1(n19187), .B2(n19265), .C1(
        n19190), .C2(n19180), .ZN(P3_U3059) );
  OAI222_X1 U22310 ( .A1(n19180), .A2(n19194), .B1(n19191), .B2(n19265), .C1(
        n19190), .C2(n19189), .ZN(P3_U3060) );
  INV_X1 U22311 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19193) );
  OAI222_X1 U22312 ( .A1(n19195), .A2(n19194), .B1(n19193), .B2(n19265), .C1(
        n19192), .C2(n19180), .ZN(P3_U3061) );
  OAI22_X1 U22313 ( .A1(n19266), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19265), .ZN(n19196) );
  INV_X1 U22314 ( .A(n19196), .ZN(P3_U3274) );
  OAI22_X1 U22315 ( .A1(n19266), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19265), .ZN(n19197) );
  INV_X1 U22316 ( .A(n19197), .ZN(P3_U3275) );
  OAI22_X1 U22317 ( .A1(n19266), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19265), .ZN(n19198) );
  INV_X1 U22318 ( .A(n19198), .ZN(P3_U3276) );
  OAI22_X1 U22319 ( .A1(n19266), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19265), .ZN(n19199) );
  INV_X1 U22320 ( .A(n19199), .ZN(P3_U3277) );
  OAI21_X1 U22321 ( .B1(n19203), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19201), 
        .ZN(n19200) );
  INV_X1 U22322 ( .A(n19200), .ZN(P3_U3280) );
  OAI21_X1 U22323 ( .B1(n19203), .B2(n19202), .A(n19201), .ZN(P3_U3281) );
  OAI221_X1 U22324 ( .B1(n19206), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19206), 
        .C2(n19205), .A(n19204), .ZN(P3_U3282) );
  INV_X1 U22325 ( .A(n19212), .ZN(n19269) );
  NOR2_X1 U22326 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19207), .ZN(
        n19210) );
  INV_X1 U22327 ( .A(n19208), .ZN(n19209) );
  AOI22_X1 U22328 ( .A1(n19269), .A2(n19210), .B1(n19230), .B2(n19209), .ZN(
        n19215) );
  INV_X1 U22329 ( .A(n19236), .ZN(n19233) );
  OAI21_X1 U22330 ( .B1(n19212), .B2(n19211), .A(n19233), .ZN(n19213) );
  INV_X1 U22331 ( .A(n19213), .ZN(n19214) );
  OAI22_X1 U22332 ( .A1(n19236), .A2(n19215), .B1(n19214), .B2(n9869), .ZN(
        P3_U3285) );
  NOR2_X1 U22333 ( .A1(n19216), .A2(n19232), .ZN(n19224) );
  OAI22_X1 U22334 ( .A1(n19218), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19217), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19223) );
  AOI222_X1 U22335 ( .A1(n19220), .A2(n19269), .B1(n19224), .B2(n19223), .C1(
        n19230), .C2(n19219), .ZN(n19221) );
  AOI22_X1 U22336 ( .A1(n19236), .A2(n9868), .B1(n19221), .B2(n19233), .ZN(
        P3_U3288) );
  INV_X1 U22337 ( .A(n19222), .ZN(n19226) );
  INV_X1 U22338 ( .A(n19223), .ZN(n19225) );
  AOI222_X1 U22339 ( .A1(n19227), .A2(n19269), .B1(n19230), .B2(n19226), .C1(
        n19225), .C2(n19224), .ZN(n19228) );
  AOI22_X1 U22340 ( .A1(n19236), .A2(n19229), .B1(n19228), .B2(n19233), .ZN(
        P3_U3289) );
  AOI222_X1 U22341 ( .A1(n19232), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19269), 
        .B2(n19231), .C1(n19235), .C2(n19230), .ZN(n19234) );
  AOI22_X1 U22342 ( .A1(n19236), .A2(n19235), .B1(n19234), .B2(n19233), .ZN(
        P3_U3290) );
  AOI21_X1 U22343 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19238) );
  AOI22_X1 U22344 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19238), .B2(n19237), .ZN(n19240) );
  INV_X1 U22345 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19239) );
  AOI22_X1 U22346 ( .A1(n19241), .A2(n19240), .B1(n19239), .B2(n19244), .ZN(
        P3_U3292) );
  INV_X1 U22347 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19245) );
  NOR2_X1 U22348 ( .A1(n19244), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19242) );
  AOI22_X1 U22349 ( .A1(n19245), .A2(n19244), .B1(n19243), .B2(n19242), .ZN(
        P3_U3293) );
  INV_X1 U22350 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19270) );
  OAI22_X1 U22351 ( .A1(n19266), .A2(n19270), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19265), .ZN(n19246) );
  INV_X1 U22352 ( .A(n19246), .ZN(P3_U3294) );
  MUX2_X1 U22353 ( .A(P3_MORE_REG_SCAN_IN), .B(n19248), .S(n19247), .Z(
        P3_U3295) );
  OAI21_X1 U22354 ( .B1(n19251), .B2(n19250), .A(n19249), .ZN(n19252) );
  AOI21_X1 U22355 ( .B1(n19253), .B2(n19257), .A(n19252), .ZN(n19264) );
  AOI21_X1 U22356 ( .B1(n19256), .B2(n19255), .A(n19254), .ZN(n19259) );
  OAI211_X1 U22357 ( .C1(n19259), .C2(n19258), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19257), .ZN(n19261) );
  AOI21_X1 U22358 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19261), .A(n19260), 
        .ZN(n19263) );
  NAND2_X1 U22359 ( .A1(n19264), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19262) );
  OAI21_X1 U22360 ( .B1(n19264), .B2(n19263), .A(n19262), .ZN(P3_U3296) );
  OAI22_X1 U22361 ( .A1(n19266), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19265), .ZN(n19267) );
  INV_X1 U22362 ( .A(n19267), .ZN(P3_U3297) );
  AOI21_X1 U22363 ( .B1(n19269), .B2(n19268), .A(n19271), .ZN(n19275) );
  AOI22_X1 U22364 ( .A1(n19272), .A2(n19271), .B1(n19275), .B2(n19270), .ZN(
        P3_U3298) );
  INV_X1 U22365 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19274) );
  AOI21_X1 U22366 ( .B1(n19275), .B2(n19274), .A(n19273), .ZN(P3_U3299) );
  AOI21_X1 U22367 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n19277), .A(n19276), 
        .ZN(n19278) );
  INV_X1 U22368 ( .A(n19278), .ZN(P2_U2814) );
  INV_X1 U22369 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19284) );
  NAND2_X1 U22370 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20183), .ZN(n20172) );
  NAND2_X1 U22371 ( .A1(n19284), .A2(n19279), .ZN(n20169) );
  OAI21_X1 U22372 ( .B1(n19284), .B2(n20172), .A(n20169), .ZN(n20239) );
  AOI21_X1 U22373 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20239), .ZN(n19280) );
  INV_X1 U22374 ( .A(n19280), .ZN(P2_U2815) );
  NAND2_X1 U22375 ( .A1(n19955), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20156) );
  INV_X1 U22376 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19281) );
  OAI22_X1 U22377 ( .A1(n19283), .A2(n20156), .B1(n19282), .B2(n19281), .ZN(
        P2_U2816) );
  NAND2_X1 U22378 ( .A1(n19284), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20293) );
  INV_X2 U22379 ( .A(n20293), .ZN(n20229) );
  AOI21_X1 U22380 ( .B1(n19284), .B2(n20183), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19285) );
  AOI22_X1 U22381 ( .A1(n20229), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19285), 
        .B2(n20293), .ZN(P2_U2817) );
  OAI21_X1 U22382 ( .B1(n20176), .B2(BS16), .A(n20239), .ZN(n20237) );
  OAI21_X1 U22383 ( .B1(n20239), .B2(n20049), .A(n20237), .ZN(P2_U2818) );
  NOR2_X1 U22384 ( .A1(n19287), .A2(n19286), .ZN(n20283) );
  OAI21_X1 U22385 ( .B1(n20283), .B2(n19289), .A(n19288), .ZN(P2_U2819) );
  NOR4_X1 U22386 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19293) );
  NOR4_X1 U22387 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19292) );
  NOR4_X1 U22388 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19291) );
  NOR4_X1 U22389 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19290) );
  NAND4_X1 U22390 ( .A1(n19293), .A2(n19292), .A3(n19291), .A4(n19290), .ZN(
        n19299) );
  NOR4_X1 U22391 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19297) );
  AOI211_X1 U22392 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19296) );
  NOR4_X1 U22393 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19295) );
  NOR4_X1 U22394 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19294) );
  NAND4_X1 U22395 ( .A1(n19297), .A2(n19296), .A3(n19295), .A4(n19294), .ZN(
        n19298) );
  NOR2_X1 U22396 ( .A1(n19299), .A2(n19298), .ZN(n19310) );
  INV_X1 U22397 ( .A(n19310), .ZN(n19308) );
  NOR2_X1 U22398 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19308), .ZN(n19302) );
  INV_X1 U22399 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19300) );
  AOI22_X1 U22400 ( .A1(n19302), .A2(n19303), .B1(n19308), .B2(n19300), .ZN(
        P2_U2820) );
  OR3_X1 U22401 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19307) );
  INV_X1 U22402 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22403 ( .A1(n19302), .A2(n19307), .B1(n19308), .B2(n19301), .ZN(
        P2_U2821) );
  INV_X1 U22404 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20238) );
  NAND2_X1 U22405 ( .A1(n19302), .A2(n20238), .ZN(n19306) );
  OAI21_X1 U22406 ( .B1(n19303), .B2(n20184), .A(n19310), .ZN(n19304) );
  OAI21_X1 U22407 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19310), .A(n19304), 
        .ZN(n19305) );
  OAI221_X1 U22408 ( .B1(n19306), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19306), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19305), .ZN(P2_U2822) );
  INV_X1 U22409 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19309) );
  OAI221_X1 U22410 ( .B1(n19310), .B2(n19309), .C1(n19308), .C2(n19307), .A(
        n19306), .ZN(P2_U2823) );
  AOI22_X1 U22411 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19443), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19444), .ZN(n19320) );
  AOI22_X1 U22412 ( .A1(n19311), .A2(n19448), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19459), .ZN(n19319) );
  AOI22_X1 U22413 ( .A1(n19313), .A2(n19437), .B1(n19450), .B2(n19312), .ZN(
        n19318) );
  OAI211_X1 U22414 ( .C1(n19316), .C2(n19315), .A(n19420), .B(n19314), .ZN(
        n19317) );
  NAND4_X1 U22415 ( .A1(n19320), .A2(n19319), .A3(n19318), .A4(n19317), .ZN(
        P2_U2834) );
  INV_X1 U22416 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20209) );
  OAI21_X1 U22417 ( .B1(n20209), .B2(n19425), .A(n19424), .ZN(n19325) );
  INV_X1 U22418 ( .A(n19321), .ZN(n19323) );
  OAI22_X1 U22419 ( .A1(n19323), .A2(n19427), .B1(n19390), .B2(n19322), .ZN(
        n19324) );
  AOI211_X1 U22420 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19443), .A(n19325), .B(
        n19324), .ZN(n19334) );
  OAI22_X1 U22421 ( .A1(n19327), .A2(n19453), .B1(n19326), .B2(n19442), .ZN(
        n19328) );
  INV_X1 U22422 ( .A(n19328), .ZN(n19333) );
  OAI211_X1 U22423 ( .C1(n19331), .C2(n19330), .A(n19420), .B(n19329), .ZN(
        n19332) );
  NAND3_X1 U22424 ( .A1(n19334), .A2(n19333), .A3(n19332), .ZN(P2_U2836) );
  OAI21_X1 U22425 ( .B1(n20206), .B2(n19425), .A(n19424), .ZN(n19338) );
  OAI22_X1 U22426 ( .A1(n19336), .A2(n19427), .B1(n19390), .B2(n19335), .ZN(
        n19337) );
  AOI211_X1 U22427 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19443), .A(n19338), .B(
        n19337), .ZN(n19345) );
  NAND2_X1 U22428 ( .A1(n9647), .A2(n19339), .ZN(n19340) );
  XOR2_X1 U22429 ( .A(n19341), .B(n19340), .Z(n19343) );
  AOI22_X1 U22430 ( .A1(n19343), .A2(n19438), .B1(n19342), .B2(n19437), .ZN(
        n19344) );
  OAI211_X1 U22431 ( .C1(n19346), .C2(n19442), .A(n19345), .B(n19344), .ZN(
        P2_U2838) );
  AOI211_X1 U22432 ( .C1(n19354), .C2(n19348), .A(n20159), .B(n19347), .ZN(
        n19349) );
  INV_X1 U22433 ( .A(n19349), .ZN(n19351) );
  AOI22_X1 U22434 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19459), .ZN(n19350) );
  OAI211_X1 U22435 ( .C1(n19427), .C2(n19352), .A(n19351), .B(n19350), .ZN(
        n19353) );
  AOI211_X1 U22436 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19444), .A(n19592), 
        .B(n19353), .ZN(n19357) );
  AOI22_X1 U22437 ( .A1(n19355), .A2(n19437), .B1(n19354), .B2(n19458), .ZN(
        n19356) );
  OAI211_X1 U22438 ( .C1(n19506), .C2(n19442), .A(n19357), .B(n19356), .ZN(
        P2_U2840) );
  NOR2_X1 U22439 ( .A1(n19416), .A2(n19358), .ZN(n19360) );
  XOR2_X1 U22440 ( .A(n19360), .B(n19359), .Z(n19368) );
  AOI22_X1 U22441 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19459), .ZN(n19361) );
  OAI21_X1 U22442 ( .B1(n19362), .B2(n19427), .A(n19361), .ZN(n19363) );
  AOI211_X1 U22443 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19444), .A(n19592), 
        .B(n19363), .ZN(n19367) );
  INV_X1 U22444 ( .A(n19513), .ZN(n19364) );
  OAI22_X1 U22445 ( .A1(n19475), .A2(n19453), .B1(n19364), .B2(n19442), .ZN(
        n19365) );
  INV_X1 U22446 ( .A(n19365), .ZN(n19366) );
  OAI211_X1 U22447 ( .C1(n20159), .C2(n19368), .A(n19367), .B(n19366), .ZN(
        P2_U2843) );
  AOI22_X1 U22448 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19443), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19459), .ZN(n19369) );
  OAI21_X1 U22449 ( .B1(n19370), .B2(n19427), .A(n19369), .ZN(n19371) );
  AOI211_X1 U22450 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19444), .A(n19592), 
        .B(n19371), .ZN(n19378) );
  NAND2_X1 U22451 ( .A1(n9647), .A2(n19372), .ZN(n19374) );
  XNOR2_X1 U22452 ( .A(n19374), .B(n19373), .ZN(n19376) );
  AOI22_X1 U22453 ( .A1(n19376), .A2(n19420), .B1(n19375), .B2(n19437), .ZN(
        n19377) );
  OAI211_X1 U22454 ( .C1(n19516), .C2(n19442), .A(n19378), .B(n19377), .ZN(
        P2_U2844) );
  NOR2_X1 U22455 ( .A1(n19416), .A2(n19379), .ZN(n19380) );
  XOR2_X1 U22456 ( .A(n19381), .B(n19380), .Z(n19387) );
  AOI22_X1 U22457 ( .A1(n19382), .A2(n19448), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19459), .ZN(n19383) );
  OAI211_X1 U22458 ( .C1(n12603), .C2(n19425), .A(n19383), .B(n19424), .ZN(
        n19385) );
  OAI22_X1 U22459 ( .A1(n19478), .A2(n19453), .B1(n19442), .B2(n19519), .ZN(
        n19384) );
  AOI211_X1 U22460 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19443), .A(n19385), .B(
        n19384), .ZN(n19386) );
  OAI21_X1 U22461 ( .B1(n20159), .B2(n19387), .A(n19386), .ZN(P2_U2845) );
  OAI21_X1 U22462 ( .B1(n12600), .B2(n19425), .A(n19424), .ZN(n19393) );
  INV_X1 U22463 ( .A(n19388), .ZN(n19391) );
  OAI22_X1 U22464 ( .A1(n19391), .A2(n19427), .B1(n19390), .B2(n19389), .ZN(
        n19392) );
  AOI211_X1 U22465 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19443), .A(n19393), .B(
        n19392), .ZN(n19400) );
  NAND2_X1 U22466 ( .A1(n9647), .A2(n19394), .ZN(n19395) );
  XNOR2_X1 U22467 ( .A(n19396), .B(n19395), .ZN(n19398) );
  AOI22_X1 U22468 ( .A1(n19398), .A2(n19420), .B1(n19397), .B2(n19437), .ZN(
        n19399) );
  OAI211_X1 U22469 ( .C1(n19521), .C2(n19442), .A(n19400), .B(n19399), .ZN(
        P2_U2846) );
  NAND2_X1 U22470 ( .A1(n9647), .A2(n19401), .ZN(n19403) );
  XOR2_X1 U22471 ( .A(n19403), .B(n19402), .Z(n19410) );
  AOI22_X1 U22472 ( .A1(n19404), .A2(n19448), .B1(n19443), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n19405) );
  OAI211_X1 U22473 ( .C1(n20194), .C2(n19425), .A(n19405), .B(n19424), .ZN(
        n19408) );
  OAI22_X1 U22474 ( .A1(n19527), .A2(n19442), .B1(n19453), .B2(n19406), .ZN(
        n19407) );
  AOI211_X1 U22475 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19459), .A(
        n19408), .B(n19407), .ZN(n19409) );
  OAI21_X1 U22476 ( .B1(n19410), .B2(n20159), .A(n19409), .ZN(P2_U2848) );
  OAI21_X1 U22477 ( .B1(n20192), .B2(n19425), .A(n19424), .ZN(n19414) );
  OAI22_X1 U22478 ( .A1(n19429), .A2(n19412), .B1(n19427), .B2(n19411), .ZN(
        n19413) );
  AOI211_X1 U22479 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19459), .A(
        n19414), .B(n19413), .ZN(n19423) );
  NOR2_X1 U22480 ( .A1(n19416), .A2(n19415), .ZN(n19418) );
  XNOR2_X1 U22481 ( .A(n19418), .B(n19417), .ZN(n19421) );
  AOI22_X1 U22482 ( .A1(n19421), .A2(n19420), .B1(n19437), .B2(n19419), .ZN(
        n19422) );
  OAI211_X1 U22483 ( .C1(n19442), .C2(n19530), .A(n19423), .B(n19422), .ZN(
        P2_U2849) );
  OAI21_X1 U22484 ( .B1(n20190), .B2(n19425), .A(n19424), .ZN(n19431) );
  OAI22_X1 U22485 ( .A1(n19429), .A2(n19428), .B1(n19427), .B2(n19426), .ZN(
        n19430) );
  AOI211_X1 U22486 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19459), .A(
        n19431), .B(n19430), .ZN(n19441) );
  NAND2_X1 U22487 ( .A1(n9647), .A2(n19432), .ZN(n19434) );
  XNOR2_X1 U22488 ( .A(n19435), .B(n19434), .ZN(n19439) );
  AOI22_X1 U22489 ( .A1(n19439), .A2(n19438), .B1(n19437), .B2(n19436), .ZN(
        n19440) );
  OAI211_X1 U22490 ( .C1(n19442), .C2(n19531), .A(n19441), .B(n19440), .ZN(
        P2_U2850) );
  AOI22_X1 U22491 ( .A1(n19444), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19443), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19452) );
  INV_X1 U22492 ( .A(n19445), .ZN(n19449) );
  INV_X1 U22493 ( .A(n19446), .ZN(n19447) );
  AOI22_X1 U22494 ( .A1(n19450), .A2(n19449), .B1(n19448), .B2(n19447), .ZN(
        n19451) );
  OAI211_X1 U22495 ( .C1(n19454), .C2(n19453), .A(n19452), .B(n19451), .ZN(
        n19455) );
  AOI21_X1 U22496 ( .B1(n19457), .B2(n19456), .A(n19455), .ZN(n19461) );
  OAI21_X1 U22497 ( .B1(n19459), .B2(n19458), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19460) );
  OAI211_X1 U22498 ( .C1(n19462), .C2(n20159), .A(n19461), .B(n19460), .ZN(
        P2_U2855) );
  AND2_X1 U22499 ( .A1(n19464), .A2(n19463), .ZN(n19466) );
  OR2_X1 U22500 ( .A1(n19466), .A2(n19465), .ZN(n19500) );
  OAI22_X1 U22501 ( .A1(n19500), .A2(n19481), .B1(n19490), .B2(n19467), .ZN(
        n19468) );
  INV_X1 U22502 ( .A(n19468), .ZN(n19469) );
  OAI21_X1 U22503 ( .B1(n19484), .B2(n19470), .A(n19469), .ZN(P2_U2871) );
  XOR2_X1 U22504 ( .A(n19472), .B(n19471), .Z(n19473) );
  AOI22_X1 U22505 ( .A1(n19473), .A2(n19487), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19484), .ZN(n19474) );
  OAI21_X1 U22506 ( .B1(n19475), .B2(n19484), .A(n19474), .ZN(P2_U2875) );
  XNOR2_X1 U22507 ( .A(n13486), .B(n9753), .ZN(n19476) );
  AOI22_X1 U22508 ( .A1(n19476), .A2(n19487), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19484), .ZN(n19477) );
  OAI21_X1 U22509 ( .B1(n19478), .B2(n19484), .A(n19477), .ZN(P2_U2877) );
  AOI21_X1 U22510 ( .B1(n19480), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n19479), .ZN(n19482) );
  NOR3_X1 U22511 ( .A1(n19482), .A2(n10051), .A3(n19481), .ZN(n19483) );
  AOI21_X1 U22512 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19484), .A(n19483), .ZN(
        n19485) );
  OAI21_X1 U22513 ( .B1(n19486), .B2(n19484), .A(n19485), .ZN(P2_U2879) );
  AOI22_X1 U22514 ( .A1(n19488), .A2(n19487), .B1(n19490), .B2(n19596), .ZN(
        n19489) );
  OAI21_X1 U22515 ( .B1(n19490), .B2(n12803), .A(n19489), .ZN(P2_U2883) );
  AOI22_X1 U22516 ( .A1(n19491), .A2(n19547), .B1(n19497), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19493) );
  AOI22_X1 U22517 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19546), .B1(n19496), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19492) );
  NAND2_X1 U22518 ( .A1(n19493), .A2(n19492), .ZN(P2_U2888) );
  AOI22_X1 U22519 ( .A1(n19495), .A2(n19494), .B1(n19546), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19504) );
  AOI22_X1 U22520 ( .A1(n19497), .A2(BUF2_REG_16__SCAN_IN), .B1(n19496), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19503) );
  INV_X1 U22521 ( .A(n19498), .ZN(n19499) );
  OAI22_X1 U22522 ( .A1(n19500), .A2(n19551), .B1(n19538), .B2(n19499), .ZN(
        n19501) );
  INV_X1 U22523 ( .A(n19501), .ZN(n19502) );
  NAND3_X1 U22524 ( .A1(n19504), .A2(n19503), .A3(n19502), .ZN(P2_U2903) );
  OAI222_X1 U22525 ( .A1(n19506), .A2(n19529), .B1(n12958), .B2(n19537), .C1(
        n19505), .C2(n19555), .ZN(P2_U2904) );
  INV_X1 U22526 ( .A(n19529), .ZN(n19534) );
  AOI22_X1 U22527 ( .A1(n19508), .A2(n19534), .B1(n19507), .B2(n19522), .ZN(
        n19509) );
  OAI21_X1 U22528 ( .B1(n19537), .B2(n19561), .A(n19509), .ZN(P2_U2905) );
  INV_X1 U22529 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19563) );
  OAI222_X1 U22530 ( .A1(n19511), .A2(n19529), .B1(n19563), .B2(n19537), .C1(
        n19555), .C2(n19510), .ZN(P2_U2906) );
  AOI22_X1 U22531 ( .A1(n19513), .A2(n19534), .B1(n19512), .B2(n19522), .ZN(
        n19514) );
  OAI21_X1 U22532 ( .B1(n19537), .B2(n19565), .A(n19514), .ZN(P2_U2907) );
  INV_X1 U22533 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19567) );
  OAI222_X1 U22534 ( .A1(n19516), .A2(n19529), .B1(n19567), .B2(n19537), .C1(
        n19555), .C2(n19515), .ZN(P2_U2908) );
  AOI22_X1 U22535 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19546), .B1(n19517), 
        .B2(n19522), .ZN(n19518) );
  OAI21_X1 U22536 ( .B1(n19529), .B2(n19519), .A(n19518), .ZN(P2_U2909) );
  INV_X1 U22537 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19571) );
  OAI222_X1 U22538 ( .A1(n19521), .A2(n19529), .B1(n19571), .B2(n19537), .C1(
        n19555), .C2(n19520), .ZN(P2_U2910) );
  AOI22_X1 U22539 ( .A1(n19524), .A2(n19534), .B1(n19523), .B2(n19522), .ZN(
        n19525) );
  OAI21_X1 U22540 ( .B1(n19537), .B2(n19574), .A(n19525), .ZN(P2_U2911) );
  OAI222_X1 U22541 ( .A1(n19527), .A2(n19529), .B1(n19576), .B2(n19537), .C1(
        n19555), .C2(n19526), .ZN(P2_U2912) );
  INV_X1 U22542 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19578) );
  OAI222_X1 U22543 ( .A1(n19530), .A2(n19529), .B1(n19578), .B2(n19537), .C1(
        n19555), .C2(n19528), .ZN(P2_U2913) );
  OAI21_X1 U22544 ( .B1(n19532), .B2(n19551), .A(n19531), .ZN(n19533) );
  AOI22_X1 U22545 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19546), .B1(n19534), .B2(
        n19533), .ZN(n19535) );
  OAI21_X1 U22546 ( .B1(n19651), .B2(n19555), .A(n19535), .ZN(P2_U2914) );
  INV_X1 U22547 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19536) );
  OAI22_X1 U22548 ( .A1(n20240), .A2(n19538), .B1(n19537), .B2(n19536), .ZN(
        n19539) );
  INV_X1 U22549 ( .A(n19539), .ZN(n19545) );
  AOI21_X1 U22550 ( .B1(n19542), .B2(n19541), .A(n19540), .ZN(n19543) );
  OR2_X1 U22551 ( .A1(n19543), .A2(n19551), .ZN(n19544) );
  OAI211_X1 U22552 ( .C1(n19643), .C2(n19555), .A(n19545), .B(n19544), .ZN(
        P2_U2916) );
  AOI22_X1 U22553 ( .A1(n19547), .A2(n20270), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19546), .ZN(n19554) );
  AOI21_X1 U22554 ( .B1(n19550), .B2(n19549), .A(n19548), .ZN(n19552) );
  OR2_X1 U22555 ( .A1(n19552), .A2(n19551), .ZN(n19553) );
  OAI211_X1 U22556 ( .C1(n19556), .C2(n19555), .A(n19554), .B(n19553), .ZN(
        P2_U2918) );
  AND2_X1 U22557 ( .A1(n19557), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22558 ( .A1(n19572), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19559) );
  OAI21_X1 U22559 ( .B1(n12958), .B2(n19591), .A(n19559), .ZN(P2_U2936) );
  AOI22_X1 U22560 ( .A1(n19572), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19560) );
  OAI21_X1 U22561 ( .B1(n19561), .B2(n19591), .A(n19560), .ZN(P2_U2937) );
  AOI22_X1 U22562 ( .A1(n19572), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19562) );
  OAI21_X1 U22563 ( .B1(n19563), .B2(n19591), .A(n19562), .ZN(P2_U2938) );
  AOI22_X1 U22564 ( .A1(n19572), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19564) );
  OAI21_X1 U22565 ( .B1(n19565), .B2(n19591), .A(n19564), .ZN(P2_U2939) );
  AOI22_X1 U22566 ( .A1(n19572), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19566) );
  OAI21_X1 U22567 ( .B1(n19567), .B2(n19591), .A(n19566), .ZN(P2_U2940) );
  AOI22_X1 U22568 ( .A1(n19572), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19568) );
  OAI21_X1 U22569 ( .B1(n19569), .B2(n19591), .A(n19568), .ZN(P2_U2941) );
  AOI22_X1 U22570 ( .A1(n19572), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19570) );
  OAI21_X1 U22571 ( .B1(n19571), .B2(n19591), .A(n19570), .ZN(P2_U2942) );
  AOI22_X1 U22572 ( .A1(n19572), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19573) );
  OAI21_X1 U22573 ( .B1(n19574), .B2(n19591), .A(n19573), .ZN(P2_U2943) );
  AOI22_X1 U22574 ( .A1(n19589), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19575) );
  OAI21_X1 U22575 ( .B1(n19576), .B2(n19591), .A(n19575), .ZN(P2_U2944) );
  AOI22_X1 U22576 ( .A1(n19589), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19577) );
  OAI21_X1 U22577 ( .B1(n19578), .B2(n19591), .A(n19577), .ZN(P2_U2945) );
  INV_X1 U22578 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U22579 ( .A1(n19589), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19579) );
  OAI21_X1 U22580 ( .B1(n19580), .B2(n19591), .A(n19579), .ZN(P2_U2946) );
  INV_X1 U22581 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19582) );
  AOI22_X1 U22582 ( .A1(n19589), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19581) );
  OAI21_X1 U22583 ( .B1(n19582), .B2(n19591), .A(n19581), .ZN(P2_U2947) );
  AOI22_X1 U22584 ( .A1(n19589), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19583) );
  OAI21_X1 U22585 ( .B1(n19536), .B2(n19591), .A(n19583), .ZN(P2_U2948) );
  INV_X1 U22586 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19585) );
  AOI22_X1 U22587 ( .A1(n19589), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19584) );
  OAI21_X1 U22588 ( .B1(n19585), .B2(n19591), .A(n19584), .ZN(P2_U2949) );
  INV_X1 U22589 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19587) );
  AOI22_X1 U22590 ( .A1(n19589), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19586) );
  OAI21_X1 U22591 ( .B1(n19587), .B2(n19591), .A(n19586), .ZN(P2_U2950) );
  AOI22_X1 U22592 ( .A1(n19589), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19588), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19590) );
  OAI21_X1 U22593 ( .B1(n13061), .B2(n19591), .A(n19590), .ZN(P2_U2951) );
  AOI22_X1 U22594 ( .A1(n19593), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19592), .ZN(n19601) );
  AOI222_X1 U22595 ( .A1(n19599), .A2(n19598), .B1(n19597), .B2(n19596), .C1(
        n19595), .C2(n19594), .ZN(n19600) );
  OAI211_X1 U22596 ( .C1(n19603), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P2_U3010) );
  AOI22_X1 U22597 ( .A1(n19606), .A2(n19605), .B1(n19604), .B2(n20270), .ZN(
        n19621) );
  AOI21_X1 U22598 ( .B1(n19608), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19607), .ZN(n19616) );
  INV_X1 U22599 ( .A(n19609), .ZN(n19610) );
  NAND2_X1 U22600 ( .A1(n19611), .A2(n19610), .ZN(n19615) );
  NAND2_X1 U22601 ( .A1(n19613), .A2(n19612), .ZN(n19614) );
  AND3_X1 U22602 ( .A1(n19616), .A2(n19615), .A3(n19614), .ZN(n19620) );
  OAI211_X1 U22603 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19618), .B(n19617), .ZN(n19619) );
  NAND3_X1 U22604 ( .A1(n19621), .A2(n19620), .A3(n19619), .ZN(P2_U3045) );
  NAND2_X1 U22605 ( .A1(n19731), .A2(n20272), .ZN(n19670) );
  NOR2_X1 U22606 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19670), .ZN(
        n19660) );
  AOI22_X1 U22607 ( .A1(n20147), .A2(n20100), .B1(n20092), .B2(n19660), .ZN(
        n19633) );
  INV_X1 U22608 ( .A(n19628), .ZN(n19622) );
  AOI21_X1 U22609 ( .B1(n19622), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19626) );
  AOI21_X1 U22610 ( .B1(n20134), .B2(n19690), .A(n20049), .ZN(n19623) );
  NOR2_X1 U22611 ( .A1(n19623), .A2(n20245), .ZN(n19627) );
  NOR2_X1 U22612 ( .A1(n20254), .A2(n19624), .ZN(n20142) );
  NOR2_X1 U22613 ( .A1(n20142), .A2(n19660), .ZN(n19630) );
  NAND2_X1 U22614 ( .A1(n19627), .A2(n19630), .ZN(n19625) );
  OAI211_X1 U22615 ( .C1(n19660), .C2(n19626), .A(n19625), .B(n20098), .ZN(
        n19663) );
  INV_X1 U22616 ( .A(n19627), .ZN(n19631) );
  OAI21_X1 U22617 ( .B1(n19628), .B2(n19660), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19629) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19663), .B1(
        n16038), .B2(n19662), .ZN(n19632) );
  OAI211_X1 U22619 ( .C1(n20103), .C2(n19690), .A(n19633), .B(n19632), .ZN(
        P2_U3048) );
  INV_X1 U22620 ( .A(n19660), .ZN(n19641) );
  OAI22_X1 U22621 ( .A1(n20134), .A2(n20109), .B1(n20062), .B2(n19641), .ZN(
        n19634) );
  INV_X1 U22622 ( .A(n19634), .ZN(n19636) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19663), .B1(
        n20105), .B2(n19662), .ZN(n19635) );
  OAI211_X1 U22624 ( .C1(n20066), .C2(n19690), .A(n19636), .B(n19635), .ZN(
        P2_U3049) );
  AOI22_X1 U22625 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19656), .ZN(n20115) );
  AOI22_X1 U22626 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19656), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19657), .ZN(n20070) );
  NOR2_X2 U22627 ( .A1(n11915), .A2(n19637), .ZN(n20110) );
  AOI22_X1 U22628 ( .A1(n20147), .A2(n20112), .B1(n20110), .B2(n19660), .ZN(
        n19640) );
  NOR2_X2 U22629 ( .A1(n19638), .A2(n19782), .ZN(n20111) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19663), .B1(
        n20111), .B2(n19662), .ZN(n19639) );
  OAI211_X1 U22631 ( .C1(n20115), .C2(n19690), .A(n19640), .B(n19639), .ZN(
        P2_U3050) );
  AOI22_X1 U22632 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19656), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19657), .ZN(n20073) );
  AND2_X1 U22633 ( .A1(n11914), .A2(n19658), .ZN(n20116) );
  INV_X1 U22634 ( .A(n20116), .ZN(n20072) );
  OAI22_X1 U22635 ( .A1(n20134), .A2(n20073), .B1(n20072), .B2(n19641), .ZN(
        n19642) );
  INV_X1 U22636 ( .A(n19642), .ZN(n19645) );
  NOR2_X2 U22637 ( .A1(n19643), .A2(n19782), .ZN(n20117) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19663), .B1(
        n20117), .B2(n19662), .ZN(n19644) );
  OAI211_X1 U22639 ( .C1(n20121), .C2(n19690), .A(n19645), .B(n19644), .ZN(
        P2_U3051) );
  AOI22_X1 U22640 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19656), .ZN(n20034) );
  AOI22_X1 U22641 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19656), .ZN(n20127) );
  AOI22_X1 U22642 ( .A1(n20147), .A2(n20031), .B1(n20122), .B2(n19660), .ZN(
        n19649) );
  NOR2_X2 U22643 ( .A1(n19647), .A2(n19782), .ZN(n20123) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19663), .B1(
        n20123), .B2(n19662), .ZN(n19648) );
  OAI211_X1 U22645 ( .C1(n20034), .C2(n19690), .A(n19649), .B(n19648), .ZN(
        P2_U3052) );
  AOI22_X1 U22646 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19656), .ZN(n20135) );
  AOI22_X1 U22647 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19656), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19657), .ZN(n20082) );
  INV_X1 U22648 ( .A(n20082), .ZN(n20130) );
  AOI22_X1 U22649 ( .A1(n20147), .A2(n20130), .B1(n20128), .B2(n19660), .ZN(
        n19653) );
  NOR2_X2 U22650 ( .A1(n19651), .A2(n19782), .ZN(n20129) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19663), .B1(
        n20129), .B2(n19662), .ZN(n19652) );
  OAI211_X1 U22652 ( .C1(n20135), .C2(n19690), .A(n19653), .B(n19652), .ZN(
        P2_U3053) );
  AOI22_X1 U22653 ( .A1(n20147), .A2(n20009), .B1(n20136), .B2(n19660), .ZN(
        n19655) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19663), .B1(
        n20137), .B2(n19662), .ZN(n19654) );
  OAI211_X1 U22655 ( .C1(n20012), .C2(n19690), .A(n19655), .B(n19654), .ZN(
        P2_U3054) );
  AOI22_X1 U22656 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19656), .ZN(n20044) );
  AOI22_X1 U22657 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19657), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19656), .ZN(n20152) );
  INV_X1 U22658 ( .A(n20152), .ZN(n20039) );
  AND2_X1 U22659 ( .A1(n19659), .A2(n19658), .ZN(n20143) );
  AOI22_X1 U22660 ( .A1(n20147), .A2(n20039), .B1(n20143), .B2(n19660), .ZN(
        n19665) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19663), .B1(
        n20144), .B2(n19662), .ZN(n19664) );
  OAI211_X1 U22662 ( .C1(n20044), .C2(n19690), .A(n19665), .B(n19664), .ZN(
        P2_U3055) );
  NAND2_X1 U22663 ( .A1(n19667), .A2(n19666), .ZN(n19704) );
  NOR2_X1 U22664 ( .A1(n19668), .A2(n19730), .ZN(n19691) );
  OAI21_X1 U22665 ( .B1(n14235), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19669) );
  OAI21_X1 U22666 ( .B1(n19670), .B2(n20245), .A(n19669), .ZN(n19692) );
  AOI22_X1 U22667 ( .A1(n19692), .A2(n16038), .B1(n20092), .B2(n19691), .ZN(
        n19677) );
  NAND2_X1 U22668 ( .A1(n20248), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20242) );
  OAI21_X1 U22669 ( .B1(n19671), .B2(n20242), .A(n19670), .ZN(n19675) );
  INV_X1 U22670 ( .A(n14235), .ZN(n19673) );
  INV_X1 U22671 ( .A(n19691), .ZN(n19672) );
  OAI211_X1 U22672 ( .C1(n19673), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19672), 
        .B(n20245), .ZN(n19674) );
  NAND3_X1 U22673 ( .A1(n19675), .A2(n20098), .A3(n19674), .ZN(n19694) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20100), .ZN(n19676) );
  OAI211_X1 U22675 ( .C1(n20103), .C2(n19704), .A(n19677), .B(n19676), .ZN(
        P2_U3056) );
  AOI22_X1 U22676 ( .A1(n19692), .A2(n20105), .B1(n20104), .B2(n19691), .ZN(
        n19679) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19694), .B1(
        n19726), .B2(n20106), .ZN(n19678) );
  OAI211_X1 U22678 ( .C1(n20109), .C2(n19690), .A(n19679), .B(n19678), .ZN(
        P2_U3057) );
  AOI22_X1 U22679 ( .A1(n19692), .A2(n20111), .B1(n20110), .B2(n19691), .ZN(
        n19681) );
  INV_X1 U22680 ( .A(n20115), .ZN(n20067) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19694), .B1(
        n19726), .B2(n20067), .ZN(n19680) );
  OAI211_X1 U22682 ( .C1(n20070), .C2(n19690), .A(n19681), .B(n19680), .ZN(
        P2_U3058) );
  AOI22_X1 U22683 ( .A1(n19692), .A2(n20117), .B1(n20116), .B2(n19691), .ZN(
        n19683) );
  INV_X1 U22684 ( .A(n20121), .ZN(n19884) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19694), .B1(
        n19726), .B2(n19884), .ZN(n19682) );
  OAI211_X1 U22686 ( .C1(n20073), .C2(n19690), .A(n19683), .B(n19682), .ZN(
        P2_U3059) );
  AOI22_X1 U22687 ( .A1(n19692), .A2(n20123), .B1(n20122), .B2(n19691), .ZN(
        n19685) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20031), .ZN(n19684) );
  OAI211_X1 U22689 ( .C1(n20034), .C2(n19704), .A(n19685), .B(n19684), .ZN(
        P2_U3060) );
  AOI22_X1 U22690 ( .A1(n19692), .A2(n20129), .B1(n20128), .B2(n19691), .ZN(
        n19687) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19694), .B1(
        n19726), .B2(n20079), .ZN(n19686) );
  OAI211_X1 U22692 ( .C1(n20082), .C2(n19690), .A(n19687), .B(n19686), .ZN(
        P2_U3061) );
  AOI22_X1 U22693 ( .A1(n19692), .A2(n20137), .B1(n20136), .B2(n19691), .ZN(
        n19689) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19694), .B1(
        n19726), .B2(n20138), .ZN(n19688) );
  OAI211_X1 U22695 ( .C1(n20141), .C2(n19690), .A(n19689), .B(n19688), .ZN(
        P2_U3062) );
  AOI22_X1 U22696 ( .A1(n19692), .A2(n20144), .B1(n20143), .B2(n19691), .ZN(
        n19696) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20039), .ZN(n19695) );
  OAI211_X1 U22698 ( .C1(n20044), .C2(n19704), .A(n19696), .B(n19695), .ZN(
        P2_U3063) );
  INV_X1 U22699 ( .A(n19698), .ZN(n19703) );
  AND2_X1 U22700 ( .A1(n19699), .A2(n19731), .ZN(n19724) );
  OAI21_X1 U22701 ( .B1(n19703), .B2(n19724), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19702) );
  NOR2_X1 U22702 ( .A1(n19700), .A2(n19730), .ZN(n19705) );
  INV_X1 U22703 ( .A(n19705), .ZN(n19701) );
  NAND2_X1 U22704 ( .A1(n19702), .A2(n19701), .ZN(n19725) );
  AOI22_X1 U22705 ( .A1(n19725), .A2(n16038), .B1(n20092), .B2(n19724), .ZN(
        n19711) );
  AOI21_X1 U22706 ( .B1(n19703), .B2(n20153), .A(n19724), .ZN(n19708) );
  NAND2_X1 U22707 ( .A1(n19753), .A2(n19704), .ZN(n19706) );
  AOI21_X1 U22708 ( .B1(n19706), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19705), 
        .ZN(n19707) );
  MUX2_X1 U22709 ( .A(n19708), .B(n19707), .S(n20243), .Z(n19709) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20100), .ZN(n19710) );
  OAI211_X1 U22711 ( .C1(n20103), .C2(n19753), .A(n19711), .B(n19710), .ZN(
        P2_U3064) );
  AOI22_X1 U22712 ( .A1(n19725), .A2(n20105), .B1(n20104), .B2(n19724), .ZN(
        n19713) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20023), .ZN(n19712) );
  OAI211_X1 U22714 ( .C1(n20066), .C2(n19753), .A(n19713), .B(n19712), .ZN(
        P2_U3065) );
  AOI22_X1 U22715 ( .A1(n19725), .A2(n20111), .B1(n20110), .B2(n19724), .ZN(
        n19715) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20112), .ZN(n19714) );
  OAI211_X1 U22717 ( .C1(n20115), .C2(n19753), .A(n19715), .B(n19714), .ZN(
        P2_U3066) );
  AOI22_X1 U22718 ( .A1(n19725), .A2(n20117), .B1(n20116), .B2(n19724), .ZN(
        n19717) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20118), .ZN(n19716) );
  OAI211_X1 U22720 ( .C1(n20121), .C2(n19753), .A(n19717), .B(n19716), .ZN(
        P2_U3067) );
  AOI22_X1 U22721 ( .A1(n19725), .A2(n20123), .B1(n20122), .B2(n19724), .ZN(
        n19719) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20031), .ZN(n19718) );
  OAI211_X1 U22723 ( .C1(n20034), .C2(n19753), .A(n19719), .B(n19718), .ZN(
        P2_U3068) );
  AOI22_X1 U22724 ( .A1(n19725), .A2(n20129), .B1(n20128), .B2(n19724), .ZN(
        n19721) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20130), .ZN(n19720) );
  OAI211_X1 U22726 ( .C1(n20135), .C2(n19753), .A(n19721), .B(n19720), .ZN(
        P2_U3069) );
  AOI22_X1 U22727 ( .A1(n19725), .A2(n20137), .B1(n20136), .B2(n19724), .ZN(
        n19723) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20009), .ZN(n19722) );
  OAI211_X1 U22729 ( .C1(n20012), .C2(n19753), .A(n19723), .B(n19722), .ZN(
        P2_U3070) );
  AOI22_X1 U22730 ( .A1(n19725), .A2(n20144), .B1(n20143), .B2(n19724), .ZN(
        n19729) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19727), .B1(
        n19726), .B2(n20039), .ZN(n19728) );
  OAI211_X1 U22732 ( .C1(n20044), .C2(n19753), .A(n19729), .B(n19728), .ZN(
        P2_U3071) );
  INV_X1 U22733 ( .A(n19753), .ZN(n19755) );
  NOR2_X1 U22734 ( .A1(n19949), .A2(n19730), .ZN(n19754) );
  AOI22_X1 U22735 ( .A1(n19755), .A2(n20100), .B1(n20092), .B2(n19754), .ZN(
        n19740) );
  OAI21_X1 U22736 ( .B1(n20244), .B2(n20242), .A(n20243), .ZN(n19738) );
  NAND2_X1 U22737 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19731), .ZN(
        n19737) );
  INV_X1 U22738 ( .A(n19737), .ZN(n19735) );
  INV_X1 U22739 ( .A(n14234), .ZN(n19733) );
  INV_X1 U22740 ( .A(n19754), .ZN(n19732) );
  OAI211_X1 U22741 ( .C1(n19733), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19732), 
        .B(n20245), .ZN(n19734) );
  OAI211_X1 U22742 ( .C1(n19738), .C2(n19735), .A(n20098), .B(n19734), .ZN(
        n19757) );
  OAI21_X1 U22743 ( .B1(n14234), .B2(n19754), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19736) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19757), .B1(
        n16038), .B2(n19756), .ZN(n19739) );
  OAI211_X1 U22745 ( .C1(n20103), .C2(n19780), .A(n19740), .B(n19739), .ZN(
        P2_U3072) );
  AOI22_X1 U22746 ( .A1(n19755), .A2(n20023), .B1(n20104), .B2(n19754), .ZN(
        n19742) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19757), .B1(
        n20105), .B2(n19756), .ZN(n19741) );
  OAI211_X1 U22748 ( .C1(n20066), .C2(n19780), .A(n19742), .B(n19741), .ZN(
        P2_U3073) );
  AOI22_X1 U22749 ( .A1(n19755), .A2(n20112), .B1(n19754), .B2(n20110), .ZN(
        n19744) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19757), .B1(
        n20111), .B2(n19756), .ZN(n19743) );
  OAI211_X1 U22751 ( .C1(n20115), .C2(n19780), .A(n19744), .B(n19743), .ZN(
        P2_U3074) );
  AOI22_X1 U22752 ( .A1(n19884), .A2(n19760), .B1(n19754), .B2(n20116), .ZN(
        n19746) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19757), .B1(
        n20117), .B2(n19756), .ZN(n19745) );
  OAI211_X1 U22754 ( .C1(n20073), .C2(n19753), .A(n19746), .B(n19745), .ZN(
        P2_U3075) );
  INV_X1 U22755 ( .A(n20034), .ZN(n20124) );
  AOI22_X1 U22756 ( .A1(n19760), .A2(n20124), .B1(n19754), .B2(n20122), .ZN(
        n19748) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19757), .B1(
        n20123), .B2(n19756), .ZN(n19747) );
  OAI211_X1 U22758 ( .C1(n20127), .C2(n19753), .A(n19748), .B(n19747), .ZN(
        P2_U3076) );
  AOI22_X1 U22759 ( .A1(n19760), .A2(n20079), .B1(n19754), .B2(n20128), .ZN(
        n19750) );
  AOI22_X1 U22760 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19757), .B1(
        n20129), .B2(n19756), .ZN(n19749) );
  OAI211_X1 U22761 ( .C1(n20082), .C2(n19753), .A(n19750), .B(n19749), .ZN(
        P2_U3077) );
  AOI22_X1 U22762 ( .A1(n20138), .A2(n19760), .B1(n20136), .B2(n19754), .ZN(
        n19752) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19757), .B1(
        n20137), .B2(n19756), .ZN(n19751) );
  OAI211_X1 U22764 ( .C1(n20141), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P2_U3078) );
  AOI22_X1 U22765 ( .A1(n19755), .A2(n20039), .B1(n19754), .B2(n20143), .ZN(
        n19759) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19757), .B1(
        n20144), .B2(n19756), .ZN(n19758) );
  OAI211_X1 U22767 ( .C1(n20044), .C2(n19780), .A(n19759), .B(n19758), .ZN(
        P2_U3079) );
  INV_X1 U22768 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U22769 ( .A1(n19776), .A2(n20105), .B1(n20104), .B2(n19775), .ZN(
        n19762) );
  AOI22_X1 U22770 ( .A1(n19760), .A2(n20023), .B1(n19800), .B2(n20106), .ZN(
        n19761) );
  OAI211_X1 U22771 ( .C1(n19764), .C2(n19763), .A(n19762), .B(n19761), .ZN(
        P2_U3081) );
  AOI22_X1 U22772 ( .A1(n19776), .A2(n20111), .B1(n20110), .B2(n19775), .ZN(
        n19766) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n20067), .ZN(n19765) );
  OAI211_X1 U22774 ( .C1(n20070), .C2(n19780), .A(n19766), .B(n19765), .ZN(
        P2_U3082) );
  AOI22_X1 U22775 ( .A1(n19776), .A2(n20117), .B1(n20116), .B2(n19775), .ZN(
        n19768) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n19884), .ZN(n19767) );
  OAI211_X1 U22777 ( .C1(n20073), .C2(n19780), .A(n19768), .B(n19767), .ZN(
        P2_U3083) );
  AOI22_X1 U22778 ( .A1(n19776), .A2(n20123), .B1(n20122), .B2(n19775), .ZN(
        n19770) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n20124), .ZN(n19769) );
  OAI211_X1 U22780 ( .C1(n20127), .C2(n19780), .A(n19770), .B(n19769), .ZN(
        P2_U3084) );
  AOI22_X1 U22781 ( .A1(n19776), .A2(n20129), .B1(n20128), .B2(n19775), .ZN(
        n19772) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n20079), .ZN(n19771) );
  OAI211_X1 U22783 ( .C1(n20082), .C2(n19780), .A(n19772), .B(n19771), .ZN(
        P2_U3085) );
  AOI22_X1 U22784 ( .A1(n19776), .A2(n20137), .B1(n20136), .B2(n19775), .ZN(
        n19774) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n20138), .ZN(n19773) );
  OAI211_X1 U22786 ( .C1(n20141), .C2(n19780), .A(n19774), .B(n19773), .ZN(
        P2_U3086) );
  AOI22_X1 U22787 ( .A1(n19776), .A2(n20144), .B1(n20143), .B2(n19775), .ZN(
        n19779) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19777), .B1(
        n19800), .B2(n20146), .ZN(n19778) );
  OAI211_X1 U22789 ( .C1(n20152), .C2(n19780), .A(n19779), .B(n19778), .ZN(
        P2_U3087) );
  AOI22_X1 U22790 ( .A1(n19800), .A2(n20100), .B1(n20092), .B2(n9772), .ZN(
        n19791) );
  OAI21_X1 U22791 ( .B1(n20242), .B2(n19781), .A(n20243), .ZN(n19789) );
  OAI21_X1 U22792 ( .B1(n14236), .B2(n19955), .A(n20153), .ZN(n19784) );
  INV_X1 U22793 ( .A(n19805), .ZN(n19783) );
  AOI21_X1 U22794 ( .B1(n19784), .B2(n19783), .A(n19782), .ZN(n19785) );
  OAI21_X1 U22795 ( .B1(n19789), .B2(n19786), .A(n19785), .ZN(n19807) );
  OAI21_X1 U22796 ( .B1(n14236), .B2(n9772), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19787) );
  OAI21_X1 U22797 ( .B1(n19789), .B2(n19788), .A(n19787), .ZN(n19806) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19807), .B1(
        n16038), .B2(n19806), .ZN(n19790) );
  OAI211_X1 U22799 ( .C1(n20103), .C2(n19829), .A(n19791), .B(n19790), .ZN(
        P2_U3088) );
  AOI22_X1 U22800 ( .A1(n19817), .A2(n20106), .B1(n20104), .B2(n9772), .ZN(
        n19793) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19807), .B1(
        n20105), .B2(n19806), .ZN(n19792) );
  OAI211_X1 U22802 ( .C1(n20109), .C2(n19810), .A(n19793), .B(n19792), .ZN(
        P2_U3089) );
  AOI22_X1 U22803 ( .A1(n19817), .A2(n20067), .B1(n20110), .B2(n9772), .ZN(
        n19795) );
  AOI22_X1 U22804 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19807), .B1(
        n20111), .B2(n19806), .ZN(n19794) );
  OAI211_X1 U22805 ( .C1(n20070), .C2(n19810), .A(n19795), .B(n19794), .ZN(
        P2_U3090) );
  AOI22_X1 U22806 ( .A1(n19884), .A2(n19817), .B1(n9772), .B2(n20116), .ZN(
        n19797) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19807), .B1(
        n20117), .B2(n19806), .ZN(n19796) );
  OAI211_X1 U22808 ( .C1(n20073), .C2(n19810), .A(n19797), .B(n19796), .ZN(
        P2_U3091) );
  AOI22_X1 U22809 ( .A1(n19800), .A2(n20031), .B1(n9772), .B2(n20122), .ZN(
        n19799) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19807), .B1(
        n20123), .B2(n19806), .ZN(n19798) );
  OAI211_X1 U22811 ( .C1(n20034), .C2(n19829), .A(n19799), .B(n19798), .ZN(
        P2_U3092) );
  AOI22_X1 U22812 ( .A1(n19800), .A2(n20130), .B1(n9772), .B2(n20128), .ZN(
        n19802) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19807), .B1(
        n20129), .B2(n19806), .ZN(n19801) );
  OAI211_X1 U22814 ( .C1(n20135), .C2(n19829), .A(n19802), .B(n19801), .ZN(
        P2_U3093) );
  AOI22_X1 U22815 ( .A1(n20138), .A2(n19817), .B1(n20136), .B2(n9772), .ZN(
        n19804) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19807), .B1(
        n20137), .B2(n19806), .ZN(n19803) );
  OAI211_X1 U22817 ( .C1(n20141), .C2(n19810), .A(n19804), .B(n19803), .ZN(
        P2_U3094) );
  AOI22_X1 U22818 ( .A1(n19817), .A2(n20146), .B1(n20143), .B2(n9772), .ZN(
        n19809) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19807), .B1(
        n20144), .B2(n19806), .ZN(n19808) );
  OAI211_X1 U22820 ( .C1(n20152), .C2(n19810), .A(n19809), .B(n19808), .ZN(
        P2_U3095) );
  AOI22_X1 U22821 ( .A1(n19825), .A2(n20105), .B1(n19824), .B2(n20104), .ZN(
        n19812) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19826), .B1(
        n19817), .B2(n20023), .ZN(n19811) );
  OAI211_X1 U22823 ( .C1(n20066), .C2(n19880), .A(n19812), .B(n19811), .ZN(
        P2_U3097) );
  AOI22_X1 U22824 ( .A1(n19825), .A2(n20111), .B1(n19824), .B2(n20110), .ZN(
        n19814) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19826), .B1(
        n19868), .B2(n20067), .ZN(n19813) );
  OAI211_X1 U22826 ( .C1(n20070), .C2(n19829), .A(n19814), .B(n19813), .ZN(
        P2_U3098) );
  AOI22_X1 U22827 ( .A1(n19825), .A2(n20117), .B1(n19824), .B2(n20116), .ZN(
        n19816) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19826), .B1(
        n19817), .B2(n20118), .ZN(n19815) );
  OAI211_X1 U22829 ( .C1(n20121), .C2(n19880), .A(n19816), .B(n19815), .ZN(
        P2_U3099) );
  AOI22_X1 U22830 ( .A1(n19825), .A2(n20123), .B1(n19824), .B2(n20122), .ZN(
        n19819) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19826), .B1(
        n19817), .B2(n20031), .ZN(n19818) );
  OAI211_X1 U22832 ( .C1(n20034), .C2(n19880), .A(n19819), .B(n19818), .ZN(
        P2_U3100) );
  AOI22_X1 U22833 ( .A1(n19825), .A2(n20129), .B1(n19824), .B2(n20128), .ZN(
        n19821) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19826), .B1(
        n19868), .B2(n20079), .ZN(n19820) );
  OAI211_X1 U22835 ( .C1(n20082), .C2(n19829), .A(n19821), .B(n19820), .ZN(
        P2_U3101) );
  AOI22_X1 U22836 ( .A1(n19825), .A2(n20137), .B1(n19824), .B2(n20136), .ZN(
        n19823) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19826), .B1(
        n19868), .B2(n20138), .ZN(n19822) );
  OAI211_X1 U22838 ( .C1(n20141), .C2(n19829), .A(n19823), .B(n19822), .ZN(
        P2_U3102) );
  AOI22_X1 U22839 ( .A1(n19825), .A2(n20144), .B1(n19824), .B2(n20143), .ZN(
        n19828) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19826), .B1(
        n19868), .B2(n20146), .ZN(n19827) );
  OAI211_X1 U22841 ( .C1(n20152), .C2(n19829), .A(n19828), .B(n19827), .ZN(
        P2_U3103) );
  NOR2_X1 U22842 ( .A1(n19839), .A2(n19955), .ZN(n19830) );
  NAND2_X1 U22843 ( .A1(n14237), .A2(n19830), .ZN(n19836) );
  OAI21_X1 U22844 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19835), .A(n19955), 
        .ZN(n19831) );
  NAND2_X1 U22845 ( .A1(n19836), .A2(n19831), .ZN(n19875) );
  INV_X1 U22846 ( .A(n16038), .ZN(n19833) );
  OAI22_X1 U22847 ( .A1(n19875), .A2(n19833), .B1(n19873), .B2(n19832), .ZN(
        n19834) );
  INV_X1 U22848 ( .A(n19834), .ZN(n19841) );
  OAI21_X1 U22849 ( .B1(n20242), .B2(n20241), .A(n19835), .ZN(n19837) );
  AND3_X1 U22850 ( .A1(n19837), .A2(n20098), .A3(n19836), .ZN(n19838) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19877), .B1(
        n19868), .B2(n20100), .ZN(n19840) );
  OAI211_X1 U22852 ( .C1(n20103), .C2(n19871), .A(n19841), .B(n19840), .ZN(
        P2_U3104) );
  INV_X1 U22853 ( .A(n20105), .ZN(n19842) );
  OAI22_X1 U22854 ( .A1(n19875), .A2(n19842), .B1(n19873), .B2(n20062), .ZN(
        n19843) );
  INV_X1 U22855 ( .A(n19843), .ZN(n19845) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19877), .B1(
        n19868), .B2(n20023), .ZN(n19844) );
  OAI211_X1 U22857 ( .C1(n20066), .C2(n19871), .A(n19845), .B(n19844), .ZN(
        P2_U3105) );
  INV_X1 U22858 ( .A(n20111), .ZN(n19847) );
  INV_X1 U22859 ( .A(n20110), .ZN(n19846) );
  OAI22_X1 U22860 ( .A1(n19875), .A2(n19847), .B1(n19873), .B2(n19846), .ZN(
        n19848) );
  INV_X1 U22861 ( .A(n19848), .ZN(n19850) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19877), .B1(
        n19868), .B2(n20112), .ZN(n19849) );
  OAI211_X1 U22863 ( .C1(n20115), .C2(n19871), .A(n19850), .B(n19849), .ZN(
        P2_U3106) );
  INV_X1 U22864 ( .A(n20117), .ZN(n19851) );
  OAI22_X1 U22865 ( .A1(n19875), .A2(n19851), .B1(n19873), .B2(n20072), .ZN(
        n19852) );
  INV_X1 U22866 ( .A(n19852), .ZN(n19854) );
  AOI22_X1 U22867 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19877), .B1(
        n19868), .B2(n20118), .ZN(n19853) );
  OAI211_X1 U22868 ( .C1(n20121), .C2(n19871), .A(n19854), .B(n19853), .ZN(
        P2_U3107) );
  INV_X1 U22869 ( .A(n20123), .ZN(n19856) );
  INV_X1 U22870 ( .A(n20122), .ZN(n19855) );
  OAI22_X1 U22871 ( .A1(n19875), .A2(n19856), .B1(n19873), .B2(n19855), .ZN(
        n19857) );
  INV_X1 U22872 ( .A(n19857), .ZN(n19859) );
  AOI22_X1 U22873 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19877), .B1(
        n19896), .B2(n20124), .ZN(n19858) );
  OAI211_X1 U22874 ( .C1(n20127), .C2(n19880), .A(n19859), .B(n19858), .ZN(
        P2_U3108) );
  INV_X1 U22875 ( .A(n20129), .ZN(n19861) );
  INV_X1 U22876 ( .A(n20128), .ZN(n19860) );
  OAI22_X1 U22877 ( .A1(n19875), .A2(n19861), .B1(n19873), .B2(n19860), .ZN(
        n19862) );
  INV_X1 U22878 ( .A(n19862), .ZN(n19864) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19877), .B1(
        n19896), .B2(n20079), .ZN(n19863) );
  OAI211_X1 U22880 ( .C1(n20082), .C2(n19880), .A(n19864), .B(n19863), .ZN(
        P2_U3109) );
  INV_X1 U22881 ( .A(n20137), .ZN(n19866) );
  INV_X1 U22882 ( .A(n20136), .ZN(n19865) );
  OAI22_X1 U22883 ( .A1(n19875), .A2(n19866), .B1(n19873), .B2(n19865), .ZN(
        n19867) );
  INV_X1 U22884 ( .A(n19867), .ZN(n19870) );
  AOI22_X1 U22885 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19877), .B1(
        n19868), .B2(n20009), .ZN(n19869) );
  OAI211_X1 U22886 ( .C1(n20012), .C2(n19871), .A(n19870), .B(n19869), .ZN(
        P2_U3110) );
  INV_X1 U22887 ( .A(n20144), .ZN(n19874) );
  INV_X1 U22888 ( .A(n20143), .ZN(n19872) );
  OAI22_X1 U22889 ( .A1(n19875), .A2(n19874), .B1(n19873), .B2(n19872), .ZN(
        n19876) );
  INV_X1 U22890 ( .A(n19876), .ZN(n19879) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19877), .B1(
        n19896), .B2(n20146), .ZN(n19878) );
  OAI211_X1 U22892 ( .C1(n20152), .C2(n19880), .A(n19879), .B(n19878), .ZN(
        P2_U3111) );
  INV_X1 U22893 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U22894 ( .A1(n19914), .A2(n20067), .B1(n19895), .B2(n20110), .ZN(
        n19882) );
  AOI22_X1 U22895 ( .A1(n20111), .A2(n19897), .B1(n19896), .B2(n20112), .ZN(
        n19881) );
  OAI211_X1 U22896 ( .C1(n19901), .C2(n19883), .A(n19882), .B(n19881), .ZN(
        P2_U3114) );
  AOI22_X1 U22897 ( .A1(n19914), .A2(n19884), .B1(n19895), .B2(n20116), .ZN(
        n19886) );
  AOI22_X1 U22898 ( .A1(n20117), .A2(n19897), .B1(n19896), .B2(n20118), .ZN(
        n19885) );
  OAI211_X1 U22899 ( .C1(n19901), .C2(n12287), .A(n19886), .B(n19885), .ZN(
        P2_U3115) );
  INV_X1 U22900 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U22901 ( .A1(n19914), .A2(n20124), .B1(n19895), .B2(n20122), .ZN(
        n19888) );
  AOI22_X1 U22902 ( .A1(n20123), .A2(n19897), .B1(n19896), .B2(n20031), .ZN(
        n19887) );
  OAI211_X1 U22903 ( .C1(n19901), .C2(n19889), .A(n19888), .B(n19887), .ZN(
        P2_U3116) );
  AOI22_X1 U22904 ( .A1(n19914), .A2(n20079), .B1(n19895), .B2(n20128), .ZN(
        n19891) );
  AOI22_X1 U22905 ( .A1(n20129), .A2(n19897), .B1(n19896), .B2(n20130), .ZN(
        n19890) );
  OAI211_X1 U22906 ( .C1(n19901), .C2(n12338), .A(n19891), .B(n19890), .ZN(
        P2_U3117) );
  INV_X1 U22907 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U22908 ( .A1(n19914), .A2(n20138), .B1(n20136), .B2(n19895), .ZN(
        n19893) );
  AOI22_X1 U22909 ( .A1(n20137), .A2(n19897), .B1(n19896), .B2(n20009), .ZN(
        n19892) );
  OAI211_X1 U22910 ( .C1(n19901), .C2(n19894), .A(n19893), .B(n19892), .ZN(
        P2_U3118) );
  INV_X1 U22911 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U22912 ( .A1(n19914), .A2(n20146), .B1(n19895), .B2(n20143), .ZN(
        n19899) );
  AOI22_X1 U22913 ( .A1(n20144), .A2(n19897), .B1(n19896), .B2(n20039), .ZN(
        n19898) );
  OAI211_X1 U22914 ( .C1(n19901), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        P2_U3119) );
  AOI22_X1 U22915 ( .A1(n19942), .A2(n20019), .B1(n20092), .B2(n19920), .ZN(
        n19903) );
  AOI22_X1 U22916 ( .A1(n16038), .A2(n19921), .B1(n19914), .B2(n20100), .ZN(
        n19902) );
  OAI211_X1 U22917 ( .C1(n19907), .C2(n12205), .A(n19903), .B(n19902), .ZN(
        P2_U3120) );
  INV_X1 U22918 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U22919 ( .A1(n19942), .A2(n20067), .B1(n19920), .B2(n20110), .ZN(
        n19905) );
  AOI22_X1 U22920 ( .A1(n20111), .A2(n19921), .B1(n19914), .B2(n20112), .ZN(
        n19904) );
  OAI211_X1 U22921 ( .C1(n19907), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P2_U3122) );
  INV_X1 U22922 ( .A(n19942), .ZN(n19917) );
  OAI22_X1 U22923 ( .A1(n19925), .A2(n20073), .B1(n19908), .B2(n20072), .ZN(
        n19909) );
  INV_X1 U22924 ( .A(n19909), .ZN(n19911) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19922), .B1(
        n20117), .B2(n19921), .ZN(n19910) );
  OAI211_X1 U22926 ( .C1(n20121), .C2(n19917), .A(n19911), .B(n19910), .ZN(
        P2_U3123) );
  AOI22_X1 U22927 ( .A1(n19914), .A2(n20031), .B1(n19920), .B2(n20122), .ZN(
        n19913) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19922), .B1(
        n20123), .B2(n19921), .ZN(n19912) );
  OAI211_X1 U22929 ( .C1(n20034), .C2(n19917), .A(n19913), .B(n19912), .ZN(
        P2_U3124) );
  AOI22_X1 U22930 ( .A1(n19914), .A2(n20130), .B1(n19920), .B2(n20128), .ZN(
        n19916) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19922), .B1(
        n20129), .B2(n19921), .ZN(n19915) );
  OAI211_X1 U22932 ( .C1(n20135), .C2(n19917), .A(n19916), .B(n19915), .ZN(
        P2_U3125) );
  AOI22_X1 U22933 ( .A1(n19942), .A2(n20138), .B1(n20136), .B2(n19920), .ZN(
        n19919) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19922), .B1(
        n20137), .B2(n19921), .ZN(n19918) );
  OAI211_X1 U22935 ( .C1(n20141), .C2(n19925), .A(n19919), .B(n19918), .ZN(
        P2_U3126) );
  AOI22_X1 U22936 ( .A1(n19942), .A2(n20146), .B1(n19920), .B2(n20143), .ZN(
        n19924) );
  AOI22_X1 U22937 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19922), .B1(
        n20144), .B2(n19921), .ZN(n19923) );
  OAI211_X1 U22938 ( .C1(n20152), .C2(n19925), .A(n19924), .B(n19923), .ZN(
        P2_U3127) );
  AOI22_X1 U22939 ( .A1(n19941), .A2(n20105), .B1(n19940), .B2(n20104), .ZN(
        n19927) );
  AOI22_X1 U22940 ( .A1(n19942), .A2(n20023), .B1(n19975), .B2(n20106), .ZN(
        n19926) );
  OAI211_X1 U22941 ( .C1(n19931), .C2(n19928), .A(n19927), .B(n19926), .ZN(
        P2_U3129) );
  AOI22_X1 U22942 ( .A1(n19941), .A2(n20111), .B1(n19940), .B2(n20110), .ZN(
        n19930) );
  AOI22_X1 U22943 ( .A1(n19942), .A2(n20112), .B1(n19975), .B2(n20067), .ZN(
        n19929) );
  OAI211_X1 U22944 ( .C1(n19931), .C2(n12252), .A(n19930), .B(n19929), .ZN(
        P2_U3130) );
  AOI22_X1 U22945 ( .A1(n19941), .A2(n20117), .B1(n19940), .B2(n20116), .ZN(
        n19933) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n20118), .ZN(n19932) );
  OAI211_X1 U22947 ( .C1(n20121), .C2(n19983), .A(n19933), .B(n19932), .ZN(
        P2_U3131) );
  AOI22_X1 U22948 ( .A1(n19941), .A2(n20123), .B1(n19940), .B2(n20122), .ZN(
        n19935) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n20031), .ZN(n19934) );
  OAI211_X1 U22950 ( .C1(n20034), .C2(n19983), .A(n19935), .B(n19934), .ZN(
        P2_U3132) );
  AOI22_X1 U22951 ( .A1(n19941), .A2(n20129), .B1(n19940), .B2(n20128), .ZN(
        n19937) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n20130), .ZN(n19936) );
  OAI211_X1 U22953 ( .C1(n20135), .C2(n19983), .A(n19937), .B(n19936), .ZN(
        P2_U3133) );
  AOI22_X1 U22954 ( .A1(n19941), .A2(n20137), .B1(n19940), .B2(n20136), .ZN(
        n19939) );
  AOI22_X1 U22955 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n20009), .ZN(n19938) );
  OAI211_X1 U22956 ( .C1(n20012), .C2(n19983), .A(n19939), .B(n19938), .ZN(
        P2_U3134) );
  AOI22_X1 U22957 ( .A1(n19941), .A2(n20144), .B1(n19940), .B2(n20143), .ZN(
        n19945) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19943), .B1(
        n19942), .B2(n20039), .ZN(n19944) );
  OAI211_X1 U22959 ( .C1(n20044), .C2(n19983), .A(n19945), .B(n19944), .ZN(
        P2_U3135) );
  NOR2_X1 U22960 ( .A1(n20272), .A2(n19947), .ZN(n19962) );
  INV_X1 U22961 ( .A(n19962), .ZN(n19948) );
  OR2_X1 U22962 ( .A1(n19948), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19954) );
  INV_X1 U22963 ( .A(n19949), .ZN(n19951) );
  NAND2_X1 U22964 ( .A1(n19951), .A2(n19950), .ZN(n19956) );
  NAND2_X1 U22965 ( .A1(n19956), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19952) );
  NOR2_X1 U22966 ( .A1(n19953), .A2(n19952), .ZN(n19958) );
  AOI21_X1 U22967 ( .B1(n19955), .B2(n19954), .A(n19958), .ZN(n19979) );
  INV_X1 U22968 ( .A(n19956), .ZN(n19978) );
  AOI22_X1 U22969 ( .A1(n19979), .A2(n16038), .B1(n20092), .B2(n19978), .ZN(
        n19964) );
  INV_X1 U22970 ( .A(n20094), .ZN(n19960) );
  OAI21_X1 U22971 ( .B1(n19978), .B2(n20153), .A(n20098), .ZN(n19957) );
  NOR2_X1 U22972 ( .A1(n19958), .A2(n19957), .ZN(n19959) );
  OAI221_X1 U22973 ( .B1(n19962), .B2(n19961), .C1(n19962), .C2(n19960), .A(
        n19959), .ZN(n19980) );
  AOI22_X1 U22974 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19980), .B1(
        n19975), .B2(n20100), .ZN(n19963) );
  OAI211_X1 U22975 ( .C1(n20103), .C2(n19990), .A(n19964), .B(n19963), .ZN(
        P2_U3136) );
  AOI22_X1 U22976 ( .A1(n19979), .A2(n20105), .B1(n20104), .B2(n19978), .ZN(
        n19966) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19980), .B1(
        n19975), .B2(n20023), .ZN(n19965) );
  OAI211_X1 U22978 ( .C1(n20066), .C2(n19990), .A(n19966), .B(n19965), .ZN(
        P2_U3137) );
  AOI22_X1 U22979 ( .A1(n19979), .A2(n20111), .B1(n20110), .B2(n19978), .ZN(
        n19968) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19980), .B1(
        n19975), .B2(n20112), .ZN(n19967) );
  OAI211_X1 U22981 ( .C1(n20115), .C2(n19990), .A(n19968), .B(n19967), .ZN(
        P2_U3138) );
  AOI22_X1 U22982 ( .A1(n19979), .A2(n20117), .B1(n20116), .B2(n19978), .ZN(
        n19970) );
  AOI22_X1 U22983 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19980), .B1(
        n19975), .B2(n20118), .ZN(n19969) );
  OAI211_X1 U22984 ( .C1(n20121), .C2(n19990), .A(n19970), .B(n19969), .ZN(
        P2_U3139) );
  AOI22_X1 U22985 ( .A1(n19979), .A2(n20123), .B1(n20122), .B2(n19978), .ZN(
        n19972) );
  AOI22_X1 U22986 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19980), .B1(
        n20015), .B2(n20124), .ZN(n19971) );
  OAI211_X1 U22987 ( .C1(n20127), .C2(n19983), .A(n19972), .B(n19971), .ZN(
        P2_U3140) );
  AOI22_X1 U22988 ( .A1(n19979), .A2(n20129), .B1(n20128), .B2(n19978), .ZN(
        n19974) );
  AOI22_X1 U22989 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19980), .B1(
        n20015), .B2(n20079), .ZN(n19973) );
  OAI211_X1 U22990 ( .C1(n20082), .C2(n19983), .A(n19974), .B(n19973), .ZN(
        P2_U3141) );
  AOI22_X1 U22991 ( .A1(n19979), .A2(n20137), .B1(n20136), .B2(n19978), .ZN(
        n19977) );
  AOI22_X1 U22992 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19980), .B1(
        n19975), .B2(n20009), .ZN(n19976) );
  OAI211_X1 U22993 ( .C1(n20012), .C2(n19990), .A(n19977), .B(n19976), .ZN(
        P2_U3142) );
  AOI22_X1 U22994 ( .A1(n19979), .A2(n20144), .B1(n20143), .B2(n19978), .ZN(
        n19982) );
  AOI22_X1 U22995 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19980), .B1(
        n20015), .B2(n20146), .ZN(n19981) );
  OAI211_X1 U22996 ( .C1(n20152), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        P2_U3143) );
  NOR2_X1 U22997 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19984), .ZN(
        n20013) );
  OAI21_X1 U22998 ( .B1(n14287), .B2(n20013), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19989) );
  NAND3_X1 U22999 ( .A1(n19987), .A2(n19986), .A3(n19985), .ZN(n19988) );
  NAND2_X1 U23000 ( .A1(n19989), .A2(n19988), .ZN(n20014) );
  AOI22_X1 U23001 ( .A1(n20014), .A2(n16038), .B1(n20092), .B2(n20013), .ZN(
        n19998) );
  AOI21_X1 U23002 ( .B1(n19990), .B2(n20037), .A(n20049), .ZN(n19996) );
  INV_X1 U23003 ( .A(n14287), .ZN(n19992) );
  INV_X1 U23004 ( .A(n20013), .ZN(n19991) );
  OAI211_X1 U23005 ( .C1(n19992), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19991), 
        .B(n20245), .ZN(n19993) );
  AND2_X1 U23006 ( .A1(n19993), .A2(n20098), .ZN(n19994) );
  OAI211_X1 U23007 ( .C1(n19996), .C2(n19995), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19994), .ZN(n20016) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20100), .ZN(n19997) );
  OAI211_X1 U23009 ( .C1(n20103), .C2(n20037), .A(n19998), .B(n19997), .ZN(
        P2_U3144) );
  AOI22_X1 U23010 ( .A1(n20014), .A2(n20105), .B1(n20104), .B2(n20013), .ZN(
        n20000) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20023), .ZN(n19999) );
  OAI211_X1 U23012 ( .C1(n20066), .C2(n20037), .A(n20000), .B(n19999), .ZN(
        P2_U3145) );
  AOI22_X1 U23013 ( .A1(n20014), .A2(n20111), .B1(n20110), .B2(n20013), .ZN(
        n20002) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20112), .ZN(n20001) );
  OAI211_X1 U23015 ( .C1(n20115), .C2(n20037), .A(n20002), .B(n20001), .ZN(
        P2_U3146) );
  AOI22_X1 U23016 ( .A1(n20014), .A2(n20117), .B1(n20116), .B2(n20013), .ZN(
        n20004) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20118), .ZN(n20003) );
  OAI211_X1 U23018 ( .C1(n20121), .C2(n20037), .A(n20004), .B(n20003), .ZN(
        P2_U3147) );
  AOI22_X1 U23019 ( .A1(n20014), .A2(n20123), .B1(n20122), .B2(n20013), .ZN(
        n20006) );
  AOI22_X1 U23020 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20031), .ZN(n20005) );
  OAI211_X1 U23021 ( .C1(n20034), .C2(n20037), .A(n20006), .B(n20005), .ZN(
        P2_U3148) );
  AOI22_X1 U23022 ( .A1(n20014), .A2(n20129), .B1(n20128), .B2(n20013), .ZN(
        n20008) );
  AOI22_X1 U23023 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20130), .ZN(n20007) );
  OAI211_X1 U23024 ( .C1(n20135), .C2(n20037), .A(n20008), .B(n20007), .ZN(
        P2_U3149) );
  AOI22_X1 U23025 ( .A1(n20014), .A2(n20137), .B1(n20136), .B2(n20013), .ZN(
        n20011) );
  AOI22_X1 U23026 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20009), .ZN(n20010) );
  OAI211_X1 U23027 ( .C1(n20012), .C2(n20037), .A(n20011), .B(n20010), .ZN(
        P2_U3150) );
  AOI22_X1 U23028 ( .A1(n20014), .A2(n20144), .B1(n20143), .B2(n20013), .ZN(
        n20018) );
  AOI22_X1 U23029 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20016), .B1(
        n20015), .B2(n20039), .ZN(n20017) );
  OAI211_X1 U23030 ( .C1(n20044), .C2(n20037), .A(n20018), .B(n20017), .ZN(
        P2_U3151) );
  AOI22_X1 U23031 ( .A1(n20038), .A2(n16038), .B1(n20092), .B2(n20051), .ZN(
        n20021) );
  AOI22_X1 U23032 ( .A1(n20040), .A2(n20100), .B1(n20048), .B2(n20019), .ZN(
        n20020) );
  OAI211_X1 U23033 ( .C1(n20026), .C2(n20022), .A(n20021), .B(n20020), .ZN(
        P2_U3152) );
  AOI22_X1 U23034 ( .A1(n20038), .A2(n20105), .B1(n20051), .B2(n20104), .ZN(
        n20025) );
  AOI22_X1 U23035 ( .A1(n20040), .A2(n20023), .B1(n20048), .B2(n20106), .ZN(
        n20024) );
  OAI211_X1 U23036 ( .C1(n20026), .C2(n13740), .A(n20025), .B(n20024), .ZN(
        P2_U3153) );
  AOI22_X1 U23037 ( .A1(n20038), .A2(n20111), .B1(n20051), .B2(n20110), .ZN(
        n20028) );
  AOI22_X1 U23038 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20041), .B1(
        n20040), .B2(n20112), .ZN(n20027) );
  OAI211_X1 U23039 ( .C1(n20115), .C2(n20090), .A(n20028), .B(n20027), .ZN(
        P2_U3154) );
  AOI22_X1 U23040 ( .A1(n20038), .A2(n20117), .B1(n20051), .B2(n20116), .ZN(
        n20030) );
  AOI22_X1 U23041 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20041), .B1(
        n20040), .B2(n20118), .ZN(n20029) );
  OAI211_X1 U23042 ( .C1(n20121), .C2(n20090), .A(n20030), .B(n20029), .ZN(
        P2_U3155) );
  AOI22_X1 U23043 ( .A1(n20038), .A2(n20123), .B1(n20051), .B2(n20122), .ZN(
        n20033) );
  AOI22_X1 U23044 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20041), .B1(
        n20040), .B2(n20031), .ZN(n20032) );
  OAI211_X1 U23045 ( .C1(n20034), .C2(n20090), .A(n20033), .B(n20032), .ZN(
        P2_U3156) );
  AOI22_X1 U23046 ( .A1(n20038), .A2(n20129), .B1(n20051), .B2(n20128), .ZN(
        n20036) );
  AOI22_X1 U23047 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20041), .B1(
        n20048), .B2(n20079), .ZN(n20035) );
  OAI211_X1 U23048 ( .C1(n20082), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        P2_U3157) );
  AOI22_X1 U23049 ( .A1(n20038), .A2(n20144), .B1(n20051), .B2(n20143), .ZN(
        n20043) );
  AOI22_X1 U23050 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20041), .B1(
        n20040), .B2(n20039), .ZN(n20042) );
  OAI211_X1 U23051 ( .C1(n20044), .C2(n20090), .A(n20043), .B(n20042), .ZN(
        P2_U3159) );
  NAND2_X1 U23052 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20047), .ZN(
        n20093) );
  NOR2_X1 U23053 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20093), .ZN(
        n20085) );
  AOI22_X1 U23054 ( .A1(n20048), .A2(n20100), .B1(n20092), .B2(n20085), .ZN(
        n20061) );
  AOI21_X1 U23055 ( .B1(n20055), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20053) );
  AOI21_X1 U23056 ( .B1(n20151), .B2(n20090), .A(n20049), .ZN(n20050) );
  NOR2_X1 U23057 ( .A1(n20050), .A2(n20245), .ZN(n20054) );
  NOR2_X1 U23058 ( .A1(n20085), .A2(n20051), .ZN(n20058) );
  NAND2_X1 U23059 ( .A1(n20054), .A2(n20058), .ZN(n20052) );
  OAI211_X1 U23060 ( .C1(n20085), .C2(n20053), .A(n20052), .B(n20098), .ZN(
        n20087) );
  INV_X1 U23061 ( .A(n20054), .ZN(n20059) );
  INV_X1 U23062 ( .A(n20055), .ZN(n20056) );
  OAI21_X1 U23063 ( .B1(n20056), .B2(n20085), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20057) );
  AOI22_X1 U23064 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20087), .B1(
        n16038), .B2(n20086), .ZN(n20060) );
  OAI211_X1 U23065 ( .C1(n20103), .C2(n20151), .A(n20061), .B(n20060), .ZN(
        P2_U3160) );
  INV_X1 U23066 ( .A(n20085), .ZN(n20071) );
  OAI22_X1 U23067 ( .A1(n20090), .A2(n20109), .B1(n20062), .B2(n20071), .ZN(
        n20063) );
  INV_X1 U23068 ( .A(n20063), .ZN(n20065) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20087), .B1(
        n20105), .B2(n20086), .ZN(n20064) );
  OAI211_X1 U23070 ( .C1(n20066), .C2(n20151), .A(n20065), .B(n20064), .ZN(
        P2_U3161) );
  AOI22_X1 U23071 ( .A1(n20131), .A2(n20067), .B1(n20110), .B2(n20085), .ZN(
        n20069) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20087), .B1(
        n20111), .B2(n20086), .ZN(n20068) );
  OAI211_X1 U23073 ( .C1(n20070), .C2(n20090), .A(n20069), .B(n20068), .ZN(
        P2_U3162) );
  OAI22_X1 U23074 ( .A1(n20090), .A2(n20073), .B1(n20072), .B2(n20071), .ZN(
        n20074) );
  INV_X1 U23075 ( .A(n20074), .ZN(n20076) );
  AOI22_X1 U23076 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20087), .B1(
        n20117), .B2(n20086), .ZN(n20075) );
  OAI211_X1 U23077 ( .C1(n20121), .C2(n20151), .A(n20076), .B(n20075), .ZN(
        P2_U3163) );
  AOI22_X1 U23078 ( .A1(n20131), .A2(n20124), .B1(n20122), .B2(n20085), .ZN(
        n20078) );
  AOI22_X1 U23079 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20087), .B1(
        n20123), .B2(n20086), .ZN(n20077) );
  OAI211_X1 U23080 ( .C1(n20127), .C2(n20090), .A(n20078), .B(n20077), .ZN(
        P2_U3164) );
  AOI22_X1 U23081 ( .A1(n20131), .A2(n20079), .B1(n20128), .B2(n20085), .ZN(
        n20081) );
  AOI22_X1 U23082 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20087), .B1(
        n20129), .B2(n20086), .ZN(n20080) );
  OAI211_X1 U23083 ( .C1(n20082), .C2(n20090), .A(n20081), .B(n20080), .ZN(
        P2_U3165) );
  AOI22_X1 U23084 ( .A1(n20131), .A2(n20138), .B1(n20136), .B2(n20085), .ZN(
        n20084) );
  AOI22_X1 U23085 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20087), .B1(
        n20137), .B2(n20086), .ZN(n20083) );
  OAI211_X1 U23086 ( .C1(n20141), .C2(n20090), .A(n20084), .B(n20083), .ZN(
        P2_U3166) );
  AOI22_X1 U23087 ( .A1(n20131), .A2(n20146), .B1(n20143), .B2(n20085), .ZN(
        n20089) );
  AOI22_X1 U23088 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20087), .B1(
        n20144), .B2(n20086), .ZN(n20088) );
  OAI211_X1 U23089 ( .C1(n20152), .C2(n20090), .A(n20089), .B(n20088), .ZN(
        P2_U3167) );
  OAI21_X1 U23090 ( .B1(n14295), .B2(n20142), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20091) );
  OAI21_X1 U23091 ( .B1(n20093), .B2(n20245), .A(n20091), .ZN(n20145) );
  AOI22_X1 U23092 ( .A1(n20145), .A2(n16038), .B1(n20092), .B2(n20142), .ZN(
        n20102) );
  OAI21_X1 U23093 ( .B1(n20094), .B2(n20241), .A(n20093), .ZN(n20099) );
  INV_X1 U23094 ( .A(n20142), .ZN(n20095) );
  OAI211_X1 U23095 ( .C1(n20096), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20095), 
        .B(n20245), .ZN(n20097) );
  NAND3_X1 U23096 ( .A1(n20099), .A2(n20098), .A3(n20097), .ZN(n20148) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20148), .B1(
        n20131), .B2(n20100), .ZN(n20101) );
  OAI211_X1 U23098 ( .C1(n20103), .C2(n20134), .A(n20102), .B(n20101), .ZN(
        P2_U3168) );
  AOI22_X1 U23099 ( .A1(n20145), .A2(n20105), .B1(n20104), .B2(n20142), .ZN(
        n20108) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20106), .ZN(n20107) );
  OAI211_X1 U23101 ( .C1(n20109), .C2(n20151), .A(n20108), .B(n20107), .ZN(
        P2_U3169) );
  AOI22_X1 U23102 ( .A1(n20145), .A2(n20111), .B1(n20110), .B2(n20142), .ZN(
        n20114) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20148), .B1(
        n20131), .B2(n20112), .ZN(n20113) );
  OAI211_X1 U23104 ( .C1(n20115), .C2(n20134), .A(n20114), .B(n20113), .ZN(
        P2_U3170) );
  AOI22_X1 U23105 ( .A1(n20145), .A2(n20117), .B1(n20116), .B2(n20142), .ZN(
        n20120) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20148), .B1(
        n20131), .B2(n20118), .ZN(n20119) );
  OAI211_X1 U23107 ( .C1(n20121), .C2(n20134), .A(n20120), .B(n20119), .ZN(
        P2_U3171) );
  AOI22_X1 U23108 ( .A1(n20145), .A2(n20123), .B1(n20122), .B2(n20142), .ZN(
        n20126) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20124), .ZN(n20125) );
  OAI211_X1 U23110 ( .C1(n20127), .C2(n20151), .A(n20126), .B(n20125), .ZN(
        P2_U3172) );
  AOI22_X1 U23111 ( .A1(n20145), .A2(n20129), .B1(n20128), .B2(n20142), .ZN(
        n20133) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20148), .B1(
        n20131), .B2(n20130), .ZN(n20132) );
  OAI211_X1 U23113 ( .C1(n20135), .C2(n20134), .A(n20133), .B(n20132), .ZN(
        P2_U3173) );
  AOI22_X1 U23114 ( .A1(n20145), .A2(n20137), .B1(n20136), .B2(n20142), .ZN(
        n20140) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20138), .ZN(n20139) );
  OAI211_X1 U23116 ( .C1(n20141), .C2(n20151), .A(n20140), .B(n20139), .ZN(
        P2_U3174) );
  AOI22_X1 U23117 ( .A1(n20145), .A2(n20144), .B1(n20143), .B2(n20142), .ZN(
        n20150) );
  AOI22_X1 U23118 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20146), .ZN(n20149) );
  OAI211_X1 U23119 ( .C1(n20152), .C2(n20151), .A(n20150), .B(n20149), .ZN(
        P2_U3175) );
  OAI221_X1 U23120 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20153), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n20155), .A(n20157), .ZN(n20161) );
  AOI211_X1 U23121 ( .C1(n20157), .C2(n20156), .A(n20155), .B(n20154), .ZN(
        n20158) );
  INV_X1 U23122 ( .A(n20158), .ZN(n20160) );
  OAI211_X1 U23123 ( .C1(n20162), .C2(n20161), .A(n20160), .B(n20159), .ZN(
        P2_U3177) );
  AND2_X1 U23124 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20163), .ZN(
        P2_U3179) );
  AND2_X1 U23125 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20163), .ZN(
        P2_U3180) );
  AND2_X1 U23126 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20163), .ZN(
        P2_U3181) );
  AND2_X1 U23127 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20163), .ZN(
        P2_U3182) );
  AND2_X1 U23128 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20163), .ZN(
        P2_U3183) );
  AND2_X1 U23129 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20163), .ZN(
        P2_U3184) );
  AND2_X1 U23130 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20163), .ZN(
        P2_U3185) );
  AND2_X1 U23131 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20163), .ZN(
        P2_U3186) );
  AND2_X1 U23132 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20163), .ZN(
        P2_U3187) );
  AND2_X1 U23133 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20163), .ZN(
        P2_U3188) );
  AND2_X1 U23134 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20163), .ZN(
        P2_U3189) );
  AND2_X1 U23135 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20163), .ZN(
        P2_U3190) );
  AND2_X1 U23136 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20163), .ZN(
        P2_U3191) );
  AND2_X1 U23137 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20163), .ZN(
        P2_U3192) );
  AND2_X1 U23138 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20163), .ZN(
        P2_U3193) );
  AND2_X1 U23139 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20163), .ZN(
        P2_U3194) );
  AND2_X1 U23140 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20163), .ZN(
        P2_U3195) );
  AND2_X1 U23141 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20163), .ZN(
        P2_U3196) );
  AND2_X1 U23142 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20163), .ZN(
        P2_U3197) );
  AND2_X1 U23143 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20163), .ZN(
        P2_U3198) );
  AND2_X1 U23144 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20163), .ZN(
        P2_U3199) );
  AND2_X1 U23145 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20163), .ZN(
        P2_U3200) );
  AND2_X1 U23146 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20163), .ZN(P2_U3201) );
  AND2_X1 U23147 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20163), .ZN(P2_U3202) );
  AND2_X1 U23148 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20163), .ZN(P2_U3203) );
  AND2_X1 U23149 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20163), .ZN(P2_U3204) );
  AND2_X1 U23150 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20163), .ZN(P2_U3205) );
  AND2_X1 U23151 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20163), .ZN(P2_U3206) );
  AND2_X1 U23152 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20163), .ZN(P2_U3207) );
  AND2_X1 U23153 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20163), .ZN(P2_U3208) );
  NAND2_X1 U23154 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20175), .ZN(n20177) );
  NAND3_X1 U23155 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20177), .ZN(n20165) );
  AOI211_X1 U23156 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20966), .A(
        n20176), .B(n20229), .ZN(n20164) );
  INV_X1 U23157 ( .A(NA), .ZN(n20970) );
  NOR2_X1 U23158 ( .A1(n20970), .A2(n20169), .ZN(n20182) );
  AOI211_X1 U23159 ( .C1(n20183), .C2(n20165), .A(n20164), .B(n20182), .ZN(
        n20166) );
  INV_X1 U23160 ( .A(n20166), .ZN(P2_U3209) );
  INV_X1 U23161 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20167) );
  AOI21_X1 U23162 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20966), .A(n20183), 
        .ZN(n20173) );
  NOR2_X1 U23163 ( .A1(n20167), .A2(n20173), .ZN(n20170) );
  AOI21_X1 U23164 ( .B1(n20170), .B2(n20169), .A(n20168), .ZN(n20171) );
  OAI211_X1 U23165 ( .C1(n20966), .C2(n20172), .A(n20171), .B(n20177), .ZN(
        P2_U3210) );
  AOI21_X1 U23166 ( .B1(n20175), .B2(n20174), .A(n20173), .ZN(n20181) );
  INV_X1 U23167 ( .A(n20176), .ZN(n20178) );
  OAI22_X1 U23168 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20178), .B1(NA), 
        .B2(n20177), .ZN(n20179) );
  OAI211_X1 U23169 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20179), .ZN(n20180) );
  OAI21_X1 U23170 ( .B1(n20182), .B2(n20181), .A(n20180), .ZN(P2_U3211) );
  OAI222_X1 U23171 ( .A1(n20232), .A2(n20187), .B1(n20185), .B2(n20229), .C1(
        n20184), .C2(n20228), .ZN(P2_U3212) );
  OAI222_X1 U23172 ( .A1(n20228), .A2(n20187), .B1(n20186), .B2(n20229), .C1(
        n13782), .C2(n20232), .ZN(P2_U3213) );
  OAI222_X1 U23173 ( .A1(n20228), .A2(n13782), .B1(n20188), .B2(n20229), .C1(
        n12535), .C2(n20232), .ZN(P2_U3214) );
  OAI222_X1 U23174 ( .A1(n20232), .A2(n20190), .B1(n20189), .B2(n20229), .C1(
        n12535), .C2(n20228), .ZN(P2_U3215) );
  OAI222_X1 U23175 ( .A1(n20232), .A2(n20192), .B1(n20191), .B2(n20229), .C1(
        n20190), .C2(n20228), .ZN(P2_U3216) );
  OAI222_X1 U23176 ( .A1(n20232), .A2(n20194), .B1(n20193), .B2(n20229), .C1(
        n20192), .C2(n20228), .ZN(P2_U3217) );
  OAI222_X1 U23177 ( .A1(n20232), .A2(n13870), .B1(n20195), .B2(n20229), .C1(
        n20194), .C2(n20228), .ZN(P2_U3218) );
  OAI222_X1 U23178 ( .A1(n20232), .A2(n12600), .B1(n20196), .B2(n20229), .C1(
        n13870), .C2(n20228), .ZN(P2_U3219) );
  OAI222_X1 U23179 ( .A1(n20232), .A2(n12603), .B1(n20197), .B2(n20229), .C1(
        n12600), .C2(n20228), .ZN(P2_U3220) );
  OAI222_X1 U23180 ( .A1(n20232), .A2(n12606), .B1(n20198), .B2(n20229), .C1(
        n12603), .C2(n20228), .ZN(P2_U3221) );
  OAI222_X1 U23181 ( .A1(n20232), .A2(n15607), .B1(n20199), .B2(n20229), .C1(
        n12606), .C2(n20228), .ZN(P2_U3222) );
  OAI222_X1 U23182 ( .A1(n20232), .A2(n15589), .B1(n20200), .B2(n20229), .C1(
        n15607), .C2(n20228), .ZN(P2_U3223) );
  OAI222_X1 U23183 ( .A1(n20232), .A2(n15576), .B1(n20201), .B2(n20229), .C1(
        n15589), .C2(n20228), .ZN(P2_U3224) );
  OAI222_X1 U23184 ( .A1(n20232), .A2(n20203), .B1(n20202), .B2(n20229), .C1(
        n15576), .C2(n20228), .ZN(P2_U3225) );
  OAI222_X1 U23185 ( .A1(n20232), .A2(n15552), .B1(n20204), .B2(n20229), .C1(
        n20203), .C2(n20228), .ZN(P2_U3226) );
  OAI222_X1 U23186 ( .A1(n20232), .A2(n20206), .B1(n20205), .B2(n20229), .C1(
        n15552), .C2(n20228), .ZN(P2_U3227) );
  OAI222_X1 U23187 ( .A1(n20232), .A2(n15535), .B1(n20207), .B2(n20229), .C1(
        n20206), .C2(n20228), .ZN(P2_U3228) );
  OAI222_X1 U23188 ( .A1(n20232), .A2(n20209), .B1(n20208), .B2(n20229), .C1(
        n15535), .C2(n20228), .ZN(P2_U3229) );
  OAI222_X1 U23189 ( .A1(n20232), .A2(n15510), .B1(n20210), .B2(n20229), .C1(
        n20209), .C2(n20228), .ZN(P2_U3230) );
  INV_X1 U23190 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20212) );
  OAI222_X1 U23191 ( .A1(n20232), .A2(n20212), .B1(n20211), .B2(n20229), .C1(
        n15510), .C2(n20228), .ZN(P2_U3231) );
  OAI222_X1 U23192 ( .A1(n20232), .A2(n15482), .B1(n20213), .B2(n20229), .C1(
        n20212), .C2(n20228), .ZN(P2_U3232) );
  OAI222_X1 U23193 ( .A1(n20232), .A2(n20215), .B1(n20214), .B2(n20229), .C1(
        n15482), .C2(n20228), .ZN(P2_U3233) );
  OAI222_X1 U23194 ( .A1(n20232), .A2(n20217), .B1(n20216), .B2(n20229), .C1(
        n20215), .C2(n20228), .ZN(P2_U3234) );
  OAI222_X1 U23195 ( .A1(n20232), .A2(n20219), .B1(n20218), .B2(n20229), .C1(
        n20217), .C2(n20228), .ZN(P2_U3235) );
  OAI222_X1 U23196 ( .A1(n20232), .A2(n20221), .B1(n20220), .B2(n20229), .C1(
        n20219), .C2(n20228), .ZN(P2_U3236) );
  OAI222_X1 U23197 ( .A1(n20232), .A2(n20224), .B1(n20222), .B2(n20229), .C1(
        n20221), .C2(n20228), .ZN(P2_U3237) );
  OAI222_X1 U23198 ( .A1(n20228), .A2(n20224), .B1(n20223), .B2(n20229), .C1(
        n14444), .C2(n20232), .ZN(P2_U3238) );
  OAI222_X1 U23199 ( .A1(n20232), .A2(n20226), .B1(n20225), .B2(n20229), .C1(
        n14444), .C2(n20228), .ZN(P2_U3239) );
  OAI222_X1 U23200 ( .A1(n20232), .A2(n12647), .B1(n20227), .B2(n20229), .C1(
        n20226), .C2(n20228), .ZN(P2_U3240) );
  INV_X1 U23201 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20231) );
  INV_X1 U23202 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20230) );
  OAI222_X1 U23203 ( .A1(n20232), .A2(n20231), .B1(n20230), .B2(n20229), .C1(
        n12647), .C2(n20228), .ZN(P2_U3241) );
  OAI22_X1 U23204 ( .A1(n20293), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20229), .ZN(n20233) );
  INV_X1 U23205 ( .A(n20233), .ZN(P2_U3585) );
  MUX2_X1 U23206 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20293), .Z(P2_U3586) );
  OAI22_X1 U23207 ( .A1(n20293), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20229), .ZN(n20234) );
  INV_X1 U23208 ( .A(n20234), .ZN(P2_U3587) );
  OAI22_X1 U23209 ( .A1(n20293), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20229), .ZN(n20235) );
  INV_X1 U23210 ( .A(n20235), .ZN(P2_U3588) );
  OAI21_X1 U23211 ( .B1(n20239), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20237), 
        .ZN(n20236) );
  INV_X1 U23212 ( .A(n20236), .ZN(P2_U3591) );
  OAI21_X1 U23213 ( .B1(n20239), .B2(n20238), .A(n20237), .ZN(P2_U3592) );
  INV_X1 U23214 ( .A(n20240), .ZN(n20252) );
  NOR3_X1 U23215 ( .A1(n20242), .A2(n20241), .A3(n20245), .ZN(n20251) );
  NAND2_X1 U23216 ( .A1(n20243), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20268) );
  NOR2_X1 U23217 ( .A1(n20244), .A2(n20268), .ZN(n20259) );
  INV_X1 U23218 ( .A(n20259), .ZN(n20249) );
  AOI21_X1 U23219 ( .B1(n20267), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20245), 
        .ZN(n20247) );
  NOR2_X1 U23220 ( .A1(n20247), .A2(n20246), .ZN(n20255) );
  AOI21_X1 U23221 ( .B1(n20249), .B2(n20255), .A(n20248), .ZN(n20250) );
  AOI211_X1 U23222 ( .C1(n20252), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20251), 
        .B(n20250), .ZN(n20253) );
  AOI22_X1 U23223 ( .A1(n20279), .A2(n20254), .B1(n20253), .B2(n20280), .ZN(
        P2_U3602) );
  INV_X1 U23224 ( .A(n20255), .ZN(n20257) );
  AOI22_X1 U23225 ( .A1(n20258), .A2(n20257), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20256), .ZN(n20261) );
  NOR2_X1 U23226 ( .A1(n20279), .A2(n20259), .ZN(n20260) );
  AOI22_X1 U23227 ( .A1(n20262), .A2(n20279), .B1(n20261), .B2(n20260), .ZN(
        P2_U3603) );
  INV_X1 U23228 ( .A(n20263), .ZN(n20275) );
  OR3_X1 U23229 ( .A1(n20265), .A2(n20275), .A3(n20264), .ZN(n20266) );
  OAI21_X1 U23230 ( .B1(n20268), .B2(n20267), .A(n20266), .ZN(n20269) );
  AOI21_X1 U23231 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20270), .A(n20269), 
        .ZN(n20271) );
  AOI22_X1 U23232 ( .A1(n20279), .A2(n20272), .B1(n20271), .B2(n20280), .ZN(
        P2_U3604) );
  NAND3_X1 U23233 ( .A1(n20273), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20274) );
  OAI21_X1 U23234 ( .B1(n20276), .B2(n20275), .A(n20274), .ZN(n20277) );
  AOI21_X1 U23235 ( .B1(n20281), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20277), 
        .ZN(n20278) );
  OAI22_X1 U23236 ( .A1(n20281), .A2(n20280), .B1(n20279), .B2(n20278), .ZN(
        P2_U3605) );
  INV_X1 U23237 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20282) );
  AOI22_X1 U23238 ( .A1(n20229), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20282), 
        .B2(n20293), .ZN(P2_U3608) );
  INV_X1 U23239 ( .A(n20283), .ZN(n20292) );
  NOR2_X1 U23240 ( .A1(n20285), .A2(n20284), .ZN(n20287) );
  AOI211_X1 U23241 ( .C1(n20289), .C2(n20288), .A(n20287), .B(n20286), .ZN(
        n20291) );
  NAND2_X1 U23242 ( .A1(n20292), .A2(P2_MORE_REG_SCAN_IN), .ZN(n20290) );
  OAI21_X1 U23243 ( .B1(n20292), .B2(n20291), .A(n20290), .ZN(P2_U3609) );
  MUX2_X1 U23244 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n20293), .Z(P2_U3611) );
  AOI21_X1 U23245 ( .B1(n20979), .B2(P1_STATE_REG_1__SCAN_IN), .A(n20971), 
        .ZN(n20973) );
  INV_X1 U23246 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21165) );
  NAND2_X1 U23247 ( .A1(n20971), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21073) );
  AOI21_X1 U23248 ( .B1(n20973), .B2(n21165), .A(n21031), .ZN(P1_U2802) );
  NAND2_X1 U23249 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21040), .ZN(n20297) );
  OAI21_X1 U23250 ( .B1(n20295), .B2(n20294), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20296) );
  OAI21_X1 U23251 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20297), .A(n20296), 
        .ZN(P1_U2803) );
  NOR2_X1 U23252 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20299) );
  OAI21_X1 U23253 ( .B1(n20299), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21073), .ZN(
        n20298) );
  OAI21_X1 U23254 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21073), .A(n20298), 
        .ZN(P1_U2804) );
  NOR2_X1 U23255 ( .A1(n20973), .A2(n21031), .ZN(n21037) );
  OAI21_X1 U23256 ( .B1(BS16), .B2(n20299), .A(n21037), .ZN(n21035) );
  OAI21_X1 U23257 ( .B1(n21037), .B2(n21129), .A(n21035), .ZN(P1_U2805) );
  AND2_X1 U23258 ( .A1(n20301), .A2(n20300), .ZN(n21058) );
  INV_X1 U23259 ( .A(n21058), .ZN(n21056) );
  AOI21_X1 U23260 ( .B1(n21056), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20302), .ZN(
        n20303) );
  INV_X1 U23261 ( .A(n20303), .ZN(P1_U2806) );
  NOR4_X1 U23262 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20307) );
  NOR4_X1 U23263 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20306) );
  NOR4_X1 U23264 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20305) );
  NOR4_X1 U23265 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20304) );
  NAND4_X1 U23266 ( .A1(n20307), .A2(n20306), .A3(n20305), .A4(n20304), .ZN(
        n20313) );
  NOR4_X1 U23267 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20311) );
  AOI211_X1 U23268 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20310) );
  NOR4_X1 U23269 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20309) );
  NOR4_X1 U23270 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20308) );
  NAND4_X1 U23271 ( .A1(n20311), .A2(n20310), .A3(n20309), .A4(n20308), .ZN(
        n20312) );
  NOR2_X1 U23272 ( .A1(n20313), .A2(n20312), .ZN(n21051) );
  INV_X1 U23273 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21117) );
  NOR3_X1 U23274 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20315) );
  OAI21_X1 U23275 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20315), .A(n21051), .ZN(
        n20314) );
  OAI21_X1 U23276 ( .B1(n21051), .B2(n21117), .A(n20314), .ZN(P1_U2807) );
  INV_X1 U23277 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21036) );
  AOI21_X1 U23278 ( .B1(n21047), .B2(n21036), .A(n20315), .ZN(n20317) );
  INV_X1 U23279 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20316) );
  INV_X1 U23280 ( .A(n21051), .ZN(n21054) );
  AOI22_X1 U23281 ( .A1(n21051), .A2(n20317), .B1(n20316), .B2(n21054), .ZN(
        P1_U2808) );
  AOI22_X1 U23282 ( .A1(n20320), .A2(n20319), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20318), .ZN(n20331) );
  OAI22_X1 U23283 ( .A1(n20363), .A2(n20323), .B1(n20322), .B2(n20321), .ZN(
        n20324) );
  AOI211_X1 U23284 ( .C1(n20345), .C2(n20325), .A(n20334), .B(n20324), .ZN(
        n20330) );
  AOI22_X1 U23285 ( .A1(n20328), .A2(n20327), .B1(n20995), .B2(n20326), .ZN(
        n20329) );
  NAND3_X1 U23286 ( .A1(n20331), .A2(n20330), .A3(n20329), .ZN(P1_U2831) );
  INV_X1 U23287 ( .A(n20332), .ZN(n20342) );
  INV_X1 U23288 ( .A(n20333), .ZN(n20340) );
  AOI21_X1 U23289 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20334), .ZN(n20335) );
  OAI21_X1 U23290 ( .B1(n20336), .B2(n20361), .A(n20335), .ZN(n20337) );
  AOI21_X1 U23291 ( .B1(n20346), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20337), .ZN(
        n20339) );
  NAND3_X1 U23292 ( .A1(n20352), .A2(n20351), .A3(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20338) );
  OAI211_X1 U23293 ( .C1(n20340), .C2(n20377), .A(n20339), .B(n20338), .ZN(
        n20341) );
  AOI21_X1 U23294 ( .B1(n20342), .B2(n20372), .A(n20341), .ZN(n20343) );
  OAI21_X1 U23295 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20344), .A(n20343), .ZN(
        P1_U2835) );
  AOI22_X1 U23296 ( .A1(n20346), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20345), .B2(
        n20428), .ZN(n20359) );
  INV_X1 U23297 ( .A(n20367), .ZN(n20349) );
  NAND3_X1 U23298 ( .A1(n20366), .A2(P1_REIP_REG_3__SCAN_IN), .A3(n20984), 
        .ZN(n20348) );
  OAI211_X1 U23299 ( .C1(n20350), .C2(n20349), .A(n20348), .B(n20347), .ZN(
        n20357) );
  NAND3_X1 U23300 ( .A1(n20352), .A2(n20351), .A3(P1_REIP_REG_4__SCAN_IN), 
        .ZN(n20353) );
  OAI21_X1 U23301 ( .B1(n20355), .B2(n20354), .A(n20353), .ZN(n20356) );
  AOI211_X1 U23302 ( .C1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n20365), .A(
        n20357), .B(n20356), .ZN(n20358) );
  OAI211_X1 U23303 ( .C1(n20360), .C2(n20361), .A(n20359), .B(n20358), .ZN(
        P1_U2836) );
  OAI22_X1 U23304 ( .A1(n20363), .A2(n13340), .B1(n20362), .B2(n20361), .ZN(
        n20364) );
  INV_X1 U23305 ( .A(n20364), .ZN(n20375) );
  AOI22_X1 U23306 ( .A1(n20366), .A2(n13373), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20365), .ZN(n20369) );
  NAND2_X1 U23307 ( .A1(n20663), .A2(n20367), .ZN(n20368) );
  OAI211_X1 U23308 ( .C1(n20370), .C2(n13373), .A(n20369), .B(n20368), .ZN(
        n20371) );
  AOI21_X1 U23309 ( .B1(n20373), .B2(n20372), .A(n20371), .ZN(n20374) );
  OAI211_X1 U23310 ( .C1(n20377), .C2(n20376), .A(n20375), .B(n20374), .ZN(
        P1_U2837) );
  AOI22_X1 U23311 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20381), .B1(n20391), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20378) );
  OAI21_X1 U23312 ( .B1(n20380), .B2(n20379), .A(n20378), .ZN(P1_U2921) );
  INV_X1 U23313 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20383) );
  AOI22_X1 U23314 ( .A1(n20394), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20382) );
  OAI21_X1 U23315 ( .B1(n20383), .B2(n20408), .A(n20382), .ZN(P1_U2922) );
  AOI22_X1 U23316 ( .A1(n20394), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20384) );
  OAI21_X1 U23317 ( .B1(n14859), .B2(n20408), .A(n20384), .ZN(P1_U2923) );
  AOI22_X1 U23318 ( .A1(n20394), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20385) );
  OAI21_X1 U23319 ( .B1(n14862), .B2(n20408), .A(n20385), .ZN(P1_U2924) );
  AOI22_X1 U23320 ( .A1(n20394), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20386) );
  OAI21_X1 U23321 ( .B1(n14866), .B2(n20408), .A(n20386), .ZN(P1_U2925) );
  INV_X1 U23322 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20388) );
  AOI22_X1 U23323 ( .A1(n20394), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20387) );
  OAI21_X1 U23324 ( .B1(n20388), .B2(n20408), .A(n20387), .ZN(P1_U2926) );
  INV_X1 U23325 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20390) );
  AOI22_X1 U23326 ( .A1(n20394), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20389) );
  OAI21_X1 U23327 ( .B1(n20390), .B2(n20408), .A(n20389), .ZN(P1_U2927) );
  AOI22_X1 U23328 ( .A1(n20394), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20392) );
  OAI21_X1 U23329 ( .B1(n20393), .B2(n20408), .A(n20392), .ZN(P1_U2928) );
  AOI22_X1 U23330 ( .A1(n20394), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20395) );
  OAI21_X1 U23331 ( .B1(n10861), .B2(n20408), .A(n20395), .ZN(P1_U2929) );
  AOI22_X1 U23332 ( .A1(n20394), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20396) );
  OAI21_X1 U23333 ( .B1(n20397), .B2(n20408), .A(n20396), .ZN(P1_U2930) );
  AOI22_X1 U23334 ( .A1(n20394), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20398) );
  OAI21_X1 U23335 ( .B1(n13593), .B2(n20408), .A(n20398), .ZN(P1_U2931) );
  AOI22_X1 U23336 ( .A1(n20394), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20399) );
  OAI21_X1 U23337 ( .B1(n20400), .B2(n20408), .A(n20399), .ZN(P1_U2932) );
  AOI22_X1 U23338 ( .A1(n20394), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20401) );
  OAI21_X1 U23339 ( .B1(n20402), .B2(n20408), .A(n20401), .ZN(P1_U2933) );
  AOI22_X1 U23340 ( .A1(n20394), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20403) );
  OAI21_X1 U23341 ( .B1(n20404), .B2(n20408), .A(n20403), .ZN(P1_U2934) );
  AOI22_X1 U23342 ( .A1(n20394), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20405) );
  OAI21_X1 U23343 ( .B1(n20406), .B2(n20408), .A(n20405), .ZN(P1_U2935) );
  AOI22_X1 U23344 ( .A1(n20394), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20391), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20407) );
  OAI21_X1 U23345 ( .B1(n20409), .B2(n20408), .A(n20407), .ZN(P1_U2936) );
  AOI22_X1 U23346 ( .A1(n20421), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20412), .ZN(n20411) );
  NAND2_X1 U23347 ( .A1(n20411), .A2(n20410), .ZN(P1_U2961) );
  AOI22_X1 U23348 ( .A1(n20421), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20412), .ZN(n20414) );
  NAND2_X1 U23349 ( .A1(n20414), .A2(n20413), .ZN(P1_U2962) );
  AOI22_X1 U23350 ( .A1(n20421), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20412), .ZN(n20416) );
  NAND2_X1 U23351 ( .A1(n20416), .A2(n20415), .ZN(P1_U2963) );
  AOI22_X1 U23352 ( .A1(n20421), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20412), .ZN(n20418) );
  NAND2_X1 U23353 ( .A1(n20418), .A2(n20417), .ZN(P1_U2964) );
  AOI22_X1 U23354 ( .A1(n20421), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20412), .ZN(n20420) );
  NAND2_X1 U23355 ( .A1(n20420), .A2(n20419), .ZN(P1_U2965) );
  AOI22_X1 U23356 ( .A1(n20421), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20412), .ZN(n20423) );
  NAND2_X1 U23357 ( .A1(n20423), .A2(n20422), .ZN(P1_U2966) );
  OAI21_X1 U23358 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20424), .ZN(n20435) );
  OR2_X1 U23359 ( .A1(n20426), .A2(n20425), .ZN(n20430) );
  AOI21_X1 U23360 ( .B1(n20438), .B2(n20428), .A(n20427), .ZN(n20429) );
  OAI211_X1 U23361 ( .C1(n20432), .C2(n20431), .A(n20430), .B(n20429), .ZN(
        n20433) );
  INV_X1 U23362 ( .A(n20433), .ZN(n20434) );
  OAI21_X1 U23363 ( .B1(n20436), .B2(n20435), .A(n20434), .ZN(P1_U3027) );
  INV_X1 U23364 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U23365 ( .A1(n20440), .A2(n20439), .B1(n20438), .B2(n20437), .ZN(
        n20449) );
  INV_X1 U23366 ( .A(n20441), .ZN(n20444) );
  NAND3_X1 U23367 ( .A1(n20444), .A2(n20443), .A3(n20442), .ZN(n20445) );
  OAI21_X1 U23368 ( .B1(n20447), .B2(n20446), .A(n20445), .ZN(n20448) );
  OAI211_X1 U23369 ( .C1(n21053), .C2(n20347), .A(n20449), .B(n20448), .ZN(
        P1_U3031) );
  NOR2_X1 U23370 ( .A1(n20451), .A2(n20450), .ZN(P1_U3032) );
  INV_X1 U23371 ( .A(n20777), .ZN(n20455) );
  NOR3_X1 U23372 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20497) );
  NAND2_X1 U23373 ( .A1(n20690), .A2(n20497), .ZN(n20487) );
  OAI22_X1 U23374 ( .A1(n20959), .A2(n20781), .B1(n20723), .B2(n20487), .ZN(
        n20456) );
  INV_X1 U23375 ( .A(n20456), .ZN(n20468) );
  INV_X1 U23376 ( .A(n20519), .ZN(n20457) );
  OAI21_X1 U23377 ( .B1(n20457), .B2(n20945), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20458) );
  NAND2_X1 U23378 ( .A1(n20458), .A2(n20907), .ZN(n20466) );
  OR2_X1 U23379 ( .A1(n20663), .A2(n20459), .ZN(n20548) );
  NOR2_X1 U23380 ( .A1(n20548), .A2(n20866), .ZN(n20463) );
  INV_X1 U23381 ( .A(n20464), .ZN(n20460) );
  NOR2_X1 U23382 ( .A1(n20460), .A2(n20769), .ZN(n20807) );
  INV_X1 U23383 ( .A(n20664), .ZN(n20461) );
  NAND2_X1 U23384 ( .A1(n20461), .A2(n20864), .ZN(n20578) );
  AOI22_X1 U23385 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20578), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20487), .ZN(n20462) );
  OAI211_X1 U23386 ( .C1(n20466), .C2(n20463), .A(n20725), .B(n20462), .ZN(
        n20490) );
  INV_X1 U23387 ( .A(n20463), .ZN(n20465) );
  NOR2_X1 U23388 ( .A1(n20464), .A2(n20769), .ZN(n20719) );
  INV_X1 U23389 ( .A(n20719), .ZN(n20665) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20490), .B1(
        n20898), .B2(n20489), .ZN(n20467) );
  OAI211_X1 U23391 ( .C1(n9777), .C2(n20519), .A(n20468), .B(n20467), .ZN(
        P1_U3033) );
  INV_X1 U23392 ( .A(n20823), .ZN(n20917) );
  OAI22_X1 U23393 ( .A1(n20959), .A2(n20821), .B1(n20820), .B2(n20487), .ZN(
        n20469) );
  INV_X1 U23394 ( .A(n20469), .ZN(n20471) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20490), .B1(
        n20912), .B2(n20489), .ZN(n20470) );
  OAI211_X1 U23396 ( .C1(n20917), .C2(n20519), .A(n20471), .B(n20470), .ZN(
        P1_U3034) );
  OAI22_X1 U23397 ( .A1(n20959), .A2(n20923), .B1(n20827), .B2(n20487), .ZN(
        n20472) );
  INV_X1 U23398 ( .A(n20472), .ZN(n20474) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20490), .B1(
        n20918), .B2(n20489), .ZN(n20473) );
  OAI211_X1 U23400 ( .C1(n9773), .C2(n20519), .A(n20474), .B(n20473), .ZN(
        P1_U3035) );
  INV_X1 U23401 ( .A(n20832), .ZN(n20929) );
  OAI22_X1 U23402 ( .A1(n20959), .A2(n20788), .B1(n20739), .B2(n20487), .ZN(
        n20475) );
  INV_X1 U23403 ( .A(n20475), .ZN(n20477) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20490), .B1(
        n20924), .B2(n20489), .ZN(n20476) );
  OAI211_X1 U23405 ( .C1(n20929), .C2(n20519), .A(n20477), .B(n20476), .ZN(
        P1_U3036) );
  INV_X1 U23406 ( .A(n20836), .ZN(n20935) );
  OAI22_X1 U23407 ( .A1(n20959), .A2(n20791), .B1(n20743), .B2(n20487), .ZN(
        n20478) );
  INV_X1 U23408 ( .A(n20478), .ZN(n20480) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20490), .B1(
        n20930), .B2(n20489), .ZN(n20479) );
  OAI211_X1 U23410 ( .C1(n20935), .C2(n20519), .A(n20480), .B(n20479), .ZN(
        P1_U3037) );
  INV_X1 U23411 ( .A(n20840), .ZN(n20941) );
  OAI22_X1 U23412 ( .A1(n20959), .A2(n20794), .B1(n20747), .B2(n20487), .ZN(
        n20481) );
  INV_X1 U23413 ( .A(n20481), .ZN(n20483) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20490), .B1(
        n20936), .B2(n20489), .ZN(n20482) );
  OAI211_X1 U23415 ( .C1(n20941), .C2(n20519), .A(n20483), .B(n20482), .ZN(
        P1_U3038) );
  OAI22_X1 U23416 ( .A1(n20959), .A2(n20949), .B1(n20845), .B2(n20487), .ZN(
        n20484) );
  INV_X1 U23417 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20490), .B1(
        n20942), .B2(n20489), .ZN(n20485) );
  OAI211_X1 U23419 ( .C1(n9775), .C2(n20519), .A(n20486), .B(n20485), .ZN(
        P1_U3039) );
  INV_X1 U23420 ( .A(n20852), .ZN(n20960) );
  OAI22_X1 U23421 ( .A1(n20959), .A2(n20803), .B1(n20756), .B2(n20487), .ZN(
        n20488) );
  INV_X1 U23422 ( .A(n20488), .ZN(n20492) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20490), .B1(
        n20951), .B2(n20489), .ZN(n20491) );
  OAI211_X1 U23424 ( .C1(n20960), .C2(n20519), .A(n20492), .B(n20491), .ZN(
        P1_U3040) );
  INV_X1 U23425 ( .A(n20497), .ZN(n20494) );
  NOR2_X1 U23426 ( .A1(n20690), .A2(n20494), .ZN(n20515) );
  INV_X1 U23427 ( .A(n20548), .ZN(n20493) );
  INV_X1 U23428 ( .A(n13548), .ZN(n20691) );
  AOI21_X1 U23429 ( .B1(n20493), .B2(n20691), .A(n20515), .ZN(n20495) );
  OAI22_X1 U23430 ( .A1(n20495), .A2(n20901), .B1(n20494), .B2(n20769), .ZN(
        n20514) );
  AOI22_X1 U23431 ( .A1(n20899), .A2(n20515), .B1(n20514), .B2(n20898), .ZN(
        n20501) );
  OAI211_X1 U23432 ( .C1(n20555), .C2(n21129), .A(n20907), .B(n20495), .ZN(
        n20496) );
  OAI211_X1 U23433 ( .C1(n20907), .C2(n20497), .A(n20496), .B(n20906), .ZN(
        n20516) );
  INV_X1 U23434 ( .A(n20697), .ZN(n20498) );
  AOI22_X1 U23435 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20542), .B2(n9778), .ZN(n20500) );
  OAI211_X1 U23436 ( .C1(n20781), .C2(n20519), .A(n20501), .B(n20500), .ZN(
        P1_U3041) );
  AOI22_X1 U23437 ( .A1(n20913), .A2(n20515), .B1(n20514), .B2(n20912), .ZN(
        n20503) );
  AOI22_X1 U23438 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20542), .B2(n20823), .ZN(n20502) );
  OAI211_X1 U23439 ( .C1(n20821), .C2(n20519), .A(n20503), .B(n20502), .ZN(
        P1_U3042) );
  AOI22_X1 U23440 ( .A1(n20919), .A2(n20515), .B1(n20514), .B2(n20918), .ZN(
        n20505) );
  AOI22_X1 U23441 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20542), .B2(n9774), .ZN(n20504) );
  OAI211_X1 U23442 ( .C1(n20923), .C2(n20519), .A(n20505), .B(n20504), .ZN(
        P1_U3043) );
  AOI22_X1 U23443 ( .A1(n20925), .A2(n20515), .B1(n20514), .B2(n20924), .ZN(
        n20507) );
  AOI22_X1 U23444 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20542), .B2(n20832), .ZN(n20506) );
  OAI211_X1 U23445 ( .C1(n20788), .C2(n20519), .A(n20507), .B(n20506), .ZN(
        P1_U3044) );
  AOI22_X1 U23446 ( .A1(n20931), .A2(n20515), .B1(n20514), .B2(n20930), .ZN(
        n20509) );
  AOI22_X1 U23447 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20542), .B2(n20836), .ZN(n20508) );
  OAI211_X1 U23448 ( .C1(n20791), .C2(n20519), .A(n20509), .B(n20508), .ZN(
        P1_U3045) );
  AOI22_X1 U23449 ( .A1(n20937), .A2(n20515), .B1(n20514), .B2(n20936), .ZN(
        n20511) );
  AOI22_X1 U23450 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20542), .B2(n20840), .ZN(n20510) );
  OAI211_X1 U23451 ( .C1(n20794), .C2(n20519), .A(n20511), .B(n20510), .ZN(
        P1_U3046) );
  AOI22_X1 U23452 ( .A1(n20943), .A2(n20515), .B1(n20514), .B2(n20942), .ZN(
        n20513) );
  AOI22_X1 U23453 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20542), .B2(n9776), .ZN(n20512) );
  OAI211_X1 U23454 ( .C1(n20949), .C2(n20519), .A(n20513), .B(n20512), .ZN(
        P1_U3047) );
  AOI22_X1 U23455 ( .A1(n20953), .A2(n20515), .B1(n20514), .B2(n20951), .ZN(
        n20518) );
  AOI22_X1 U23456 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20542), .B2(n20852), .ZN(n20517) );
  OAI211_X1 U23457 ( .C1(n20803), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P1_U3048) );
  NOR3_X1 U23458 ( .A1(n20571), .A2(n20542), .A3(n20901), .ZN(n20520) );
  NOR2_X1 U23459 ( .A1(n20520), .A2(n20804), .ZN(n20526) );
  INV_X1 U23460 ( .A(n20526), .ZN(n20521) );
  NOR2_X1 U23461 ( .A1(n20548), .A2(n9669), .ZN(n20525) );
  NOR3_X1 U23462 ( .A1(n20522), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20550) );
  NAND2_X1 U23463 ( .A1(n20690), .A2(n20550), .ZN(n20523) );
  INV_X1 U23464 ( .A(n20523), .ZN(n20541) );
  AOI22_X1 U23465 ( .A1(n20571), .A2(n9778), .B1(n20899), .B2(n20541), .ZN(
        n20528) );
  NOR2_X1 U23466 ( .A1(n10212), .A2(n20769), .ZN(n20635) );
  AOI21_X1 U23467 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20523), .A(n20635), 
        .ZN(n20524) );
  OAI211_X1 U23468 ( .C1(n20526), .C2(n20525), .A(n20725), .B(n20524), .ZN(
        n20543) );
  AOI22_X1 U23469 ( .A1(n20543), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n20909), .B2(n20542), .ZN(n20527) );
  OAI211_X1 U23470 ( .C1(n20546), .C2(n20819), .A(n20528), .B(n20527), .ZN(
        P1_U3049) );
  AOI22_X1 U23471 ( .A1(n20542), .A2(n20914), .B1(n20913), .B2(n20541), .ZN(
        n20530) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20543), .B1(
        n20571), .B2(n20823), .ZN(n20529) );
  OAI211_X1 U23473 ( .C1(n20546), .C2(n20826), .A(n20530), .B(n20529), .ZN(
        P1_U3050) );
  AOI22_X1 U23474 ( .A1(n20542), .A2(n20876), .B1(n20919), .B2(n20541), .ZN(
        n20532) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20543), .B1(
        n20571), .B2(n9774), .ZN(n20531) );
  OAI211_X1 U23476 ( .C1(n20546), .C2(n20831), .A(n20532), .B(n20531), .ZN(
        P1_U3051) );
  AOI22_X1 U23477 ( .A1(n20571), .A2(n20832), .B1(n20925), .B2(n20541), .ZN(
        n20534) );
  AOI22_X1 U23478 ( .A1(n20543), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n20542), .B2(n20926), .ZN(n20533) );
  OAI211_X1 U23479 ( .C1(n20546), .C2(n20835), .A(n20534), .B(n20533), .ZN(
        P1_U3052) );
  AOI22_X1 U23480 ( .A1(n20571), .A2(n20836), .B1(n20931), .B2(n20541), .ZN(
        n20536) );
  AOI22_X1 U23481 ( .A1(n20543), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n20542), .B2(n20932), .ZN(n20535) );
  OAI211_X1 U23482 ( .C1(n20546), .C2(n20839), .A(n20536), .B(n20535), .ZN(
        P1_U3053) );
  AOI22_X1 U23483 ( .A1(n20571), .A2(n20840), .B1(n20937), .B2(n20541), .ZN(
        n20538) );
  AOI22_X1 U23484 ( .A1(n20543), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n20542), .B2(n20938), .ZN(n20537) );
  OAI211_X1 U23485 ( .C1(n20546), .C2(n20843), .A(n20538), .B(n20537), .ZN(
        P1_U3054) );
  AOI22_X1 U23486 ( .A1(n20542), .A2(n20885), .B1(n20943), .B2(n20541), .ZN(
        n20540) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20543), .B1(
        n20571), .B2(n9776), .ZN(n20539) );
  OAI211_X1 U23488 ( .C1(n20546), .C2(n20850), .A(n20540), .B(n20539), .ZN(
        P1_U3055) );
  AOI22_X1 U23489 ( .A1(n20542), .A2(n20954), .B1(n20953), .B2(n20541), .ZN(
        n20545) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20543), .B1(
        n20571), .B2(n20852), .ZN(n20544) );
  OAI211_X1 U23491 ( .C1(n20546), .C2(n20858), .A(n20545), .B(n20544), .ZN(
        P1_U3056) );
  NOR2_X1 U23492 ( .A1(n20764), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20570) );
  INV_X1 U23493 ( .A(n20570), .ZN(n20547) );
  OAI21_X1 U23494 ( .B1(n20548), .B2(n20767), .A(n20547), .ZN(n20553) );
  AOI21_X1 U23495 ( .B1(n20555), .B2(n20907), .A(n20771), .ZN(n20554) );
  INV_X1 U23496 ( .A(n20554), .ZN(n20549) );
  AOI22_X1 U23497 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20550), .B1(n20553), 
        .B2(n20549), .ZN(n20575) );
  AOI22_X1 U23498 ( .A1(n20571), .A2(n20909), .B1(n20899), .B2(n20570), .ZN(
        n20557) );
  INV_X1 U23499 ( .A(n20550), .ZN(n20551) );
  AOI21_X1 U23500 ( .B1(n20901), .B2(n20551), .A(n20772), .ZN(n20552) );
  OAI21_X1 U23501 ( .B1(n20554), .B2(n20553), .A(n20552), .ZN(n20572) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n9778), .ZN(n20556) );
  OAI211_X1 U23503 ( .C1(n20575), .C2(n20819), .A(n20557), .B(n20556), .ZN(
        P1_U3057) );
  AOI22_X1 U23504 ( .A1(n20571), .A2(n20914), .B1(n20913), .B2(n20570), .ZN(
        n20559) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n20823), .ZN(n20558) );
  OAI211_X1 U23506 ( .C1(n20575), .C2(n20826), .A(n20559), .B(n20558), .ZN(
        P1_U3058) );
  AOI22_X1 U23507 ( .A1(n20571), .A2(n20876), .B1(n20919), .B2(n20570), .ZN(
        n20561) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n9774), .ZN(n20560) );
  OAI211_X1 U23509 ( .C1(n20575), .C2(n20831), .A(n20561), .B(n20560), .ZN(
        P1_U3059) );
  AOI22_X1 U23510 ( .A1(n20571), .A2(n20926), .B1(n20925), .B2(n20570), .ZN(
        n20563) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n20832), .ZN(n20562) );
  OAI211_X1 U23512 ( .C1(n20575), .C2(n20835), .A(n20563), .B(n20562), .ZN(
        P1_U3060) );
  AOI22_X1 U23513 ( .A1(n20571), .A2(n20932), .B1(n20931), .B2(n20570), .ZN(
        n20565) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n20836), .ZN(n20564) );
  OAI211_X1 U23515 ( .C1(n20575), .C2(n20839), .A(n20565), .B(n20564), .ZN(
        P1_U3061) );
  AOI22_X1 U23516 ( .A1(n20571), .A2(n20938), .B1(n20937), .B2(n20570), .ZN(
        n20567) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n20840), .ZN(n20566) );
  OAI211_X1 U23518 ( .C1(n20575), .C2(n20843), .A(n20567), .B(n20566), .ZN(
        P1_U3062) );
  AOI22_X1 U23519 ( .A1(n20571), .A2(n20885), .B1(n20943), .B2(n20570), .ZN(
        n20569) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n9776), .ZN(n20568) );
  OAI211_X1 U23521 ( .C1(n20575), .C2(n20850), .A(n20569), .B(n20568), .ZN(
        P1_U3063) );
  AOI22_X1 U23522 ( .A1(n20571), .A2(n20954), .B1(n20953), .B2(n20570), .ZN(
        n20574) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20572), .B1(
        n20600), .B2(n20852), .ZN(n20573) );
  OAI211_X1 U23524 ( .C1(n20575), .C2(n20858), .A(n20574), .B(n20573), .ZN(
        P1_U3064) );
  NOR3_X1 U23525 ( .A1(n20722), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20608) );
  INV_X1 U23526 ( .A(n20608), .ZN(n20605) );
  NOR2_X1 U23527 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20605), .ZN(
        n20599) );
  INV_X1 U23528 ( .A(n20807), .ZN(n20863) );
  NAND3_X1 U23529 ( .A1(n20604), .A2(n20907), .A3(n9669), .ZN(n20577) );
  OAI21_X1 U23530 ( .B1(n20863), .B2(n20578), .A(n20577), .ZN(n20598) );
  AOI22_X1 U23531 ( .A1(n20899), .A2(n20599), .B1(n20898), .B2(n20598), .ZN(
        n20585) );
  INV_X1 U23532 ( .A(n20600), .ZN(n20579) );
  AOI21_X1 U23533 ( .B1(n20579), .B2(n20629), .A(n21129), .ZN(n20580) );
  AOI21_X1 U23534 ( .B1(n20604), .B2(n9669), .A(n20580), .ZN(n20581) );
  NOR2_X1 U23535 ( .A1(n20581), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20909), .ZN(n20584) );
  OAI211_X1 U23537 ( .C1(n9777), .C2(n20629), .A(n20585), .B(n20584), .ZN(
        P1_U3065) );
  AOI22_X1 U23538 ( .A1(n20913), .A2(n20599), .B1(n20912), .B2(n20598), .ZN(
        n20587) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20914), .ZN(n20586) );
  OAI211_X1 U23540 ( .C1(n20917), .C2(n20629), .A(n20587), .B(n20586), .ZN(
        P1_U3066) );
  AOI22_X1 U23541 ( .A1(n20919), .A2(n20599), .B1(n20918), .B2(n20598), .ZN(
        n20589) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20876), .ZN(n20588) );
  OAI211_X1 U23543 ( .C1(n9773), .C2(n20629), .A(n20589), .B(n20588), .ZN(
        P1_U3067) );
  AOI22_X1 U23544 ( .A1(n20925), .A2(n20599), .B1(n20924), .B2(n20598), .ZN(
        n20591) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20926), .ZN(n20590) );
  OAI211_X1 U23546 ( .C1(n20929), .C2(n20629), .A(n20591), .B(n20590), .ZN(
        P1_U3068) );
  AOI22_X1 U23547 ( .A1(n20931), .A2(n20599), .B1(n20930), .B2(n20598), .ZN(
        n20593) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20932), .ZN(n20592) );
  OAI211_X1 U23549 ( .C1(n20935), .C2(n20629), .A(n20593), .B(n20592), .ZN(
        P1_U3069) );
  AOI22_X1 U23550 ( .A1(n20937), .A2(n20599), .B1(n20936), .B2(n20598), .ZN(
        n20595) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20938), .ZN(n20594) );
  OAI211_X1 U23552 ( .C1(n20941), .C2(n20629), .A(n20595), .B(n20594), .ZN(
        P1_U3070) );
  AOI22_X1 U23553 ( .A1(n20943), .A2(n20599), .B1(n20942), .B2(n20598), .ZN(
        n20597) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20885), .ZN(n20596) );
  OAI211_X1 U23555 ( .C1(n9775), .C2(n20629), .A(n20597), .B(n20596), .ZN(
        P1_U3071) );
  AOI22_X1 U23556 ( .A1(n20953), .A2(n20599), .B1(n20951), .B2(n20598), .ZN(
        n20603) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20601), .B1(
        n20600), .B2(n20954), .ZN(n20602) );
  OAI211_X1 U23558 ( .C1(n20960), .C2(n20629), .A(n20603), .B(n20602), .ZN(
        P1_U3072) );
  NOR2_X1 U23559 ( .A1(n20690), .A2(n20605), .ZN(n20625) );
  AOI21_X1 U23560 ( .B1(n20604), .B2(n20691), .A(n20625), .ZN(n20606) );
  OAI22_X1 U23561 ( .A1(n20606), .A2(n20901), .B1(n20605), .B2(n20769), .ZN(
        n20624) );
  AOI22_X1 U23562 ( .A1(n20899), .A2(n20625), .B1(n20898), .B2(n20624), .ZN(
        n20611) );
  OAI211_X1 U23563 ( .C1(n20609), .C2(n21129), .A(n20907), .B(n20606), .ZN(
        n20607) );
  OAI211_X1 U23564 ( .C1(n20907), .C2(n20608), .A(n20607), .B(n20906), .ZN(
        n20626) );
  AOI22_X1 U23565 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9778), .B2(n20655), .ZN(n20610) );
  OAI211_X1 U23566 ( .C1(n20781), .C2(n20629), .A(n20611), .B(n20610), .ZN(
        P1_U3073) );
  AOI22_X1 U23567 ( .A1(n20913), .A2(n20625), .B1(n20912), .B2(n20624), .ZN(
        n20613) );
  AOI22_X1 U23568 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n20823), .B2(n20655), .ZN(n20612) );
  OAI211_X1 U23569 ( .C1(n20821), .C2(n20629), .A(n20613), .B(n20612), .ZN(
        P1_U3074) );
  AOI22_X1 U23570 ( .A1(n20919), .A2(n20625), .B1(n20918), .B2(n20624), .ZN(
        n20615) );
  AOI22_X1 U23571 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9774), .B2(n20655), .ZN(n20614) );
  OAI211_X1 U23572 ( .C1(n20923), .C2(n20629), .A(n20615), .B(n20614), .ZN(
        P1_U3075) );
  AOI22_X1 U23573 ( .A1(n20925), .A2(n20625), .B1(n20924), .B2(n20624), .ZN(
        n20617) );
  AOI22_X1 U23574 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n20655), .B2(n20832), .ZN(n20616) );
  OAI211_X1 U23575 ( .C1(n20788), .C2(n20629), .A(n20617), .B(n20616), .ZN(
        P1_U3076) );
  AOI22_X1 U23576 ( .A1(n20931), .A2(n20625), .B1(n20930), .B2(n20624), .ZN(
        n20619) );
  AOI22_X1 U23577 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n20655), .B2(n20836), .ZN(n20618) );
  OAI211_X1 U23578 ( .C1(n20791), .C2(n20629), .A(n20619), .B(n20618), .ZN(
        P1_U3077) );
  AOI22_X1 U23579 ( .A1(n20937), .A2(n20625), .B1(n20936), .B2(n20624), .ZN(
        n20621) );
  AOI22_X1 U23580 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n20655), .B2(n20840), .ZN(n20620) );
  OAI211_X1 U23581 ( .C1(n20794), .C2(n20629), .A(n20621), .B(n20620), .ZN(
        P1_U3078) );
  AOI22_X1 U23582 ( .A1(n20943), .A2(n20625), .B1(n20942), .B2(n20624), .ZN(
        n20623) );
  AOI22_X1 U23583 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9776), .B2(n20655), .ZN(n20622) );
  OAI211_X1 U23584 ( .C1(n20949), .C2(n20629), .A(n20623), .B(n20622), .ZN(
        P1_U3079) );
  AOI22_X1 U23585 ( .A1(n20953), .A2(n20625), .B1(n20951), .B2(n20624), .ZN(
        n20628) );
  AOI22_X1 U23586 ( .A1(n20626), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n20655), .B2(n20852), .ZN(n20627) );
  OAI211_X1 U23587 ( .C1(n20803), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        P1_U3080) );
  NOR3_X1 U23588 ( .A1(n20656), .A2(n20655), .A3(n20901), .ZN(n20630) );
  NOR2_X1 U23589 ( .A1(n20630), .A2(n20804), .ZN(n20639) );
  INV_X1 U23590 ( .A(n20639), .ZN(n20632) );
  NOR2_X1 U23591 ( .A1(n20631), .A2(n9669), .ZN(n20638) );
  NOR2_X1 U23592 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20633), .ZN(
        n20654) );
  AOI22_X1 U23593 ( .A1(n20655), .A2(n20909), .B1(n20899), .B2(n20654), .ZN(
        n20641) );
  INV_X1 U23594 ( .A(n20654), .ZN(n20636) );
  INV_X1 U23595 ( .A(n20869), .ZN(n20634) );
  AOI211_X1 U23596 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20636), .A(n20635), 
        .B(n20634), .ZN(n20637) );
  AOI22_X1 U23597 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20656), .B2(n9778), .ZN(n20640) );
  OAI211_X1 U23598 ( .C1(n20660), .C2(n20819), .A(n20641), .B(n20640), .ZN(
        P1_U3081) );
  AOI22_X1 U23599 ( .A1(n20655), .A2(n20914), .B1(n20913), .B2(n20654), .ZN(
        n20643) );
  AOI22_X1 U23600 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20823), .B2(n20656), .ZN(n20642) );
  OAI211_X1 U23601 ( .C1(n20660), .C2(n20826), .A(n20643), .B(n20642), .ZN(
        P1_U3082) );
  AOI22_X1 U23602 ( .A1(n20655), .A2(n20876), .B1(n20919), .B2(n20654), .ZN(
        n20645) );
  AOI22_X1 U23603 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9774), .B2(n20656), .ZN(n20644) );
  OAI211_X1 U23604 ( .C1(n20660), .C2(n20831), .A(n20645), .B(n20644), .ZN(
        P1_U3083) );
  AOI22_X1 U23605 ( .A1(n20655), .A2(n20926), .B1(n20925), .B2(n20654), .ZN(
        n20647) );
  AOI22_X1 U23606 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20656), .B2(n20832), .ZN(n20646) );
  OAI211_X1 U23607 ( .C1(n20660), .C2(n20835), .A(n20647), .B(n20646), .ZN(
        P1_U3084) );
  AOI22_X1 U23608 ( .A1(n20655), .A2(n20932), .B1(n20931), .B2(n20654), .ZN(
        n20649) );
  AOI22_X1 U23609 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20656), .B2(n20836), .ZN(n20648) );
  OAI211_X1 U23610 ( .C1(n20660), .C2(n20839), .A(n20649), .B(n20648), .ZN(
        P1_U3085) );
  AOI22_X1 U23611 ( .A1(n20655), .A2(n20938), .B1(n20937), .B2(n20654), .ZN(
        n20651) );
  AOI22_X1 U23612 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20656), .B2(n20840), .ZN(n20650) );
  OAI211_X1 U23613 ( .C1(n20660), .C2(n20843), .A(n20651), .B(n20650), .ZN(
        P1_U3086) );
  AOI22_X1 U23614 ( .A1(n20655), .A2(n20885), .B1(n20943), .B2(n20654), .ZN(
        n20653) );
  AOI22_X1 U23615 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9776), .B2(n20656), .ZN(n20652) );
  OAI211_X1 U23616 ( .C1(n20660), .C2(n20850), .A(n20653), .B(n20652), .ZN(
        P1_U3087) );
  AOI22_X1 U23617 ( .A1(n20655), .A2(n20954), .B1(n20953), .B2(n20654), .ZN(
        n20659) );
  AOI22_X1 U23618 ( .A1(n20657), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20656), .B2(n20852), .ZN(n20658) );
  OAI211_X1 U23619 ( .C1(n20660), .C2(n20858), .A(n20659), .B(n20658), .ZN(
        P1_U3088) );
  INV_X1 U23620 ( .A(n20778), .ZN(n20662) );
  NOR3_X1 U23621 ( .A1(n20862), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20696) );
  INV_X1 U23622 ( .A(n20696), .ZN(n20693) );
  NOR2_X1 U23623 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20693), .ZN(
        n20685) );
  NAND2_X1 U23624 ( .A1(n20663), .A2(n13257), .ZN(n20768) );
  INV_X1 U23625 ( .A(n20768), .ZN(n20692) );
  AOI21_X1 U23626 ( .B1(n20692), .B2(n9669), .A(n20685), .ZN(n20667) );
  NAND2_X1 U23627 ( .A1(n20664), .A2(n20864), .ZN(n20813) );
  OAI22_X1 U23628 ( .A1(n20667), .A2(n20901), .B1(n20813), .B2(n20665), .ZN(
        n20684) );
  AOI22_X1 U23629 ( .A1(n20899), .A2(n20685), .B1(n20684), .B2(n20898), .ZN(
        n20671) );
  INV_X1 U23630 ( .A(n20717), .ZN(n20666) );
  OAI21_X1 U23631 ( .B1(n20666), .B2(n20686), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20668) );
  NAND2_X1 U23632 ( .A1(n20668), .A2(n20667), .ZN(n20669) );
  AOI22_X1 U23633 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20909), .B2(n20686), .ZN(n20670) );
  OAI211_X1 U23634 ( .C1(n9777), .C2(n20717), .A(n20671), .B(n20670), .ZN(
        P1_U3097) );
  AOI22_X1 U23635 ( .A1(n20913), .A2(n20685), .B1(n20684), .B2(n20912), .ZN(
        n20673) );
  AOI22_X1 U23636 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20914), .B2(n20686), .ZN(n20672) );
  OAI211_X1 U23637 ( .C1(n20917), .C2(n20717), .A(n20673), .B(n20672), .ZN(
        P1_U3098) );
  AOI22_X1 U23638 ( .A1(n20919), .A2(n20685), .B1(n20684), .B2(n20918), .ZN(
        n20675) );
  AOI22_X1 U23639 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20876), .B2(n20686), .ZN(n20674) );
  OAI211_X1 U23640 ( .C1(n9773), .C2(n20717), .A(n20675), .B(n20674), .ZN(
        P1_U3099) );
  AOI22_X1 U23641 ( .A1(n20925), .A2(n20685), .B1(n20684), .B2(n20924), .ZN(
        n20677) );
  AOI22_X1 U23642 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20926), .B2(n20686), .ZN(n20676) );
  OAI211_X1 U23643 ( .C1(n20929), .C2(n20717), .A(n20677), .B(n20676), .ZN(
        P1_U3100) );
  AOI22_X1 U23644 ( .A1(n20931), .A2(n20685), .B1(n20684), .B2(n20930), .ZN(
        n20679) );
  AOI22_X1 U23645 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20932), .B2(n20686), .ZN(n20678) );
  OAI211_X1 U23646 ( .C1(n20935), .C2(n20717), .A(n20679), .B(n20678), .ZN(
        P1_U3101) );
  AOI22_X1 U23647 ( .A1(n20937), .A2(n20685), .B1(n20684), .B2(n20936), .ZN(
        n20681) );
  AOI22_X1 U23648 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20938), .B2(n20686), .ZN(n20680) );
  OAI211_X1 U23649 ( .C1(n20941), .C2(n20717), .A(n20681), .B(n20680), .ZN(
        P1_U3102) );
  AOI22_X1 U23650 ( .A1(n20943), .A2(n20685), .B1(n20684), .B2(n20942), .ZN(
        n20683) );
  AOI22_X1 U23651 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20885), .B2(n20686), .ZN(n20682) );
  OAI211_X1 U23652 ( .C1(n9775), .C2(n20717), .A(n20683), .B(n20682), .ZN(
        P1_U3103) );
  AOI22_X1 U23653 ( .A1(n20953), .A2(n20685), .B1(n20684), .B2(n20951), .ZN(
        n20689) );
  AOI22_X1 U23654 ( .A1(n20687), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20954), .B2(n20686), .ZN(n20688) );
  OAI211_X1 U23655 ( .C1(n20960), .C2(n20717), .A(n20689), .B(n20688), .ZN(
        P1_U3104) );
  NOR2_X1 U23656 ( .A1(n20690), .A2(n20693), .ZN(n20713) );
  AOI21_X1 U23657 ( .B1(n20692), .B2(n20691), .A(n20713), .ZN(n20694) );
  OAI22_X1 U23658 ( .A1(n20694), .A2(n20901), .B1(n20693), .B2(n20769), .ZN(
        n20712) );
  AOI22_X1 U23659 ( .A1(n20899), .A2(n20713), .B1(n20712), .B2(n20898), .ZN(
        n20699) );
  OAI211_X1 U23660 ( .C1(n20778), .C2(n21129), .A(n20907), .B(n20694), .ZN(
        n20695) );
  OAI211_X1 U23661 ( .C1(n20907), .C2(n20696), .A(n20695), .B(n20906), .ZN(
        n20714) );
  AOI22_X1 U23662 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n20752), .B2(n9778), .ZN(n20698) );
  OAI211_X1 U23663 ( .C1(n20781), .C2(n20717), .A(n20699), .B(n20698), .ZN(
        P1_U3105) );
  AOI22_X1 U23664 ( .A1(n20913), .A2(n20713), .B1(n20712), .B2(n20912), .ZN(
        n20701) );
  AOI22_X1 U23665 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n20752), .B2(n20823), .ZN(n20700) );
  OAI211_X1 U23666 ( .C1(n20821), .C2(n20717), .A(n20701), .B(n20700), .ZN(
        P1_U3106) );
  AOI22_X1 U23667 ( .A1(n20919), .A2(n20713), .B1(n20712), .B2(n20918), .ZN(
        n20703) );
  AOI22_X1 U23668 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n20752), .B2(n9774), .ZN(n20702) );
  OAI211_X1 U23669 ( .C1(n20923), .C2(n20717), .A(n20703), .B(n20702), .ZN(
        P1_U3107) );
  AOI22_X1 U23670 ( .A1(n20925), .A2(n20713), .B1(n20712), .B2(n20924), .ZN(
        n20705) );
  AOI22_X1 U23671 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n20752), .B2(n20832), .ZN(n20704) );
  OAI211_X1 U23672 ( .C1(n20788), .C2(n20717), .A(n20705), .B(n20704), .ZN(
        P1_U3108) );
  AOI22_X1 U23673 ( .A1(n20931), .A2(n20713), .B1(n20712), .B2(n20930), .ZN(
        n20707) );
  AOI22_X1 U23674 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n20752), .B2(n20836), .ZN(n20706) );
  OAI211_X1 U23675 ( .C1(n20791), .C2(n20717), .A(n20707), .B(n20706), .ZN(
        P1_U3109) );
  AOI22_X1 U23676 ( .A1(n20937), .A2(n20713), .B1(n20712), .B2(n20936), .ZN(
        n20709) );
  AOI22_X1 U23677 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n20752), .B2(n20840), .ZN(n20708) );
  OAI211_X1 U23678 ( .C1(n20794), .C2(n20717), .A(n20709), .B(n20708), .ZN(
        P1_U3110) );
  AOI22_X1 U23679 ( .A1(n20943), .A2(n20713), .B1(n20712), .B2(n20942), .ZN(
        n20711) );
  AOI22_X1 U23680 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n20752), .B2(n9776), .ZN(n20710) );
  OAI211_X1 U23681 ( .C1(n20949), .C2(n20717), .A(n20711), .B(n20710), .ZN(
        P1_U3111) );
  AOI22_X1 U23682 ( .A1(n20953), .A2(n20713), .B1(n20712), .B2(n20951), .ZN(
        n20716) );
  AOI22_X1 U23683 ( .A1(n20714), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n20752), .B2(n20852), .ZN(n20715) );
  OAI211_X1 U23684 ( .C1(n20803), .C2(n20717), .A(n20716), .B(n20715), .ZN(
        P1_U3112) );
  NOR3_X1 U23685 ( .A1(n20759), .A2(n20752), .A3(n20901), .ZN(n20718) );
  NOR2_X1 U23686 ( .A1(n20718), .A2(n20804), .ZN(n20730) );
  INV_X1 U23687 ( .A(n20730), .ZN(n20721) );
  NOR2_X1 U23688 ( .A1(n20768), .A2(n9669), .ZN(n20729) );
  NOR2_X1 U23689 ( .A1(n20864), .A2(n20862), .ZN(n20720) );
  NAND3_X1 U23690 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20722), .ZN(n20773) );
  OR2_X1 U23691 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20773), .ZN(
        n20755) );
  OAI22_X1 U23692 ( .A1(n20757), .A2(n20781), .B1(n20723), .B2(n20755), .ZN(
        n20724) );
  INV_X1 U23693 ( .A(n20724), .ZN(n20732) );
  INV_X1 U23694 ( .A(n20725), .ZN(n20727) );
  OAI21_X1 U23695 ( .B1(n20862), .B2(n20864), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20870) );
  INV_X1 U23696 ( .A(n20870), .ZN(n20726) );
  AOI211_X1 U23697 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20755), .A(n20727), 
        .B(n20726), .ZN(n20728) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20760), .B1(
        n20759), .B2(n9778), .ZN(n20731) );
  OAI211_X1 U23699 ( .C1(n20763), .C2(n20819), .A(n20732), .B(n20731), .ZN(
        P1_U3113) );
  OAI22_X1 U23700 ( .A1(n20802), .A2(n20917), .B1(n20820), .B2(n20755), .ZN(
        n20733) );
  INV_X1 U23701 ( .A(n20733), .ZN(n20735) );
  AOI22_X1 U23702 ( .A1(n20760), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n20752), .B2(n20914), .ZN(n20734) );
  OAI211_X1 U23703 ( .C1(n20763), .C2(n20826), .A(n20735), .B(n20734), .ZN(
        P1_U3114) );
  OAI22_X1 U23704 ( .A1(n20802), .A2(n9773), .B1(n20827), .B2(n20755), .ZN(
        n20736) );
  INV_X1 U23705 ( .A(n20736), .ZN(n20738) );
  AOI22_X1 U23706 ( .A1(n20760), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20752), .B2(n20876), .ZN(n20737) );
  OAI211_X1 U23707 ( .C1(n20763), .C2(n20831), .A(n20738), .B(n20737), .ZN(
        P1_U3115) );
  OAI22_X1 U23708 ( .A1(n20802), .A2(n20929), .B1(n20739), .B2(n20755), .ZN(
        n20740) );
  INV_X1 U23709 ( .A(n20740), .ZN(n20742) );
  AOI22_X1 U23710 ( .A1(n20760), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20926), .B2(n20752), .ZN(n20741) );
  OAI211_X1 U23711 ( .C1(n20763), .C2(n20835), .A(n20742), .B(n20741), .ZN(
        P1_U3116) );
  OAI22_X1 U23712 ( .A1(n20757), .A2(n20791), .B1(n20743), .B2(n20755), .ZN(
        n20744) );
  INV_X1 U23713 ( .A(n20744), .ZN(n20746) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20760), .B1(
        n20759), .B2(n20836), .ZN(n20745) );
  OAI211_X1 U23715 ( .C1(n20763), .C2(n20839), .A(n20746), .B(n20745), .ZN(
        P1_U3117) );
  OAI22_X1 U23716 ( .A1(n20802), .A2(n20941), .B1(n20747), .B2(n20755), .ZN(
        n20748) );
  INV_X1 U23717 ( .A(n20748), .ZN(n20750) );
  AOI22_X1 U23718 ( .A1(n20760), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n20938), .B2(n20752), .ZN(n20749) );
  OAI211_X1 U23719 ( .C1(n20763), .C2(n20843), .A(n20750), .B(n20749), .ZN(
        P1_U3118) );
  OAI22_X1 U23720 ( .A1(n20802), .A2(n9775), .B1(n20845), .B2(n20755), .ZN(
        n20751) );
  INV_X1 U23721 ( .A(n20751), .ZN(n20754) );
  AOI22_X1 U23722 ( .A1(n20760), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n20752), .B2(n20885), .ZN(n20753) );
  OAI211_X1 U23723 ( .C1(n20763), .C2(n20850), .A(n20754), .B(n20753), .ZN(
        P1_U3119) );
  OAI22_X1 U23724 ( .A1(n20757), .A2(n20803), .B1(n20756), .B2(n20755), .ZN(
        n20758) );
  INV_X1 U23725 ( .A(n20758), .ZN(n20762) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20760), .B1(
        n20759), .B2(n20852), .ZN(n20761) );
  OAI211_X1 U23727 ( .C1(n20763), .C2(n20858), .A(n20762), .B(n20761), .ZN(
        P1_U3120) );
  INV_X1 U23728 ( .A(n20764), .ZN(n20765) );
  NAND2_X1 U23729 ( .A1(n20765), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20766) );
  INV_X1 U23730 ( .A(n20766), .ZN(n20798) );
  OAI21_X1 U23731 ( .B1(n20768), .B2(n20767), .A(n20766), .ZN(n20775) );
  INV_X1 U23732 ( .A(n20775), .ZN(n20770) );
  OAI22_X1 U23733 ( .A1(n20770), .A2(n20901), .B1(n20773), .B2(n20769), .ZN(
        n20797) );
  AOI22_X1 U23734 ( .A1(n20899), .A2(n20798), .B1(n20797), .B2(n20898), .ZN(
        n20780) );
  AOI21_X1 U23735 ( .B1(n20778), .B2(n20907), .A(n20771), .ZN(n20776) );
  AOI21_X1 U23736 ( .B1(n20901), .B2(n20773), .A(n20772), .ZN(n20774) );
  OAI21_X1 U23737 ( .B1(n20776), .B2(n20775), .A(n20774), .ZN(n20799) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n9778), .ZN(n20779) );
  OAI211_X1 U23739 ( .C1(n20781), .C2(n20802), .A(n20780), .B(n20779), .ZN(
        P1_U3121) );
  AOI22_X1 U23740 ( .A1(n20913), .A2(n20798), .B1(n20797), .B2(n20912), .ZN(
        n20783) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n20823), .ZN(n20782) );
  OAI211_X1 U23742 ( .C1(n20821), .C2(n20802), .A(n20783), .B(n20782), .ZN(
        P1_U3122) );
  AOI22_X1 U23743 ( .A1(n20919), .A2(n20798), .B1(n20797), .B2(n20918), .ZN(
        n20785) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n9774), .ZN(n20784) );
  OAI211_X1 U23745 ( .C1(n20923), .C2(n20802), .A(n20785), .B(n20784), .ZN(
        P1_U3123) );
  AOI22_X1 U23746 ( .A1(n20925), .A2(n20798), .B1(n20797), .B2(n20924), .ZN(
        n20787) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n20832), .ZN(n20786) );
  OAI211_X1 U23748 ( .C1(n20788), .C2(n20802), .A(n20787), .B(n20786), .ZN(
        P1_U3124) );
  AOI22_X1 U23749 ( .A1(n20931), .A2(n20798), .B1(n20797), .B2(n20930), .ZN(
        n20790) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n20836), .ZN(n20789) );
  OAI211_X1 U23751 ( .C1(n20791), .C2(n20802), .A(n20790), .B(n20789), .ZN(
        P1_U3125) );
  AOI22_X1 U23752 ( .A1(n20937), .A2(n20798), .B1(n20797), .B2(n20936), .ZN(
        n20793) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n20840), .ZN(n20792) );
  OAI211_X1 U23754 ( .C1(n20794), .C2(n20802), .A(n20793), .B(n20792), .ZN(
        P1_U3126) );
  AOI22_X1 U23755 ( .A1(n20943), .A2(n20798), .B1(n20797), .B2(n20942), .ZN(
        n20796) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n9776), .ZN(n20795) );
  OAI211_X1 U23757 ( .C1(n20949), .C2(n20802), .A(n20796), .B(n20795), .ZN(
        P1_U3127) );
  AOI22_X1 U23758 ( .A1(n20953), .A2(n20798), .B1(n20797), .B2(n20951), .ZN(
        n20801) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20799), .B1(
        n20854), .B2(n20852), .ZN(n20800) );
  OAI211_X1 U23760 ( .C1(n20803), .C2(n20802), .A(n20801), .B(n20800), .ZN(
        P1_U3128) );
  NOR3_X1 U23761 ( .A1(n20854), .A2(n20853), .A3(n20901), .ZN(n20805) );
  NOR2_X1 U23762 ( .A1(n20805), .A2(n20804), .ZN(n20816) );
  INV_X1 U23763 ( .A(n20816), .ZN(n20808) );
  NOR2_X1 U23764 ( .A1(n20865), .A2(n20866), .ZN(n20815) );
  INV_X1 U23765 ( .A(n20813), .ZN(n20806) );
  NOR2_X1 U23766 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20809), .ZN(
        n20851) );
  AOI22_X1 U23767 ( .A1(n20853), .A2(n9778), .B1(n20899), .B2(n20851), .ZN(
        n20818) );
  OAI21_X1 U23768 ( .B1(n20811), .B2(n20851), .A(n20869), .ZN(n20812) );
  AOI21_X1 U23769 ( .B1(n20813), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n20812), 
        .ZN(n20814) );
  AOI22_X1 U23770 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n20909), .ZN(n20817) );
  OAI211_X1 U23771 ( .C1(n20859), .C2(n20819), .A(n20818), .B(n20817), .ZN(
        P1_U3129) );
  INV_X1 U23772 ( .A(n20851), .ZN(n20844) );
  OAI22_X1 U23773 ( .A1(n20846), .A2(n20821), .B1(n20820), .B2(n20844), .ZN(
        n20822) );
  INV_X1 U23774 ( .A(n20822), .ZN(n20825) );
  AOI22_X1 U23775 ( .A1(n20855), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20853), .B2(n20823), .ZN(n20824) );
  OAI211_X1 U23776 ( .C1(n20859), .C2(n20826), .A(n20825), .B(n20824), .ZN(
        P1_U3130) );
  OAI22_X1 U23777 ( .A1(n20846), .A2(n20923), .B1(n20827), .B2(n20844), .ZN(
        n20828) );
  INV_X1 U23778 ( .A(n20828), .ZN(n20830) );
  AOI22_X1 U23779 ( .A1(n20855), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20853), .B2(n9774), .ZN(n20829) );
  OAI211_X1 U23780 ( .C1(n20859), .C2(n20831), .A(n20830), .B(n20829), .ZN(
        P1_U3131) );
  AOI22_X1 U23781 ( .A1(n20853), .A2(n20832), .B1(n20925), .B2(n20851), .ZN(
        n20834) );
  AOI22_X1 U23782 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n20926), .ZN(n20833) );
  OAI211_X1 U23783 ( .C1(n20859), .C2(n20835), .A(n20834), .B(n20833), .ZN(
        P1_U3132) );
  AOI22_X1 U23784 ( .A1(n20853), .A2(n20836), .B1(n20931), .B2(n20851), .ZN(
        n20838) );
  AOI22_X1 U23785 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n20932), .ZN(n20837) );
  OAI211_X1 U23786 ( .C1(n20859), .C2(n20839), .A(n20838), .B(n20837), .ZN(
        P1_U3133) );
  AOI22_X1 U23787 ( .A1(n20853), .A2(n20840), .B1(n20937), .B2(n20851), .ZN(
        n20842) );
  AOI22_X1 U23788 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n20938), .ZN(n20841) );
  OAI211_X1 U23789 ( .C1(n20859), .C2(n20843), .A(n20842), .B(n20841), .ZN(
        P1_U3134) );
  OAI22_X1 U23790 ( .A1(n20846), .A2(n20949), .B1(n20845), .B2(n20844), .ZN(
        n20847) );
  INV_X1 U23791 ( .A(n20847), .ZN(n20849) );
  AOI22_X1 U23792 ( .A1(n20855), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20853), .B2(n9776), .ZN(n20848) );
  OAI211_X1 U23793 ( .C1(n20859), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        P1_U3135) );
  AOI22_X1 U23794 ( .A1(n20853), .A2(n20852), .B1(n20953), .B2(n20851), .ZN(
        n20857) );
  AOI22_X1 U23795 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20855), .B1(
        n20854), .B2(n20954), .ZN(n20856) );
  OAI211_X1 U23796 ( .C1(n20859), .C2(n20858), .A(n20857), .B(n20856), .ZN(
        P1_U3136) );
  INV_X1 U23797 ( .A(n20860), .ZN(n20861) );
  INV_X1 U23798 ( .A(n20908), .ZN(n20897) );
  NOR2_X1 U23799 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20897), .ZN(
        n20889) );
  OAI33_X1 U23800 ( .A1(n9669), .A2(n20865), .A3(n20901), .B1(n20864), .B2(
        n20863), .B3(n20862), .ZN(n20888) );
  AOI22_X1 U23801 ( .A1(n20899), .A2(n20889), .B1(n9780), .B2(n20898), .ZN(
        n20873) );
  OAI21_X1 U23802 ( .B1(n20955), .B2(n20890), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20868) );
  INV_X1 U23803 ( .A(n20865), .ZN(n20896) );
  NAND2_X1 U23804 ( .A1(n20896), .A2(n20866), .ZN(n20867) );
  AOI21_X1 U23805 ( .B1(n20868), .B2(n20867), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20871) );
  AOI22_X1 U23806 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20909), .B2(n20890), .ZN(n20872) );
  OAI211_X1 U23807 ( .C1(n9777), .C2(n20948), .A(n20873), .B(n20872), .ZN(
        P1_U3145) );
  AOI22_X1 U23808 ( .A1(n20913), .A2(n20889), .B1(n9780), .B2(n20912), .ZN(
        n20875) );
  AOI22_X1 U23809 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20914), .B2(n20890), .ZN(n20874) );
  OAI211_X1 U23810 ( .C1(n20917), .C2(n20948), .A(n20875), .B(n20874), .ZN(
        P1_U3146) );
  AOI22_X1 U23811 ( .A1(n20919), .A2(n20889), .B1(n9780), .B2(n20918), .ZN(
        n20878) );
  AOI22_X1 U23812 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20876), .B2(n20890), .ZN(n20877) );
  OAI211_X1 U23813 ( .C1(n9773), .C2(n20948), .A(n20878), .B(n20877), .ZN(
        P1_U3147) );
  AOI22_X1 U23814 ( .A1(n20925), .A2(n20889), .B1(n9780), .B2(n20924), .ZN(
        n20880) );
  AOI22_X1 U23815 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n20926), .B2(n20890), .ZN(n20879) );
  OAI211_X1 U23816 ( .C1(n20929), .C2(n20948), .A(n20880), .B(n20879), .ZN(
        P1_U3148) );
  AOI22_X1 U23817 ( .A1(n20931), .A2(n20889), .B1(n9780), .B2(n20930), .ZN(
        n20882) );
  AOI22_X1 U23818 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n20932), .B2(n20890), .ZN(n20881) );
  OAI211_X1 U23819 ( .C1(n20935), .C2(n20948), .A(n20882), .B(n20881), .ZN(
        P1_U3149) );
  AOI22_X1 U23820 ( .A1(n20937), .A2(n20889), .B1(n9780), .B2(n20936), .ZN(
        n20884) );
  AOI22_X1 U23821 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20938), .B2(n20890), .ZN(n20883) );
  OAI211_X1 U23822 ( .C1(n20941), .C2(n20948), .A(n20884), .B(n20883), .ZN(
        P1_U3150) );
  AOI22_X1 U23823 ( .A1(n20943), .A2(n20889), .B1(n9780), .B2(n20942), .ZN(
        n20887) );
  AOI22_X1 U23824 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20885), .B2(n20890), .ZN(n20886) );
  OAI211_X1 U23825 ( .C1(n9775), .C2(n20948), .A(n20887), .B(n20886), .ZN(
        P1_U3151) );
  AOI22_X1 U23826 ( .A1(n20953), .A2(n20889), .B1(n9780), .B2(n20951), .ZN(
        n20893) );
  AOI22_X1 U23827 ( .A1(n20891), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20890), .B2(n20954), .ZN(n20892) );
  OAI211_X1 U23828 ( .C1(n20960), .C2(n20948), .A(n20893), .B(n20892), .ZN(
        P1_U3152) );
  INV_X1 U23829 ( .A(n20894), .ZN(n20952) );
  AOI21_X1 U23830 ( .B1(n20896), .B2(n20895), .A(n20952), .ZN(n20903) );
  OAI22_X1 U23831 ( .A1(n20903), .A2(n20901), .B1(n20769), .B2(n20897), .ZN(
        n20950) );
  AOI22_X1 U23832 ( .A1(n20899), .A2(n20952), .B1(n20898), .B2(n20950), .ZN(
        n20911) );
  OAI21_X1 U23833 ( .B1(n20902), .B2(n20901), .A(n20900), .ZN(n20904) );
  NAND2_X1 U23834 ( .A1(n20904), .A2(n20903), .ZN(n20905) );
  OAI211_X1 U23835 ( .C1(n20908), .C2(n20907), .A(n20906), .B(n20905), .ZN(
        n20956) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20909), .ZN(n20910) );
  OAI211_X1 U23837 ( .C1(n9777), .C2(n20959), .A(n20911), .B(n20910), .ZN(
        P1_U3153) );
  AOI22_X1 U23838 ( .A1(n20913), .A2(n20952), .B1(n20912), .B2(n20950), .ZN(
        n20916) );
  AOI22_X1 U23839 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20914), .ZN(n20915) );
  OAI211_X1 U23840 ( .C1(n20917), .C2(n20959), .A(n20916), .B(n20915), .ZN(
        P1_U3154) );
  AOI22_X1 U23841 ( .A1(n20919), .A2(n20952), .B1(n20918), .B2(n20950), .ZN(
        n20922) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20956), .B1(
        n20945), .B2(n9774), .ZN(n20921) );
  OAI211_X1 U23843 ( .C1(n20923), .C2(n20948), .A(n20922), .B(n20921), .ZN(
        P1_U3155) );
  AOI22_X1 U23844 ( .A1(n20925), .A2(n20952), .B1(n20924), .B2(n20950), .ZN(
        n20928) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20926), .ZN(n20927) );
  OAI211_X1 U23846 ( .C1(n20929), .C2(n20959), .A(n20928), .B(n20927), .ZN(
        P1_U3156) );
  AOI22_X1 U23847 ( .A1(n20931), .A2(n20952), .B1(n20930), .B2(n20950), .ZN(
        n20934) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20932), .ZN(n20933) );
  OAI211_X1 U23849 ( .C1(n20935), .C2(n20959), .A(n20934), .B(n20933), .ZN(
        P1_U3157) );
  AOI22_X1 U23850 ( .A1(n20937), .A2(n20952), .B1(n20936), .B2(n20950), .ZN(
        n20940) );
  AOI22_X1 U23851 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20938), .ZN(n20939) );
  OAI211_X1 U23852 ( .C1(n20941), .C2(n20959), .A(n20940), .B(n20939), .ZN(
        P1_U3158) );
  AOI22_X1 U23853 ( .A1(n20943), .A2(n20952), .B1(n20942), .B2(n20950), .ZN(
        n20947) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20956), .B1(
        n20945), .B2(n9776), .ZN(n20946) );
  OAI211_X1 U23855 ( .C1(n20949), .C2(n20948), .A(n20947), .B(n20946), .ZN(
        P1_U3159) );
  AOI22_X1 U23856 ( .A1(n20953), .A2(n20952), .B1(n20951), .B2(n20950), .ZN(
        n20958) );
  AOI22_X1 U23857 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20956), .B1(
        n20955), .B2(n20954), .ZN(n20957) );
  OAI211_X1 U23858 ( .C1(n20960), .C2(n20959), .A(n20958), .B(n20957), .ZN(
        P1_U3160) );
  OAI221_X1 U23859 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20963), .C1(n20769), 
        .C2(n20962), .A(n20961), .ZN(P1_U3163) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20964), .ZN(
        P1_U3164) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20964), .ZN(
        P1_U3165) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20964), .ZN(
        P1_U3166) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20964), .ZN(
        P1_U3167) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20964), .ZN(
        P1_U3168) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20964), .ZN(
        P1_U3169) );
  AND2_X1 U23866 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20964), .ZN(
        P1_U3170) );
  AND2_X1 U23867 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20964), .ZN(
        P1_U3171) );
  AND2_X1 U23868 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20964), .ZN(
        P1_U3172) );
  AND2_X1 U23869 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20964), .ZN(
        P1_U3173) );
  AND2_X1 U23870 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20964), .ZN(
        P1_U3174) );
  AND2_X1 U23871 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20964), .ZN(
        P1_U3175) );
  AND2_X1 U23872 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20964), .ZN(
        P1_U3176) );
  AND2_X1 U23873 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20964), .ZN(
        P1_U3177) );
  AND2_X1 U23874 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20964), .ZN(
        P1_U3178) );
  AND2_X1 U23875 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20964), .ZN(
        P1_U3179) );
  AND2_X1 U23876 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20964), .ZN(
        P1_U3180) );
  AND2_X1 U23877 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20964), .ZN(
        P1_U3181) );
  AND2_X1 U23878 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20964), .ZN(
        P1_U3182) );
  AND2_X1 U23879 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20964), .ZN(
        P1_U3183) );
  AND2_X1 U23880 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20964), .ZN(
        P1_U3184) );
  AND2_X1 U23881 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20964), .ZN(
        P1_U3185) );
  AND2_X1 U23882 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20964), .ZN(P1_U3186) );
  AND2_X1 U23883 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20964), .ZN(P1_U3187) );
  AND2_X1 U23884 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20964), .ZN(P1_U3188) );
  AND2_X1 U23885 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20964), .ZN(P1_U3189) );
  AND2_X1 U23886 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20964), .ZN(P1_U3190) );
  AND2_X1 U23887 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20964), .ZN(P1_U3191) );
  AND2_X1 U23888 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20964), .ZN(P1_U3192) );
  AND2_X1 U23889 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20964), .ZN(P1_U3193) );
  AOI21_X1 U23890 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20965), .A(n20971), 
        .ZN(n20978) );
  INV_X1 U23891 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21072) );
  NOR2_X1 U23892 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20967) );
  OAI22_X1 U23893 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20970), .B1(n20967), 
        .B2(n20966), .ZN(n20968) );
  NOR2_X1 U23894 ( .A1(n21072), .A2(n20968), .ZN(n20969) );
  OAI22_X1 U23895 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20978), .B1(n21031), 
        .B2(n20969), .ZN(P1_U3194) );
  OAI21_X1 U23896 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20970), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20977) );
  NOR3_X1 U23897 ( .A1(NA), .A2(n20971), .A3(n21064), .ZN(n20972) );
  NAND3_X1 U23898 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .A3(n20972), .ZN(n20976) );
  OR2_X1 U23899 ( .A1(n20973), .A2(n20972), .ZN(n20974) );
  OAI211_X1 U23900 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21072), .A(HOLD), .B(
        n20974), .ZN(n20975) );
  OAI211_X1 U23901 ( .C1(n20978), .C2(n20977), .A(n20976), .B(n20975), .ZN(
        P1_U3196) );
  INV_X1 U23902 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20980) );
  OAI222_X1 U23903 ( .A1(n21025), .A2(n20981), .B1(n20980), .B2(n21031), .C1(
        n21047), .C2(n21028), .ZN(P1_U3197) );
  INV_X1 U23904 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20982) );
  OAI222_X1 U23905 ( .A1(n21025), .A2(n13373), .B1(n20982), .B2(n21031), .C1(
        n20981), .C2(n21028), .ZN(P1_U3198) );
  OAI222_X1 U23906 ( .A1(n21028), .A2(n13373), .B1(n20983), .B2(n21031), .C1(
        n20984), .C2(n21025), .ZN(P1_U3199) );
  INV_X1 U23907 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20985) );
  OAI222_X1 U23908 ( .A1(n21025), .A2(n20987), .B1(n20985), .B2(n21031), .C1(
        n20984), .C2(n21028), .ZN(P1_U3200) );
  INV_X1 U23909 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20986) );
  OAI222_X1 U23910 ( .A1(n21028), .A2(n20987), .B1(n20986), .B2(n21031), .C1(
        n20989), .C2(n21025), .ZN(P1_U3201) );
  INV_X1 U23911 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20988) );
  OAI222_X1 U23912 ( .A1(n21028), .A2(n20989), .B1(n20988), .B2(n21031), .C1(
        n20991), .C2(n21025), .ZN(P1_U3202) );
  INV_X1 U23913 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20990) );
  OAI222_X1 U23914 ( .A1(n21028), .A2(n20991), .B1(n20990), .B2(n21031), .C1(
        n20992), .C2(n21025), .ZN(P1_U3203) );
  INV_X1 U23915 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20993) );
  OAI222_X1 U23916 ( .A1(n21025), .A2(n20995), .B1(n20993), .B2(n21031), .C1(
        n20992), .C2(n21028), .ZN(P1_U3204) );
  INV_X1 U23917 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20994) );
  OAI222_X1 U23918 ( .A1(n21028), .A2(n20995), .B1(n20994), .B2(n21031), .C1(
        n20996), .C2(n21025), .ZN(P1_U3205) );
  INV_X1 U23919 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20997) );
  OAI222_X1 U23920 ( .A1(n21025), .A2(n20999), .B1(n20997), .B2(n21031), .C1(
        n20996), .C2(n21028), .ZN(P1_U3206) );
  INV_X1 U23921 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20998) );
  OAI222_X1 U23922 ( .A1(n21028), .A2(n20999), .B1(n20998), .B2(n21031), .C1(
        n21001), .C2(n21025), .ZN(P1_U3207) );
  INV_X1 U23923 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21000) );
  OAI222_X1 U23924 ( .A1(n21028), .A2(n21001), .B1(n21000), .B2(n21031), .C1(
        n21003), .C2(n21025), .ZN(P1_U3208) );
  INV_X1 U23925 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21002) );
  OAI222_X1 U23926 ( .A1(n21028), .A2(n21003), .B1(n21002), .B2(n21031), .C1(
        n21004), .C2(n21025), .ZN(P1_U3209) );
  INV_X1 U23927 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21005) );
  OAI222_X1 U23928 ( .A1(n21025), .A2(n21007), .B1(n21005), .B2(n21031), .C1(
        n21004), .C2(n21028), .ZN(P1_U3210) );
  INV_X1 U23929 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21006) );
  OAI222_X1 U23930 ( .A1(n21028), .A2(n21007), .B1(n21006), .B2(n21031), .C1(
        n21009), .C2(n21025), .ZN(P1_U3211) );
  INV_X1 U23931 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21008) );
  OAI222_X1 U23932 ( .A1(n21028), .A2(n21009), .B1(n21008), .B2(n21031), .C1(
        n21010), .C2(n21025), .ZN(P1_U3212) );
  INV_X1 U23933 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21011) );
  OAI222_X1 U23934 ( .A1(n21025), .A2(n14971), .B1(n21011), .B2(n21031), .C1(
        n21010), .C2(n21028), .ZN(P1_U3213) );
  INV_X1 U23935 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21012) );
  OAI222_X1 U23936 ( .A1(n21028), .A2(n14971), .B1(n21012), .B2(n21031), .C1(
        n21014), .C2(n21025), .ZN(P1_U3214) );
  INV_X1 U23937 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21013) );
  OAI222_X1 U23938 ( .A1(n21028), .A2(n21014), .B1(n21013), .B2(n21031), .C1(
        n21164), .C2(n21025), .ZN(P1_U3215) );
  INV_X1 U23939 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21015) );
  OAI222_X1 U23940 ( .A1(n21025), .A2(n21131), .B1(n21015), .B2(n21031), .C1(
        n21164), .C2(n21028), .ZN(P1_U3216) );
  INV_X1 U23941 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21016) );
  OAI222_X1 U23942 ( .A1(n21028), .A2(n21131), .B1(n21016), .B2(n21031), .C1(
        n21168), .C2(n21025), .ZN(P1_U3217) );
  INV_X1 U23943 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21017) );
  OAI222_X1 U23944 ( .A1(n21028), .A2(n21168), .B1(n21017), .B2(n21031), .C1(
        n21018), .C2(n21025), .ZN(P1_U3218) );
  INV_X1 U23945 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21019) );
  OAI222_X1 U23946 ( .A1(n21025), .A2(n21095), .B1(n21019), .B2(n21031), .C1(
        n21018), .C2(n21028), .ZN(P1_U3219) );
  INV_X1 U23947 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21020) );
  INV_X1 U23948 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21235) );
  OAI222_X1 U23949 ( .A1(n21028), .A2(n21095), .B1(n21020), .B2(n21031), .C1(
        n21235), .C2(n21025), .ZN(P1_U3220) );
  INV_X1 U23950 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21021) );
  OAI222_X1 U23951 ( .A1(n21028), .A2(n21235), .B1(n21021), .B2(n21031), .C1(
        n21173), .C2(n21025), .ZN(P1_U3221) );
  INV_X1 U23952 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21022) );
  OAI222_X1 U23953 ( .A1(n21028), .A2(n21173), .B1(n21022), .B2(n21031), .C1(
        n21185), .C2(n21025), .ZN(P1_U3222) );
  INV_X1 U23954 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21023) );
  OAI222_X1 U23955 ( .A1(n21028), .A2(n21185), .B1(n21023), .B2(n21031), .C1(
        n21138), .C2(n21025), .ZN(P1_U3223) );
  INV_X1 U23956 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21024) );
  OAI222_X1 U23957 ( .A1(n21025), .A2(n21182), .B1(n21024), .B2(n21031), .C1(
        n21138), .C2(n21028), .ZN(P1_U3224) );
  INV_X1 U23958 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21026) );
  OAI222_X1 U23959 ( .A1(n21025), .A2(n21201), .B1(n21026), .B2(n21031), .C1(
        n21182), .C2(n21028), .ZN(P1_U3225) );
  INV_X1 U23960 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21027) );
  OAI222_X1 U23961 ( .A1(n21028), .A2(n21201), .B1(n21027), .B2(n21031), .C1(
        n21197), .C2(n21025), .ZN(P1_U3226) );
  OAI22_X1 U23962 ( .A1(n21073), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21031), .ZN(n21029) );
  INV_X1 U23963 ( .A(n21029), .ZN(P1_U3458) );
  OAI22_X1 U23964 ( .A1(n21073), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21031), .ZN(n21030) );
  INV_X1 U23965 ( .A(n21030), .ZN(P1_U3459) );
  OAI22_X1 U23966 ( .A1(n21073), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21031), .ZN(n21032) );
  INV_X1 U23967 ( .A(n21032), .ZN(P1_U3460) );
  OAI22_X1 U23968 ( .A1(n21073), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21031), .ZN(n21033) );
  INV_X1 U23969 ( .A(n21033), .ZN(P1_U3461) );
  OAI21_X1 U23970 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21037), .A(n21035), 
        .ZN(n21034) );
  INV_X1 U23971 ( .A(n21034), .ZN(P1_U3464) );
  OAI21_X1 U23972 ( .B1(n21037), .B2(n21036), .A(n21035), .ZN(P1_U3465) );
  AOI22_X1 U23973 ( .A1(n21041), .A2(n21040), .B1(n21039), .B2(n21038), .ZN(
        n21042) );
  INV_X1 U23974 ( .A(n21042), .ZN(n21044) );
  OAI22_X1 U23975 ( .A1(n21045), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21044), .B2(n21043), .ZN(n21046) );
  INV_X1 U23976 ( .A(n21046), .ZN(P1_U3469) );
  AOI21_X1 U23977 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21048) );
  AOI22_X1 U23978 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21048), .B2(n21047), .ZN(n21050) );
  INV_X1 U23979 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U23980 ( .A1(n21051), .A2(n21050), .B1(n21049), .B2(n21054), .ZN(
        P1_U3481) );
  INV_X1 U23981 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21179) );
  NOR2_X1 U23982 ( .A1(n21054), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21052) );
  AOI22_X1 U23983 ( .A1(n21179), .A2(n21054), .B1(n21053), .B2(n21052), .ZN(
        P1_U3482) );
  AOI22_X1 U23984 ( .A1(n21031), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21055), 
        .B2(n21073), .ZN(P1_U3483) );
  AOI22_X1 U23985 ( .A1(n21058), .A2(n21057), .B1(n16262), .B2(n21056), .ZN(
        P1_U3484) );
  AOI211_X1 U23986 ( .C1(n20394), .C2(n21064), .A(n21060), .B(n21059), .ZN(
        n21071) );
  AOI21_X1 U23987 ( .B1(n21062), .B2(n21129), .A(n21061), .ZN(n21066) );
  INV_X1 U23988 ( .A(n21063), .ZN(n21065) );
  OAI211_X1 U23989 ( .C1(n21066), .C2(n21065), .A(n21064), .B(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21067) );
  NAND2_X1 U23990 ( .A1(n21067), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21070) );
  NOR2_X1 U23991 ( .A1(n21071), .A2(n21068), .ZN(n21069) );
  AOI22_X1 U23992 ( .A1(n21072), .A2(n21071), .B1(n21070), .B2(n21069), .ZN(
        P1_U3485) );
  INV_X1 U23993 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21082) );
  AOI22_X1 U23994 ( .A1(n21031), .A2(n21167), .B1(n21082), .B2(n21073), .ZN(
        P1_U3486) );
  AOI22_X1 U23995 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_f46), .B1(
        DATAI_18_), .B2(keyinput_f14), .ZN(n21074) );
  OAI221_X1 U23996 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .C1(
        DATAI_18_), .C2(keyinput_f14), .A(n21074), .ZN(n21081) );
  AOI22_X1 U23997 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f0), .B1(
        READY1), .B2(keyinput_f36), .ZN(n21075) );
  OAI221_X1 U23998 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .C1(
        READY1), .C2(keyinput_f36), .A(n21075), .ZN(n21080) );
  AOI22_X1 U23999 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(DATAI_5_), .B2(keyinput_f27), .ZN(n21076) );
  OAI221_X1 U24000 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        DATAI_5_), .C2(keyinput_f27), .A(n21076), .ZN(n21079) );
  AOI22_X1 U24001 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n21077) );
  OAI221_X1 U24002 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n21077), .ZN(n21078)
         );
  NOR4_X1 U24003 ( .A1(n21081), .A2(n21080), .A3(n21079), .A4(n21078), .ZN(
        n21111) );
  XNOR2_X1 U24004 ( .A(keyinput_f41), .B(n21082), .ZN(n21089) );
  AOI22_X1 U24005 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n21083) );
  OAI221_X1 U24006 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n21083), .ZN(n21088)
         );
  AOI22_X1 U24007 ( .A1(DATAI_22_), .A2(keyinput_f10), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .ZN(n21084) );
  OAI221_X1 U24008 ( .B1(DATAI_22_), .B2(keyinput_f10), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_f61), .A(n21084), .ZN(n21087)
         );
  AOI22_X1 U24009 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(DATAI_20_), .B2(
        keyinput_f12), .ZN(n21085) );
  OAI221_X1 U24010 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(DATAI_20_), .C2(
        keyinput_f12), .A(n21085), .ZN(n21086) );
  NOR4_X1 U24011 ( .A1(n21089), .A2(n21088), .A3(n21087), .A4(n21086), .ZN(
        n21110) );
  AOI22_X1 U24012 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n21090) );
  OAI221_X1 U24013 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f43), .A(n21090), 
        .ZN(n21099) );
  AOI22_X1 U24014 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_2_), .B2(
        keyinput_f30), .ZN(n21091) );
  OAI221_X1 U24015 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_2_), .C2(
        keyinput_f30), .A(n21091), .ZN(n21098) );
  INV_X1 U24016 ( .A(DATAI_0_), .ZN(n21093) );
  AOI22_X1 U24017 ( .A1(n21093), .A2(keyinput_f32), .B1(n21170), .B2(
        keyinput_f3), .ZN(n21092) );
  OAI221_X1 U24018 ( .B1(n21093), .B2(keyinput_f32), .C1(n21170), .C2(
        keyinput_f3), .A(n21092), .ZN(n21097) );
  AOI22_X1 U24019 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_f54), .B1(
        n21095), .B2(keyinput_f59), .ZN(n21094) );
  OAI221_X1 U24020 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .C1(
        n21095), .C2(keyinput_f59), .A(n21094), .ZN(n21096) );
  NOR4_X1 U24021 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21109) );
  AOI22_X1 U24022 ( .A1(keyinput_f50), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        DATAI_10_), .B2(keyinput_f22), .ZN(n21100) );
  OAI221_X1 U24023 ( .B1(keyinput_f50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), 
        .C1(DATAI_10_), .C2(keyinput_f22), .A(n21100), .ZN(n21107) );
  AOI22_X1 U24024 ( .A1(DATAI_6_), .A2(keyinput_f26), .B1(DATAI_7_), .B2(
        keyinput_f25), .ZN(n21101) );
  OAI221_X1 U24025 ( .B1(DATAI_6_), .B2(keyinput_f26), .C1(DATAI_7_), .C2(
        keyinput_f25), .A(n21101), .ZN(n21106) );
  AOI22_X1 U24026 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n21102) );
  OAI221_X1 U24027 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_f58), .A(n21102), .ZN(n21105)
         );
  AOI22_X1 U24028 ( .A1(DATAI_3_), .A2(keyinput_f29), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .ZN(n21103) );
  OAI221_X1 U24029 ( .B1(DATAI_3_), .B2(keyinput_f29), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21103), .ZN(n21104)
         );
  NOR4_X1 U24030 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21108) );
  NAND4_X1 U24031 ( .A1(n21111), .A2(n21110), .A3(n21109), .A4(n21108), .ZN(
        n21161) );
  INV_X1 U24032 ( .A(keyinput_f35), .ZN(n21113) );
  AOI22_X1 U24033 ( .A1(n21173), .A2(keyinput_f57), .B1(BS16), .B2(n21113), 
        .ZN(n21112) );
  OAI221_X1 U24034 ( .B1(n21173), .B2(keyinput_f57), .C1(n21113), .C2(BS16), 
        .A(n21112), .ZN(n21123) );
  AOI22_X1 U24035 ( .A1(n21115), .A2(keyinput_f2), .B1(keyinput_f20), .B2(
        n21203), .ZN(n21114) );
  OAI221_X1 U24036 ( .B1(n21115), .B2(keyinput_f2), .C1(n21203), .C2(
        keyinput_f20), .A(n21114), .ZN(n21122) );
  AOI22_X1 U24037 ( .A1(n21214), .A2(keyinput_f13), .B1(keyinput_f49), .B2(
        n21117), .ZN(n21116) );
  OAI221_X1 U24038 ( .B1(n21214), .B2(keyinput_f13), .C1(n21117), .C2(
        keyinput_f49), .A(n21116), .ZN(n21121) );
  AOI22_X1 U24039 ( .A1(n21119), .A2(keyinput_f4), .B1(keyinput_f21), .B2(
        n21212), .ZN(n21118) );
  OAI221_X1 U24040 ( .B1(n21119), .B2(keyinput_f4), .C1(n21212), .C2(
        keyinput_f21), .A(n21118), .ZN(n21120) );
  NOR4_X1 U24041 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21159) );
  INV_X1 U24042 ( .A(keyinput_f47), .ZN(n21125) );
  AOI22_X1 U24043 ( .A1(n21237), .A2(keyinput_f6), .B1(P1_W_R_N_REG_SCAN_IN), 
        .B2(n21125), .ZN(n21124) );
  OAI221_X1 U24044 ( .B1(n21237), .B2(keyinput_f6), .C1(n21125), .C2(
        P1_W_R_N_REG_SCAN_IN), .A(n21124), .ZN(n21135) );
  AOI22_X1 U24045 ( .A1(n21195), .A2(keyinput_f8), .B1(n21180), .B2(
        keyinput_f18), .ZN(n21126) );
  OAI221_X1 U24046 ( .B1(n21195), .B2(keyinput_f8), .C1(n21180), .C2(
        keyinput_f18), .A(n21126), .ZN(n21134) );
  INV_X1 U24047 ( .A(keyinput_f33), .ZN(n21128) );
  AOI22_X1 U24048 ( .A1(n21129), .A2(keyinput_f44), .B1(HOLD), .B2(n21128), 
        .ZN(n21127) );
  OAI221_X1 U24049 ( .B1(n21129), .B2(keyinput_f44), .C1(n21128), .C2(HOLD), 
        .A(n21127), .ZN(n21133) );
  AOI22_X1 U24050 ( .A1(n21131), .A2(keyinput_f62), .B1(keyinput_f45), .B2(
        n16262), .ZN(n21130) );
  OAI221_X1 U24051 ( .B1(n21131), .B2(keyinput_f62), .C1(n16262), .C2(
        keyinput_f45), .A(n21130), .ZN(n21132) );
  NOR4_X1 U24052 ( .A1(n21135), .A2(n21134), .A3(n21133), .A4(n21132), .ZN(
        n21158) );
  INV_X1 U24053 ( .A(DATAI_1_), .ZN(n21188) );
  AOI22_X1 U24054 ( .A1(n21165), .A2(keyinput_f39), .B1(n21188), .B2(
        keyinput_f31), .ZN(n21136) );
  OAI221_X1 U24055 ( .B1(n21165), .B2(keyinput_f39), .C1(n21188), .C2(
        keyinput_f31), .A(n21136), .ZN(n21144) );
  AOI22_X1 U24056 ( .A1(n21198), .A2(keyinput_f24), .B1(n21138), .B2(
        keyinput_f55), .ZN(n21137) );
  OAI221_X1 U24057 ( .B1(n21198), .B2(keyinput_f24), .C1(n21138), .C2(
        keyinput_f55), .A(n21137), .ZN(n21143) );
  AOI22_X1 U24058 ( .A1(n21185), .A2(keyinput_f56), .B1(keyinput_f9), .B2(
        n21218), .ZN(n21139) );
  OAI221_X1 U24059 ( .B1(n21185), .B2(keyinput_f56), .C1(n21218), .C2(
        keyinput_f9), .A(n21139), .ZN(n21142) );
  AOI22_X1 U24060 ( .A1(n21200), .A2(keyinput_f19), .B1(keyinput_f48), .B2(
        n21179), .ZN(n21140) );
  OAI221_X1 U24061 ( .B1(n21200), .B2(keyinput_f19), .C1(n21179), .C2(
        keyinput_f48), .A(n21140), .ZN(n21141) );
  NOR4_X1 U24062 ( .A1(n21144), .A2(n21143), .A3(n21142), .A4(n21141), .ZN(
        n21157) );
  AOI22_X1 U24063 ( .A1(n21210), .A2(keyinput_f7), .B1(keyinput_f38), .B2(
        n21187), .ZN(n21145) );
  OAI221_X1 U24064 ( .B1(n21210), .B2(keyinput_f7), .C1(n21187), .C2(
        keyinput_f38), .A(n21145), .ZN(n21155) );
  AOI22_X1 U24065 ( .A1(n21147), .A2(keyinput_f15), .B1(keyinput_f16), .B2(
        n21171), .ZN(n21146) );
  OAI221_X1 U24066 ( .B1(n21147), .B2(keyinput_f15), .C1(n21171), .C2(
        keyinput_f16), .A(n21146), .ZN(n21154) );
  INV_X1 U24067 ( .A(READY2), .ZN(n21184) );
  AOI22_X1 U24068 ( .A1(n21149), .A2(keyinput_f5), .B1(keyinput_f37), .B2(
        n21184), .ZN(n21148) );
  OAI221_X1 U24069 ( .B1(n21149), .B2(keyinput_f5), .C1(n21184), .C2(
        keyinput_f37), .A(n21148), .ZN(n21153) );
  AOI22_X1 U24070 ( .A1(n21201), .A2(keyinput_f53), .B1(n21151), .B2(
        keyinput_f1), .ZN(n21150) );
  OAI221_X1 U24071 ( .B1(n21201), .B2(keyinput_f53), .C1(n21151), .C2(
        keyinput_f1), .A(n21150), .ZN(n21152) );
  NOR4_X1 U24072 ( .A1(n21155), .A2(n21154), .A3(n21153), .A4(n21152), .ZN(
        n21156) );
  NAND4_X1 U24073 ( .A1(n21159), .A2(n21158), .A3(n21157), .A4(n21156), .ZN(
        n21160) );
  OAI22_X1 U24074 ( .A1(n21161), .A2(n21160), .B1(keyinput_f28), .B2(DATAI_4_), 
        .ZN(n21162) );
  AOI21_X1 U24075 ( .B1(keyinput_f28), .B2(DATAI_4_), .A(n21162), .ZN(n21267)
         );
  AOI22_X1 U24076 ( .A1(n21165), .A2(keyinput_g39), .B1(n21164), .B2(
        keyinput_g63), .ZN(n21163) );
  OAI221_X1 U24077 ( .B1(n21165), .B2(keyinput_g39), .C1(n21164), .C2(
        keyinput_g63), .A(n21163), .ZN(n21177) );
  AOI22_X1 U24078 ( .A1(n21168), .A2(keyinput_g61), .B1(keyinput_g0), .B2(
        n21167), .ZN(n21166) );
  OAI221_X1 U24079 ( .B1(n21168), .B2(keyinput_g61), .C1(n21167), .C2(
        keyinput_g0), .A(n21166), .ZN(n21176) );
  AOI22_X1 U24080 ( .A1(n21171), .A2(keyinput_g16), .B1(n21170), .B2(
        keyinput_g3), .ZN(n21169) );
  OAI221_X1 U24081 ( .B1(n21171), .B2(keyinput_g16), .C1(n21170), .C2(
        keyinput_g3), .A(n21169), .ZN(n21175) );
  AOI22_X1 U24082 ( .A1(n13400), .A2(keyinput_g25), .B1(n21173), .B2(
        keyinput_g57), .ZN(n21172) );
  OAI221_X1 U24083 ( .B1(n13400), .B2(keyinput_g25), .C1(n21173), .C2(
        keyinput_g57), .A(n21172), .ZN(n21174) );
  NOR4_X1 U24084 ( .A1(n21177), .A2(n21176), .A3(n21175), .A4(n21174), .ZN(
        n21226) );
  AOI22_X1 U24085 ( .A1(n21180), .A2(keyinput_g18), .B1(keyinput_g48), .B2(
        n21179), .ZN(n21178) );
  OAI221_X1 U24086 ( .B1(n21180), .B2(keyinput_g18), .C1(n21179), .C2(
        keyinput_g48), .A(n21178), .ZN(n21192) );
  AOI22_X1 U24087 ( .A1(n16262), .A2(keyinput_g45), .B1(n21182), .B2(
        keyinput_g54), .ZN(n21181) );
  OAI221_X1 U24088 ( .B1(n16262), .B2(keyinput_g45), .C1(n21182), .C2(
        keyinput_g54), .A(n21181), .ZN(n21191) );
  AOI22_X1 U24089 ( .A1(n21185), .A2(keyinput_g56), .B1(keyinput_g37), .B2(
        n21184), .ZN(n21183) );
  OAI221_X1 U24090 ( .B1(n21185), .B2(keyinput_g56), .C1(n21184), .C2(
        keyinput_g37), .A(n21183), .ZN(n21190) );
  AOI22_X1 U24091 ( .A1(n21188), .A2(keyinput_g31), .B1(keyinput_g38), .B2(
        n21187), .ZN(n21186) );
  OAI221_X1 U24092 ( .B1(n21188), .B2(keyinput_g31), .C1(n21187), .C2(
        keyinput_g38), .A(n21186), .ZN(n21189) );
  NOR4_X1 U24093 ( .A1(n21192), .A2(n21191), .A3(n21190), .A4(n21189), .ZN(
        n21225) );
  INV_X1 U24094 ( .A(BS16), .ZN(n21194) );
  AOI22_X1 U24095 ( .A1(n21195), .A2(keyinput_g8), .B1(keyinput_g35), .B2(
        n21194), .ZN(n21193) );
  OAI221_X1 U24096 ( .B1(n21195), .B2(keyinput_g8), .C1(n21194), .C2(
        keyinput_g35), .A(n21193), .ZN(n21207) );
  AOI22_X1 U24097 ( .A1(n21198), .A2(keyinput_g24), .B1(n21197), .B2(
        keyinput_g52), .ZN(n21196) );
  OAI221_X1 U24098 ( .B1(n21198), .B2(keyinput_g24), .C1(n21197), .C2(
        keyinput_g52), .A(n21196), .ZN(n21206) );
  AOI22_X1 U24099 ( .A1(n21201), .A2(keyinput_g53), .B1(keyinput_g19), .B2(
        n21200), .ZN(n21199) );
  OAI221_X1 U24100 ( .B1(n21201), .B2(keyinput_g53), .C1(n21200), .C2(
        keyinput_g19), .A(n21199), .ZN(n21205) );
  AOI22_X1 U24101 ( .A1(n13424), .A2(keyinput_g27), .B1(n21203), .B2(
        keyinput_g20), .ZN(n21202) );
  OAI221_X1 U24102 ( .B1(n13424), .B2(keyinput_g27), .C1(n21203), .C2(
        keyinput_g20), .A(n21202), .ZN(n21204) );
  NOR4_X1 U24103 ( .A1(n21207), .A2(n21206), .A3(n21205), .A4(n21204), .ZN(
        n21224) );
  INV_X1 U24104 ( .A(DATAI_3_), .ZN(n21209) );
  AOI22_X1 U24105 ( .A1(n21210), .A2(keyinput_g7), .B1(keyinput_g29), .B2(
        n21209), .ZN(n21208) );
  OAI221_X1 U24106 ( .B1(n21210), .B2(keyinput_g7), .C1(n21209), .C2(
        keyinput_g29), .A(n21208), .ZN(n21222) );
  AOI22_X1 U24107 ( .A1(n21212), .A2(keyinput_g21), .B1(keyinput_g26), .B2(
        n13431), .ZN(n21211) );
  OAI221_X1 U24108 ( .B1(n21212), .B2(keyinput_g21), .C1(n13431), .C2(
        keyinput_g26), .A(n21211), .ZN(n21221) );
  INV_X1 U24109 ( .A(DATAI_2_), .ZN(n21215) );
  AOI22_X1 U24110 ( .A1(n21215), .A2(keyinput_g30), .B1(n21214), .B2(
        keyinput_g13), .ZN(n21213) );
  OAI221_X1 U24111 ( .B1(n21215), .B2(keyinput_g30), .C1(n21214), .C2(
        keyinput_g13), .A(n21213), .ZN(n21220) );
  AOI22_X1 U24112 ( .A1(n21218), .A2(keyinput_g9), .B1(keyinput_g10), .B2(
        n21217), .ZN(n21216) );
  OAI221_X1 U24113 ( .B1(n21218), .B2(keyinput_g9), .C1(n21217), .C2(
        keyinput_g10), .A(n21216), .ZN(n21219) );
  NOR4_X1 U24114 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        n21223) );
  NAND4_X1 U24115 ( .A1(n21226), .A2(n21225), .A3(n21224), .A4(n21223), .ZN(
        n21265) );
  AOI22_X1 U24116 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_30_), .B2(keyinput_g2), .ZN(n21227) );
  OAI221_X1 U24117 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(DATAI_30_), .C2(keyinput_g2), .A(n21227), .ZN(n21234) );
  AOI22_X1 U24118 ( .A1(NA), .A2(keyinput_g34), .B1(P1_STATEBS16_REG_SCAN_IN), 
        .B2(keyinput_g44), .ZN(n21228) );
  OAI221_X1 U24119 ( .B1(NA), .B2(keyinput_g34), .C1(P1_STATEBS16_REG_SCAN_IN), 
        .C2(keyinput_g44), .A(n21228), .ZN(n21233) );
  AOI22_X1 U24120 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g51), .B1(
        P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n21229) );
  OAI221_X1 U24121 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), 
        .C1(P1_D_C_N_REG_SCAN_IN), .C2(keyinput_g42), .A(n21229), .ZN(n21232)
         );
  AOI22_X1 U24122 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        DATAI_18_), .B2(keyinput_g14), .ZN(n21230) );
  OAI221_X1 U24123 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        DATAI_18_), .C2(keyinput_g14), .A(n21230), .ZN(n21231) );
  NOR4_X1 U24124 ( .A1(n21234), .A2(n21233), .A3(n21232), .A4(n21231), .ZN(
        n21263) );
  XOR2_X1 U24125 ( .A(n21235), .B(keyinput_g58), .Z(n21243) );
  AOI22_X1 U24126 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(n21237), .B2(
        keyinput_g6), .ZN(n21236) );
  OAI221_X1 U24127 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(n21237), .C2(
        keyinput_g6), .A(n21236), .ZN(n21242) );
  AOI22_X1 U24128 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        DATAI_31_), .B2(keyinput_g1), .ZN(n21238) );
  OAI221_X1 U24129 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        DATAI_31_), .C2(keyinput_g1), .A(n21238), .ZN(n21241) );
  AOI22_X1 U24130 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g43), 
        .B1(READY1), .B2(keyinput_g36), .ZN(n21239) );
  OAI221_X1 U24131 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g43), 
        .C1(READY1), .C2(keyinput_g36), .A(n21239), .ZN(n21240) );
  NOR4_X1 U24132 ( .A1(n21243), .A2(n21242), .A3(n21241), .A4(n21240), .ZN(
        n21262) );
  AOI22_X1 U24133 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        DATAI_20_), .B2(keyinput_g12), .ZN(n21244) );
  OAI221_X1 U24134 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        DATAI_20_), .C2(keyinput_g12), .A(n21244), .ZN(n21251) );
  AOI22_X1 U24135 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .ZN(n21245) );
  OAI221_X1 U24136 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_g55), .A(n21245), .ZN(n21250)
         );
  AOI22_X1 U24137 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(DATAI_10_), .B2(
        keyinput_g22), .ZN(n21246) );
  OAI221_X1 U24138 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(DATAI_10_), .C2(
        keyinput_g22), .A(n21246), .ZN(n21249) );
  AOI22_X1 U24139 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(DATAI_28_), .B2(
        keyinput_g4), .ZN(n21247) );
  OAI221_X1 U24140 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(DATAI_28_), .C2(
        keyinput_g4), .A(n21247), .ZN(n21248) );
  NOR4_X1 U24141 ( .A1(n21251), .A2(n21250), .A3(n21249), .A4(n21248), .ZN(
        n21261) );
  AOI22_X1 U24142 ( .A1(HOLD), .A2(keyinput_g33), .B1(P1_W_R_N_REG_SCAN_IN), 
        .B2(keyinput_g47), .ZN(n21252) );
  OAI221_X1 U24143 ( .B1(HOLD), .B2(keyinput_g33), .C1(P1_W_R_N_REG_SCAN_IN), 
        .C2(keyinput_g47), .A(n21252), .ZN(n21259) );
  AOI22_X1 U24144 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        DATAI_21_), .B2(keyinput_g11), .ZN(n21253) );
  OAI221_X1 U24145 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(DATAI_21_), .C2(keyinput_g11), .A(n21253), .ZN(n21258) );
  AOI22_X1 U24146 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(DATAI_27_), .B2(
        keyinput_g5), .ZN(n21254) );
  OAI221_X1 U24147 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(DATAI_27_), .C2(
        keyinput_g5), .A(n21254), .ZN(n21257) );
  AOI22_X1 U24148 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n21255) );
  OAI221_X1 U24149 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n21255), .ZN(n21256)
         );
  NOR4_X1 U24150 ( .A1(n21259), .A2(n21258), .A3(n21257), .A4(n21256), .ZN(
        n21260) );
  NAND4_X1 U24151 ( .A1(n21263), .A2(n21262), .A3(n21261), .A4(n21260), .ZN(
        n21264) );
  OAI22_X1 U24152 ( .A1(keyinput_g28), .A2(n13411), .B1(n21265), .B2(n21264), 
        .ZN(n21266) );
  AOI211_X1 U24153 ( .C1(keyinput_g28), .C2(n13411), .A(n21267), .B(n21266), 
        .ZN(n21269) );
  AOI22_X1 U24154 ( .A1(n16906), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16908), .ZN(n21268) );
  XNOR2_X1 U24155 ( .A(n21269), .B(n21268), .ZN(U355) );
  AND2_X1 U11164 ( .A1(n15992), .A2(n16709), .ZN(n9640) );
  AND3_X1 U11179 ( .A1(n12397), .A2(n16709), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9644) );
  NOR2_X1 U15930 ( .A1(n13756), .A2(n13755), .ZN(n13898) );
  AND2_X2 U12552 ( .A1(n11824), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12478) );
  AND2_X2 U14978 ( .A1(n12383), .A2(n12026), .ZN(n12167) );
  NAND2_X1 U15937 ( .A1(n14406), .A2(n9633), .ZN(n14335) );
  NAND2_X1 U17622 ( .A1(n14390), .A2(n14406), .ZN(n14371) );
  CLKBUF_X1 U11091 ( .A(n10551), .Z(n10511) );
  INV_X1 U11106 ( .A(n11925), .ZN(n11926) );
  CLKBUF_X2 U11126 ( .A(n13702), .Z(n16001) );
  CLKBUF_X1 U11141 ( .A(n13238), .Z(n9669) );
  CLKBUF_X1 U11158 ( .A(n19589), .Z(n19572) );
  CLKBUF_X1 U11163 ( .A(n11933), .Z(n15993) );
  CLKBUF_X1 U11171 ( .A(n11638), .Z(n17466) );
  OR3_X1 U11209 ( .A1(n14847), .A2(n13623), .A3(n12862), .ZN(n21270) );
endmodule

