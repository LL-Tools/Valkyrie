

module b15_C_gen_AntiSAT_k_256_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031;

  INV_X2 U3597 ( .A(n5065), .ZN(n5448) );
  INV_X2 U3598 ( .A(n3636), .ZN(n5065) );
  NAND2_X1 U3599 ( .A1(n4358), .A2(n4357), .ZN(n5263) );
  NAND2_X1 U3600 ( .A1(n4523), .A2(n4334), .ZN(n4621) );
  NAND2_X1 U3601 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  MUX2_X1 U3602 ( .A(n3501), .B(n3500), .S(n3499), .Z(n6361) );
  BUF_X1 U3603 ( .A(n3340), .Z(n4544) );
  CLKBUF_X2 U3604 ( .A(n4211), .Z(n4116) );
  INV_X1 U3605 ( .A(n4528), .ZN(n4653) );
  CLKBUF_X2 U3606 ( .A(n3415), .Z(n4208) );
  CLKBUF_X2 U3607 ( .A(n3305), .Z(n4217) );
  AND2_X4 U3608 ( .A1(n4582), .A2(n3213), .ZN(n3314) );
  OR2_X1 U3609 ( .A1(n3692), .A2(n3691), .ZN(n3696) );
  AND2_X1 U3610 ( .A1(n3288), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3235) );
  AOI21_X1 U3611 ( .B1(n3150), .B2(INSTQUEUE_REG_14__6__SCAN_IN), .A(n3235), 
        .ZN(n3239) );
  CLKBUF_X2 U3612 ( .A(n3416), .Z(n3393) );
  BUF_X1 U3613 ( .A(n4289), .Z(n4335) );
  NAND2_X2 U3614 ( .A1(n4738), .A2(n4528), .ZN(n4350) );
  INV_X1 U3615 ( .A(n4335), .ZN(n5316) );
  CLKBUF_X2 U3616 ( .A(n3402), .Z(n4563) );
  NOR2_X2 U3617 ( .A1(n3152), .A2(n5312), .ZN(n5311) );
  NOR2_X1 U3619 ( .A1(n5102), .A2(n5293), .ZN(n5662) );
  INV_X1 U3620 ( .A(n5821), .ZN(n5813) );
  OAI21_X2 U3621 ( .B1(n5004), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5065), 
        .ZN(n3639) );
  NAND2_X2 U3622 ( .A1(n4202), .A2(n3659), .ZN(n5393) );
  NAND2_X2 U3623 ( .A1(n3658), .A2(n3657), .ZN(n4202) );
  NOR2_X2 U3624 ( .A1(n4623), .A2(n4715), .ZN(n4709) );
  OAI21_X2 U3625 ( .B1(n4251), .B2(n5463), .A(n4204), .ZN(n4205) );
  OAI22_X2 U3626 ( .A1(n4570), .A2(STATE2_REG_0__SCAN_IN), .B1(n3536), .B2(
        n3471), .ZN(n3476) );
  NAND2_X2 U3627 ( .A1(n3447), .A2(n3366), .ZN(n3445) );
  AND2_X2 U3628 ( .A1(n3386), .A2(n3721), .ZN(n3446) );
  OAI21_X2 U3629 ( .B1(n3643), .B2(n3194), .A(n3192), .ZN(n5051) );
  NAND2_X2 U3630 ( .A1(n5682), .A2(n5683), .ZN(n3643) );
  OR2_X2 U3631 ( .A1(n3370), .A2(n3369), .ZN(n3373) );
  NAND2_X2 U3632 ( .A1(n4256), .A2(n3355), .ZN(n4285) );
  NAND2_X2 U3633 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  XNOR2_X2 U3634 ( .A(n3542), .B(n5988), .ZN(n5900) );
  NAND2_X2 U3635 ( .A1(n3541), .A2(n3540), .ZN(n3542) );
  CLKBUF_X1 U3636 ( .A(n3447), .Z(n3448) );
  AND2_X1 U3637 ( .A1(n4799), .A2(n4514), .ZN(n4494) );
  NOR2_X1 U3638 ( .A1(n4290), .A2(n3350), .ZN(n3374) );
  OAI21_X1 U3639 ( .B1(n3368), .B2(n4512), .A(n3283), .ZN(n4290) );
  AND2_X1 U3641 ( .A1(n3260), .A2(n3357), .ZN(n3283) );
  CLKBUF_X2 U3642 ( .A(n3332), .Z(n4512) );
  CLKBUF_X1 U3643 ( .A(n3357), .Z(n5349) );
  INV_X2 U3644 ( .A(n4291), .ZN(n4649) );
  BUF_X1 U3645 ( .A(n3282), .Z(n4422) );
  BUF_X2 U3646 ( .A(n4220), .Z(n4117) );
  CLKBUF_X2 U3647 ( .A(n3458), .Z(n4219) );
  CLKBUF_X2 U3648 ( .A(n6628), .Z(n6534) );
  CLKBUF_X2 U3649 ( .A(n3408), .Z(n4209) );
  CLKBUF_X2 U3650 ( .A(n3459), .Z(n3388) );
  NOR2_X4 U3651 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U3652 ( .A1(n5059), .A2(n3650), .ZN(n5427) );
  INV_X1 U3653 ( .A(n5189), .ZN(n5283) );
  OR2_X1 U3654 ( .A1(n3735), .A2(n4522), .ZN(n4602) );
  OAI21_X1 U3655 ( .B1(n3716), .B2(n3901), .A(n3758), .ZN(n3735) );
  CLKBUF_X1 U3656 ( .A(n4593), .Z(n6202) );
  NAND2_X1 U3657 ( .A1(n3477), .A2(n3478), .ZN(n3544) );
  NAND2_X1 U3658 ( .A1(n5369), .A2(n4616), .ZN(n5653) );
  NOR2_X1 U3659 ( .A1(n6534), .A2(n4529), .ZN(n5883) );
  AND2_X2 U3660 ( .A1(n5918), .A2(n4192), .ZN(n5921) );
  CLKBUF_X1 U3661 ( .A(n4552), .Z(n6392) );
  OR2_X1 U3662 ( .A1(n3439), .A2(n3438), .ZN(n3444) );
  NAND3_X1 U3663 ( .A1(n3448), .A2(n3168), .A3(n3456), .ZN(n4585) );
  NAND2_X1 U3664 ( .A1(n3449), .A2(n3726), .ZN(n3168) );
  NAND2_X1 U3665 ( .A1(n4341), .A2(n3202), .ZN(n4717) );
  NOR2_X1 U3666 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  INV_X1 U3667 ( .A(n4621), .ZN(n4341) );
  AND2_X1 U3668 ( .A1(n3373), .A2(n3372), .ZN(n4297) );
  INV_X2 U3669 ( .A(n6361), .ZN(n6611) );
  AND2_X1 U3670 ( .A1(n3157), .A2(n3371), .ZN(n3372) );
  NAND2_X1 U3671 ( .A1(n4494), .A2(n4276), .ZN(n4423) );
  AND2_X1 U3672 ( .A1(n3374), .A2(n3351), .ZN(n4273) );
  NOR2_X1 U3673 ( .A1(n4290), .A2(n3491), .ZN(n3715) );
  INV_X1 U3674 ( .A(n3380), .ZN(n4799) );
  CLKBUF_X1 U3675 ( .A(n3482), .Z(n4443) );
  CLKBUF_X1 U3677 ( .A(n3377), .Z(n4790) );
  OR2_X1 U3678 ( .A1(n3426), .A2(n3425), .ZN(n3504) );
  INV_X2 U3679 ( .A(n3340), .ZN(n4733) );
  INV_X1 U3680 ( .A(n3368), .ZN(n3149) );
  INV_X1 U3681 ( .A(n4422), .ZN(n4782) );
  NAND2_X1 U3682 ( .A1(n3245), .A2(n3244), .ZN(n3332) );
  CLKBUF_X1 U3683 ( .A(n3341), .Z(n5350) );
  NAND2_X1 U3684 ( .A1(n3259), .A2(n3258), .ZN(n3357) );
  OR2_X1 U3685 ( .A1(n3414), .A2(n3413), .ZN(n3620) );
  NAND3_X1 U3686 ( .A1(n3155), .A2(n3269), .A3(n3268), .ZN(n4291) );
  NAND4_X2 U3687 ( .A1(n3249), .A2(n3248), .A3(n3246), .A4(n3247), .ZN(n3492)
         );
  AND4_X1 U3688 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3301)
         );
  AND4_X1 U3689 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3303)
         );
  NAND2_X1 U3690 ( .A1(n3153), .A2(n3218), .ZN(n3282) );
  AND3_X1 U3691 ( .A1(n3267), .A2(n3266), .A3(n3265), .ZN(n3268) );
  AND4_X1 U3692 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3341)
         );
  AND4_X1 U3693 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3248)
         );
  AND4_X1 U3694 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3249)
         );
  AND4_X1 U3695 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3246)
         );
  AND4_X1 U3696 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3218)
         );
  NAND2_X2 U3697 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7027), .ZN(n6598) );
  AND2_X2 U3698 ( .A1(n4560), .A2(n4555), .ZN(n4123) );
  AND2_X2 U3699 ( .A1(n4560), .A2(n5583), .ZN(n4220) );
  BUF_X4 U3700 ( .A(n3274), .Z(n3150) );
  AND2_X2 U3701 ( .A1(n3208), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4560)
         );
  AND2_X2 U3702 ( .A1(n3367), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5583)
         );
  AND2_X2 U3703 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4555) );
  INV_X1 U3704 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3367) );
  NOR2_X2 U3705 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4556) );
  NOR2_X4 U3706 ( .A1(n3203), .A2(n5238), .ZN(n5240) );
  NOR2_X2 U3707 ( .A1(n4825), .A2(n4826), .ZN(n4824) );
  NOR3_X4 U3708 ( .A1(n5179), .A2(n5120), .A3(n4415), .ZN(n4420) );
  NOR2_X2 U3709 ( .A1(n5263), .A2(n4367), .ZN(n4943) );
  AOI21_X2 U3710 ( .B1(n5125), .B2(n5168), .A(n5124), .ZN(n5129) );
  OR2_X1 U3711 ( .A1(n3604), .A2(n3603), .ZN(n3630) );
  AND2_X1 U3712 ( .A1(n3345), .A2(n4295), .ZN(n3346) );
  NAND2_X2 U3713 ( .A1(n4501), .A2(n6548), .ZN(n4605) );
  NAND2_X1 U3714 ( .A1(n3630), .A2(n3629), .ZN(n3636) );
  AND2_X1 U3715 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  CLKBUF_X1 U3716 ( .A(n3314), .Z(n4016) );
  CLKBUF_X1 U3717 ( .A(n4145), .Z(n4060) );
  AND2_X2 U3718 ( .A1(n4557), .A2(n4555), .ZN(n3403) );
  NAND2_X1 U3719 ( .A1(n5310), .A2(n3176), .ZN(n3175) );
  INV_X1 U3720 ( .A(n3177), .ZN(n3176) );
  INV_X1 U3721 ( .A(n4233), .ZN(n4183) );
  NAND2_X1 U3722 ( .A1(n4790), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3901) );
  XNOR2_X1 U3723 ( .A(n3630), .B(n3616), .ZN(n3766) );
  INV_X1 U3724 ( .A(n3901), .ZN(n3871) );
  NOR2_X1 U3725 ( .A1(n5393), .A2(n3200), .ZN(n5373) );
  OR2_X1 U3726 ( .A1(n3450), .A2(n4562), .ZN(n3522) );
  XNOR2_X1 U3727 ( .A(n4585), .B(n4584), .ZN(n4552) );
  NAND2_X1 U3728 ( .A1(n5142), .A2(n4441), .ZN(n5140) );
  NOR2_X1 U3729 ( .A1(n5085), .A2(n3171), .ZN(n3170) );
  INV_X1 U3730 ( .A(n4190), .ZN(n3171) );
  INV_X1 U3731 ( .A(n5051), .ZN(n3648) );
  NAND2_X1 U3732 ( .A1(n5065), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5063) );
  AND2_X1 U3733 ( .A1(n4280), .A2(n4279), .ZN(n4426) );
  OR2_X1 U3734 ( .A1(n4605), .A2(n4278), .ZN(n4279) );
  XNOR2_X1 U3735 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U3736 ( .A1(n3158), .A2(n3644), .ZN(n3194) );
  OAI21_X1 U3737 ( .B1(n3352), .B2(n3339), .A(n4653), .ZN(n3370) );
  NAND2_X1 U3738 ( .A1(n4220), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3296)
         );
  AND4_X1 U3739 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3247)
         );
  AND4_X1 U3740 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  AND4_X1 U3741 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3245)
         );
  AOI22_X1 U3742 ( .A1(n3387), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3241) );
  CLKBUF_X1 U3743 ( .A(n3349), .Z(n4615) );
  OR2_X1 U3744 ( .A1(n5099), .A2(n5078), .ZN(n5101) );
  NOR2_X1 U3745 ( .A1(n4430), .A2(n3175), .ZN(n5189) );
  NAND2_X1 U3746 ( .A1(n5321), .A2(n3178), .ZN(n3177) );
  INV_X1 U3747 ( .A(n5324), .ZN(n3178) );
  NAND2_X1 U3748 ( .A1(n3904), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4233) );
  NOR2_X1 U3749 ( .A1(n4980), .A2(n4991), .ZN(n3858) );
  INV_X1 U3750 ( .A(n3732), .ZN(n4186) );
  AND2_X1 U3751 ( .A1(n3470), .A2(n3620), .ZN(n3628) );
  AND2_X1 U3752 ( .A1(n5415), .A2(n5406), .ZN(n3188) );
  XNOR2_X1 U3753 ( .A(n3476), .B(n3475), .ZN(n3478) );
  OR2_X1 U3754 ( .A1(n3450), .A2(n5117), .ZN(n3455) );
  NAND2_X1 U3755 ( .A1(n3328), .A2(n3149), .ZN(n4496) );
  INV_X1 U3756 ( .A(n6202), .ZN(n6238) );
  NAND2_X1 U3757 ( .A1(n6436), .A2(n6793), .ZN(n4236) );
  CLKBUF_X1 U3758 ( .A(n4273), .Z(n4274) );
  AND4_X1 U3759 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3258)
         );
  AND4_X1 U3760 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3259)
         );
  AND4_X1 U3761 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3324)
         );
  AND4_X1 U3762 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3323)
         );
  AND4_X1 U3763 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3326)
         );
  INV_X1 U3764 ( .A(n3175), .ZN(n3174) );
  CLKBUF_X1 U3765 ( .A(n5374), .Z(n5399) );
  NOR2_X1 U3766 ( .A1(n5283), .A2(n5101), .ZN(n5293) );
  OR2_X1 U3767 ( .A1(n5283), .A2(n5078), .ZN(n5100) );
  AND2_X1 U3768 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3985), .ZN(n3986)
         );
  OR2_X1 U3769 ( .A1(n5047), .A2(n3179), .ZN(n4432) );
  OR2_X1 U3770 ( .A1(n3181), .A2(n3180), .ZN(n3179) );
  INV_X1 U3771 ( .A(n5224), .ZN(n3180) );
  AND2_X1 U3772 ( .A1(n3871), .A2(n3870), .ZN(n5042) );
  AND2_X1 U3773 ( .A1(n3785), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3790)
         );
  NOR2_X1 U3774 ( .A1(n5262), .A2(n5260), .ZN(n3773) );
  INV_X1 U3775 ( .A(n5415), .ZN(n3184) );
  NOR2_X1 U3776 ( .A1(n3190), .A2(n5091), .ZN(n3187) );
  NOR2_X1 U3777 ( .A1(n5448), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5406)
         );
  AOI21_X1 U3778 ( .B1(n5420), .B2(n3199), .A(n3161), .ZN(n5413) );
  INV_X1 U3779 ( .A(n5430), .ZN(n5062) );
  NOR2_X1 U3780 ( .A1(n3645), .A2(n3196), .ZN(n3195) );
  INV_X1 U3781 ( .A(n3642), .ZN(n3196) );
  MUX2_X1 U3782 ( .A(n3711), .B(n4197), .S(n6619), .Z(n3723) );
  NAND2_X1 U3783 ( .A1(n3486), .A2(n3489), .ZN(n4593) );
  CLKBUF_X1 U3784 ( .A(n3738), .Z(n4594) );
  NOR2_X1 U3785 ( .A1(n6030), .A2(n6029), .ZN(n6434) );
  NAND2_X1 U3786 ( .A1(n3535), .A2(n3534), .ZN(n6383) );
  NAND2_X1 U3787 ( .A1(n4552), .A2(n6542), .ZN(n3535) );
  NOR2_X1 U3788 ( .A1(n6027), .A2(n6238), .ZN(n6384) );
  AND2_X1 U3789 ( .A1(n5587), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3711) );
  OR2_X1 U3790 ( .A1(n5634), .A2(n5136), .ZN(n5617) );
  NAND2_X1 U3791 ( .A1(n4708), .A2(n4614), .ZN(n5369) );
  AOI21_X1 U3792 ( .B1(n4613), .B2(n4612), .A(n4611), .ZN(n4614) );
  XNOR2_X1 U3793 ( .A(n4243), .B(n5144), .ZN(n4447) );
  XNOR2_X1 U3794 ( .A(n3173), .B(n3172), .ZN(n5345) );
  OR2_X2 U3795 ( .A1(n4605), .A2(n4281), .ZN(n5918) );
  OR2_X1 U3796 ( .A1(n4426), .A2(n4288), .ZN(n6018) );
  INV_X1 U3797 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6619) );
  CLKBUF_X1 U3798 ( .A(n4570), .Z(n6030) );
  INV_X1 U3799 ( .A(n6612), .ZN(n6438) );
  AND2_X1 U3800 ( .A1(n3711), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6548) );
  OR2_X1 U3801 ( .A1(n3681), .A2(n3682), .ZN(n3664) );
  CLKBUF_X1 U3802 ( .A(n4122), .Z(n4017) );
  INV_X1 U3803 ( .A(n3566), .ZN(n3590) );
  NAND2_X1 U3804 ( .A1(n3590), .A2(n3589), .ZN(n3604) );
  AND2_X1 U3805 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  AND2_X1 U3806 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  OR2_X1 U3807 ( .A1(n3576), .A2(n3575), .ZN(n3606) );
  OR2_X1 U3808 ( .A1(n3556), .A2(n3555), .ZN(n3605) );
  OR2_X1 U3809 ( .A1(n3399), .A2(n3398), .ZN(n3490) );
  OR2_X1 U3810 ( .A1(n3469), .A2(n3468), .ZN(n3473) );
  NAND2_X1 U3811 ( .A1(n3348), .A2(n3160), .ZN(n3169) );
  AND2_X2 U3812 ( .A1(n3207), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3213)
         );
  NAND2_X1 U3813 ( .A1(n3344), .A2(n3343), .ZN(n4295) );
  NAND2_X1 U3814 ( .A1(n3348), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U3815 ( .A1(n3431), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3670) );
  NOR2_X1 U3816 ( .A1(n3679), .A2(n3678), .ZN(n4265) );
  AND2_X1 U3817 ( .A1(n3673), .A2(n5736), .ZN(n3679) );
  NAND2_X1 U3818 ( .A1(n3354), .A2(n4733), .ZN(n3380) );
  NAND2_X1 U3819 ( .A1(n3403), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U3820 ( .A1(n4123), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3316)
         );
  OR2_X1 U3821 ( .A1(n5250), .A2(n5056), .ZN(n3181) );
  NOR2_X1 U3822 ( .A1(n3835), .A2(n5784), .ZN(n3853) );
  AND2_X1 U3823 ( .A1(n4940), .A2(n4931), .ZN(n3182) );
  INV_X1 U3824 ( .A(n5401), .ZN(n3657) );
  INV_X1 U3825 ( .A(n3193), .ZN(n3192) );
  OAI21_X1 U3826 ( .B1(n3195), .B2(n3194), .A(n3646), .ZN(n3193) );
  NAND2_X1 U3827 ( .A1(n4957), .A2(n4954), .ZN(n3197) );
  NAND2_X1 U3828 ( .A1(n3492), .A2(n4544), .ZN(n3669) );
  INV_X1 U3829 ( .A(n3669), .ZN(n3627) );
  OR2_X1 U3830 ( .A1(n4426), .A2(n4299), .ZN(n5709) );
  CLKBUF_X1 U3831 ( .A(n3374), .Z(n3375) );
  NAND2_X1 U3832 ( .A1(n3439), .A2(n3438), .ZN(n3198) );
  INV_X1 U3833 ( .A(n4649), .ZN(n4267) );
  AND2_X1 U3834 ( .A1(n6030), .A2(n5586), .ZN(n4871) );
  AND2_X1 U3835 ( .A1(n3518), .A2(n6433), .ZN(n6203) );
  INV_X1 U3836 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U3837 ( .A1(n6027), .A2(n6202), .ZN(n4747) );
  AND2_X1 U3838 ( .A1(n3429), .A2(n3428), .ZN(n3500) );
  OR2_X1 U3839 ( .A1(n3440), .A2(n3427), .ZN(n3429) );
  INV_X1 U3840 ( .A(n3504), .ZN(n3427) );
  AND4_X1 U3841 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3304)
         );
  AND4_X1 U3842 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3302)
         );
  OR2_X1 U3843 ( .A1(n3533), .A2(n3532), .ZN(n3559) );
  AND2_X1 U3844 ( .A1(n3523), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3707) );
  INV_X1 U3845 ( .A(n3670), .ZN(n3702) );
  AOI21_X1 U3846 ( .B1(n6555), .B2(n6530), .A(n5590), .ZN(n4636) );
  NOR2_X1 U3847 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4636), .ZN(n6101) );
  INV_X1 U3848 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6517) );
  AND2_X1 U3849 ( .A1(n4473), .A2(n4434), .ZN(n4469) );
  INV_X1 U3850 ( .A(n3482), .ZN(n6630) );
  NOR2_X1 U3851 ( .A1(n6969), .A2(n5229), .ZN(n5147) );
  AND2_X1 U3852 ( .A1(n4409), .A2(n4408), .ZN(n5288) );
  AND2_X1 U3853 ( .A1(n4381), .A2(n4380), .ZN(n5238) );
  INV_X1 U3854 ( .A(n5885), .ZN(n4529) );
  NOR2_X1 U3855 ( .A1(n4543), .A2(READY_N), .ZN(n4545) );
  OR2_X1 U3856 ( .A1(n4206), .A2(n5170), .ZN(n4241) );
  NOR2_X1 U3857 ( .A1(n4163), .A2(n4162), .ZN(n4164) );
  OR2_X1 U3858 ( .A1(n4168), .A2(n4167), .ZN(n5178) );
  NAND2_X1 U3859 ( .A1(n4084), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4163)
         );
  AND2_X1 U3860 ( .A1(n4136), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4103)
         );
  NOR2_X1 U3861 ( .A1(n4074), .A2(n5627), .ZN(n4134) );
  AND2_X1 U3862 ( .A1(n4134), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4136)
         );
  AND2_X1 U3863 ( .A1(n5625), .A2(n4436), .ZN(n4003) );
  AND2_X1 U3864 ( .A1(n3988), .A2(n3987), .ZN(n5321) );
  NOR2_X1 U3865 ( .A1(n3935), .A2(n3934), .ZN(n3936) );
  INV_X1 U3866 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U3867 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3984)
         );
  INV_X1 U3868 ( .A(n4432), .ZN(n3953) );
  NAND2_X1 U3869 ( .A1(n3919), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3935)
         );
  NOR2_X1 U3870 ( .A1(n3903), .A2(n5255), .ZN(n3919) );
  CLKBUF_X1 U3871 ( .A(n5051), .Z(n5052) );
  NOR2_X1 U3872 ( .A1(n5047), .A2(n3181), .ZN(n5223) );
  NAND2_X1 U3873 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3903)
         );
  INV_X1 U3874 ( .A(n3886), .ZN(n3887) );
  OR2_X1 U3875 ( .A1(n5047), .A2(n5250), .ZN(n5248) );
  AND2_X1 U3876 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3854)
         );
  NAND2_X1 U3877 ( .A1(n3818), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3835)
         );
  NOR2_X1 U3878 ( .A1(n3814), .A2(n5793), .ZN(n3818) );
  NAND2_X1 U3879 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3814)
         );
  AND4_X1 U3880 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n4826)
         );
  AOI21_X1 U3881 ( .B1(n3766), .B2(n3871), .A(n3765), .ZN(n5262) );
  NAND2_X1 U3882 ( .A1(n3762), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3767)
         );
  INV_X1 U3883 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3769) );
  NOR2_X1 U3884 ( .A1(n3767), .A2(n3769), .ZN(n3785) );
  NAND2_X1 U3885 ( .A1(n4913), .A2(n4912), .ZN(n4911) );
  AND2_X1 U3886 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3751), .ZN(n3762)
         );
  INV_X1 U3887 ( .A(n3739), .ZN(n3740) );
  AND2_X1 U3888 ( .A1(n4520), .A2(n4519), .ZN(n4522) );
  OR2_X1 U3889 ( .A1(n4282), .A2(n3368), .ZN(n4281) );
  NOR2_X2 U3890 ( .A1(n5300), .A2(n5288), .ZN(n5287) );
  AND2_X1 U3891 ( .A1(n4385), .A2(n4384), .ZN(n5225) );
  NOR2_X2 U3892 ( .A1(n5725), .A2(n5724), .ZN(n5727) );
  INV_X1 U3893 ( .A(n5266), .ZN(n4357) );
  INV_X1 U3894 ( .A(n5265), .ZN(n4358) );
  NAND2_X1 U3895 ( .A1(n4809), .A2(n4808), .ZN(n5265) );
  AND2_X1 U3896 ( .A1(n4719), .A2(n4712), .ZN(n4809) );
  NOR2_X2 U3897 ( .A1(n4717), .A2(n4716), .ZN(n4719) );
  AND2_X1 U3898 ( .A1(n6025), .A2(n5709), .ZN(n5927) );
  AOI21_X1 U3899 ( .B1(n4904), .B2(n4903), .A(n3512), .ZN(n5906) );
  OR2_X1 U3900 ( .A1(n4426), .A2(n4554), .ZN(n5708) );
  CLKBUF_X1 U3901 ( .A(n4283), .Z(n4284) );
  NAND2_X1 U3902 ( .A1(n3168), .A2(n3448), .ZN(n3167) );
  CLKBUF_X1 U3903 ( .A(n4638), .Z(n5586) );
  CLKBUF_X1 U3904 ( .A(n3712), .Z(n3713) );
  INV_X1 U3905 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3208) );
  INV_X1 U3906 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4562) );
  NOR2_X1 U3907 ( .A1(n4594), .A2(n6028), .ZN(n6063) );
  NOR2_X1 U3908 ( .A1(n6030), .A2(n5586), .ZN(n6353) );
  NOR2_X1 U3909 ( .A1(n6240), .A2(n6202), .ZN(n6233) );
  OAI21_X1 U3910 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6609), .A(n6101), 
        .ZN(n6129) );
  AND2_X1 U3911 ( .A1(n4747), .A2(n6383), .ZN(n6360) );
  OR2_X1 U3912 ( .A1(n6607), .A2(n4636), .ZN(n4791) );
  INV_X1 U3913 ( .A(n6101), .ZN(n6208) );
  INV_X1 U3914 ( .A(n6129), .ZN(n6446) );
  AND2_X1 U3915 ( .A1(n4589), .A2(n4588), .ZN(n6532) );
  NAND2_X1 U3916 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n6530) );
  AND2_X1 U3917 ( .A1(n5133), .A2(n5138), .ZN(n5634) );
  AND2_X1 U3918 ( .A1(n4922), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5820) );
  INV_X1 U3919 ( .A(n5646), .ZN(n5810) );
  AND2_X1 U3920 ( .A1(n4841), .A2(n4449), .ZN(n4802) );
  AND2_X1 U3921 ( .A1(n4922), .A2(n4448), .ZN(n5821) );
  AND2_X1 U3922 ( .A1(n4447), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4448) );
  INV_X1 U3923 ( .A(n5140), .ZN(n4841) );
  INV_X1 U3924 ( .A(n5820), .ZN(n5794) );
  OR2_X1 U3925 ( .A1(n5286), .A2(n5285), .ZN(n5394) );
  INV_X1 U3926 ( .A(n5336), .ZN(n5836) );
  NAND2_X2 U3927 ( .A1(n4516), .A2(n4515), .ZN(n5840) );
  OR2_X1 U3928 ( .A1(n4607), .A2(n5126), .ZN(n4515) );
  OR2_X1 U3929 ( .A1(n5295), .A2(n5294), .ZN(n5658) );
  INV_X1 U3930 ( .A(n5653), .ZN(n5848) );
  AND2_X1 U3931 ( .A1(n5369), .A2(n5351), .ZN(n5847) );
  NOR2_X2 U3932 ( .A1(n5850), .A2(n5346), .ZN(n5851) );
  NAND2_X1 U3933 ( .A1(n5369), .A2(n4617), .ZN(n5371) );
  AOI21_X1 U3935 ( .B1(n5085), .B2(n4237), .A(n5084), .ZN(n5155) );
  INV_X1 U3936 ( .A(n5394), .ZN(n5654) );
  AND2_X1 U3937 ( .A1(n5100), .A2(n5080), .ZN(n5201) );
  AND2_X1 U3938 ( .A1(n5045), .A2(n5044), .ZN(n5832) );
  OR2_X1 U3939 ( .A1(n5168), .A2(n5167), .ZN(n5472) );
  AOI22_X1 U3940 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n3156), .B2(n5492), .ZN(n5377) );
  INV_X1 U3941 ( .A(n3187), .ZN(n3186) );
  CLKBUF_X1 U3942 ( .A(n5059), .Z(n5060) );
  NAND2_X1 U3943 ( .A1(n5414), .A2(n3189), .ZN(n5408) );
  INV_X1 U3944 ( .A(n5420), .ZN(n5422) );
  NAND2_X1 U3945 ( .A1(n3191), .A2(n3644), .ZN(n5439) );
  NAND2_X1 U3946 ( .A1(n3643), .A2(n3195), .ZN(n3191) );
  CLKBUF_X1 U3947 ( .A(n4961), .Z(n4962) );
  CLKBUF_X1 U3948 ( .A(n4963), .Z(n4964) );
  INV_X1 U3949 ( .A(n5708), .ZN(n5992) );
  AND2_X1 U3950 ( .A1(n6025), .A2(n4308), .ZN(n6004) );
  INV_X1 U3951 ( .A(n6018), .ZN(n6012) );
  AND2_X1 U3952 ( .A1(n3726), .A2(n3725), .ZN(n6614) );
  INV_X1 U3953 ( .A(n5586), .ZN(n6029) );
  NOR2_X2 U3954 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6612) );
  INV_X1 U3955 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6525) );
  INV_X1 U3956 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5117) );
  INV_X1 U3957 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5587) );
  INV_X1 U3958 ( .A(n6543), .ZN(n5590) );
  INV_X1 U3959 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5736) );
  NOR2_X1 U3960 ( .A1(n4870), .A2(n6361), .ZN(n4899) );
  NOR2_X2 U3961 ( .A1(n6240), .A2(n4728), .ZN(n6349) );
  OAI211_X1 U3962 ( .C1(n6426), .C2(n6609), .A(n6396), .B(n6395), .ZN(n6429)
         );
  OR2_X1 U3963 ( .A1(n6441), .A2(n6611), .ZN(n6497) );
  AND2_X1 U3964 ( .A1(n6384), .A2(n6033), .ZN(n6492) );
  INV_X1 U3965 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U3966 ( .A1(n5587), .A2(n6436), .ZN(n6555) );
  NAND2_X1 U3967 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4501), .ZN(n6543) );
  AND2_X1 U3968 ( .A1(n6540), .A2(n6539), .ZN(n6554) );
  INV_X1 U3969 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6609) );
  INV_X1 U3970 ( .A(n6554), .ZN(n6608) );
  AOI21_X1 U3971 ( .B1(n5345), .B2(n5910), .A(n4245), .ZN(n4246) );
  NAND2_X1 U3972 ( .A1(n4191), .A2(n5910), .ZN(n4201) );
  AND2_X1 U3973 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  OR2_X1 U3974 ( .A1(n4430), .A2(n3154), .ZN(n5177) );
  NOR2_X1 U3975 ( .A1(n4430), .A2(n5324), .ZN(n5320) );
  AND2_X1 U3976 ( .A1(n4955), .A2(n5935), .ZN(n3151) );
  OR2_X2 U3977 ( .A1(n5315), .A2(n4396), .ZN(n3152) );
  NAND2_X1 U3978 ( .A1(n3149), .A2(n4512), .ZN(n3353) );
  NOR2_X1 U3979 ( .A1(n4430), .A2(n3177), .ZN(n5309) );
  AND4_X1 U3980 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3153)
         );
  NAND2_X1 U3981 ( .A1(n4142), .A2(n3174), .ZN(n3154) );
  AND4_X1 U3982 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3155)
         );
  NAND2_X1 U3983 ( .A1(n3643), .A2(n3642), .ZN(n5446) );
  NOR3_X1 U3984 ( .A1(n5399), .A2(n5448), .A3(n5501), .ZN(n3156) );
  AND2_X2 U3985 ( .A1(n3213), .A2(n4555), .ZN(n3402) );
  OR2_X1 U3986 ( .A1(n6630), .A2(n4615), .ZN(n3157) );
  NAND2_X1 U3987 ( .A1(n3444), .A2(n3198), .ZN(n3487) );
  OR2_X1 U3988 ( .A1(n5448), .A2(n5706), .ZN(n3158) );
  NOR2_X1 U3989 ( .A1(n5177), .A2(n5178), .ZN(n4189) );
  NAND2_X1 U3990 ( .A1(n4824), .A2(n3182), .ZN(n4939) );
  INV_X1 U3991 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3661) );
  AND2_X1 U3992 ( .A1(n4824), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U3993 ( .A1(n3636), .A2(n3647), .ZN(n3159) );
  INV_X1 U3994 ( .A(n3190), .ZN(n3189) );
  NOR2_X1 U3995 ( .A1(n5065), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3190)
         );
  AND2_X1 U3996 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3160) );
  AND2_X1 U3997 ( .A1(n5065), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3161)
         );
  AND2_X1 U3998 ( .A1(n3182), .A2(n3834), .ZN(n3162) );
  AND2_X1 U3999 ( .A1(n3188), .A2(n3653), .ZN(n3163) );
  AND2_X1 U4000 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3164) );
  AND2_X2 U4001 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4557) );
  CLKBUF_X1 U4002 ( .A(n6182), .Z(n3165) );
  NAND2_X1 U4003 ( .A1(n3167), .A2(n3166), .ZN(n3457) );
  INV_X1 U4004 ( .A(n3456), .ZN(n3166) );
  NAND2_X1 U4005 ( .A1(n3348), .A2(n3164), .ZN(n3722) );
  NAND3_X1 U4006 ( .A1(n3169), .A2(n3364), .A3(n3361), .ZN(n3447) );
  NAND2_X1 U4007 ( .A1(n4189), .A2(n3170), .ZN(n3173) );
  NAND2_X1 U4008 ( .A1(n4189), .A2(n4190), .ZN(n4237) );
  INV_X1 U4009 ( .A(n3173), .ZN(n5084) );
  INV_X1 U4010 ( .A(n4240), .ZN(n3172) );
  NAND2_X1 U4011 ( .A1(n4824), .A2(n3162), .ZN(n4980) );
  NAND2_X1 U4012 ( .A1(n5413), .A2(n3188), .ZN(n5092) );
  NAND2_X1 U4013 ( .A1(n5413), .A2(n5415), .ZN(n5414) );
  OAI211_X1 U4014 ( .C1(n5413), .C2(n3186), .A(n3185), .B(n3183), .ZN(n5093)
         );
  NAND2_X1 U4015 ( .A1(n3184), .A2(n3187), .ZN(n3183) );
  NAND2_X1 U4016 ( .A1(n5413), .A2(n3163), .ZN(n3185) );
  NAND2_X1 U4017 ( .A1(n3197), .A2(n4955), .ZN(n3637) );
  NAND2_X1 U4018 ( .A1(n3197), .A2(n3151), .ZN(n5004) );
  NAND3_X1 U4019 ( .A1(n3444), .A2(n3443), .A3(n3198), .ZN(n3486) );
  NAND2_X1 U4020 ( .A1(n5428), .A2(n5063), .ZN(n5420) );
  NAND2_X1 U4021 ( .A1(n5427), .A2(n5062), .ZN(n5428) );
  NOR2_X1 U4022 ( .A1(n4249), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4255)
         );
  CLKBUF_X1 U4023 ( .A(n3367), .Z(n6508) );
  CLKBUF_X1 U4024 ( .A(n5373), .Z(n5383) );
  NAND2_X1 U4025 ( .A1(n5373), .A2(n4322), .ZN(n4251) );
  CLKBUF_X1 U4026 ( .A(n3716), .Z(n6027) );
  CLKBUF_X2 U4027 ( .A(n4218), .Z(n4146) );
  AOI22_X1 U4028 ( .A1(n4218), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3211) );
  INV_X1 U4029 ( .A(n5427), .ZN(n5431) );
  NAND2_X1 U4030 ( .A1(n4649), .A2(n3483), .ZN(n3491) );
  NAND2_X1 U4032 ( .A1(n3774), .A2(n3773), .ZN(n4825) );
  NAND2_X1 U4033 ( .A1(n4422), .A2(n4528), .ZN(n3523) );
  NOR2_X1 U4034 ( .A1(n4422), .A2(n6542), .ZN(n3470) );
  XNOR2_X1 U4035 ( .A(n3566), .B(n3587), .ZN(n3756) );
  NAND2_X1 U4036 ( .A1(n3545), .A2(n6383), .ZN(n3566) );
  AND2_X1 U4037 ( .A1(n3349), .A2(n4422), .ZN(n3350) );
  AND2_X1 U4038 ( .A1(n3349), .A2(n4528), .ZN(n3344) );
  INV_X1 U4039 ( .A(n3445), .ZN(n3449) );
  INV_X1 U4040 ( .A(n3282), .ZN(n3333) );
  NAND2_X1 U4041 ( .A1(n3636), .A2(n5064), .ZN(n3199) );
  OR2_X1 U4042 ( .A1(n5065), .A2(n5391), .ZN(n3200) );
  INV_X1 U4043 ( .A(n5428), .ZN(n5429) );
  OR2_X1 U4044 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6965), .ZN(n7026) );
  INV_X1 U4045 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5793) );
  INV_X1 U4046 ( .A(READY_N), .ZN(n6627) );
  OR2_X1 U4047 ( .A1(n6556), .A2(n6438), .ZN(n4644) );
  NOR2_X1 U4048 ( .A1(n4809), .A2(n4713), .ZN(n3201) );
  NOR2_X1 U4049 ( .A1(n5349), .A2(n6436), .ZN(n4239) );
  AND2_X1 U4050 ( .A1(n4340), .A2(n4618), .ZN(n3202) );
  NAND2_X1 U4051 ( .A1(n3377), .A2(n3492), .ZN(n3349) );
  INV_X1 U4052 ( .A(n3332), .ZN(n3377) );
  OR2_X2 U4053 ( .A1(n5252), .A2(n5251), .ZN(n3203) );
  AND2_X1 U4054 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3204) );
  NOR2_X4 U4055 ( .A1(n4605), .A2(n6538), .ZN(n3205) );
  INV_X1 U4056 ( .A(n3859), .ZN(n5041) );
  OR2_X1 U4057 ( .A1(n5146), .A2(n5145), .ZN(n3206) );
  NAND2_X1 U4058 ( .A1(n4512), .A2(n3492), .ZN(n3334) );
  NAND2_X1 U4059 ( .A1(n6517), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3667) );
  OAI21_X1 U4060 ( .B1(n4512), .B2(n3282), .A(n3334), .ZN(n3335) );
  BUF_X2 U4061 ( .A(n3403), .Z(n4171) );
  AND2_X1 U4062 ( .A1(n3676), .A2(n3677), .ZN(n3674) );
  NOR2_X1 U4063 ( .A1(n3491), .A2(n3492), .ZN(n3351) );
  OR2_X1 U4064 ( .A1(n4101), .A2(n4048), .ZN(n4092) );
  INV_X1 U4065 ( .A(n4431), .ZN(n3952) );
  INV_X1 U4066 ( .A(n4982), .ZN(n3834) );
  OR2_X1 U4067 ( .A1(n3600), .A2(n3599), .ZN(n3618) );
  INV_X1 U4068 ( .A(n3544), .ZN(n3545) );
  INV_X1 U4069 ( .A(n3473), .ZN(n3536) );
  INV_X1 U4070 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3207) );
  BUF_X4 U4071 ( .A(n4123), .Z(n4212) );
  AOI21_X1 U4072 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6525), .A(n3674), 
        .ZN(n3672) );
  NAND2_X1 U4073 ( .A1(n3340), .A2(n3483), .ZN(n4289) );
  INV_X1 U4074 ( .A(n4239), .ZN(n3732) );
  NAND2_X1 U4075 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4096)
         );
  INV_X1 U4076 ( .A(n3620), .ZN(n3631) );
  NAND2_X1 U4077 ( .A1(n3558), .A2(n3557), .ZN(n3587) );
  NAND2_X1 U4078 ( .A1(n3455), .A2(n3454), .ZN(n3456) );
  NAND2_X1 U4079 ( .A1(n3522), .A2(n3521), .ZN(n4584) );
  AND2_X1 U4080 ( .A1(n3327), .A2(n4528), .ZN(n3482) );
  INV_X1 U4081 ( .A(n4096), .ZN(n4075) );
  INV_X1 U4082 ( .A(n3758), .ZN(n4238) );
  NAND2_X1 U4083 ( .A1(n4164), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4206)
         );
  OR2_X1 U4084 ( .A1(n5079), .A2(n5213), .ZN(n5078) );
  INV_X1 U4085 ( .A(n3750), .ZN(n3751) );
  NAND2_X1 U4086 ( .A1(n4524), .A2(n4335), .ZN(n5121) );
  NAND2_X1 U4087 ( .A1(n4350), .A2(n4289), .ZN(n5127) );
  AND2_X1 U4088 ( .A1(n4297), .A2(n4296), .ZN(n4499) );
  AND2_X1 U4089 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3451) );
  AND2_X1 U4090 ( .A1(n4493), .A2(n4492), .ZN(n6515) );
  AND2_X1 U4091 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4075), .ZN(n4084)
         );
  INV_X1 U4092 ( .A(n3984), .ZN(n3985) );
  INV_X1 U4093 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5255) );
  INV_X1 U4094 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U4095 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4802), .ZN(n5272) );
  INV_X1 U4096 ( .A(n5790), .ZN(n5825) );
  BUF_X1 U4097 ( .A(n4289), .Z(n5119) );
  OR2_X1 U4098 ( .A1(n4140), .A2(n5101), .ZN(n5282) );
  AND2_X1 U4099 ( .A1(n4373), .A2(n4372), .ZN(n4992) );
  AND2_X1 U4100 ( .A1(n4499), .A2(n4300), .ZN(n4510) );
  INV_X1 U4101 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5627) );
  AOI21_X1 U4102 ( .B1(n3772), .B2(n3871), .A(n3771), .ZN(n5260) );
  NAND2_X1 U4103 ( .A1(n4251), .A2(n4316), .ZN(n4252) );
  NAND2_X1 U4104 ( .A1(n5448), .A2(n5375), .ZN(n3659) );
  AND2_X1 U4105 ( .A1(n4303), .A2(n6026), .ZN(n5011) );
  AND2_X1 U4106 ( .A1(n4256), .A2(n4257), .ZN(n4434) );
  INV_X1 U4107 ( .A(n6515), .ZN(n4578) );
  AND2_X1 U4108 ( .A1(n4874), .A2(n4873), .ZN(n4881) );
  AND2_X1 U4109 ( .A1(n4754), .A2(n4753), .ZN(n4793) );
  INV_X2 U4110 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U4111 ( .A1(n4543), .A2(n4466), .ZN(n6625) );
  AND2_X1 U4112 ( .A1(n5610), .A2(REIP_REG_24__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U4113 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4074)
         );
  AND2_X1 U4114 ( .A1(n5142), .A2(n4459), .ZN(n5790) );
  OR3_X1 U4115 ( .A1(n6625), .A2(n6541), .A3(n4437), .ZN(n4922) );
  INV_X1 U4116 ( .A(n5840), .ZN(n5341) );
  INV_X1 U4117 ( .A(n5369), .ZN(n5850) );
  NOR2_X1 U4118 ( .A1(n6530), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U4119 ( .A1(n4545), .A2(n3205), .ZN(n4665) );
  INV_X1 U4120 ( .A(n4708), .ZN(n4684) );
  AOI21_X1 U4121 ( .B1(n4005), .B2(n4004), .A(n4003), .ZN(n5310) );
  NAND2_X1 U4122 ( .A1(n3854), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3886)
         );
  INV_X1 U4123 ( .A(n5915), .ZN(n5888) );
  INV_X1 U4124 ( .A(n5918), .ZN(n5909) );
  OR2_X1 U4125 ( .A1(n5686), .A2(n4313), .ZN(n5494) );
  AND2_X1 U4126 ( .A1(n5326), .A2(n4456), .ZN(n5548) );
  OAI21_X1 U4127 ( .B1(n6025), .B2(n5014), .A(n5714), .ZN(n5722) );
  NOR2_X1 U4128 ( .A1(n5927), .A2(n6004), .ZN(n5998) );
  INV_X1 U4129 ( .A(n6009), .ZN(n6023) );
  NOR2_X1 U4130 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5113) );
  OAI221_X1 U4131 ( .B1(n6118), .B2(n6609), .C1(n6118), .C2(n6102), .A(n6285), 
        .ZN(n6120) );
  OAI21_X1 U4132 ( .B1(n4879), .B2(n4880), .A(n4878), .ZN(n4897) );
  NAND2_X1 U4133 ( .A1(n4752), .A2(n4751), .ZN(n4789) );
  INV_X1 U4134 ( .A(n6205), .ZN(n6229) );
  OAI21_X1 U4135 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6307) );
  INV_X1 U4136 ( .A(n6321), .ZN(n6306) );
  NAND2_X1 U4137 ( .A1(n4594), .A2(n6027), .ZN(n6240) );
  NOR2_X2 U4138 ( .A1(n6362), .A2(n6361), .ZN(n6427) );
  INV_X1 U4139 ( .A(n4236), .ZN(n4436) );
  INV_X1 U4140 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6575) );
  OR2_X1 U4141 ( .A1(n4605), .A2(n4284), .ZN(n4543) );
  INV_X1 U4142 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6793) );
  NAND2_X1 U4143 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4856), .ZN(n5802) );
  NAND2_X1 U4144 ( .A1(n4922), .A2(n4438), .ZN(n5646) );
  AND2_X1 U4145 ( .A1(n4800), .A2(n5646), .ZN(n5817) );
  NAND2_X1 U4146 ( .A1(n5840), .A2(n5344), .ZN(n5336) );
  INV_X1 U4147 ( .A(n5201), .ZN(n5365) );
  INV_X1 U4148 ( .A(n4988), .ZN(n4951) );
  OR3_X1 U4149 ( .A1(n4605), .A2(n4527), .A3(n6564), .ZN(n5885) );
  NAND2_X1 U4150 ( .A1(n4545), .A2(n4544), .ZN(n4708) );
  INV_X1 U4151 ( .A(n4199), .ZN(n4200) );
  OR2_X1 U4152 ( .A1(n5921), .A2(n4195), .ZN(n5915) );
  OR2_X1 U4153 ( .A1(n5068), .A2(n4321), .ZN(n5693) );
  OR2_X1 U4154 ( .A1(n4426), .A2(n4425), .ZN(n6009) );
  OR2_X1 U4155 ( .A1(n4197), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5721) );
  OR2_X1 U4156 ( .A1(n5931), .A2(n5977), .ZN(n5962) );
  OR2_X1 U4157 ( .A1(n4426), .A2(n6507), .ZN(n6025) );
  NAND2_X1 U4158 ( .A1(n6063), .A2(n6361), .ZN(n6090) );
  NAND2_X1 U4159 ( .A1(n6063), .A2(n6611), .ZN(n6123) );
  INV_X1 U4160 ( .A(n6119), .ZN(n4902) );
  INV_X1 U4161 ( .A(n4899), .ZN(n4798) );
  OR2_X1 U4162 ( .A1(n6124), .A2(n6611), .ZN(n6154) );
  OR2_X1 U4163 ( .A1(n4646), .A2(n6611), .ZN(n6201) );
  NAND2_X1 U4164 ( .A1(n6233), .A2(n6361), .ZN(n6280) );
  NAND2_X1 U4165 ( .A1(n6233), .A2(n6611), .ZN(n6311) );
  OR2_X1 U4166 ( .A1(n6240), .A2(n4721), .ZN(n6321) );
  NAND2_X1 U4167 ( .A1(n6360), .A2(n6361), .ZN(n6382) );
  INV_X1 U4168 ( .A(n6397), .ZN(n6451) );
  INV_X1 U4169 ( .A(n6413), .ZN(n6475) );
  AND3_X1 U4170 ( .A1(n6529), .A2(n6528), .A3(n6527), .ZN(n6547) );
  CLKBUF_X1 U4171 ( .A(n6600), .Z(n6596) );
  OR4_X1 U4172 ( .A1(n4465), .A2(n4464), .A3(n4463), .A4(n4462), .ZN(U2809) );
  OAI211_X1 U4173 ( .C1(n5481), .C2(n5918), .A(n4201), .B(n4200), .ZN(U2957)
         );
  AND2_X4 U4174 ( .A1(n5583), .A2(n3213), .ZN(n4145) );
  AND2_X2 U4175 ( .A1(n5583), .A2(n4556), .ZN(n3458) );
  AOI22_X1 U4176 ( .A1(n4145), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3212) );
  AND2_X2 U4177 ( .A1(n3661), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5582)
         );
  AND2_X4 U4178 ( .A1(n4557), .A2(n5582), .ZN(n4218) );
  AND2_X2 U4179 ( .A1(n4556), .A2(n4582), .ZN(n3408) );
  AND2_X2 U4180 ( .A1(n4556), .A2(n4555), .ZN(n3459) );
  AOI22_X1 U4181 ( .A1(n4220), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3210) );
  AND2_X2 U4182 ( .A1(n3213), .A2(n5582), .ZN(n3305) );
  AOI22_X1 U4183 ( .A1(n3402), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3209) );
  AND2_X2 U4184 ( .A1(n5582), .A2(n4560), .ZN(n3415) );
  AOI22_X1 U4185 ( .A1(n3314), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3217) );
  AND2_X2 U4186 ( .A1(n5583), .A2(n4557), .ZN(n3274) );
  AND2_X2 U4187 ( .A1(n4560), .A2(n4582), .ZN(n3416) );
  AOI22_X1 U4188 ( .A1(n3274), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3216) );
  AND2_X2 U4189 ( .A1(n5582), .A2(n4556), .ZN(n3387) );
  AND2_X2 U4190 ( .A1(n4582), .A2(n4557), .ZN(n3288) );
  AOI22_X1 U4191 ( .A1(n3387), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4192 ( .A1(n4123), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4193 ( .A1(n3458), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4194 ( .A1(n4145), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4195 ( .A1(n3402), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4196 ( .A1(n3305), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4197 ( .A1(n3387), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4198 ( .A1(n3274), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3225)
         );
  NAND2_X1 U4199 ( .A1(n3416), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4200 ( .A1(n3288), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4201 ( .A1(n4218), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3230)
         );
  NAND2_X1 U4202 ( .A1(n4220), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3229)
         );
  NAND2_X1 U4203 ( .A1(n3408), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4204 ( .A1(n3459), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4205 ( .A1(n3415), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4206 ( .A1(n3314), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4207 ( .A1(n4123), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3232)
         );
  NAND2_X1 U4208 ( .A1(n3403), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3231)
         );
  NAND2_X2 U4209 ( .A1(n3333), .A2(n3492), .ZN(n3368) );
  AOI22_X1 U4210 ( .A1(n3403), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4211 ( .A1(n4218), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4212 ( .A1(n3458), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4213 ( .A1(n4145), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4220), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4214 ( .A1(n3402), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4215 ( .A1(n3415), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4216 ( .A1(n3341), .A2(n3332), .ZN(n3260) );
  AOI22_X1 U4217 ( .A1(n3150), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4218 ( .A1(n4220), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4219 ( .A1(n3458), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4220 ( .A1(n3314), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4221 ( .A1(n4145), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4222 ( .A1(n3415), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4223 ( .A1(n4123), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4224 ( .A1(n3408), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4225 ( .A1(n4145), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4226 ( .A1(n3402), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4227 ( .A1(n4220), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4228 ( .A1(n4218), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4229 ( .A1(n4212), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4230 ( .A1(n3150), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4231 ( .A1(n3314), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3266) );
  BUF_X4 U4232 ( .A(n3387), .Z(n4211) );
  AOI22_X1 U4233 ( .A1(n4211), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4234 ( .A1(n3314), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4235 ( .A1(n3458), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4236 ( .A1(n4145), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4237 ( .A1(n4123), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3270) );
  NAND4_X1 U4238 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3280)
         );
  AOI22_X1 U4239 ( .A1(n4211), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4240 ( .A1(n3402), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4241 ( .A1(n3274), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4242 ( .A1(n4220), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3275) );
  NAND4_X1 U4243 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3279)
         );
  OR2_X2 U4244 ( .A1(n3280), .A2(n3279), .ZN(n3483) );
  INV_X1 U4245 ( .A(n3715), .ZN(n3330) );
  NAND2_X1 U4246 ( .A1(n4782), .A2(n3283), .ZN(n3343) );
  NAND2_X1 U4247 ( .A1(n4145), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4248 ( .A1(n3402), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4249 ( .A1(n3458), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U4250 ( .A1(n3415), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4251 ( .A1(n3387), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4252 ( .A1(n3314), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4253 ( .A1(n3416), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4254 ( .A1(n3288), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4255 ( .A1(n3305), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4256 ( .A1(n4218), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4257 ( .A1(n3408), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4258 ( .A1(n3150), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3300)
         );
  NAND2_X1 U4259 ( .A1(n4123), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3299)
         );
  NAND2_X1 U4260 ( .A1(n3403), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3298)
         );
  NAND2_X1 U4261 ( .A1(n3459), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3297) );
  NAND4_X4 U4262 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3340)
         );
  INV_X1 U4263 ( .A(n3340), .ZN(n3327) );
  NAND2_X1 U4264 ( .A1(n3458), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4265 ( .A1(n4145), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4266 ( .A1(n3402), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4267 ( .A1(n3305), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4268 ( .A1(n3387), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4269 ( .A1(n3150), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3312)
         );
  NAND2_X1 U4270 ( .A1(n3416), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4271 ( .A1(n3288), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3310)
         );
  AND4_X2 U4272 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3325)
         );
  NAND2_X1 U4273 ( .A1(n3415), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4274 ( .A1(n3314), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4275 ( .A1(n4218), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3322)
         );
  NAND2_X1 U4276 ( .A1(n4220), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3321)
         );
  NAND2_X1 U4277 ( .A1(n3408), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4278 ( .A1(n3459), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3319) );
  NAND4_X4 U4279 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n4528)
         );
  NAND2_X1 U4280 ( .A1(n3343), .A2(n3482), .ZN(n3329) );
  INV_X1 U4281 ( .A(n4289), .ZN(n3328) );
  NAND2_X1 U4282 ( .A1(n3329), .A2(n4496), .ZN(n3383) );
  NOR2_X1 U4283 ( .A1(n3330), .A2(n3383), .ZN(n3347) );
  INV_X1 U4284 ( .A(n3357), .ZN(n5344) );
  INV_X1 U4285 ( .A(n3349), .ZN(n3331) );
  NAND2_X1 U4286 ( .A1(n3331), .A2(n3357), .ZN(n3712) );
  OAI21_X1 U4287 ( .B1(n5344), .B2(n3483), .A(n3712), .ZN(n3337) );
  NAND2_X1 U4288 ( .A1(n3335), .A2(n4649), .ZN(n3336) );
  NAND2_X1 U4289 ( .A1(n3337), .A2(n3336), .ZN(n3352) );
  NAND2_X1 U4290 ( .A1(n3353), .A2(n4291), .ZN(n3338) );
  NAND2_X1 U4291 ( .A1(n3338), .A2(n4733), .ZN(n3339) );
  XNOR2_X1 U4292 ( .A(n6575), .B(STATE_REG_1__SCAN_IN), .ZN(n4261) );
  NOR2_X1 U4293 ( .A1(n3340), .A2(n4261), .ZN(n3358) );
  INV_X1 U4294 ( .A(n3358), .ZN(n3342) );
  NAND2_X1 U4295 ( .A1(n3342), .A2(n5350), .ZN(n3345) );
  NAND3_X1 U4296 ( .A1(n3347), .A2(n3370), .A3(n3346), .ZN(n3348) );
  NAND2_X1 U4297 ( .A1(n4273), .A2(n4528), .ZN(n4283) );
  INV_X1 U4298 ( .A(n3352), .ZN(n4256) );
  INV_X1 U4299 ( .A(n4528), .ZN(n3354) );
  NOR2_X1 U4300 ( .A1(n3353), .A2(n3380), .ZN(n3355) );
  NOR2_X1 U4301 ( .A1(n3483), .A2(n3492), .ZN(n3356) );
  AND2_X1 U4302 ( .A1(n4649), .A2(n3356), .ZN(n4514) );
  AND2_X1 U4303 ( .A1(n5349), .A2(n4512), .ZN(n4276) );
  OAI211_X1 U4304 ( .C1(n4283), .C2(n3358), .A(n4285), .B(n4423), .ZN(n3359)
         );
  NAND2_X1 U4305 ( .A1(n3359), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4306 ( .A1(n5113), .A2(n6542), .ZN(n4197) );
  INV_X1 U4307 ( .A(n4197), .ZN(n3520) );
  XNOR2_X1 U4308 ( .A(n6619), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6385)
         );
  INV_X1 U4309 ( .A(n3711), .ZN(n3519) );
  AND2_X1 U4310 ( .A1(n3519), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3360)
         );
  AOI21_X1 U4311 ( .B1(n3520), .B2(n6385), .A(n3360), .ZN(n3361) );
  INV_X1 U4312 ( .A(n3361), .ZN(n3362) );
  NOR2_X1 U4313 ( .A1(n3362), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3363)
         );
  INV_X1 U4314 ( .A(n3365), .ZN(n3366) );
  NAND2_X1 U4315 ( .A1(n3722), .A2(n3723), .ZN(n3386) );
  NOR2_X1 U4316 ( .A1(n3368), .A2(n4733), .ZN(n3369) );
  NAND2_X1 U4317 ( .A1(n4291), .A2(n4528), .ZN(n3371) );
  INV_X1 U4318 ( .A(n3375), .ZN(n3376) );
  NAND2_X1 U4319 ( .A1(n3376), .A2(n4544), .ZN(n3385) );
  AND2_X1 U4320 ( .A1(n4653), .A2(n4422), .ZN(n3379) );
  NOR2_X1 U4321 ( .A1(n4267), .A2(n3483), .ZN(n3378) );
  NAND4_X1 U4322 ( .A1(n3379), .A2(n4790), .A3(n3378), .A4(n5349), .ZN(n4571)
         );
  AND2_X1 U4323 ( .A1(n5113), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6549) );
  INV_X1 U4324 ( .A(n3483), .ZN(n4738) );
  NAND2_X1 U4325 ( .A1(n4608), .A2(n4738), .ZN(n3381) );
  NAND3_X1 U4326 ( .A1(n4571), .A2(n6549), .A3(n3381), .ZN(n3382) );
  NOR2_X1 U4327 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  NAND3_X1 U4328 ( .A1(n4297), .A2(n3385), .A3(n3384), .ZN(n3721) );
  XNOR2_X1 U4329 ( .A(n3445), .B(n3446), .ZN(n4638) );
  NAND2_X1 U4330 ( .A1(n4638), .A2(n6542), .ZN(n3401) );
  AOI22_X1 U4331 ( .A1(n4016), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4332 ( .A1(n3458), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4333 ( .A1(n4208), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4334 ( .A1(n4212), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3389) );
  NAND4_X1 U4335 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), .ZN(n3399)
         );
  AOI22_X1 U4336 ( .A1(n4563), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4337 ( .A1(n4117), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4338 ( .A1(n4145), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3395) );
  BUF_X1 U4339 ( .A(n3288), .Z(n4122) );
  AOI22_X1 U4340 ( .A1(n7031), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3394) );
  NAND4_X1 U4341 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3398)
         );
  NAND2_X1 U4342 ( .A1(n3470), .A2(n3490), .ZN(n3400) );
  NAND2_X1 U4343 ( .A1(n3401), .A2(n3400), .ZN(n3439) );
  AOI22_X1 U4344 ( .A1(n3314), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4345 ( .A1(n4117), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4346 ( .A1(n3150), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4347 ( .A1(n4212), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4348 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3414)
         );
  AOI22_X1 U4349 ( .A1(n3458), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4350 ( .A1(n4211), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4351 ( .A1(n4145), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4352 ( .A1(n4146), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3409) );
  NAND4_X1 U4353 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3413)
         );
  NAND2_X1 U4354 ( .A1(n3470), .A2(n3631), .ZN(n3440) );
  AOI22_X1 U4355 ( .A1(n3150), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4356 ( .A1(n4145), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4357 ( .A1(n4208), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4358 ( .A1(n3388), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3417) );
  NAND4_X1 U4359 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3426)
         );
  AOI22_X1 U4360 ( .A1(n3458), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4361 ( .A1(n4117), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4362 ( .A1(n4146), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4363 ( .A1(n3314), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4364 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3425)
         );
  NAND2_X1 U4365 ( .A1(n3427), .A2(n3628), .ZN(n3428) );
  NAND2_X1 U4366 ( .A1(n3723), .A2(n6542), .ZN(n3430) );
  NAND2_X1 U4367 ( .A1(n3500), .A2(n3430), .ZN(n3501) );
  INV_X1 U4368 ( .A(n3523), .ZN(n3431) );
  NAND2_X1 U4369 ( .A1(n3702), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4370 ( .A1(n4653), .A2(n3504), .ZN(n3432) );
  OAI211_X1 U4371 ( .C1(n3631), .C2(n4422), .A(STATE2_REG_0__SCAN_IN), .B(
        n3432), .ZN(n3433) );
  INV_X1 U4372 ( .A(n3433), .ZN(n3434) );
  NAND2_X1 U4373 ( .A1(n3435), .A2(n3434), .ZN(n3498) );
  NAND2_X1 U4374 ( .A1(n3501), .A2(n3498), .ZN(n3437) );
  INV_X1 U4375 ( .A(n3628), .ZN(n3436) );
  NAND2_X1 U4376 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  INV_X1 U4377 ( .A(n3490), .ZN(n3442) );
  NAND2_X1 U4378 ( .A1(n4653), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U4379 ( .A1(n3702), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3441) );
  OAI211_X1 U4380 ( .C1(n3442), .C2(n3472), .A(n3441), .B(n3440), .ZN(n3488)
         );
  INV_X1 U4381 ( .A(n3488), .ZN(n3443) );
  AND2_X2 U4382 ( .A1(n3486), .A2(n3444), .ZN(n3477) );
  INV_X1 U4383 ( .A(n3446), .ZN(n3726) );
  NAND2_X1 U4384 ( .A1(n3451), .A2(n6517), .ZN(n4872) );
  INV_X1 U4385 ( .A(n3451), .ZN(n3452) );
  NAND2_X1 U4386 ( .A1(n3452), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3453) );
  NAND2_X1 U4387 ( .A1(n4872), .A2(n3453), .ZN(n6155) );
  AOI22_X1 U4388 ( .A1(n3520), .A2(n6155), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3519), .ZN(n3454) );
  NAND2_X1 U4389 ( .A1(n4585), .A2(n3457), .ZN(n4570) );
  AOI22_X1 U4390 ( .A1(n4145), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4391 ( .A1(n4563), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4392 ( .A1(n4117), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4393 ( .A1(n4146), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3460) );
  NAND4_X1 U4394 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3469)
         );
  AOI22_X1 U4395 ( .A1(n4016), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4396 ( .A1(n7031), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4397 ( .A1(n4116), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4398 ( .A1(n4212), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U4399 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3468)
         );
  INV_X1 U4400 ( .A(n3470), .ZN(n3471) );
  INV_X1 U4401 ( .A(n3472), .ZN(n3474) );
  AOI22_X1 U4402 ( .A1(n3702), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3474), 
        .B2(n3473), .ZN(n3475) );
  INV_X1 U4403 ( .A(n3477), .ZN(n3480) );
  INV_X1 U4404 ( .A(n3478), .ZN(n3479) );
  NAND2_X1 U4405 ( .A1(n3480), .A2(n3479), .ZN(n3481) );
  NAND2_X1 U4406 ( .A1(n3544), .A2(n3481), .ZN(n3716) );
  NAND2_X1 U4407 ( .A1(n3504), .A2(n3490), .ZN(n3537) );
  XNOR2_X1 U4408 ( .A(n3537), .B(n3536), .ZN(n3484) );
  AND2_X1 U4409 ( .A1(n4653), .A2(n3483), .ZN(n3502) );
  AOI21_X1 U4410 ( .B1(n3484), .B2(n4443), .A(n3502), .ZN(n3485) );
  OAI21_X2 U4411 ( .B1(n3716), .B2(n3669), .A(n3485), .ZN(n5908) );
  NAND2_X1 U4412 ( .A1(n5908), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3513)
         );
  NAND2_X1 U4413 ( .A1(n3487), .A2(n3488), .ZN(n3489) );
  NAND2_X1 U4414 ( .A1(n4593), .A2(n4544), .ZN(n3497) );
  XNOR2_X1 U4415 ( .A(n3504), .B(n3490), .ZN(n3494) );
  INV_X1 U4416 ( .A(n3491), .ZN(n3493) );
  OAI211_X1 U4417 ( .C1(n3494), .C2(n6630), .A(n3493), .B(n3492), .ZN(n3495)
         );
  INV_X1 U4418 ( .A(n3495), .ZN(n3496) );
  NAND2_X1 U4419 ( .A1(n3497), .A2(n3496), .ZN(n4904) );
  INV_X1 U4420 ( .A(n3498), .ZN(n3499) );
  NAND2_X1 U4421 ( .A1(n6611), .A2(n3627), .ZN(n3507) );
  INV_X1 U4422 ( .A(n3502), .ZN(n3503) );
  OAI21_X1 U4423 ( .B1(n6630), .B2(n3504), .A(n3503), .ZN(n3505) );
  INV_X1 U4424 ( .A(n3505), .ZN(n3506) );
  NAND2_X1 U4425 ( .A1(n3507), .A2(n3506), .ZN(n5916) );
  NAND2_X1 U4426 ( .A1(n5916), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3508)
         );
  INV_X1 U4427 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U4428 ( .A1(n3508), .A2(n6015), .ZN(n3510) );
  AND2_X1 U4429 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4430 ( .A1(n5916), .A2(n3509), .ZN(n3511) );
  AND2_X1 U4431 ( .A1(n3510), .A2(n3511), .ZN(n4903) );
  INV_X1 U4432 ( .A(n3511), .ZN(n3512) );
  NAND2_X1 U4433 ( .A1(n3513), .A2(n5906), .ZN(n3516) );
  INV_X1 U4434 ( .A(n5908), .ZN(n3514) );
  INV_X1 U4435 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U4436 ( .A1(n3514), .A2(n5997), .ZN(n3515) );
  AND2_X1 U4437 ( .A1(n3516), .A2(n3515), .ZN(n5898) );
  NAND3_X1 U4438 ( .A1(n6525), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6159) );
  INV_X1 U4439 ( .A(n6159), .ZN(n3517) );
  NAND2_X1 U4440 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3517), .ZN(n6187) );
  NAND2_X1 U4441 ( .A1(n6525), .A2(n6187), .ZN(n3518) );
  NAND3_X1 U4442 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6437) );
  INV_X1 U4443 ( .A(n6437), .ZN(n6447) );
  NAND2_X1 U4444 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6447), .ZN(n6433) );
  AOI22_X1 U4445 ( .A1(n3520), .A2(n6203), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3519), .ZN(n3521) );
  AOI22_X1 U4446 ( .A1(n4016), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4447 ( .A1(n4117), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4448 ( .A1(n4208), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4449 ( .A1(n4116), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3524) );
  NAND4_X1 U4450 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n3533)
         );
  AOI22_X1 U4451 ( .A1(n4145), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4452 ( .A1(n7031), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4453 ( .A1(n4219), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4454 ( .A1(n4563), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3528) );
  NAND4_X1 U4455 ( .A1(n3531), .A2(n3530), .A3(n3529), .A4(n3528), .ZN(n3532)
         );
  AOI22_X1 U4456 ( .A1(n3702), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3707), 
        .B2(n3559), .ZN(n3534) );
  XNOR2_X1 U4457 ( .A(n3544), .B(n6383), .ZN(n3738) );
  NAND2_X1 U4458 ( .A1(n3738), .A2(n3627), .ZN(n3541) );
  NAND2_X1 U4459 ( .A1(n3537), .A2(n3536), .ZN(n3560) );
  INV_X1 U4460 ( .A(n3559), .ZN(n3538) );
  XNOR2_X1 U4461 ( .A(n3560), .B(n3538), .ZN(n3539) );
  NAND2_X1 U4462 ( .A1(n3539), .A2(n4443), .ZN(n3540) );
  INV_X1 U4463 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U4464 ( .A1(n5898), .A2(n5900), .ZN(n5899) );
  NAND2_X1 U4465 ( .A1(n3542), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3543)
         );
  NAND2_X1 U4466 ( .A1(n5899), .A2(n3543), .ZN(n4961) );
  INV_X1 U4467 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3546) );
  OR2_X1 U4468 ( .A1(n3670), .A2(n3546), .ZN(n3558) );
  AOI22_X1 U4469 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4563), .B1(n4219), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4470 ( .A1(n4016), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4471 ( .A1(n4116), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4472 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4146), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4473 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3556)
         );
  AOI22_X1 U4474 ( .A1(n4060), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4475 ( .A1(n7031), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4476 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4117), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4477 ( .A1(n4212), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4478 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  NAND2_X1 U4479 ( .A1(n3707), .A2(n3605), .ZN(n3557) );
  NAND2_X1 U4480 ( .A1(n3756), .A2(n3627), .ZN(n3563) );
  NAND2_X1 U4481 ( .A1(n3560), .A2(n3559), .ZN(n3608) );
  XNOR2_X1 U4482 ( .A(n3608), .B(n3605), .ZN(n3561) );
  NAND2_X1 U4483 ( .A1(n3561), .A2(n4443), .ZN(n3562) );
  INV_X1 U4484 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U4485 ( .A(n3564), .B(n5981), .ZN(n4965) );
  NAND2_X1 U4486 ( .A1(n4961), .A2(n4965), .ZN(n4963) );
  NAND2_X1 U4487 ( .A1(n3564), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3565)
         );
  NAND2_X1 U4488 ( .A1(n4963), .A2(n3565), .ZN(n4913) );
  NAND2_X1 U4489 ( .A1(n3590), .A2(n3587), .ZN(n3579) );
  NAND2_X1 U4490 ( .A1(n3702), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4491 ( .A1(n4060), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4492 ( .A1(n4563), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4493 ( .A1(n4117), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4494 ( .A1(n4146), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4495 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3576)
         );
  AOI22_X1 U4496 ( .A1(n4016), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4497 ( .A1(n7031), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4498 ( .A1(n4116), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4499 ( .A1(n4212), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3571) );
  NAND4_X1 U4500 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n3575)
         );
  NAND2_X1 U4501 ( .A1(n3707), .A2(n3606), .ZN(n3577) );
  NAND2_X1 U4502 ( .A1(n3578), .A2(n3577), .ZN(n3588) );
  XNOR2_X1 U4503 ( .A(n3579), .B(n3588), .ZN(n3757) );
  NAND2_X1 U4504 ( .A1(n3757), .A2(n3627), .ZN(n3584) );
  INV_X1 U4505 ( .A(n3605), .ZN(n3580) );
  OR2_X1 U4506 ( .A1(n3608), .A2(n3580), .ZN(n3581) );
  XNOR2_X1 U4507 ( .A(n3581), .B(n3606), .ZN(n3582) );
  NAND2_X1 U4508 ( .A1(n3582), .A2(n4443), .ZN(n3583) );
  NAND2_X1 U4509 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  INV_X1 U4510 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U4511 ( .A(n3585), .B(n5963), .ZN(n4912) );
  NAND2_X1 U4512 ( .A1(n3585), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3586)
         );
  NAND2_X1 U4513 ( .A1(n4911), .A2(n3586), .ZN(n4816) );
  NAND2_X1 U4514 ( .A1(n3702), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4515 ( .A1(n4060), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4516 ( .A1(n4563), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4517 ( .A1(n4117), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4518 ( .A1(n4146), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3591) );
  NAND4_X1 U4519 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3600)
         );
  AOI22_X1 U4520 ( .A1(n4016), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4521 ( .A1(n7031), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4522 ( .A1(n4116), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4523 ( .A1(n4212), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4524 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  NAND2_X1 U4525 ( .A1(n3707), .A2(n3618), .ZN(n3601) );
  NAND2_X1 U4526 ( .A1(n3604), .A2(n3603), .ZN(n3772) );
  NAND3_X1 U4527 ( .A1(n3630), .A2(n3772), .A3(n3627), .ZN(n3611) );
  NAND2_X1 U4528 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  OR2_X1 U4529 ( .A1(n3608), .A2(n3607), .ZN(n3617) );
  XNOR2_X1 U4530 ( .A(n3617), .B(n3618), .ZN(n3609) );
  NAND2_X1 U4531 ( .A1(n3609), .A2(n4443), .ZN(n3610) );
  NAND2_X1 U4532 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  INV_X1 U4533 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4819) );
  XNOR2_X1 U4534 ( .A(n3612), .B(n4819), .ZN(n4815) );
  NAND2_X1 U4535 ( .A1(n4816), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U4536 ( .A1(n3612), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3613)
         );
  NAND2_X1 U4537 ( .A1(n4814), .A2(n3613), .ZN(n5457) );
  INV_X1 U4538 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4539 ( .A1(n3707), .A2(n3620), .ZN(n3614) );
  OAI21_X1 U4540 ( .B1(n3670), .B2(n3615), .A(n3614), .ZN(n3616) );
  NAND2_X1 U4541 ( .A1(n3766), .A2(n3627), .ZN(n3623) );
  INV_X1 U4542 ( .A(n3617), .ZN(n3619) );
  NAND2_X1 U4543 ( .A1(n3619), .A2(n3618), .ZN(n3632) );
  XNOR2_X1 U4544 ( .A(n3632), .B(n3620), .ZN(n3621) );
  NAND2_X1 U4545 ( .A1(n3621), .A2(n4443), .ZN(n3622) );
  NAND2_X1 U4546 ( .A1(n3623), .A2(n3622), .ZN(n3625) );
  INV_X1 U4547 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3624) );
  XNOR2_X1 U4548 ( .A(n3625), .B(n3624), .ZN(n5456) );
  NAND2_X1 U4549 ( .A1(n5457), .A2(n5456), .ZN(n5455) );
  NAND2_X1 U4550 ( .A1(n3625), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3626)
         );
  NAND2_X1 U4551 ( .A1(n5455), .A2(n3626), .ZN(n4974) );
  OR3_X1 U4552 ( .A1(n3632), .A2(n3631), .A3(n6630), .ZN(n3633) );
  NAND2_X1 U4553 ( .A1(n3636), .A2(n3633), .ZN(n3634) );
  INV_X1 U4554 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4361) );
  XNOR2_X1 U4555 ( .A(n3634), .B(n4361), .ZN(n4973) );
  NAND2_X1 U4556 ( .A1(n4974), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U4557 ( .A1(n3634), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3635)
         );
  NAND2_X1 U4558 ( .A1(n4972), .A2(n3635), .ZN(n4957) );
  INV_X1 U4559 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U4560 ( .A1(n3636), .A2(n5943), .ZN(n4954) );
  OR2_X1 U4561 ( .A1(n3636), .A2(n5943), .ZN(n4955) );
  NAND2_X1 U4562 ( .A1(n3637), .A2(n3204), .ZN(n3638) );
  NAND2_X1 U4563 ( .A1(n3639), .A2(n3638), .ZN(n5022) );
  INV_X1 U4564 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3640) );
  NOR2_X1 U4565 ( .A1(n5448), .A2(n3640), .ZN(n5020) );
  NAND2_X1 U4566 ( .A1(n3636), .A2(n3640), .ZN(n5018) );
  OAI21_X2 U4567 ( .B1(n5022), .B2(n5020), .A(n5018), .ZN(n5682) );
  XNOR2_X1 U4568 ( .A(n5448), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5683)
         );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4570 ( .A1(n5448), .A2(n3641), .ZN(n3642) );
  INV_X1 U4571 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5447) );
  AND2_X1 U4572 ( .A1(n3636), .A2(n5447), .ZN(n3645) );
  NAND2_X1 U4573 ( .A1(n5065), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3644) );
  INV_X1 U4574 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U4575 ( .A1(n5448), .A2(n5706), .ZN(n3646) );
  AND2_X1 U4576 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U4577 ( .A1(n5538), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3647) );
  NAND2_X1 U4578 ( .A1(n3648), .A2(n3159), .ZN(n5059) );
  INV_X1 U4579 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5560) );
  INV_X1 U4580 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5569) );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5551) );
  NAND3_X1 U4582 ( .A1(n5560), .A2(n5569), .A3(n5551), .ZN(n3649) );
  NAND2_X1 U4583 ( .A1(n5065), .A2(n3649), .ZN(n3650) );
  AND2_X1 U4584 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5512) );
  AND2_X1 U4585 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4309) );
  AND2_X1 U4586 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5540) );
  NAND3_X1 U4587 ( .A1(n5512), .A2(n4309), .A3(n5540), .ZN(n3651) );
  NAND2_X1 U4588 ( .A1(n5448), .A2(n3651), .ZN(n3652) );
  NAND2_X1 U4589 ( .A1(n5427), .A2(n3652), .ZN(n3656) );
  NOR2_X1 U4590 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5539) );
  NOR2_X1 U4591 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5511) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3653) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5096) );
  NAND4_X1 U4594 ( .A1(n5539), .A2(n5511), .A3(n3653), .A4(n5096), .ZN(n3654)
         );
  NAND2_X1 U4595 ( .A1(n5065), .A2(n3654), .ZN(n3655) );
  NAND2_X1 U4596 ( .A1(n3656), .A2(n3655), .ZN(n5374) );
  INV_X1 U4597 ( .A(n5374), .ZN(n3658) );
  INV_X1 U4598 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5375) );
  XNOR2_X1 U4599 ( .A(n5448), .B(n5375), .ZN(n5401) );
  INV_X1 U4600 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5391) );
  AND2_X1 U4601 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4322) );
  NOR4_X1 U4602 ( .A1(n5448), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A4(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n4203) );
  NAND2_X1 U4603 ( .A1(n5393), .A2(n4203), .ZN(n4250) );
  NAND2_X1 U4604 ( .A1(n4251), .A2(n4250), .ZN(n3660) );
  XNOR2_X1 U4605 ( .A(n3660), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5481)
         );
  NAND2_X1 U4606 ( .A1(n6512), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4607 ( .A1(n3661), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4608 ( .A1(n3663), .A2(n3662), .ZN(n3681) );
  NAND2_X1 U4609 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6619), .ZN(n3682) );
  NAND2_X1 U4610 ( .A1(n3664), .A2(n3663), .ZN(n3694) );
  NAND2_X1 U4611 ( .A1(n5117), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4612 ( .A1(n3667), .A2(n3665), .ZN(n3693) );
  INV_X1 U4613 ( .A(n3693), .ZN(n3666) );
  NAND2_X1 U4614 ( .A1(n3694), .A2(n3666), .ZN(n3668) );
  NAND2_X1 U4615 ( .A1(n3668), .A2(n3667), .ZN(n3676) );
  AOI222_X1 U4616 ( .A1(n3672), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3672), .B2(n5736), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n5736), 
        .ZN(n4264) );
  OR2_X2 U4617 ( .A1(n3670), .A2(n3669), .ZN(n3705) );
  INV_X1 U4618 ( .A(n3705), .ZN(n3671) );
  NAND2_X1 U4619 ( .A1(n4264), .A2(n3671), .ZN(n3710) );
  AND2_X1 U4620 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3672), .ZN(n3673)
         );
  INV_X1 U4621 ( .A(n3674), .ZN(n3675) );
  OAI21_X1 U4622 ( .B1(n3677), .B2(n3676), .A(n3675), .ZN(n3678) );
  AOI21_X1 U4623 ( .B1(n3707), .B2(n4544), .A(n5350), .ZN(n3690) );
  INV_X1 U4624 ( .A(n3682), .ZN(n3680) );
  XNOR2_X1 U4625 ( .A(n3681), .B(n3680), .ZN(n4262) );
  NAND2_X1 U4626 ( .A1(n4262), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3689) );
  AOI21_X1 U4627 ( .B1(n5350), .B2(n4528), .A(n4544), .ZN(n3697) );
  OAI21_X1 U4628 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6619), .A(n3682), 
        .ZN(n3684) );
  INV_X1 U4629 ( .A(n3684), .ZN(n3683) );
  AOI21_X1 U4630 ( .B1(n3368), .B2(n3683), .A(n4653), .ZN(n3687) );
  INV_X1 U4631 ( .A(n3707), .ZN(n3685) );
  OAI21_X1 U4632 ( .B1(n3685), .B2(n3684), .A(n3705), .ZN(n3686) );
  OAI21_X1 U4633 ( .B1(n3697), .B2(n3687), .A(n3686), .ZN(n3688) );
  AOI21_X1 U4634 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3692) );
  AOI22_X1 U4635 ( .A1(n3690), .A2(n4262), .B1(n3705), .B2(n3689), .ZN(n3691)
         );
  INV_X1 U4636 ( .A(n3696), .ZN(n3700) );
  XNOR2_X1 U4637 ( .A(n3694), .B(n3693), .ZN(n4263) );
  INV_X1 U4638 ( .A(n4263), .ZN(n3695) );
  AOI21_X1 U4639 ( .B1(n3702), .B2(n3695), .A(n3697), .ZN(n3699) );
  OAI211_X1 U4640 ( .C1(n3697), .C2(n3696), .A(n3707), .B(n4263), .ZN(n3698)
         );
  OAI21_X1 U4641 ( .B1(n3700), .B2(n3699), .A(n3698), .ZN(n3701) );
  OAI21_X1 U4642 ( .B1(n3702), .B2(n4265), .A(n3701), .ZN(n3704) );
  NAND2_X1 U4643 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6542), .ZN(n3703) );
  OAI211_X1 U4644 ( .C1(n4265), .C2(n3705), .A(n3704), .B(n3703), .ZN(n3706)
         );
  AOI21_X1 U4645 ( .B1(n3707), .B2(n4264), .A(n3706), .ZN(n3708) );
  INV_X1 U4646 ( .A(n3708), .ZN(n3709) );
  NAND2_X4 U4647 ( .A1(n3710), .A2(n3709), .ZN(n4501) );
  NAND2_X1 U4648 ( .A1(n3713), .A2(n4653), .ZN(n3714) );
  NAND2_X1 U4649 ( .A1(n3715), .A2(n3714), .ZN(n4282) );
  NAND2_X1 U4650 ( .A1(n6436), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3758) );
  NAND2_X1 U4651 ( .A1(n4593), .A2(n3871), .ZN(n3720) );
  AOI22_X1 U4652 ( .A1(n4239), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6436), .ZN(n3718) );
  AND2_X1 U4653 ( .A1(n4276), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4654 ( .A1(n3747), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3717) );
  AND2_X1 U4655 ( .A1(n3718), .A2(n3717), .ZN(n3719) );
  NAND2_X1 U4656 ( .A1(n3720), .A2(n3719), .ZN(n4520) );
  INV_X1 U4657 ( .A(n3721), .ZN(n3724) );
  NAND3_X1 U4658 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3725) );
  NAND2_X1 U4659 ( .A1(n6614), .A2(n3871), .ZN(n3730) );
  AOI22_X1 U4660 ( .A1(n4239), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6436), .ZN(n3728) );
  NAND2_X1 U4661 ( .A1(n3747), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3727) );
  AND2_X1 U4662 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  NAND2_X1 U4663 ( .A1(n3730), .A2(n3729), .ZN(n4507) );
  AOI21_X1 U4664 ( .B1(n6361), .B2(n4790), .A(n6436), .ZN(n4506) );
  NAND2_X1 U4665 ( .A1(n4507), .A2(n4506), .ZN(n4509) );
  OR2_X1 U4666 ( .A1(n4507), .A2(n4236), .ZN(n3731) );
  NAND2_X1 U4667 ( .A1(n4509), .A2(n3731), .ZN(n4519) );
  INV_X1 U4668 ( .A(n3747), .ZN(n3743) );
  NAND2_X1 U4669 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3739) );
  OAI21_X1 U4670 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3739), .ZN(n5914) );
  AOI22_X1 U4671 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4436), 
        .B2(n5914), .ZN(n3734) );
  NAND2_X1 U4672 ( .A1(n4186), .A2(EAX_REG_2__SCAN_IN), .ZN(n3733) );
  OAI211_X1 U4673 ( .C1(n3743), .C2(n5117), .A(n3734), .B(n3733), .ZN(n4601)
         );
  NAND2_X1 U4674 ( .A1(n4602), .A2(n4601), .ZN(n3737) );
  NAND2_X1 U4675 ( .A1(n3735), .A2(n4522), .ZN(n3736) );
  NAND2_X1 U4676 ( .A1(n3737), .A2(n3736), .ZN(n4600) );
  NAND2_X1 U4677 ( .A1(n4594), .A2(n3871), .ZN(n3746) );
  NAND2_X1 U4678 ( .A1(n3740), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3750)
         );
  OAI21_X1 U4679 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3740), .A(n3750), 
        .ZN(n5905) );
  AOI22_X1 U4680 ( .A1(n4436), .A2(n5905), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4681 ( .A1(n4186), .A2(EAX_REG_3__SCAN_IN), .ZN(n3741) );
  OAI211_X1 U4682 ( .C1(n3743), .C2(n4562), .A(n3742), .B(n3741), .ZN(n3744)
         );
  INV_X1 U4683 ( .A(n3744), .ZN(n3745) );
  NAND2_X1 U4684 ( .A1(n3746), .A2(n3745), .ZN(n4624) );
  NAND2_X1 U4685 ( .A1(n4600), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U4686 ( .A1(n3747), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3754) );
  INV_X1 U4687 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3748) );
  AOI21_X1 U4688 ( .B1(n3748), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3749) );
  AOI21_X1 U4689 ( .B1(n4186), .B2(EAX_REG_4__SCAN_IN), .A(n3749), .ZN(n3753)
         );
  NOR2_X1 U4690 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3751), .ZN(n3752)
         );
  NOR2_X1 U4691 ( .A1(n3762), .A2(n3752), .ZN(n4966) );
  AOI22_X1 U4692 ( .A1(n3754), .A2(n3753), .B1(n4436), .B2(n4966), .ZN(n3755)
         );
  AOI21_X1 U4693 ( .B1(n3756), .B2(n3871), .A(n3755), .ZN(n4715) );
  NAND2_X1 U4694 ( .A1(n3757), .A2(n3871), .ZN(n3761) );
  INV_X1 U4695 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4915) );
  XNOR2_X1 U4696 ( .A(n3762), .B(n4915), .ZN(n4919) );
  OAI22_X1 U4697 ( .A1(n4919), .A2(n4236), .B1(n3758), .B2(n4915), .ZN(n3759)
         );
  AOI21_X1 U4698 ( .B1(n4186), .B2(EAX_REG_5__SCAN_IN), .A(n3759), .ZN(n3760)
         );
  NAND2_X1 U4699 ( .A1(n3761), .A2(n3760), .ZN(n4711) );
  NAND2_X1 U4700 ( .A1(n4709), .A2(n4711), .ZN(n4710) );
  INV_X1 U4701 ( .A(n4710), .ZN(n3774) );
  INV_X1 U4702 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3764) );
  XNOR2_X1 U4703 ( .A(n3785), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5459) );
  AOI22_X1 U4704 ( .A1(n5459), .A2(n4436), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3763) );
  OAI21_X1 U4705 ( .B1(n3732), .B2(n3764), .A(n3763), .ZN(n3765) );
  AND2_X1 U4706 ( .A1(n3767), .A2(n3769), .ZN(n3768) );
  OR2_X1 U4707 ( .A1(n3768), .A2(n3785), .ZN(n5897) );
  OAI22_X1 U4708 ( .A1(n3732), .A2(n5871), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3769), .ZN(n3770) );
  MUX2_X1 U4709 ( .A(n5897), .B(n3770), .S(n4236), .Z(n3771) );
  AOI22_X1 U4710 ( .A1(n4219), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4711 ( .A1(n4212), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4712 ( .A1(n4060), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4713 ( .A1(n4016), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4714 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3784)
         );
  AOI22_X1 U4715 ( .A1(n7031), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4716 ( .A1(n4117), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4717 ( .A1(n4208), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4718 ( .A1(n3388), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4719 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  OAI21_X1 U4720 ( .B1(n3784), .B2(n3783), .A(n3871), .ZN(n3789) );
  NAND2_X1 U4721 ( .A1(n4186), .A2(EAX_REG_8__SCAN_IN), .ZN(n3788) );
  XNOR2_X1 U4722 ( .A(n3790), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U4723 ( .A1(n4976), .A2(n4436), .ZN(n3787) );
  NAND2_X1 U4724 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3786)
         );
  XNOR2_X1 U4725 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3814), .ZN(n5798) );
  AOI22_X1 U4726 ( .A1(n4219), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4727 ( .A1(n4016), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4728 ( .A1(n3393), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4729 ( .A1(n4146), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4730 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4731 ( .A1(n4060), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4732 ( .A1(n7031), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4733 ( .A1(n4117), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4734 ( .A1(n4212), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4735 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  OR2_X1 U4736 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  AOI22_X1 U4737 ( .A1(n3871), .A2(n3801), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4738 ( .A1(n4186), .A2(EAX_REG_9__SCAN_IN), .ZN(n3802) );
  OAI211_X1 U4739 ( .C1(n5798), .C2(n4236), .A(n3803), .B(n3802), .ZN(n4931)
         );
  AOI22_X1 U4740 ( .A1(n4208), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4741 ( .A1(n4060), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4742 ( .A1(n4117), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4743 ( .A1(n4016), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4744 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4745 ( .A1(n4563), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4747 ( .A1(n7031), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4748 ( .A1(n3393), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4749 ( .A1(n4209), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4750 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  NOR2_X1 U4751 ( .A1(n3813), .A2(n3812), .ZN(n3817) );
  XNOR2_X1 U4752 ( .A(n3818), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4986)
         );
  NAND2_X1 U4753 ( .A1(n4986), .A2(n4436), .ZN(n3816) );
  AOI22_X1 U4754 ( .A1(n4186), .A2(EAX_REG_10__SCAN_IN), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U4755 ( .C1(n3817), .C2(n3901), .A(n3816), .B(n3815), .ZN(n4940)
         );
  XNOR2_X1 U4756 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3835), .ZN(n5887)
         );
  INV_X1 U4757 ( .A(n5887), .ZN(n3833) );
  AOI22_X1 U4758 ( .A1(n4016), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4759 ( .A1(n4208), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4760 ( .A1(n4563), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4761 ( .A1(n4117), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4762 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4763 ( .A1(n4219), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4764 ( .A1(n4116), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4765 ( .A1(n4060), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4766 ( .A1(n7031), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4767 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  NOR2_X1 U4768 ( .A1(n3828), .A2(n3827), .ZN(n3831) );
  NAND2_X1 U4769 ( .A1(n4186), .A2(EAX_REG_11__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4770 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3829)
         );
  OAI211_X1 U4771 ( .C1(n3901), .C2(n3831), .A(n3830), .B(n3829), .ZN(n3832)
         );
  AOI21_X1 U4772 ( .B1(n3833), .B2(n4436), .A(n3832), .ZN(n4982) );
  INV_X1 U4773 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3836) );
  XNOR2_X1 U4774 ( .A(n3853), .B(n3836), .ZN(n4995) );
  NAND2_X1 U4775 ( .A1(n4995), .A2(n4436), .ZN(n3852) );
  INV_X1 U4776 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3838) );
  OAI21_X1 U4777 ( .B1(n6793), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6436), 
        .ZN(n3837) );
  OAI21_X1 U4778 ( .B1(n3732), .B2(n3838), .A(n3837), .ZN(n3851) );
  AOI22_X1 U4779 ( .A1(n4208), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4780 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4219), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4781 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4060), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4782 ( .A1(n3393), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4783 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4784 ( .A1(n7031), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4785 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4563), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4786 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4117), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4787 ( .A1(n4016), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4788 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4789 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  NOR2_X1 U4790 ( .A1(n3901), .A2(n3849), .ZN(n3850) );
  AOI21_X1 U4791 ( .B1(n3852), .B2(n3851), .A(n3850), .ZN(n4991) );
  NAND2_X1 U4792 ( .A1(n4186), .A2(EAX_REG_13__SCAN_IN), .ZN(n3856) );
  OAI21_X1 U4793 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3854), .A(n3886), 
        .ZN(n5780) );
  AOI22_X1 U4794 ( .A1(n4436), .A2(n5780), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U4795 ( .A1(n3856), .A2(n3855), .ZN(n3857) );
  NAND2_X1 U4796 ( .A1(n3858), .A2(n3857), .ZN(n3872) );
  OAI21_X1 U4797 ( .B1(n3858), .B2(n3857), .A(n3872), .ZN(n3859) );
  AOI22_X1 U4798 ( .A1(n4116), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4799 ( .A1(n4060), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4800 ( .A1(n4117), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4801 ( .A1(n4146), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4802 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3869)
         );
  AOI22_X1 U4803 ( .A1(n4219), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4804 ( .A1(n4016), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4805 ( .A1(n7031), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4806 ( .A1(n3388), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4807 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3868)
         );
  OR2_X1 U4808 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  NAND2_X1 U4809 ( .A1(n5041), .A2(n5042), .ZN(n5044) );
  NAND2_X1 U4810 ( .A1(n5044), .A2(n3872), .ZN(n5049) );
  AOI22_X1 U4811 ( .A1(n7031), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4812 ( .A1(n4016), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4813 ( .A1(n4219), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4814 ( .A1(n4116), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4815 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3882)
         );
  AOI22_X1 U4816 ( .A1(n4563), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4817 ( .A1(n4060), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4818 ( .A1(n4208), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4819 ( .A1(n4117), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4820 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  NOR2_X1 U4821 ( .A1(n3882), .A2(n3881), .ZN(n3885) );
  XNOR2_X1 U4822 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3886), .ZN(n5764)
         );
  INV_X1 U4823 ( .A(n5764), .ZN(n5452) );
  AOI22_X1 U4824 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4436), 
        .B2(n5452), .ZN(n3884) );
  NAND2_X1 U4825 ( .A1(n4186), .A2(EAX_REG_14__SCAN_IN), .ZN(n3883) );
  OAI211_X1 U4826 ( .C1(n3901), .C2(n3885), .A(n3884), .B(n3883), .ZN(n5048)
         );
  NAND2_X1 U4827 ( .A1(n5049), .A2(n5048), .ZN(n5047) );
  XNOR2_X1 U4828 ( .A(n3903), .B(n5255), .ZN(n5441) );
  AOI22_X1 U4829 ( .A1(n4016), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4830 ( .A1(n4060), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4831 ( .A1(n4116), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4832 ( .A1(n4117), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4833 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  AOI22_X1 U4834 ( .A1(n4563), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4835 ( .A1(n7031), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4836 ( .A1(n4219), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4837 ( .A1(n4208), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4838 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NOR2_X1 U4839 ( .A1(n3897), .A2(n3896), .ZN(n3900) );
  NAND2_X1 U4840 ( .A1(n4186), .A2(EAX_REG_15__SCAN_IN), .ZN(n3899) );
  NAND2_X1 U4841 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3898)
         );
  OAI211_X1 U4842 ( .C1(n3901), .C2(n3900), .A(n3899), .B(n3898), .ZN(n3902)
         );
  AOI21_X1 U4843 ( .B1(n5441), .B2(n4436), .A(n3902), .ZN(n5250) );
  XOR2_X1 U4844 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3919), .Z(n5241) );
  INV_X1 U4845 ( .A(n5241), .ZN(n3918) );
  INV_X1 U4846 ( .A(n3713), .ZN(n3904) );
  AOI22_X1 U4847 ( .A1(n4060), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4848 ( .A1(n4208), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4849 ( .A1(n7031), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4850 ( .A1(n4117), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4851 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3914)
         );
  AOI22_X1 U4852 ( .A1(n4219), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4853 ( .A1(n4016), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4854 ( .A1(n4146), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4855 ( .A1(n4212), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4856 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3913)
         );
  NOR2_X1 U4857 ( .A1(n3914), .A2(n3913), .ZN(n3916) );
  AOI22_X1 U4858 ( .A1(n4186), .A2(EAX_REG_16__SCAN_IN), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3915) );
  OAI21_X1 U4859 ( .B1(n4233), .B2(n3916), .A(n3915), .ZN(n3917) );
  AOI21_X1 U4860 ( .B1(n3918), .B2(n4436), .A(n3917), .ZN(n5056) );
  XNOR2_X1 U4861 ( .A(n3935), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5678)
         );
  AOI22_X1 U4862 ( .A1(n4186), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6436), .ZN(n3933) );
  AOI22_X1 U4863 ( .A1(n7031), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4864 ( .A1(n4219), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4865 ( .A1(n4116), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4866 ( .A1(n4016), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4867 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3931)
         );
  NAND2_X1 U4868 ( .A1(n4563), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3925)
         );
  NAND2_X1 U4869 ( .A1(n3393), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3924)
         );
  AND3_X1 U4870 ( .A1(n3925), .A2(n3924), .A3(n4236), .ZN(n3929) );
  AOI22_X1 U4871 ( .A1(n4060), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4872 ( .A1(n4146), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4873 ( .A1(n4217), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4874 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NAND2_X1 U4875 ( .A1(n4233), .A2(n4236), .ZN(n4002) );
  OAI21_X1 U4876 ( .B1(n3931), .B2(n3930), .A(n4002), .ZN(n3932) );
  AOI22_X1 U4877 ( .A1(n5678), .A2(n4436), .B1(n3933), .B2(n3932), .ZN(n5224)
         );
  OR2_X1 U4878 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3937)
         );
  NAND2_X1 U4879 ( .A1(n3937), .A2(n3984), .ZN(n5677) );
  AOI22_X1 U4880 ( .A1(n4016), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4881 ( .A1(n4208), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4882 ( .A1(n4219), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4883 ( .A1(n4116), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4884 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3947)
         );
  AOI22_X1 U4885 ( .A1(n4563), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4886 ( .A1(n4060), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4887 ( .A1(n7031), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4888 ( .A1(n4117), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4889 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  NOR2_X1 U4890 ( .A1(n3947), .A2(n3946), .ZN(n3950) );
  OAI21_X1 U4891 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6793), .A(n6436), 
        .ZN(n3949) );
  NAND2_X1 U4892 ( .A1(n4186), .A2(EAX_REG_18__SCAN_IN), .ZN(n3948) );
  OAI211_X1 U4893 ( .C1(n4233), .C2(n3950), .A(n3949), .B(n3948), .ZN(n3951)
         );
  OAI21_X1 U4894 ( .B1(n5677), .B2(n4236), .A(n3951), .ZN(n4431) );
  NAND2_X1 U4895 ( .A1(n3953), .A2(n3952), .ZN(n4430) );
  AOI22_X1 U4896 ( .A1(n4016), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4897 ( .A1(n7031), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4898 ( .A1(n3393), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4899 ( .A1(n4209), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4900 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3965)
         );
  NAND2_X1 U4901 ( .A1(n4217), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3959) );
  NAND2_X1 U4902 ( .A1(n4116), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3958) );
  AND3_X1 U4903 ( .A1(n3959), .A2(n3958), .A3(n4236), .ZN(n3963) );
  AOI22_X1 U4904 ( .A1(n4117), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4905 ( .A1(n4219), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4906 ( .A1(n4060), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4907 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  OAI21_X1 U4908 ( .B1(n3965), .B2(n3964), .A(n4002), .ZN(n3967) );
  AOI22_X1 U4909 ( .A1(n4239), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6436), .ZN(n3966) );
  NAND2_X1 U4910 ( .A1(n3967), .A2(n3966), .ZN(n3969) );
  XNOR2_X1 U4911 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3984), .ZN(n5642)
         );
  NAND2_X1 U4912 ( .A1(n4436), .A2(n5642), .ZN(n3968) );
  NAND2_X1 U4913 ( .A1(n3969), .A2(n3968), .ZN(n5324) );
  AOI22_X1 U4914 ( .A1(n4016), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4915 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4208), .B1(n4212), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4916 ( .A1(n4219), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4917 ( .A1(n4117), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4918 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3979)
         );
  AOI22_X1 U4919 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4217), .B1(n4563), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4920 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4060), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4921 ( .A1(n4116), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4922 ( .A1(n7031), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4923 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  NOR2_X1 U4924 ( .A1(n3979), .A2(n3978), .ZN(n3983) );
  NAND2_X1 U4925 ( .A1(n6436), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3980)
         );
  NAND2_X1 U4926 ( .A1(n4236), .A2(n3980), .ZN(n3981) );
  AOI21_X1 U4927 ( .B1(n4186), .B2(EAX_REG_20__SCAN_IN), .A(n3981), .ZN(n3982)
         );
  OAI21_X1 U4928 ( .B1(n4233), .B2(n3983), .A(n3982), .ZN(n3988) );
  OAI21_X1 U4929 ( .B1(n3986), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4074), 
        .ZN(n5641) );
  OR2_X1 U4930 ( .A1(n5641), .A2(n4236), .ZN(n3987) );
  AOI22_X1 U4931 ( .A1(n4117), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4932 ( .A1(n4563), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3990)
         );
  NAND2_X1 U4933 ( .A1(n3150), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3989) );
  AND3_X1 U4934 ( .A1(n3990), .A2(n3989), .A3(n4236), .ZN(n3993) );
  AOI22_X1 U4935 ( .A1(n4219), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4936 ( .A1(n4217), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4937 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4000)
         );
  AOI22_X1 U4938 ( .A1(n3393), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4939 ( .A1(n4208), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4940 ( .A1(n4016), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4941 ( .A1(n4060), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4942 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  OR2_X1 U4943 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  NAND2_X1 U4944 ( .A1(n4002), .A2(n4001), .ZN(n4005) );
  AOI22_X1 U4945 ( .A1(n4239), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6436), .ZN(n4004) );
  XNOR2_X1 U4946 ( .A(n4074), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5625)
         );
  AOI22_X1 U4947 ( .A1(n4219), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4948 ( .A1(n3314), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4949 ( .A1(n4116), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4950 ( .A1(n4117), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4951 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4015)
         );
  AOI22_X1 U4952 ( .A1(n4060), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4953 ( .A1(n7031), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4954 ( .A1(n4212), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4955 ( .A1(n4146), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4956 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4014)
         );
  NOR2_X1 U4957 ( .A1(n4015), .A2(n4014), .ZN(n4091) );
  AOI22_X1 U4958 ( .A1(n4016), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4959 ( .A1(n7031), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4960 ( .A1(n4211), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4017), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4961 ( .A1(n4212), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4962 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4027)
         );
  AOI22_X1 U4963 ( .A1(n4060), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4964 ( .A1(n4563), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4965 ( .A1(n4117), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4966 ( .A1(n4146), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U4967 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4026)
         );
  NOR2_X1 U4968 ( .A1(n4027), .A2(n4026), .ZN(n4109) );
  AOI22_X1 U4969 ( .A1(n3150), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4970 ( .A1(n4208), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4971 ( .A1(n4217), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4972 ( .A1(n3388), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U4973 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4037)
         );
  AOI22_X1 U4974 ( .A1(n4117), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4975 ( .A1(n4219), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4976 ( .A1(n4145), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4977 ( .A1(n3314), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U4978 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4036)
         );
  NOR2_X1 U4979 ( .A1(n4037), .A2(n4036), .ZN(n4108) );
  OR2_X1 U4980 ( .A1(n4109), .A2(n4108), .ZN(n4101) );
  AOI22_X1 U4981 ( .A1(n7031), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4982 ( .A1(n4211), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4983 ( .A1(n4145), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4984 ( .A1(n4208), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U4985 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U4986 ( .A1(n3314), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4987 ( .A1(n4212), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4988 ( .A1(n4117), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4989 ( .A1(n4219), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U4990 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  OR2_X1 U4991 ( .A1(n4047), .A2(n4046), .ZN(n4100) );
  INV_X1 U4992 ( .A(n4100), .ZN(n4048) );
  NOR2_X1 U4993 ( .A1(n4091), .A2(n4092), .ZN(n4081) );
  AOI22_X1 U4994 ( .A1(n4145), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4995 ( .A1(n4563), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4996 ( .A1(n4117), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4997 ( .A1(n4146), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U4998 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4059)
         );
  AOI22_X1 U4999 ( .A1(n3314), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5000 ( .A1(n7031), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5001 ( .A1(n4211), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5002 ( .A1(n4123), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U5003 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4058)
         );
  OR2_X1 U5004 ( .A1(n4059), .A2(n4058), .ZN(n4079) );
  NAND2_X1 U5005 ( .A1(n4081), .A2(n4079), .ZN(n4143) );
  AOI22_X1 U5006 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4060), .B1(n4117), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5007 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4217), .B1(n4563), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5008 ( .A1(n3150), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5009 ( .A1(n4208), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4061) );
  NAND4_X1 U5010 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4070)
         );
  AOI22_X1 U5011 ( .A1(n4211), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5012 ( .A1(n4219), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5013 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4146), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5014 ( .A1(n3314), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5015 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4069)
         );
  NOR2_X1 U5016 ( .A1(n4070), .A2(n4069), .ZN(n4144) );
  XOR2_X1 U5017 ( .A(n4143), .B(n4144), .Z(n4071) );
  NAND2_X1 U5018 ( .A1(n4071), .A2(n4183), .ZN(n4078) );
  NAND2_X1 U5019 ( .A1(n6436), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4072)
         );
  NAND2_X1 U5020 ( .A1(n4236), .A2(n4072), .ZN(n4073) );
  AOI21_X1 U5021 ( .B1(n4186), .B2(EAX_REG_27__SCAN_IN), .A(n4073), .ZN(n4077)
         );
  XNOR2_X1 U5022 ( .A(n4163), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5385)
         );
  AND2_X1 U5023 ( .A1(n5385), .A2(n4436), .ZN(n4076) );
  AOI21_X1 U5024 ( .B1(n4078), .B2(n4077), .A(n4076), .ZN(n5190) );
  INV_X1 U5025 ( .A(n4079), .ZN(n4080) );
  XNOR2_X1 U5026 ( .A(n4081), .B(n4080), .ZN(n4082) );
  NAND2_X1 U5027 ( .A1(n4082), .A2(n4183), .ZN(n4090) );
  INV_X1 U5028 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4086) );
  AOI21_X1 U5029 ( .B1(n4086), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4083) );
  AOI21_X1 U5030 ( .B1(n4186), .B2(EAX_REG_26__SCAN_IN), .A(n4083), .ZN(n4089)
         );
  INV_X1 U5031 ( .A(n4084), .ZN(n4085) );
  NAND2_X1 U5032 ( .A1(n4086), .A2(n4085), .ZN(n4087) );
  NAND2_X1 U5033 ( .A1(n4163), .A2(n4087), .ZN(n5605) );
  NOR2_X1 U5034 ( .A1(n5605), .A2(n4236), .ZN(n4088) );
  AOI21_X1 U5035 ( .B1(n4090), .B2(n4089), .A(n4088), .ZN(n5284) );
  INV_X1 U5036 ( .A(n5284), .ZN(n4141) );
  XOR2_X1 U5037 ( .A(n4092), .B(n4091), .Z(n4093) );
  NAND2_X1 U5038 ( .A1(n4093), .A2(n4183), .ZN(n4099) );
  NAND2_X1 U5039 ( .A1(n6436), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4094)
         );
  NAND2_X1 U5040 ( .A1(n4236), .A2(n4094), .ZN(n4095) );
  AOI21_X1 U5041 ( .B1(n4186), .B2(EAX_REG_25__SCAN_IN), .A(n4095), .ZN(n4098)
         );
  XNOR2_X1 U5042 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4096), .ZN(n5402)
         );
  AND2_X1 U5043 ( .A1(n4436), .A2(n5402), .ZN(n4097) );
  AOI21_X1 U5044 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(n5292) );
  INV_X1 U5045 ( .A(n5292), .ZN(n4140) );
  XNOR2_X1 U5046 ( .A(n4101), .B(n4100), .ZN(n4107) );
  INV_X1 U5047 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4102) );
  XNOR2_X1 U5048 ( .A(n4103), .B(n4102), .ZN(n5616) );
  NAND2_X1 U5049 ( .A1(n4186), .A2(EAX_REG_24__SCAN_IN), .ZN(n4105) );
  NAND2_X1 U5050 ( .A1(n4238), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4104)
         );
  OAI211_X1 U5051 ( .C1(n5616), .C2(n4236), .A(n4105), .B(n4104), .ZN(n4106)
         );
  AOI21_X1 U5052 ( .B1(n4107), .B2(n4183), .A(n4106), .ZN(n5099) );
  XOR2_X1 U5053 ( .A(n4109), .B(n4108), .Z(n4110) );
  NAND2_X1 U5054 ( .A1(n4110), .A2(n4183), .ZN(n4113) );
  INV_X1 U5055 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5075) );
  AOI21_X1 U5056 ( .B1(n5075), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4111) );
  AOI21_X1 U5057 ( .B1(n4186), .B2(EAX_REG_23__SCAN_IN), .A(n4111), .ZN(n4112)
         );
  NAND2_X1 U5058 ( .A1(n4113), .A2(n4112), .ZN(n4115) );
  XNOR2_X1 U5059 ( .A(n4136), .B(n5075), .ZN(n5205) );
  NAND2_X1 U5060 ( .A1(n5205), .A2(n4436), .ZN(n4114) );
  NAND2_X1 U5061 ( .A1(n4115), .A2(n4114), .ZN(n5079) );
  AOI22_X1 U5062 ( .A1(n7031), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5063 ( .A1(n4145), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5064 ( .A1(n4016), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5065 ( .A1(n4117), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4118) );
  NAND4_X1 U5066 ( .A1(n4121), .A2(n4120), .A3(n4119), .A4(n4118), .ZN(n4129)
         );
  AOI22_X1 U5067 ( .A1(n4219), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4563), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5068 ( .A1(n4208), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5069 ( .A1(n4146), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5070 ( .A1(n4123), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5071 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4128)
         );
  NOR2_X1 U5072 ( .A1(n4129), .A2(n4128), .ZN(n4133) );
  NAND2_X1 U5073 ( .A1(n6436), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4130)
         );
  NAND2_X1 U5074 ( .A1(n4236), .A2(n4130), .ZN(n4131) );
  AOI21_X1 U5075 ( .B1(n4186), .B2(EAX_REG_22__SCAN_IN), .A(n4131), .ZN(n4132)
         );
  OAI21_X1 U5076 ( .B1(n4233), .B2(n4133), .A(n4132), .ZN(n4139) );
  NOR2_X1 U5077 ( .A1(n4134), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4135)
         );
  OR2_X1 U5078 ( .A1(n4136), .A2(n4135), .ZN(n5410) );
  INV_X1 U5079 ( .A(n5410), .ZN(n4137) );
  NAND2_X1 U5080 ( .A1(n4137), .A2(n4436), .ZN(n4138) );
  NAND2_X1 U5081 ( .A1(n4139), .A2(n4138), .ZN(n5213) );
  NOR2_X1 U5082 ( .A1(n4141), .A2(n5282), .ZN(n5188) );
  AND2_X1 U5083 ( .A1(n5190), .A2(n5188), .ZN(n4142) );
  NOR2_X1 U5084 ( .A1(n4144), .A2(n4143), .ZN(n4170) );
  AOI22_X1 U5085 ( .A1(n4145), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4219), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5086 ( .A1(n4563), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5087 ( .A1(n4220), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5088 ( .A1(n4146), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5089 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4156)
         );
  AOI22_X1 U5090 ( .A1(n3314), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5091 ( .A1(n3150), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5092 ( .A1(n4211), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5093 ( .A1(n4212), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U5094 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4155)
         );
  OR2_X1 U5095 ( .A1(n4156), .A2(n4155), .ZN(n4169) );
  INV_X1 U5096 ( .A(n4169), .ZN(n4157) );
  XNOR2_X1 U5097 ( .A(n4170), .B(n4157), .ZN(n4161) );
  INV_X1 U5098 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U5099 ( .A1(n6436), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4158)
         );
  OAI211_X1 U5100 ( .C1(n3732), .C2(n4159), .A(n4236), .B(n4158), .ZN(n4160)
         );
  AOI21_X1 U5101 ( .B1(n4161), .B2(n4183), .A(n4160), .ZN(n4168) );
  INV_X1 U5102 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4162) );
  INV_X1 U5103 ( .A(n4164), .ZN(n4165) );
  INV_X1 U5104 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U5105 ( .A1(n4165), .A2(n5181), .ZN(n4166) );
  NAND2_X1 U5106 ( .A1(n4206), .A2(n4166), .ZN(n5379) );
  NOR2_X1 U5107 ( .A1(n5379), .A2(n4236), .ZN(n4167) );
  NAND2_X1 U5108 ( .A1(n4170), .A2(n4169), .ZN(n4227) );
  AOI22_X1 U5109 ( .A1(n4219), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5110 ( .A1(n3150), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5111 ( .A1(n3314), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5112 ( .A1(n4145), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U5113 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4182)
         );
  AOI22_X1 U5114 ( .A1(n4208), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4212), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5115 ( .A1(n4220), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5116 ( .A1(n4563), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5117 ( .A1(n4211), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4177) );
  NAND4_X1 U5118 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), .ZN(n4181)
         );
  NOR2_X1 U5119 ( .A1(n4182), .A2(n4181), .ZN(n4228) );
  XOR2_X1 U5120 ( .A(n4227), .B(n4228), .Z(n4184) );
  NAND2_X1 U5121 ( .A1(n4184), .A2(n4183), .ZN(n4188) );
  INV_X1 U5122 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5170) );
  NOR2_X1 U5123 ( .A1(n5170), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4185) );
  AOI211_X1 U5124 ( .C1(n4186), .C2(EAX_REG_29__SCAN_IN), .A(n4436), .B(n4185), 
        .ZN(n4187) );
  XNOR2_X1 U5125 ( .A(n4206), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4196)
         );
  AOI22_X1 U5126 ( .A1(n4188), .A2(n4187), .B1(n4436), .B2(n4196), .ZN(n4190)
         );
  OAI21_X1 U5127 ( .B1(n4189), .B2(n4190), .A(n4237), .ZN(n5165) );
  INV_X1 U5128 ( .A(n5165), .ZN(n4191) );
  AND2_X1 U5129 ( .A1(n6542), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4435) );
  NAND2_X1 U5130 ( .A1(n4435), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6556) );
  INV_X2 U5131 ( .A(n4644), .ZN(n5910) );
  NAND2_X1 U5132 ( .A1(n6438), .A2(n4197), .ZN(n6626) );
  NAND2_X1 U5133 ( .A1(n6626), .A2(n6542), .ZN(n4192) );
  NAND2_X1 U5134 ( .A1(n6542), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5135 ( .A1(n6793), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U5136 ( .A1(n4194), .A2(n4193), .ZN(n5920) );
  INV_X1 U5137 ( .A(n5920), .ZN(n4195) );
  INV_X1 U5138 ( .A(n4196), .ZN(n5169) );
  INV_X1 U5139 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6597) );
  NOR2_X1 U5140 ( .A1(n5721), .A2(n6597), .ZN(n5473) );
  AOI21_X1 U5141 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5473), 
        .ZN(n4198) );
  OAI21_X1 U5142 ( .B1(n5915), .B2(n5169), .A(n4198), .ZN(n4199) );
  NAND2_X1 U5143 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5463) );
  INV_X1 U5144 ( .A(n4202), .ZN(n5400) );
  INV_X1 U5145 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5476) );
  INV_X1 U5146 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U5147 ( .A1(n5400), .A2(n4203), .A3(n5476), .A4(n4323), .ZN(n4204)
         );
  XNOR2_X1 U5148 ( .A(n4205), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5471)
         );
  INV_X1 U5149 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4207) );
  XNOR2_X1 U5150 ( .A(n4241), .B(n4207), .ZN(n5157) );
  AOI22_X1 U5151 ( .A1(n3150), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4208), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5152 ( .A1(n4145), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5153 ( .A1(n4211), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5154 ( .A1(n4212), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4171), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U5155 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4226)
         );
  AOI22_X1 U5156 ( .A1(n4016), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5157 ( .A1(n4563), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4217), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5158 ( .A1(n4219), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5159 ( .A1(n4220), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4221) );
  NAND4_X1 U5160 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  NOR2_X1 U5161 ( .A1(n4226), .A2(n4225), .ZN(n4230) );
  NOR2_X1 U5162 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  XOR2_X1 U5163 ( .A(n4230), .B(n4229), .Z(n4234) );
  AOI21_X1 U5164 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6436), .A(n4436), 
        .ZN(n4232) );
  NAND2_X1 U5165 ( .A1(n4239), .A2(EAX_REG_30__SCAN_IN), .ZN(n4231) );
  OAI211_X1 U5166 ( .C1(n4234), .C2(n4233), .A(n4232), .B(n4231), .ZN(n4235)
         );
  OAI21_X1 U5167 ( .B1(n4236), .B2(n5157), .A(n4235), .ZN(n5085) );
  AOI22_X1 U5168 ( .A1(n4239), .A2(EAX_REG_31__SCAN_IN), .B1(n4238), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4240) );
  INV_X1 U5169 ( .A(n4241), .ZN(n4242) );
  NAND2_X1 U5170 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4243)
         );
  INV_X1 U5171 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5144) );
  INV_X1 U5172 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U5173 ( .A1(n5721), .A2(n6786), .ZN(n5466) );
  AOI21_X1 U5174 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5466), 
        .ZN(n4244) );
  OAI21_X1 U5175 ( .B1(n5915), .B2(n4447), .A(n4244), .ZN(n4245) );
  OAI21_X1 U5176 ( .B1(n5918), .B2(n5471), .A(n4246), .ZN(U2955) );
  NAND2_X1 U5177 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U5178 ( .A1(n4250), .A2(n5476), .ZN(n4247) );
  NAND2_X1 U5179 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  NAND3_X1 U5180 ( .A1(n4250), .A2(n5476), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4253) );
  INV_X1 U5181 ( .A(n5463), .ZN(n4316) );
  NAND2_X1 U5182 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  NOR2_X1 U5183 ( .A1(n4255), .A2(n4254), .ZN(n5090) );
  NOR2_X1 U5184 ( .A1(n3713), .A2(n4733), .ZN(n4300) );
  INV_X1 U5185 ( .A(n4300), .ZN(n4271) );
  NOR2_X1 U5186 ( .A1(n3353), .A2(n4528), .ZN(n4257) );
  INV_X1 U5187 ( .A(n4434), .ZN(n4472) );
  NAND2_X1 U5188 ( .A1(n4295), .A2(n3157), .ZN(n4258) );
  OR2_X1 U5189 ( .A1(n4282), .A2(n4258), .ZN(n4259) );
  NAND2_X1 U5190 ( .A1(n4472), .A2(n4259), .ZN(n4489) );
  INV_X1 U5191 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U5192 ( .A1(n4261), .A2(n4260), .ZN(n6564) );
  INV_X1 U5193 ( .A(n6564), .ZN(n4269) );
  AND2_X1 U5194 ( .A1(n4263), .A2(n4262), .ZN(n4266) );
  AOI21_X1 U5195 ( .B1(n4266), .B2(n4265), .A(n4264), .ZN(n4473) );
  NAND2_X1 U5196 ( .A1(n4473), .A2(n6627), .ZN(n4610) );
  INV_X1 U5197 ( .A(n4610), .ZN(n4268) );
  OAI211_X1 U5198 ( .C1(n4733), .C2(n4269), .A(n4268), .B(n4267), .ZN(n4270)
         );
  OAI211_X1 U5199 ( .C1(n4501), .C2(n4271), .A(n4489), .B(n4270), .ZN(n4272)
         );
  NAND2_X1 U5200 ( .A1(n4272), .A2(n6548), .ZN(n4280) );
  NAND2_X1 U5201 ( .A1(n4733), .A2(n6564), .ZN(n4440) );
  AND2_X1 U5202 ( .A1(n4440), .A2(n6627), .ZN(n4275) );
  NAND2_X1 U5203 ( .A1(n4274), .A2(n4275), .ZN(n4483) );
  INV_X1 U5204 ( .A(n4276), .ZN(n5346) );
  NAND3_X1 U5205 ( .A1(n4483), .A2(n4528), .A3(n5346), .ZN(n4277) );
  NAND2_X1 U5206 ( .A1(n4277), .A2(n4649), .ZN(n4278) );
  INV_X1 U5207 ( .A(n4281), .ZN(n6500) );
  NOR2_X1 U5208 ( .A1(n4282), .A2(n4608), .ZN(n4612) );
  OR2_X1 U5209 ( .A1(n6500), .A2(n4612), .ZN(n4471) );
  NOR2_X1 U5210 ( .A1(n4284), .A2(n4733), .ZN(n4287) );
  OAI21_X1 U5211 ( .B1(n4782), .B2(n4423), .A(n4285), .ZN(n4286) );
  NOR3_X1 U5212 ( .A1(n4471), .A2(n4287), .A3(n4286), .ZN(n4288) );
  NAND2_X1 U5213 ( .A1(n4434), .A2(n4544), .ZN(n6507) );
  NAND2_X1 U5214 ( .A1(n4653), .A2(n4544), .ZN(n4828) );
  NOR2_X1 U5215 ( .A1(n4828), .A2(n4291), .ZN(n4487) );
  OAI21_X1 U5216 ( .B1(n4487), .B2(n5127), .A(n3491), .ZN(n4294) );
  NAND2_X1 U5217 ( .A1(n4290), .A2(n5316), .ZN(n4293) );
  NAND2_X1 U5218 ( .A1(n5346), .A2(n4291), .ZN(n4292) );
  AND4_X1 U5219 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4296)
         );
  OAI211_X1 U5220 ( .C1(n4496), .C2(n4528), .A(n4499), .B(n4571), .ZN(n4298)
         );
  INV_X1 U5221 ( .A(n4298), .ZN(n4299) );
  INV_X1 U5222 ( .A(n4510), .ZN(n4554) );
  NAND2_X1 U5223 ( .A1(n5927), .A2(n5708), .ZN(n5928) );
  INV_X1 U5224 ( .A(n5928), .ZN(n6005) );
  INV_X1 U5225 ( .A(n5512), .ZN(n4301) );
  AND2_X1 U5226 ( .A1(n5928), .A2(n4301), .ZN(n4307) );
  NOR2_X1 U5227 ( .A1(n5997), .A2(n6015), .ZN(n5993) );
  NAND3_X1 U5228 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n5993), .ZN(n5965) );
  NOR3_X1 U5229 ( .A1(n5963), .A2(n4819), .A3(n5965), .ZN(n5926) );
  NAND2_X1 U5230 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5231 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5932) );
  NOR2_X1 U5232 ( .A1(n5945), .A2(n5932), .ZN(n4304) );
  NAND2_X1 U5233 ( .A1(n5926), .A2(n4304), .ZN(n5014) );
  NAND2_X1 U5234 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5712) );
  NOR2_X1 U5235 ( .A1(n3641), .A2(n5712), .ZN(n5718) );
  NAND2_X1 U5236 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5718), .ZN(n5564) );
  NAND2_X1 U5237 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5573) );
  NOR2_X1 U5238 ( .A1(n5564), .A2(n5573), .ZN(n5533) );
  NAND4_X1 U5239 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5533), .A4(n5538), .ZN(n4305)
         );
  NOR2_X1 U5240 ( .A1(n5014), .A2(n4305), .ZN(n4318) );
  INV_X1 U5241 ( .A(n5709), .ZN(n4302) );
  INV_X1 U5242 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4308) );
  NAND2_X1 U5243 ( .A1(n4302), .A2(n4308), .ZN(n4303) );
  NAND2_X1 U5244 ( .A1(n4426), .A2(n5721), .ZN(n6026) );
  AOI21_X1 U5245 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5994) );
  NAND2_X1 U5246 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U5247 ( .A1(n5994), .A2(n5978), .ZN(n5967) );
  NAND2_X1 U5248 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5967), .ZN(n4818)
         );
  NOR2_X1 U5249 ( .A1(n4819), .A2(n4818), .ZN(n5923) );
  NAND2_X1 U5250 ( .A1(n4304), .A2(n5923), .ZN(n5530) );
  NOR2_X1 U5251 ( .A1(n4305), .A2(n5530), .ZN(n4317) );
  OR2_X1 U5252 ( .A1(n4317), .A2(n5708), .ZN(n4306) );
  OAI211_X1 U5253 ( .C1(n5927), .C2(n4318), .A(n5011), .B(n4306), .ZN(n5524)
         );
  OR2_X1 U5254 ( .A1(n4307), .A2(n5524), .ZN(n5070) );
  INV_X1 U5255 ( .A(n5070), .ZN(n4312) );
  INV_X1 U5256 ( .A(n5998), .ZN(n5964) );
  NAND2_X1 U5257 ( .A1(n5708), .A2(n5964), .ZN(n4310) );
  INV_X1 U5258 ( .A(n4309), .ZN(n4321) );
  NAND2_X1 U5259 ( .A1(n4310), .A2(n4321), .ZN(n4311) );
  NAND2_X1 U5260 ( .A1(n4312), .A2(n4311), .ZN(n5686) );
  NAND2_X1 U5261 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5502) );
  AND2_X1 U5262 ( .A1(n5928), .A2(n5502), .ZN(n4313) );
  INV_X1 U5263 ( .A(n4322), .ZN(n4314) );
  AND2_X1 U5264 ( .A1(n5928), .A2(n4314), .ZN(n4315) );
  NOR2_X1 U5265 ( .A1(n5494), .A2(n4315), .ZN(n5477) );
  OAI21_X1 U5266 ( .B1(n4316), .B2(n6005), .A(n5477), .ZN(n5467) );
  INV_X1 U5267 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U5268 ( .A1(n5721), .A2(n6599), .ZN(n5086) );
  INV_X1 U5269 ( .A(n4317), .ZN(n4320) );
  NAND2_X1 U5270 ( .A1(n4318), .A2(n5998), .ZN(n4319) );
  OAI21_X1 U5271 ( .B1(n5708), .B2(n4320), .A(n4319), .ZN(n5510) );
  NAND2_X1 U5272 ( .A1(n5510), .A2(n5512), .ZN(n5068) );
  NOR2_X1 U5273 ( .A1(n5693), .A2(n5502), .ZN(n5493) );
  NAND2_X1 U5274 ( .A1(n5493), .A2(n4322), .ZN(n5464) );
  INV_X1 U5275 ( .A(n5464), .ZN(n5474) );
  AND3_X1 U5276 ( .A1(n5474), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4323), 
        .ZN(n4324) );
  AOI211_X1 U5277 ( .C1(n5467), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5086), .B(n4324), .ZN(n4428) );
  NAND2_X1 U5278 ( .A1(n4350), .A2(n6015), .ZN(n4326) );
  AND2_X2 U5279 ( .A1(n4528), .A2(n3340), .ZN(n4524) );
  INV_X1 U5280 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4327) );
  NAND2_X1 U5281 ( .A1(n4524), .A2(n4327), .ZN(n4325) );
  NAND3_X1 U5282 ( .A1(n4326), .A2(n4335), .A3(n4325), .ZN(n4329) );
  NAND2_X1 U5283 ( .A1(n5316), .A2(n4327), .ZN(n4328) );
  NAND2_X1 U5284 ( .A1(n4329), .A2(n4328), .ZN(n4333) );
  NAND2_X1 U5285 ( .A1(n4350), .A2(EBX_REG_0__SCAN_IN), .ZN(n4331) );
  INV_X1 U5286 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U5287 ( .A1(n4335), .A2(n4865), .ZN(n4330) );
  NAND2_X1 U5288 ( .A1(n4331), .A2(n4330), .ZN(n4517) );
  XNOR2_X1 U5289 ( .A(n4333), .B(n4517), .ZN(n4525) );
  INV_X1 U5290 ( .A(n4517), .ZN(n4332) );
  OR2_X1 U5291 ( .A1(n4333), .A2(n4332), .ZN(n4334) );
  MUX2_X1 U5292 ( .A(n5121), .B(n4335), .S(EBX_REG_3__SCAN_IN), .Z(n4337) );
  OR2_X1 U5293 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4336)
         );
  NAND2_X1 U5294 ( .A1(n4337), .A2(n4336), .ZN(n4619) );
  INV_X1 U5295 ( .A(n4619), .ZN(n4340) );
  MUX2_X1 U5296 ( .A(n4335), .B(n4350), .S(EBX_REG_2__SCAN_IN), .Z(n4339) );
  NAND2_X1 U5297 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4338)
         );
  NAND2_X1 U5298 ( .A1(n4339), .A2(n4338), .ZN(n4618) );
  NAND2_X1 U5299 ( .A1(n4350), .A2(n5981), .ZN(n4343) );
  INV_X1 U5300 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U5301 ( .A1(n4524), .A2(n4344), .ZN(n4342) );
  NAND3_X1 U5302 ( .A1(n4343), .A2(n5119), .A3(n4342), .ZN(n4346) );
  NAND2_X1 U5303 ( .A1(n5316), .A2(n4344), .ZN(n4345) );
  AND2_X1 U5304 ( .A1(n4346), .A2(n4345), .ZN(n4716) );
  INV_X1 U5305 ( .A(n5121), .ZN(n4382) );
  INV_X1 U5306 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5307 ( .A1(n4382), .A2(n4804), .ZN(n4349) );
  NAND2_X1 U5308 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4347)
         );
  OAI211_X1 U5309 ( .C1(n5126), .C2(EBX_REG_5__SCAN_IN), .A(n4350), .B(n4347), 
        .ZN(n4348) );
  AND2_X1 U5310 ( .A1(n4349), .A2(n4348), .ZN(n4712) );
  NAND2_X1 U5311 ( .A1(n4350), .A2(n4819), .ZN(n4352) );
  INV_X1 U5312 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4811) );
  NAND2_X1 U5313 ( .A1(n4524), .A2(n4811), .ZN(n4351) );
  NAND3_X1 U5314 ( .A1(n4352), .A2(n5119), .A3(n4351), .ZN(n4354) );
  NAND2_X1 U5315 ( .A1(n5316), .A2(n4811), .ZN(n4353) );
  NAND2_X1 U5316 ( .A1(n4354), .A2(n4353), .ZN(n4808) );
  NAND2_X1 U5317 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4355)
         );
  OAI211_X1 U5318 ( .C1(n5126), .C2(EBX_REG_7__SCAN_IN), .A(n4350), .B(n4355), 
        .ZN(n4356) );
  OAI21_X1 U5319 ( .B1(n5121), .B2(EBX_REG_7__SCAN_IN), .A(n4356), .ZN(n5266)
         );
  MUX2_X1 U5320 ( .A(n5121), .B(n5119), .S(EBX_REG_9__SCAN_IN), .Z(n4360) );
  OR2_X1 U5321 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4359)
         );
  NAND2_X1 U5322 ( .A1(n4360), .A2(n4359), .ZN(n4934) );
  INV_X1 U5323 ( .A(n4934), .ZN(n4366) );
  NAND2_X1 U5324 ( .A1(n4350), .A2(n4361), .ZN(n4363) );
  INV_X1 U5325 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U5326 ( .A1(n4524), .A2(n4858), .ZN(n4362) );
  NAND3_X1 U5327 ( .A1(n4363), .A2(n5119), .A3(n4362), .ZN(n4365) );
  NAND2_X1 U5328 ( .A1(n5316), .A2(n4858), .ZN(n4364) );
  NAND2_X1 U5329 ( .A1(n4365), .A2(n4364), .ZN(n4933) );
  NAND2_X1 U5330 ( .A1(n4366), .A2(n4933), .ZN(n4367) );
  MUX2_X1 U5331 ( .A(n5119), .B(n4350), .S(EBX_REG_10__SCAN_IN), .Z(n4369) );
  NAND2_X1 U5332 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5333 ( .A1(n4369), .A2(n4368), .ZN(n4942) );
  NAND2_X1 U5334 ( .A1(n4943), .A2(n4942), .ZN(n5009) );
  NAND2_X1 U5335 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4370) );
  OAI211_X1 U5336 ( .C1(n5126), .C2(EBX_REG_11__SCAN_IN), .A(n4350), .B(n4370), 
        .ZN(n4371) );
  OAI21_X1 U5337 ( .B1(n5121), .B2(EBX_REG_11__SCAN_IN), .A(n4371), .ZN(n5010)
         );
  OR2_X2 U5338 ( .A1(n5009), .A2(n5010), .ZN(n5007) );
  MUX2_X1 U5339 ( .A(n5119), .B(n4350), .S(EBX_REG_12__SCAN_IN), .Z(n4373) );
  NAND2_X1 U5340 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4372) );
  OR2_X2 U5341 ( .A1(n5007), .A2(n4992), .ZN(n5725) );
  NAND2_X1 U5342 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4374) );
  OAI211_X1 U5343 ( .C1(n5126), .C2(EBX_REG_13__SCAN_IN), .A(n4350), .B(n4374), 
        .ZN(n4375) );
  OAI21_X1 U5344 ( .B1(n5121), .B2(EBX_REG_13__SCAN_IN), .A(n4375), .ZN(n5724)
         );
  MUX2_X1 U5345 ( .A(n5119), .B(n4350), .S(EBX_REG_14__SCAN_IN), .Z(n4377) );
  NAND2_X1 U5346 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U5347 ( .A1(n4377), .A2(n4376), .ZN(n5050) );
  NAND2_X1 U5348 ( .A1(n5727), .A2(n5050), .ZN(n5252) );
  NAND2_X1 U5349 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U5350 ( .C1(n5126), .C2(EBX_REG_15__SCAN_IN), .A(n4350), .B(n4378), 
        .ZN(n4379) );
  OAI21_X1 U5351 ( .B1(n5121), .B2(EBX_REG_15__SCAN_IN), .A(n4379), .ZN(n5251)
         );
  MUX2_X1 U5352 ( .A(n5119), .B(n4350), .S(EBX_REG_16__SCAN_IN), .Z(n4381) );
  NAND2_X1 U5353 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4380) );
  INV_X1 U5354 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U5355 ( .A1(n4382), .A2(n5331), .ZN(n4385) );
  NAND2_X1 U5356 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4383) );
  OAI211_X1 U5357 ( .C1(n5126), .C2(EBX_REG_17__SCAN_IN), .A(n4350), .B(n4383), 
        .ZN(n4384) );
  AND2_X2 U5358 ( .A1(n5240), .A2(n5225), .ZN(n5227) );
  INV_X1 U5359 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U5360 ( .A1(n4350), .A2(n5061), .ZN(n4387) );
  INV_X1 U5361 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5362 ( .A1(n4524), .A2(n4388), .ZN(n4386) );
  NAND3_X1 U5363 ( .A1(n4387), .A2(n5119), .A3(n4386), .ZN(n4390) );
  NAND2_X1 U5364 ( .A1(n5316), .A2(n4388), .ZN(n4389) );
  NAND2_X1 U5365 ( .A1(n4390), .A2(n4389), .ZN(n5325) );
  NAND2_X1 U5366 ( .A1(n5227), .A2(n5325), .ZN(n5315) );
  INV_X1 U5367 ( .A(n5127), .ZN(n4392) );
  INV_X1 U5368 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5064) );
  NOR2_X1 U5369 ( .A1(n5126), .A2(EBX_REG_20__SCAN_IN), .ZN(n4391) );
  AOI21_X1 U5370 ( .B1(n4392), .B2(n5064), .A(n4391), .ZN(n5318) );
  OR2_X1 U5371 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4393)
         );
  INV_X1 U5372 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U5373 ( .A1(n4524), .A2(n5329), .ZN(n4453) );
  NAND2_X1 U5374 ( .A1(n4393), .A2(n4453), .ZN(n5314) );
  NAND2_X1 U5375 ( .A1(n5316), .A2(EBX_REG_20__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5376 ( .A1(n5314), .A2(n5119), .ZN(n4394) );
  OAI211_X1 U5377 ( .C1(n5318), .C2(n5314), .A(n4395), .B(n4394), .ZN(n4396)
         );
  MUX2_X1 U5378 ( .A(n5121), .B(n5119), .S(EBX_REG_21__SCAN_IN), .Z(n4397) );
  OAI21_X1 U5379 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5127), .A(n4397), 
        .ZN(n5312) );
  MUX2_X1 U5380 ( .A(n5119), .B(n4350), .S(EBX_REG_22__SCAN_IN), .Z(n4399) );
  NAND2_X1 U5381 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5382 ( .A1(n4399), .A2(n4398), .ZN(n5216) );
  NAND2_X1 U5383 ( .A1(n5311), .A2(n5216), .ZN(n5215) );
  NAND2_X1 U5384 ( .A1(n5119), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4400) );
  OAI211_X1 U5385 ( .C1(n5126), .C2(EBX_REG_23__SCAN_IN), .A(n4350), .B(n4400), 
        .ZN(n4401) );
  OAI21_X1 U5386 ( .B1(n5121), .B2(EBX_REG_23__SCAN_IN), .A(n4401), .ZN(n5072)
         );
  OR2_X2 U5387 ( .A1(n5215), .A2(n5072), .ZN(n5299) );
  MUX2_X1 U5388 ( .A(n5121), .B(n5119), .S(EBX_REG_25__SCAN_IN), .Z(n4403) );
  OR2_X1 U5389 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4402)
         );
  NAND2_X1 U5390 ( .A1(n4403), .A2(n4402), .ZN(n5297) );
  INV_X1 U5391 ( .A(n5297), .ZN(n4406) );
  MUX2_X1 U5392 ( .A(n5119), .B(n4350), .S(EBX_REG_24__SCAN_IN), .Z(n4405) );
  NAND2_X1 U5393 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5394 ( .A1(n4405), .A2(n4404), .ZN(n5296) );
  NAND2_X1 U5395 ( .A1(n4406), .A2(n5296), .ZN(n4407) );
  OR2_X2 U5396 ( .A1(n5299), .A2(n4407), .ZN(n5300) );
  MUX2_X1 U5397 ( .A(n5119), .B(n4350), .S(EBX_REG_26__SCAN_IN), .Z(n4409) );
  NAND2_X1 U5398 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4408) );
  MUX2_X1 U5399 ( .A(n5121), .B(n5119), .S(EBX_REG_27__SCAN_IN), .Z(n4411) );
  OR2_X1 U5400 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4410)
         );
  AND2_X1 U5401 ( .A1(n4411), .A2(n4410), .ZN(n5191) );
  AND2_X2 U5402 ( .A1(n5287), .A2(n5191), .ZN(n5193) );
  INV_X1 U5403 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U5404 ( .A1(n4350), .A2(n5376), .ZN(n4412) );
  OAI211_X1 U5405 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5126), .A(n4412), .B(n5119), 
        .ZN(n4414) );
  INV_X1 U5406 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U5407 ( .A1(n5316), .A2(n5280), .ZN(n4413) );
  NAND2_X1 U5408 ( .A1(n4414), .A2(n4413), .ZN(n5180) );
  NAND2_X2 U5409 ( .A1(n5193), .A2(n5180), .ZN(n5179) );
  NOR2_X1 U5410 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5120)
         );
  INV_X1 U5411 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5279) );
  AND2_X1 U5412 ( .A1(n4524), .A2(n5279), .ZN(n4415) );
  NOR2_X1 U5413 ( .A1(n4420), .A2(n5316), .ZN(n5124) );
  AND2_X1 U5414 ( .A1(n5126), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4416)
         );
  AOI21_X1 U5415 ( .B1(n5127), .B2(EBX_REG_30__SCAN_IN), .A(n4416), .ZN(n5125)
         );
  INV_X1 U5416 ( .A(n5125), .ZN(n4417) );
  OAI21_X1 U5417 ( .B1(n4420), .B2(n5179), .A(n4417), .ZN(n4421) );
  INV_X1 U5418 ( .A(n5179), .ZN(n4418) );
  OAI21_X1 U5419 ( .B1(n4418), .B2(n5119), .A(n5125), .ZN(n4419) );
  OAI22_X1 U5420 ( .A1(n5124), .A2(n4421), .B1(n4420), .B2(n4419), .ZN(n5277)
         );
  INV_X1 U5421 ( .A(n5277), .ZN(n5162) );
  NAND2_X1 U5422 ( .A1(n4274), .A2(n4443), .ZN(n6538) );
  OR2_X1 U5423 ( .A1(n4423), .A2(n4422), .ZN(n4424) );
  AND2_X1 U5424 ( .A1(n6538), .A2(n4424), .ZN(n4425) );
  NAND2_X1 U5425 ( .A1(n5162), .A2(n6023), .ZN(n4427) );
  OAI21_X1 U5426 ( .B1(n5090), .B2(n6018), .A(n4429), .ZN(U2988) );
  NAND2_X1 U5427 ( .A1(n4432), .A2(n4431), .ZN(n4433) );
  AND2_X1 U5428 ( .A1(n4430), .A2(n4433), .ZN(n5841) );
  INV_X1 U5429 ( .A(n5841), .ZN(n5328) );
  NAND2_X1 U5430 ( .A1(n4469), .A2(n6548), .ZN(n4466) );
  NOR3_X1 U5431 ( .A1(n6542), .A2(n6609), .A3(n6555), .ZN(n6541) );
  NAND2_X1 U5432 ( .A1(n4436), .A2(n4435), .ZN(n6552) );
  NAND2_X1 U5433 ( .A1(n6552), .A2(n5721), .ZN(n4437) );
  NOR2_X1 U5434 ( .A1(n4447), .A2(n5587), .ZN(n4438) );
  NOR2_X1 U5435 ( .A1(n5328), .A2(n5646), .ZN(n4465) );
  INV_X1 U5436 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6969) );
  INV_X1 U5437 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6588) );
  AND2_X2 U5438 ( .A1(n4922), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U5439 ( .A1(n6627), .A2(n6793), .ZN(n4457) );
  INV_X1 U5440 ( .A(n4457), .ZN(n4439) );
  AND3_X1 U5441 ( .A1(n4440), .A2(n4528), .A3(n4439), .ZN(n4441) );
  INV_X1 U5442 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6579) );
  NAND3_X1 U5443 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U5444 ( .A1(n6579), .A2(n4845), .ZN(n4449) );
  NAND2_X1 U5445 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n4450) );
  NOR2_X2 U5446 ( .A1(n5272), .A2(n4450), .ZN(n4856) );
  NAND3_X1 U5447 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4442) );
  NOR2_X2 U5448 ( .A1(n5802), .A2(n4442), .ZN(n5777) );
  NAND3_X1 U5449 ( .A1(n5777), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n5768) );
  NOR2_X2 U5450 ( .A1(n6588), .A2(n5768), .ZN(n5257) );
  NAND3_X1 U5451 ( .A1(n5257), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5229) );
  INV_X1 U5452 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U5453 ( .A1(n5147), .A2(n6764), .ZN(n5651) );
  INV_X1 U5454 ( .A(n5651), .ZN(n4464) );
  OR2_X1 U5455 ( .A1(n6564), .A2(n4457), .ZN(n6537) );
  AND2_X1 U5456 ( .A1(n4443), .A2(n6537), .ZN(n5141) );
  INV_X1 U5457 ( .A(n5141), .ZN(n4445) );
  INV_X1 U5458 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5275) );
  NAND3_X1 U5459 ( .A1(n4528), .A2(n4457), .A3(n5275), .ZN(n4444) );
  NAND2_X1 U5460 ( .A1(n4445), .A2(n4444), .ZN(n4446) );
  AND2_X2 U5461 ( .A1(n5142), .A2(n4446), .ZN(n5818) );
  NAND2_X1 U5462 ( .A1(n5140), .A2(n4922), .ZN(n5138) );
  NAND2_X1 U5463 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5776) );
  INV_X1 U5464 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6582) );
  NAND3_X1 U5465 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4449), .A3(n4922), .ZN(n4801) );
  NOR3_X1 U5466 ( .A1(n6582), .A2(n4450), .A3(n4801), .ZN(n4855) );
  NAND4_X1 U5467 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n4855), .ZN(n4994) );
  NOR3_X1 U5468 ( .A1(n6588), .A2(n5776), .A3(n4994), .ZN(n5235) );
  NAND4_X1 U5469 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5235), .ZN(n5130) );
  NAND2_X1 U5470 ( .A1(n5138), .A2(n5130), .ZN(n5652) );
  OAI22_X1 U5471 ( .A1(n5677), .A2(n5813), .B1(n6764), .B2(n5652), .ZN(n4451)
         );
  AOI21_X1 U5472 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5818), .A(n4451), .ZN(n4452)
         );
  INV_X1 U5473 ( .A(n4452), .ZN(n4463) );
  INV_X1 U5474 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4461) );
  MUX2_X1 U5475 ( .A(n5314), .B(n4453), .S(n5316), .Z(n4454) );
  INV_X1 U5476 ( .A(n4454), .ZN(n4455) );
  NAND2_X1 U5477 ( .A1(n5227), .A2(n4455), .ZN(n5326) );
  OR2_X1 U5478 ( .A1(n5227), .A2(n4455), .ZN(n4456) );
  NAND2_X1 U5479 ( .A1(n4457), .A2(EBX_REG_31__SCAN_IN), .ZN(n4458) );
  NOR2_X1 U5480 ( .A1(n5126), .A2(n4458), .ZN(n4459) );
  NAND2_X1 U5481 ( .A1(n5548), .A2(n5790), .ZN(n4460) );
  AND2_X1 U5482 ( .A1(n6612), .A2(n5587), .ZN(n4479) );
  NAND2_X1 U5483 ( .A1(n4922), .A2(n4479), .ZN(n5791) );
  OAI211_X1 U5484 ( .C1(n4461), .C2(n5794), .A(n4460), .B(n5791), .ZN(n4462)
         );
  INV_X1 U5485 ( .A(n4466), .ZN(n4468) );
  INV_X1 U5486 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6636) );
  INV_X1 U5487 ( .A(n4479), .ZN(n4467) );
  OAI211_X1 U5488 ( .C1(n4468), .C2(n6636), .A(n4543), .B(n4467), .ZN(U2788)
         );
  INV_X1 U5489 ( .A(n4284), .ZN(n4470) );
  OAI22_X1 U5490 ( .A1(n4501), .A2(n4799), .B1(n4469), .B2(n4470), .ZN(n5739)
         );
  AND2_X1 U5491 ( .A1(n5126), .A2(n4608), .ZN(n4481) );
  AOI21_X1 U5492 ( .B1(n4481), .B2(n6564), .A(READY_N), .ZN(n6629) );
  OR2_X1 U5493 ( .A1(n5739), .A2(n6629), .ZN(n6503) );
  AND2_X1 U5494 ( .A1(n6503), .A2(n6548), .ZN(n5744) );
  INV_X1 U5495 ( .A(MORE_REG_SCAN_IN), .ZN(n4478) );
  NOR2_X1 U5496 ( .A1(n4471), .A2(n4470), .ZN(n4476) );
  NAND2_X1 U5497 ( .A1(n4510), .A2(n4501), .ZN(n4475) );
  OR2_X1 U5498 ( .A1(n4473), .A2(n4472), .ZN(n4474) );
  OAI211_X1 U5499 ( .C1(n4476), .C2(n4501), .A(n4475), .B(n4474), .ZN(n6501)
         );
  NAND2_X1 U5500 ( .A1(n5744), .A2(n6501), .ZN(n4477) );
  OAI21_X1 U5501 ( .B1(n5744), .B2(n4478), .A(n4477), .ZN(U3471) );
  INV_X1 U5502 ( .A(n6625), .ZN(n4482) );
  OAI21_X1 U5503 ( .B1(n4479), .B2(READREQUEST_REG_SCAN_IN), .A(n4482), .ZN(
        n4480) );
  OAI21_X1 U5504 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(U3474) );
  INV_X1 U5505 ( .A(n5113), .ZN(n5732) );
  NAND2_X1 U5506 ( .A1(n6542), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6607) );
  INV_X1 U5507 ( .A(n4501), .ZN(n4511) );
  NAND2_X1 U5508 ( .A1(n4511), .A2(n4510), .ZN(n4493) );
  OAI21_X1 U5509 ( .B1(n6507), .B2(READY_N), .A(n4483), .ZN(n4485) );
  NAND2_X1 U5510 ( .A1(n4284), .A2(n6564), .ZN(n4484) );
  NAND2_X1 U5511 ( .A1(n4485), .A2(n4484), .ZN(n4486) );
  INV_X1 U5512 ( .A(n4612), .ZN(n4553) );
  NAND2_X1 U5513 ( .A1(n4486), .A2(n4553), .ZN(n4491) );
  INV_X1 U5514 ( .A(n4487), .ZN(n4488) );
  OAI211_X1 U5515 ( .C1(n4610), .C2(n4285), .A(n4489), .B(n4488), .ZN(n4490)
         );
  AOI21_X1 U5516 ( .B1(n4501), .B2(n4491), .A(n4490), .ZN(n4492) );
  OR2_X1 U5517 ( .A1(n6542), .A2(n6530), .ZN(n6606) );
  INV_X1 U5518 ( .A(n6606), .ZN(n4590) );
  AOI22_X1 U5519 ( .A1(n4578), .A2(n6548), .B1(n4590), .B2(FLUSH_REG_SCAN_IN), 
        .ZN(n5733) );
  NAND2_X1 U5520 ( .A1(n6607), .A2(n5733), .ZN(n5737) );
  OAI21_X1 U5521 ( .B1(n5732), .B2(n6507), .A(n5737), .ZN(n4504) );
  INV_X1 U5522 ( .A(n4274), .ZN(n4497) );
  INV_X1 U5523 ( .A(n4494), .ZN(n4495) );
  AND4_X1 U5524 ( .A1(n4497), .A2(n4496), .A3(n4495), .A4(n4285), .ZN(n4498)
         );
  NAND2_X1 U5525 ( .A1(n4499), .A2(n4498), .ZN(n5585) );
  NOR2_X1 U5526 ( .A1(n3713), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4500)
         );
  AOI21_X1 U5527 ( .B1(n6614), .B2(n5585), .A(n4500), .ZN(n6506) );
  AOI22_X1 U5528 ( .A1(n6508), .A2(n5590), .B1(n4308), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5529 ( .B1(n6506), .B2(n5732), .A(n4502), .ZN(n4503) );
  AOI22_X1 U5530 ( .A1(n4504), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n5737), .B2(n4503), .ZN(n4505) );
  INV_X1 U5531 ( .A(n4505), .ZN(U3461) );
  OR2_X1 U5532 ( .A1(n4507), .A2(n4506), .ZN(n4508) );
  NAND2_X1 U5533 ( .A1(n4509), .A2(n4508), .ZN(n5917) );
  NAND3_X1 U5534 ( .A1(n4511), .A2(n6548), .A3(n4510), .ZN(n4516) );
  AND4_X1 U5535 ( .A1(n4782), .A2(n5344), .A3(n6548), .A4(n4512), .ZN(n4513)
         );
  NAND2_X1 U5536 ( .A1(n4514), .A2(n4513), .ZN(n4607) );
  NAND2_X2 U5537 ( .A1(n5840), .A2(n5349), .ZN(n5343) );
  OR2_X1 U5538 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4518)
         );
  AND2_X1 U5539 ( .A1(n4518), .A2(n4517), .ZN(n6022) );
  INV_X1 U5540 ( .A(n6022), .ZN(n4864) );
  OAI222_X1 U5541 ( .A1(n5917), .A2(n5343), .B1(n5840), .B2(n4865), .C1(n4864), 
        .C2(n5336), .ZN(U2859) );
  NOR2_X1 U5542 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  NOR2_X1 U5543 ( .A1(n4522), .A2(n4521), .ZN(n4908) );
  INV_X1 U5544 ( .A(n4908), .ZN(n4929) );
  OAI21_X1 U5545 ( .B1(n4525), .B2(n4524), .A(n4523), .ZN(n6006) );
  AOI22_X1 U5546 ( .A1(n5836), .A2(n6006), .B1(n5341), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4526) );
  OAI21_X1 U5547 ( .B1(n4929), .B2(n5343), .A(n4526), .ZN(U2858) );
  INV_X1 U5548 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4531) );
  AND2_X1 U5549 ( .A1(n6538), .A2(n6507), .ZN(n4527) );
  NAND2_X1 U5550 ( .A1(n4529), .A2(n4528), .ZN(n4663) );
  AOI22_X1 U5551 ( .A1(n6534), .A2(UWORD_REG_14__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4530) );
  OAI21_X1 U5552 ( .B1(n4531), .B2(n4663), .A(n4530), .ZN(U2893) );
  INV_X1 U5553 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4533) );
  AOI22_X1 U5554 ( .A1(n6628), .A2(UWORD_REG_9__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4532) );
  OAI21_X1 U5555 ( .B1(n4533), .B2(n4663), .A(n4532), .ZN(U2898) );
  INV_X1 U5556 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5557 ( .A1(n6628), .A2(UWORD_REG_8__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4534) );
  OAI21_X1 U5558 ( .B1(n4535), .B2(n4663), .A(n4534), .ZN(U2899) );
  INV_X1 U5559 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U5560 ( .A1(n6628), .A2(UWORD_REG_10__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U5561 ( .B1(n4537), .B2(n4663), .A(n4536), .ZN(U2897) );
  INV_X1 U5562 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5563 ( .A1(n6628), .A2(UWORD_REG_11__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5564 ( .B1(n4539), .B2(n4663), .A(n4538), .ZN(U2896) );
  INV_X1 U5565 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5566 ( .A1(n6628), .A2(UWORD_REG_13__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4540) );
  OAI21_X1 U5567 ( .B1(n4541), .B2(n4663), .A(n4540), .ZN(U2894) );
  AOI22_X1 U5568 ( .A1(n6628), .A2(UWORD_REG_12__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4542) );
  OAI21_X1 U5569 ( .B1(n4159), .B2(n4663), .A(n4542), .ZN(U2895) );
  NAND2_X1 U5570 ( .A1(n4684), .A2(DATAI_5_), .ZN(n4687) );
  AOI22_X1 U5571 ( .A1(n3205), .A2(EAX_REG_5__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U5572 ( .A1(n4687), .A2(n4546), .ZN(U2944) );
  NAND2_X1 U5573 ( .A1(n4684), .A2(DATAI_10_), .ZN(n4678) );
  AOI22_X1 U5574 ( .A1(n3205), .A2(EAX_REG_10__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U5575 ( .A1(n4678), .A2(n4547), .ZN(U2949) );
  NAND2_X1 U5576 ( .A1(n4684), .A2(DATAI_12_), .ZN(n4670) );
  AOI22_X1 U5577 ( .A1(n3205), .A2(EAX_REG_12__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U5578 ( .A1(n4670), .A2(n4548), .ZN(U2951) );
  NAND2_X1 U5579 ( .A1(n4684), .A2(DATAI_11_), .ZN(n4668) );
  AOI22_X1 U5580 ( .A1(n3205), .A2(EAX_REG_11__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U5581 ( .A1(n4668), .A2(n4549), .ZN(U2950) );
  NAND2_X1 U5582 ( .A1(n4684), .A2(DATAI_9_), .ZN(n4676) );
  AOI22_X1 U5583 ( .A1(n3205), .A2(EAX_REG_9__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5584 ( .A1(n4676), .A2(n4550), .ZN(U2948) );
  NAND2_X1 U5585 ( .A1(n4684), .A2(DATAI_7_), .ZN(n4691) );
  AOI22_X1 U5586 ( .A1(n3205), .A2(EAX_REG_7__SCAN_IN), .B1(n4665), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5587 ( .A1(n4691), .A2(n4551), .ZN(U2946) );
  NAND2_X1 U5588 ( .A1(n6392), .A2(n5585), .ZN(n4569) );
  NAND2_X1 U5589 ( .A1(n4554), .A2(n4553), .ZN(n4575) );
  MUX2_X1 U5590 ( .A(n4556), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4555), 
        .Z(n4558) );
  NOR2_X1 U5591 ( .A1(n4558), .A2(n4557), .ZN(n4567) );
  NAND2_X1 U5592 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4559) );
  XNOR2_X1 U5593 ( .A(n4562), .B(n4559), .ZN(n4565) );
  INV_X1 U5594 ( .A(n4560), .ZN(n4561) );
  OAI21_X1 U5595 ( .B1(n4555), .B2(n4562), .A(n4561), .ZN(n4564) );
  NOR2_X1 U5596 ( .A1(n4564), .A2(n4563), .ZN(n5596) );
  OAI22_X1 U5597 ( .A1(n6507), .A2(n4565), .B1(n5596), .B2(n4571), .ZN(n4566)
         );
  AOI21_X1 U5598 ( .B1(n4575), .B2(n4567), .A(n4566), .ZN(n4568) );
  NAND2_X1 U5599 ( .A1(n4569), .A2(n4568), .ZN(n5595) );
  MUX2_X1 U5600 ( .A(n5595), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6515), 
        .Z(n6526) );
  INV_X1 U5601 ( .A(n5585), .ZN(n4577) );
  XNOR2_X1 U5602 ( .A(n4555), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4574)
         );
  XNOR2_X1 U5603 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4572) );
  OAI22_X1 U5604 ( .A1(n6507), .A2(n4572), .B1(n4571), .B2(n4574), .ZN(n4573)
         );
  AOI21_X1 U5605 ( .B1(n4575), .B2(n4574), .A(n4573), .ZN(n4576) );
  OAI21_X1 U5606 ( .B1(n6030), .B2(n4577), .A(n4576), .ZN(n5114) );
  MUX2_X1 U5607 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5114), .S(n4578), 
        .Z(n6520) );
  NAND3_X1 U5608 ( .A1(n6526), .A2(n6520), .A3(n5587), .ZN(n4581) );
  INV_X1 U5609 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6721) );
  AND2_X1 U5610 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6721), .ZN(n4579) );
  NAND2_X1 U5611 ( .A1(n4557), .A2(n4579), .ZN(n4580) );
  NAND2_X1 U5612 ( .A1(n4581), .A2(n4580), .ZN(n6499) );
  INV_X1 U5613 ( .A(n4582), .ZN(n4583) );
  NAND2_X1 U5614 ( .A1(n6499), .A2(n4583), .ZN(n6533) );
  INV_X1 U5615 ( .A(n4584), .ZN(n6327) );
  NOR2_X1 U5616 ( .A1(n4585), .A2(n6327), .ZN(n4586) );
  XNOR2_X1 U5617 ( .A(n4586), .B(n5736), .ZN(n4840) );
  INV_X1 U5618 ( .A(n4285), .ZN(n4606) );
  NAND2_X1 U5619 ( .A1(n4840), .A2(n4606), .ZN(n5734) );
  OR2_X1 U5620 ( .A1(n5734), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4589) );
  MUX2_X1 U5621 ( .A(n6515), .B(n6721), .S(STATE2_REG_1__SCAN_IN), .Z(n4587)
         );
  NAND2_X1 U5622 ( .A1(n4587), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4588) );
  NAND3_X1 U5623 ( .A1(n6533), .A2(n6721), .A3(n6532), .ZN(n4591) );
  NAND2_X1 U5624 ( .A1(n4591), .A2(n4590), .ZN(n4592) );
  NAND2_X1 U5625 ( .A1(n4592), .A2(n6208), .ZN(n6610) );
  NAND2_X1 U5626 ( .A1(n6360), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6356) );
  AND2_X1 U5627 ( .A1(n6356), .A2(n6240), .ZN(n4876) );
  INV_X1 U5628 ( .A(n6027), .ZN(n4596) );
  NAND2_X1 U5629 ( .A1(n6202), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5578) );
  NOR2_X1 U5630 ( .A1(n5578), .A2(n6383), .ZN(n4595) );
  NAND2_X1 U5631 ( .A1(n4596), .A2(n4595), .ZN(n4637) );
  AOI21_X1 U5632 ( .B1(n4876), .B2(n4637), .A(n6438), .ZN(n4598) );
  INV_X1 U5633 ( .A(n4594), .ZN(n4745) );
  AND2_X1 U5634 ( .A1(n6612), .A2(n6793), .ZN(n6443) );
  INV_X1 U5635 ( .A(n6443), .ZN(n6162) );
  INV_X1 U5636 ( .A(n6392), .ZN(n6207) );
  NAND2_X1 U5637 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6609), .ZN(n6613) );
  INV_X1 U5638 ( .A(n6613), .ZN(n5579) );
  OAI22_X1 U5639 ( .A1(n4745), .A2(n6162), .B1(n6207), .B2(n5579), .ZN(n4597)
         );
  OAI21_X1 U5640 ( .B1(n4598), .B2(n4597), .A(n6610), .ZN(n4599) );
  OAI21_X1 U5641 ( .B1(n6610), .B2(n6525), .A(n4599), .ZN(U3462) );
  NOR2_X1 U5642 ( .A1(n4602), .A2(n4601), .ZN(n4603) );
  NOR2_X1 U5643 ( .A1(n4600), .A2(n4603), .ZN(n5911) );
  INV_X1 U5644 ( .A(n5911), .ZN(n4839) );
  XNOR2_X1 U5645 ( .A(n4621), .B(n4618), .ZN(n5991) );
  AOI22_X1 U5646 ( .A1(n5836), .A2(n5991), .B1(n5341), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4604) );
  OAI21_X1 U5647 ( .B1(n4839), .B2(n5343), .A(n4604), .ZN(U2857) );
  INV_X1 U5648 ( .A(n4605), .ZN(n4613) );
  NAND2_X1 U5649 ( .A1(n4606), .A2(n6548), .ZN(n4609) );
  OAI22_X1 U5650 ( .A1(n4610), .A2(n4609), .B1(n4608), .B2(n4607), .ZN(n4611)
         );
  NAND2_X1 U5651 ( .A1(n4615), .A2(n5349), .ZN(n4616) );
  INV_X1 U5652 ( .A(n4616), .ZN(n4617) );
  INV_X1 U5653 ( .A(DATAI_1_), .ZN(n6859) );
  INV_X1 U5654 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5882) );
  OAI222_X1 U5655 ( .A1(n4929), .A2(n5653), .B1(n5371), .B2(n6859), .C1(n5369), 
        .C2(n5882), .ZN(U2890) );
  INV_X1 U5656 ( .A(DATAI_0_), .ZN(n6972) );
  INV_X1 U5657 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5886) );
  OAI222_X1 U5658 ( .A1(n5917), .A2(n5653), .B1(n5371), .B2(n6972), .C1(n5369), 
        .C2(n5886), .ZN(U2891) );
  INV_X1 U5659 ( .A(DATAI_2_), .ZN(n6873) );
  INV_X1 U5660 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5879) );
  OAI222_X1 U5661 ( .A1(n4839), .A2(n5653), .B1(n5371), .B2(n6873), .C1(n5369), 
        .C2(n5879), .ZN(U2889) );
  INV_X1 U5662 ( .A(n4618), .ZN(n4620) );
  OAI21_X1 U5663 ( .B1(n4621), .B2(n4620), .A(n4619), .ZN(n4622) );
  NAND2_X1 U5664 ( .A1(n4622), .A2(n4717), .ZN(n5982) );
  INV_X1 U5665 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5666 ( .B1(n4600), .B2(n4624), .A(n4623), .ZN(n5816) );
  OAI222_X1 U5667 ( .A1(n5982), .A2(n5336), .B1(n4625), .B2(n5840), .C1(n5816), 
        .C2(n5343), .ZN(U2856) );
  INV_X1 U5668 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5669 ( .A1(n6534), .A2(UWORD_REG_3__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4626) );
  OAI21_X1 U5670 ( .B1(n4627), .B2(n4663), .A(n4626), .ZN(U2904) );
  INV_X1 U5671 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5672 ( .A1(n6534), .A2(UWORD_REG_1__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U5673 ( .B1(n4629), .B2(n4663), .A(n4628), .ZN(U2906) );
  INV_X1 U5674 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4631) );
  AOI22_X1 U5675 ( .A1(n6534), .A2(UWORD_REG_4__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4630) );
  OAI21_X1 U5676 ( .B1(n4631), .B2(n4663), .A(n4630), .ZN(U2903) );
  INV_X1 U5677 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5678 ( .A1(n6534), .A2(UWORD_REG_2__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U5679 ( .B1(n4633), .B2(n4663), .A(n4632), .ZN(U2905) );
  INV_X1 U5680 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5681 ( .A1(n6534), .A2(UWORD_REG_0__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4634) );
  OAI21_X1 U5682 ( .B1(n4635), .B2(n4663), .A(n4634), .ZN(U2907) );
  NOR2_X2 U5683 ( .A1(n4791), .A2(n5344), .ZN(n6491) );
  INV_X1 U5684 ( .A(n6491), .ZN(n6274) );
  NAND2_X1 U5685 ( .A1(n6612), .A2(n4637), .ZN(n4642) );
  NAND3_X1 U5686 ( .A1(n6434), .A2(n6327), .A3(n6614), .ZN(n4639) );
  AND2_X1 U5687 ( .A1(n4639), .A2(n6187), .ZN(n4643) );
  INV_X1 U5688 ( .A(n4643), .ZN(n4641) );
  AOI21_X1 U5689 ( .B1(n6159), .B2(n6438), .A(n6129), .ZN(n4640) );
  OAI21_X1 U5690 ( .B1(n4642), .B2(n4641), .A(n4640), .ZN(n6198) );
  INV_X1 U5691 ( .A(DATAI_7_), .ZN(n5370) );
  NOR2_X2 U5692 ( .A1(n5370), .A2(n6208), .ZN(n6489) );
  OAI22_X1 U5693 ( .A1(n4643), .A2(n4642), .B1(n6436), .B2(n6159), .ZN(n6197)
         );
  AOI22_X1 U5694 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6198), .B1(n6489), 
        .B2(n6197), .ZN(n4648) );
  INV_X1 U5695 ( .A(DATAI_31_), .ZN(n4645) );
  NOR2_X1 U5696 ( .A1(n4644), .A2(n4645), .ZN(n6428) );
  INV_X1 U5697 ( .A(n6383), .ZN(n4746) );
  NAND2_X1 U5698 ( .A1(n6384), .A2(n4746), .ZN(n4646) );
  INV_X1 U5699 ( .A(n6201), .ZN(n4655) );
  OR2_X1 U5700 ( .A1(n4646), .A2(n6361), .ZN(n6205) );
  INV_X1 U5701 ( .A(DATAI_23_), .ZN(n6995) );
  NOR2_X1 U5702 ( .A1(n4644), .A2(n6995), .ZN(n6493) );
  AOI22_X1 U5703 ( .A1(n6428), .A2(n4655), .B1(n6229), .B2(n6493), .ZN(n4647)
         );
  OAI211_X1 U5704 ( .C1(n6187), .C2(n6274), .A(n4648), .B(n4647), .ZN(U3083)
         );
  NOR2_X2 U5705 ( .A1(n4791), .A2(n4649), .ZN(n6459) );
  INV_X1 U5706 ( .A(n6459), .ZN(n6253) );
  NOR2_X2 U5707 ( .A1(n6873), .A2(n6208), .ZN(n6458) );
  AOI22_X1 U5708 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6198), .B1(n6458), 
        .B2(n6197), .ZN(n4652) );
  INV_X1 U5709 ( .A(DATAI_26_), .ZN(n4650) );
  NOR2_X1 U5710 ( .A1(n4644), .A2(n4650), .ZN(n6405) );
  INV_X1 U5711 ( .A(DATAI_18_), .ZN(n6958) );
  NOR2_X1 U5712 ( .A1(n4644), .A2(n6958), .ZN(n6460) );
  AOI22_X1 U5713 ( .A1(n6405), .A2(n4655), .B1(n6229), .B2(n6460), .ZN(n4651)
         );
  OAI211_X1 U5714 ( .C1(n6187), .C2(n6253), .A(n4652), .B(n4651), .ZN(U3078)
         );
  NOR2_X2 U5715 ( .A1(n4791), .A2(n4653), .ZN(n6440) );
  INV_X1 U5716 ( .A(n6440), .ZN(n6234) );
  NOR2_X2 U5717 ( .A1(n6972), .A2(n6208), .ZN(n6439) );
  AOI22_X1 U5718 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6198), .B1(n6439), 
        .B2(n6197), .ZN(n4657) );
  INV_X1 U5719 ( .A(DATAI_24_), .ZN(n4654) );
  NOR2_X1 U5720 ( .A1(n4644), .A2(n4654), .ZN(n6397) );
  INV_X1 U5721 ( .A(DATAI_16_), .ZN(n6725) );
  NOR2_X1 U5722 ( .A1(n4644), .A2(n6725), .ZN(n6448) );
  AOI22_X1 U5723 ( .A1(n6397), .A2(n4655), .B1(n6229), .B2(n6448), .ZN(n4656)
         );
  OAI211_X1 U5724 ( .C1(n6187), .C2(n6234), .A(n4657), .B(n4656), .ZN(U3076)
         );
  INV_X1 U5725 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5726 ( .A1(n6628), .A2(UWORD_REG_7__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4658) );
  OAI21_X1 U5727 ( .B1(n4659), .B2(n4663), .A(n4658), .ZN(U2900) );
  INV_X1 U5728 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5729 ( .A1(n6628), .A2(UWORD_REG_6__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4660) );
  OAI21_X1 U5730 ( .B1(n4661), .B2(n4663), .A(n4660), .ZN(U2901) );
  INV_X1 U5731 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5732 ( .A1(n6628), .A2(UWORD_REG_5__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5733 ( .B1(n4664), .B2(n4663), .A(n4662), .ZN(U2902) );
  NAND2_X1 U5734 ( .A1(n4684), .A2(DATAI_4_), .ZN(n4699) );
  AOI22_X1 U5735 ( .A1(n3205), .A2(EAX_REG_20__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U5736 ( .A1(n4699), .A2(n4666), .ZN(U2928) );
  AOI22_X1 U5737 ( .A1(n3205), .A2(EAX_REG_27__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5738 ( .A1(n4668), .A2(n4667), .ZN(U2935) );
  AOI22_X1 U5739 ( .A1(n3205), .A2(EAX_REG_28__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5740 ( .A1(n4670), .A2(n4669), .ZN(U2936) );
  NAND2_X1 U5741 ( .A1(n4684), .A2(DATAI_2_), .ZN(n4705) );
  AOI22_X1 U5742 ( .A1(n3205), .A2(EAX_REG_18__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5743 ( .A1(n4705), .A2(n4671), .ZN(U2926) );
  NAND2_X1 U5744 ( .A1(n4684), .A2(DATAI_14_), .ZN(n4697) );
  AOI22_X1 U5745 ( .A1(n3205), .A2(EAX_REG_30__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5746 ( .A1(n4697), .A2(n4672), .ZN(U2938) );
  NAND2_X1 U5747 ( .A1(n4684), .A2(DATAI_0_), .ZN(n4680) );
  AOI22_X1 U5748 ( .A1(n3205), .A2(EAX_REG_0__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5749 ( .A1(n4680), .A2(n4673), .ZN(U2939) );
  NAND2_X1 U5750 ( .A1(n4684), .A2(DATAI_13_), .ZN(n4695) );
  AOI22_X1 U5751 ( .A1(n3205), .A2(EAX_REG_29__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5752 ( .A1(n4695), .A2(n4674), .ZN(U2937) );
  AOI22_X1 U5753 ( .A1(n3205), .A2(EAX_REG_25__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U5754 ( .A1(n4676), .A2(n4675), .ZN(U2933) );
  AOI22_X1 U5755 ( .A1(n3205), .A2(EAX_REG_26__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U5756 ( .A1(n4678), .A2(n4677), .ZN(U2934) );
  AOI22_X1 U5757 ( .A1(n3205), .A2(EAX_REG_16__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5758 ( .A1(n4680), .A2(n4679), .ZN(U2924) );
  NAND2_X1 U5759 ( .A1(n4684), .A2(DATAI_1_), .ZN(n4703) );
  AOI22_X1 U5760 ( .A1(n3205), .A2(EAX_REG_17__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U5761 ( .A1(n4703), .A2(n4681), .ZN(U2925) );
  NAND2_X1 U5762 ( .A1(n4684), .A2(DATAI_6_), .ZN(n4689) );
  AOI22_X1 U5763 ( .A1(n3205), .A2(EAX_REG_6__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5764 ( .A1(n4689), .A2(n4682), .ZN(U2945) );
  NAND2_X1 U5765 ( .A1(n4684), .A2(DATAI_3_), .ZN(n4701) );
  AOI22_X1 U5766 ( .A1(n3205), .A2(EAX_REG_19__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5767 ( .A1(n4701), .A2(n4683), .ZN(U2927) );
  NAND2_X1 U5768 ( .A1(n4684), .A2(DATAI_8_), .ZN(n4693) );
  AOI22_X1 U5769 ( .A1(n3205), .A2(EAX_REG_8__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U5770 ( .A1(n4693), .A2(n4685), .ZN(U2947) );
  AOI22_X1 U5771 ( .A1(n3205), .A2(EAX_REG_21__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U5772 ( .A1(n4687), .A2(n4686), .ZN(U2929) );
  AOI22_X1 U5773 ( .A1(n3205), .A2(EAX_REG_22__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5774 ( .A1(n4689), .A2(n4688), .ZN(U2930) );
  AOI22_X1 U5775 ( .A1(n3205), .A2(EAX_REG_23__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5776 ( .A1(n4691), .A2(n4690), .ZN(U2931) );
  AOI22_X1 U5777 ( .A1(n3205), .A2(EAX_REG_24__SCAN_IN), .B1(n4706), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U5778 ( .A1(n4693), .A2(n4692), .ZN(U2932) );
  AOI22_X1 U5779 ( .A1(n3205), .A2(EAX_REG_13__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U5780 ( .A1(n4695), .A2(n4694), .ZN(U2952) );
  AOI22_X1 U5781 ( .A1(n3205), .A2(EAX_REG_14__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U5782 ( .A1(n4697), .A2(n4696), .ZN(U2953) );
  AOI22_X1 U5783 ( .A1(n3205), .A2(EAX_REG_4__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5784 ( .A1(n4699), .A2(n4698), .ZN(U2943) );
  AOI22_X1 U5785 ( .A1(n3205), .A2(EAX_REG_3__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5786 ( .A1(n4701), .A2(n4700), .ZN(U2942) );
  AOI22_X1 U5787 ( .A1(n3205), .A2(EAX_REG_1__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5788 ( .A1(n4703), .A2(n4702), .ZN(U2940) );
  AOI22_X1 U5789 ( .A1(n3205), .A2(EAX_REG_2__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5790 ( .A1(n4705), .A2(n4704), .ZN(U2941) );
  INV_X1 U5791 ( .A(DATAI_15_), .ZN(n6927) );
  AOI22_X1 U5792 ( .A1(n3205), .A2(EAX_REG_15__SCAN_IN), .B1(n4706), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4707) );
  OAI21_X1 U5793 ( .B1(n4708), .B2(n6927), .A(n4707), .ZN(U2954) );
  OAI21_X1 U5794 ( .B1(n4709), .B2(n4711), .A(n4710), .ZN(n4916) );
  NOR2_X1 U5795 ( .A1(n4719), .A2(n4712), .ZN(n4713) );
  AOI22_X1 U5796 ( .A1(n5836), .A2(n3201), .B1(n5341), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4714) );
  OAI21_X1 U5797 ( .B1(n4916), .B2(n5343), .A(n4714), .ZN(U2854) );
  INV_X1 U5798 ( .A(DATAI_3_), .ZN(n6997) );
  INV_X1 U5799 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5877) );
  OAI222_X1 U5800 ( .A1(n5816), .A2(n5653), .B1(n5371), .B2(n6997), .C1(n5369), 
        .C2(n5877), .ZN(U2888) );
  AOI21_X1 U5801 ( .B1(n4715), .B2(n4623), .A(n4709), .ZN(n4970) );
  INV_X1 U5802 ( .A(n4970), .ZN(n4853) );
  AND2_X1 U5803 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  NOR2_X1 U5804 ( .A1(n4719), .A2(n4718), .ZN(n5976) );
  AOI22_X1 U5805 ( .A1(n5836), .A2(n5976), .B1(n5341), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4720) );
  OAI21_X1 U5806 ( .B1(n4853), .B2(n5343), .A(n4720), .ZN(U2855) );
  INV_X1 U5807 ( .A(n6428), .ZN(n6498) );
  NAND2_X1 U5808 ( .A1(n6202), .A2(n6361), .ZN(n4721) );
  NAND2_X1 U5809 ( .A1(n4871), .A2(n6392), .ZN(n6289) );
  INV_X1 U5810 ( .A(n6614), .ZN(n6125) );
  OR2_X1 U5811 ( .A1(n6289), .A2(n6125), .ZN(n4723) );
  NOR2_X1 U5812 ( .A1(n4872), .A2(n6525), .ZN(n6316) );
  INV_X1 U5813 ( .A(n6316), .ZN(n4722) );
  AND2_X1 U5814 ( .A1(n4723), .A2(n4722), .ZN(n4727) );
  INV_X1 U5815 ( .A(n4727), .ZN(n4725) );
  OAI21_X1 U5816 ( .B1(n6240), .B2(n5578), .A(n6612), .ZN(n4726) );
  NAND3_X1 U5817 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6517), .ZN(n6281) );
  AOI21_X1 U5818 ( .B1(n6438), .B2(n6281), .A(n6129), .ZN(n4724) );
  OAI21_X1 U5819 ( .B1(n4725), .B2(n4726), .A(n4724), .ZN(n6318) );
  OAI22_X1 U5820 ( .A1(n4727), .A2(n4726), .B1(n6436), .B2(n6281), .ZN(n6317)
         );
  AOI22_X1 U5821 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6318), .B1(n6489), 
        .B2(n6317), .ZN(n4730) );
  NAND2_X1 U5822 ( .A1(n6202), .A2(n6611), .ZN(n4728) );
  AOI22_X1 U5823 ( .A1(n6349), .A2(n6493), .B1(n6491), .B2(n6316), .ZN(n4729)
         );
  OAI211_X1 U5824 ( .C1(n6498), .C2(n6321), .A(n4730), .B(n4729), .ZN(U3115)
         );
  INV_X1 U5825 ( .A(DATAI_25_), .ZN(n4731) );
  NOR2_X1 U5826 ( .A1(n4644), .A2(n4731), .ZN(n6401) );
  INV_X1 U5827 ( .A(n6401), .ZN(n6457) );
  NOR2_X2 U5828 ( .A1(n6859), .A2(n6208), .ZN(n6452) );
  AOI22_X1 U5829 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6318), .B1(n6452), 
        .B2(n6317), .ZN(n4735) );
  INV_X1 U5830 ( .A(DATAI_17_), .ZN(n4732) );
  NOR2_X1 U5831 ( .A1(n4644), .A2(n4732), .ZN(n6454) );
  NOR2_X2 U5832 ( .A1(n4791), .A2(n4733), .ZN(n6453) );
  AOI22_X1 U5833 ( .A1(n6349), .A2(n6454), .B1(n6453), .B2(n6316), .ZN(n4734)
         );
  OAI211_X1 U5834 ( .C1(n6457), .C2(n6321), .A(n4735), .B(n4734), .ZN(U3109)
         );
  INV_X1 U5835 ( .A(DATAI_27_), .ZN(n4736) );
  NOR2_X1 U5836 ( .A1(n4644), .A2(n4736), .ZN(n6409) );
  INV_X1 U5837 ( .A(n6409), .ZN(n6469) );
  NOR2_X2 U5838 ( .A1(n6997), .A2(n6208), .ZN(n6464) );
  AOI22_X1 U5839 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6318), .B1(n6464), 
        .B2(n6317), .ZN(n4740) );
  INV_X1 U5840 ( .A(DATAI_19_), .ZN(n4737) );
  NOR2_X1 U5841 ( .A1(n4644), .A2(n4737), .ZN(n6466) );
  NOR2_X2 U5842 ( .A1(n4791), .A2(n4738), .ZN(n6465) );
  AOI22_X1 U5843 ( .A1(n6349), .A2(n6466), .B1(n6465), .B2(n6316), .ZN(n4739)
         );
  OAI211_X1 U5844 ( .C1(n6469), .C2(n6321), .A(n4740), .B(n4739), .ZN(U3111)
         );
  AOI22_X1 U5845 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6318), .B1(n6439), 
        .B2(n6317), .ZN(n4742) );
  AOI22_X1 U5846 ( .A1(n6349), .A2(n6448), .B1(n6440), .B2(n6316), .ZN(n4741)
         );
  OAI211_X1 U5847 ( .C1(n6451), .C2(n6321), .A(n4742), .B(n4741), .ZN(U3108)
         );
  INV_X1 U5848 ( .A(n6405), .ZN(n6463) );
  AOI22_X1 U5849 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6318), .B1(n6458), 
        .B2(n6317), .ZN(n4744) );
  AOI22_X1 U5850 ( .A1(n6349), .A2(n6460), .B1(n6459), .B2(n6316), .ZN(n4743)
         );
  OAI211_X1 U5851 ( .C1(n6463), .C2(n6321), .A(n4744), .B(n4743), .ZN(U3110)
         );
  INV_X1 U5852 ( .A(DATAI_4_), .ZN(n6790) );
  INV_X1 U5853 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5875) );
  OAI222_X1 U5854 ( .A1(n4853), .A2(n5653), .B1(n5371), .B2(n6790), .C1(n5369), 
        .C2(n5875), .ZN(U2887) );
  NAND3_X1 U5855 ( .A1(n4745), .A2(n6027), .A3(n6202), .ZN(n4870) );
  NAND2_X1 U5856 ( .A1(n4747), .A2(n4746), .ZN(n6124) );
  OR2_X1 U5857 ( .A1(n6124), .A2(n6793), .ZN(n4748) );
  NAND2_X1 U5858 ( .A1(n4748), .A2(n6612), .ZN(n6133) );
  INV_X1 U5859 ( .A(n6133), .ZN(n4749) );
  NAND2_X1 U5860 ( .A1(n6353), .A2(n6327), .ZN(n6126) );
  OAI211_X1 U5861 ( .C1(n4798), .C2(n6443), .A(n4749), .B(n6126), .ZN(n4752)
         );
  NAND2_X1 U5862 ( .A1(n6512), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6354) );
  OR2_X1 U5863 ( .A1(n6354), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6132)
         );
  NOR2_X1 U5864 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6132), .ZN(n4795)
         );
  INV_X1 U5865 ( .A(n4795), .ZN(n4750) );
  NOR2_X1 U5866 ( .A1(n6155), .A2(n6436), .ZN(n6287) );
  NOR2_X1 U5867 ( .A1(n6385), .A2(n6203), .ZN(n6031) );
  OAI21_X1 U5868 ( .B1(n6031), .B2(n6436), .A(n6101), .ZN(n6036) );
  AOI211_X1 U5869 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4750), .A(n6287), .B(
        n6036), .ZN(n4751) );
  NAND2_X1 U5870 ( .A1(n4789), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4758) );
  INV_X1 U5871 ( .A(n6466), .ZN(n6412) );
  NAND3_X1 U5872 ( .A1(n6207), .A2(n6612), .A3(n6353), .ZN(n4754) );
  AND2_X1 U5873 ( .A1(n6155), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U5874 ( .A1(n6031), .A2(n6386), .ZN(n4753) );
  INV_X1 U5875 ( .A(n6464), .ZN(n4755) );
  OAI22_X1 U5876 ( .A1(n6154), .A2(n6412), .B1(n4793), .B2(n4755), .ZN(n4756)
         );
  AOI21_X1 U5877 ( .B1(n6465), .B2(n4795), .A(n4756), .ZN(n4757) );
  OAI211_X1 U5878 ( .C1(n6469), .C2(n4798), .A(n4758), .B(n4757), .ZN(U3055)
         );
  NAND2_X1 U5879 ( .A1(n4789), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4762) );
  INV_X1 U5880 ( .A(n6448), .ZN(n6400) );
  INV_X1 U5881 ( .A(n6439), .ZN(n4759) );
  OAI22_X1 U5882 ( .A1(n6154), .A2(n6400), .B1(n4793), .B2(n4759), .ZN(n4760)
         );
  AOI21_X1 U5883 ( .B1(n6440), .B2(n4795), .A(n4760), .ZN(n4761) );
  OAI211_X1 U5884 ( .C1(n4798), .C2(n6451), .A(n4762), .B(n4761), .ZN(U3052)
         );
  INV_X1 U5885 ( .A(DATAI_29_), .ZN(n4763) );
  NOR2_X1 U5886 ( .A1(n4644), .A2(n4763), .ZN(n6417) );
  INV_X1 U5887 ( .A(n6417), .ZN(n6481) );
  NAND2_X1 U5888 ( .A1(n4789), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4768) );
  NOR2_X2 U5889 ( .A1(n4791), .A2(n5350), .ZN(n6477) );
  INV_X1 U5890 ( .A(DATAI_21_), .ZN(n4764) );
  NOR2_X1 U5891 ( .A1(n4644), .A2(n4764), .ZN(n6478) );
  INV_X1 U5892 ( .A(n6478), .ZN(n6420) );
  INV_X1 U5893 ( .A(DATAI_5_), .ZN(n6735) );
  NOR2_X2 U5894 ( .A1(n6735), .A2(n6208), .ZN(n6476) );
  INV_X1 U5895 ( .A(n6476), .ZN(n4765) );
  OAI22_X1 U5896 ( .A1(n6154), .A2(n6420), .B1(n4793), .B2(n4765), .ZN(n4766)
         );
  AOI21_X1 U5897 ( .B1(n6477), .B2(n4795), .A(n4766), .ZN(n4767) );
  OAI211_X1 U5898 ( .C1(n6481), .C2(n4798), .A(n4768), .B(n4767), .ZN(U3057)
         );
  NAND2_X1 U5899 ( .A1(n4789), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4772) );
  INV_X1 U5900 ( .A(n6460), .ZN(n6408) );
  INV_X1 U5901 ( .A(n6458), .ZN(n4769) );
  OAI22_X1 U5902 ( .A1(n6154), .A2(n6408), .B1(n4793), .B2(n4769), .ZN(n4770)
         );
  AOI21_X1 U5903 ( .B1(n6459), .B2(n4795), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5904 ( .C1(n6463), .C2(n4798), .A(n4772), .B(n4771), .ZN(U3054)
         );
  NAND2_X1 U5905 ( .A1(n4789), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4776) );
  INV_X1 U5906 ( .A(n6493), .ZN(n6432) );
  INV_X1 U5907 ( .A(n6489), .ZN(n4773) );
  OAI22_X1 U5908 ( .A1(n6154), .A2(n6432), .B1(n4793), .B2(n4773), .ZN(n4774)
         );
  AOI21_X1 U5909 ( .B1(n6491), .B2(n4795), .A(n4774), .ZN(n4775) );
  OAI211_X1 U5910 ( .C1(n6498), .C2(n4798), .A(n4776), .B(n4775), .ZN(U3059)
         );
  NAND2_X1 U5911 ( .A1(n4789), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4780) );
  INV_X1 U5912 ( .A(n6454), .ZN(n6404) );
  INV_X1 U5913 ( .A(n6452), .ZN(n4777) );
  OAI22_X1 U5914 ( .A1(n6154), .A2(n6404), .B1(n4793), .B2(n4777), .ZN(n4778)
         );
  AOI21_X1 U5915 ( .B1(n6453), .B2(n4795), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5916 ( .C1(n6457), .C2(n4798), .A(n4780), .B(n4779), .ZN(U3053)
         );
  INV_X1 U5917 ( .A(DATAI_28_), .ZN(n4781) );
  NOR2_X1 U5918 ( .A1(n4644), .A2(n4781), .ZN(n6413) );
  NAND2_X1 U5919 ( .A1(n4789), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4787) );
  NOR2_X2 U5920 ( .A1(n4791), .A2(n4782), .ZN(n6471) );
  INV_X1 U5921 ( .A(DATAI_20_), .ZN(n4783) );
  NOR2_X1 U5922 ( .A1(n4644), .A2(n4783), .ZN(n6472) );
  INV_X1 U5923 ( .A(n6472), .ZN(n6416) );
  NOR2_X2 U5924 ( .A1(n6790), .A2(n6208), .ZN(n6470) );
  INV_X1 U5925 ( .A(n6470), .ZN(n4784) );
  OAI22_X1 U5926 ( .A1(n6154), .A2(n6416), .B1(n4793), .B2(n4784), .ZN(n4785)
         );
  AOI21_X1 U5927 ( .B1(n6471), .B2(n4795), .A(n4785), .ZN(n4786) );
  OAI211_X1 U5928 ( .C1(n6475), .C2(n4798), .A(n4787), .B(n4786), .ZN(U3056)
         );
  INV_X1 U5929 ( .A(DATAI_30_), .ZN(n4788) );
  NOR2_X1 U5930 ( .A1(n4644), .A2(n4788), .ZN(n6421) );
  INV_X1 U5931 ( .A(n6421), .ZN(n6487) );
  NAND2_X1 U5932 ( .A1(n4789), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4797) );
  NOR2_X2 U5933 ( .A1(n4791), .A2(n4790), .ZN(n6483) );
  INV_X1 U5934 ( .A(DATAI_22_), .ZN(n6715) );
  NOR2_X1 U5935 ( .A1(n4644), .A2(n6715), .ZN(n6484) );
  INV_X1 U5936 ( .A(n6484), .ZN(n6424) );
  INV_X1 U5937 ( .A(DATAI_6_), .ZN(n6955) );
  NOR2_X2 U5938 ( .A1(n6955), .A2(n6208), .ZN(n6482) );
  INV_X1 U5939 ( .A(n6482), .ZN(n4792) );
  OAI22_X1 U5940 ( .A1(n6154), .A2(n6424), .B1(n4793), .B2(n4792), .ZN(n4794)
         );
  AOI21_X1 U5941 ( .B1(n6483), .B2(n4795), .A(n4794), .ZN(n4796) );
  OAI211_X1 U5942 ( .C1(n6487), .C2(n4798), .A(n4797), .B(n4796), .ZN(U3058)
         );
  INV_X1 U5943 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5873) );
  OAI222_X1 U5944 ( .A1(n4916), .A2(n5653), .B1(n5371), .B2(n6735), .C1(n5369), 
        .C2(n5873), .ZN(U2886) );
  NAND2_X1 U5945 ( .A1(n5142), .A2(n4799), .ZN(n4800) );
  AND2_X1 U5946 ( .A1(n5138), .A2(n4801), .ZN(n5809) );
  OAI21_X1 U5947 ( .B1(REIP_REG_5__SCAN_IN), .B2(n4802), .A(n5809), .ZN(n4807)
         );
  INV_X1 U5948 ( .A(n5818), .ZN(n5761) );
  AOI22_X1 U5949 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5820), .B1(n5790), 
        .B2(n3201), .ZN(n4803) );
  OAI211_X1 U5950 ( .C1(n5761), .C2(n4804), .A(n4803), .B(n5791), .ZN(n4805)
         );
  AOI21_X1 U5951 ( .B1(n5821), .B2(n4919), .A(n4805), .ZN(n4806) );
  OAI211_X1 U5952 ( .C1(n4916), .C2(n5817), .A(n4807), .B(n4806), .ZN(U2822)
         );
  XOR2_X1 U5953 ( .A(n4710), .B(n5260), .Z(n5893) );
  INV_X1 U5954 ( .A(n5343), .ZN(n5837) );
  OR2_X1 U5955 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  NAND2_X1 U5956 ( .A1(n5265), .A2(n4810), .ZN(n5806) );
  OAI22_X1 U5957 ( .A1(n5336), .A2(n5806), .B1(n4811), .B2(n5840), .ZN(n4812)
         );
  AOI21_X1 U5958 ( .B1(n5893), .B2(n5837), .A(n4812), .ZN(n4813) );
  INV_X1 U5959 ( .A(n4813), .ZN(U2853) );
  OAI21_X1 U5960 ( .B1(n4816), .B2(n4815), .A(n4814), .ZN(n4817) );
  INV_X1 U5961 ( .A(n4817), .ZN(n5894) );
  OAI22_X1 U5962 ( .A1(n6009), .A2(n5806), .B1(n5721), .B2(n6580), .ZN(n4822)
         );
  OAI21_X1 U5964 ( .B1(n5927), .B2(n5993), .A(n5011), .ZN(n5996) );
  AOI21_X1 U5965 ( .B1(n4818), .B2(n5928), .A(n5996), .ZN(n5973) );
  AOI21_X1 U5966 ( .B1(n5993), .B2(n5998), .A(n5992), .ZN(n5977) );
  OAI33_X1 U5967 ( .A1(1'b0), .A2(n5973), .A3(n4819), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4818), .B3(n5977), .ZN(n4821) );
  AOI211_X1 U5968 ( .C1(n5894), .C2(n6012), .A(n4822), .B(n4821), .ZN(n4823)
         );
  INV_X1 U5969 ( .A(n4823), .ZN(U3012) );
  AOI21_X1 U5970 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(n4978) );
  INV_X1 U5971 ( .A(n4978), .ZN(n4863) );
  XNOR2_X1 U5972 ( .A(n5263), .B(n4933), .ZN(n5948) );
  AOI22_X1 U5973 ( .A1(n5948), .A2(n5836), .B1(n5341), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4827) );
  OAI21_X1 U5974 ( .B1(n4863), .B2(n5343), .A(n4827), .ZN(U2851) );
  OR2_X1 U5975 ( .A1(n5140), .A2(REIP_REG_1__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5976 ( .A1(n4921), .A2(n4922), .ZN(n5814) );
  INV_X1 U5977 ( .A(n6030), .ZN(n4830) );
  INV_X1 U5978 ( .A(n4828), .ZN(n4829) );
  AND2_X1 U5979 ( .A1(n5142), .A2(n4829), .ZN(n5819) );
  AOI22_X1 U5980 ( .A1(n4830), .A2(n5819), .B1(n5790), .B2(n5991), .ZN(n4836)
         );
  INV_X1 U5981 ( .A(n5914), .ZN(n4831) );
  AOI22_X1 U5982 ( .A1(n5820), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5821), 
        .B2(n4831), .ZN(n4835) );
  INV_X1 U5983 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4832) );
  NAND3_X1 U5984 ( .A1(n4841), .A2(REIP_REG_1__SCAN_IN), .A3(n4832), .ZN(n4834) );
  NAND2_X1 U5985 ( .A1(n5818), .A2(EBX_REG_2__SCAN_IN), .ZN(n4833) );
  NAND4_X1 U5986 ( .A1(n4836), .A2(n4835), .A3(n4834), .A4(n4833), .ZN(n4837)
         );
  AOI21_X1 U5987 ( .B1(REIP_REG_2__SCAN_IN), .B2(n5814), .A(n4837), .ZN(n4838)
         );
  OAI21_X1 U5988 ( .B1(n4839), .B2(n5817), .A(n4838), .ZN(U2825) );
  AOI22_X1 U5989 ( .A1(n4840), .A2(n5819), .B1(n5790), .B2(n5976), .ZN(n4851)
         );
  NOR2_X1 U5990 ( .A1(REIP_REG_4__SCAN_IN), .A2(n4845), .ZN(n4842) );
  AOI22_X1 U5991 ( .A1(n4842), .A2(n4841), .B1(n5818), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4850) );
  NAND2_X1 U5992 ( .A1(n5821), .A2(n4966), .ZN(n4844) );
  NAND2_X1 U5993 ( .A1(n5820), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4843)
         );
  AND3_X1 U5994 ( .A1(n4844), .A2(n4843), .A3(n5791), .ZN(n4849) );
  INV_X1 U5995 ( .A(n4845), .ZN(n4846) );
  NAND2_X1 U5996 ( .A1(n4922), .A2(n4846), .ZN(n4847) );
  NAND2_X1 U5997 ( .A1(n5138), .A2(n4847), .ZN(n5830) );
  OR2_X1 U5998 ( .A1(n5830), .A2(n6579), .ZN(n4848) );
  AND4_X1 U5999 ( .A1(n4851), .A2(n4850), .A3(n4849), .A4(n4848), .ZN(n4852)
         );
  OAI21_X1 U6000 ( .B1(n4853), .B2(n5817), .A(n4852), .ZN(U2823) );
  INV_X1 U6001 ( .A(n5893), .ZN(n4854) );
  INV_X1 U6002 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5871) );
  OAI222_X1 U6003 ( .A1(n5653), .A2(n4854), .B1(n5371), .B2(n6955), .C1(n5369), 
        .C2(n5871), .ZN(U2885) );
  INV_X1 U6004 ( .A(n5138), .ZN(n5236) );
  NOR2_X1 U6005 ( .A1(n5236), .A2(n4855), .ZN(n5796) );
  OAI21_X1 U6006 ( .B1(REIP_REG_8__SCAN_IN), .B2(n4856), .A(n5796), .ZN(n4862)
         );
  INV_X1 U6007 ( .A(n4976), .ZN(n4860) );
  AOI22_X1 U6008 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5820), .B1(n5790), 
        .B2(n5948), .ZN(n4857) );
  OAI211_X1 U6009 ( .C1(n5761), .C2(n4858), .A(n4857), .B(n5791), .ZN(n4859)
         );
  AOI21_X1 U6010 ( .B1(n5821), .B2(n4860), .A(n4859), .ZN(n4861) );
  OAI211_X1 U6011 ( .C1(n4863), .C2(n5646), .A(n4862), .B(n4861), .ZN(U2819)
         );
  INV_X1 U6012 ( .A(DATAI_8_), .ZN(n6714) );
  INV_X1 U6013 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5868) );
  OAI222_X1 U6014 ( .A1(n4863), .A2(n5653), .B1(n5371), .B2(n6714), .C1(n5369), 
        .C2(n5868), .ZN(U2883) );
  OAI22_X1 U6015 ( .A1(n4865), .A2(n5761), .B1(n5825), .B2(n4864), .ZN(n4866)
         );
  AOI21_X1 U6016 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5138), .A(n4866), .ZN(n4869)
         );
  NAND2_X1 U6017 ( .A1(n5794), .A2(n5813), .ZN(n4867) );
  AOI22_X1 U6018 ( .A1(n4867), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n5819), 
        .B2(n6614), .ZN(n4868) );
  OAI211_X1 U6019 ( .C1(n5817), .C2(n5917), .A(n4869), .B(n4868), .ZN(U2827)
         );
  NOR2_X1 U6020 ( .A1(n4870), .A2(n6611), .ZN(n6119) );
  NAND2_X1 U6021 ( .A1(n6207), .A2(n4871), .ZN(n6099) );
  OR2_X1 U6022 ( .A1(n6099), .A2(n6125), .ZN(n4874) );
  NOR2_X1 U6023 ( .A1(n4872), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4898)
         );
  INV_X1 U6024 ( .A(n4898), .ZN(n4873) );
  INV_X1 U6025 ( .A(n4881), .ZN(n4879) );
  INV_X1 U6026 ( .A(n5578), .ZN(n4875) );
  NAND3_X1 U6027 ( .A1(n4876), .A2(n4875), .A3(n6027), .ZN(n4877) );
  NAND2_X1 U6028 ( .A1(n4877), .A2(n6612), .ZN(n4880) );
  NAND3_X1 U6029 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6525), .A3(n6517), .ZN(n6096) );
  AOI21_X1 U6030 ( .B1(n6438), .B2(n6096), .A(n6129), .ZN(n4878) );
  OAI22_X1 U6031 ( .A1(n4881), .A2(n4880), .B1(n6436), .B2(n6096), .ZN(n4896)
         );
  AOI22_X1 U6032 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4897), .B1(n6439), 
        .B2(n4896), .ZN(n4883) );
  AOI22_X1 U6033 ( .A1(n4899), .A2(n6448), .B1(n6440), .B2(n4898), .ZN(n4882)
         );
  OAI211_X1 U6034 ( .C1(n4902), .C2(n6451), .A(n4883), .B(n4882), .ZN(U3044)
         );
  AOI22_X1 U6035 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4897), .B1(n6489), 
        .B2(n4896), .ZN(n4885) );
  AOI22_X1 U6036 ( .A1(n4899), .A2(n6493), .B1(n4898), .B2(n6491), .ZN(n4884)
         );
  OAI211_X1 U6037 ( .C1(n4902), .C2(n6498), .A(n4885), .B(n4884), .ZN(U3051)
         );
  AOI22_X1 U6038 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4897), .B1(n6470), 
        .B2(n4896), .ZN(n4887) );
  AOI22_X1 U6039 ( .A1(n4899), .A2(n6472), .B1(n4898), .B2(n6471), .ZN(n4886)
         );
  OAI211_X1 U6040 ( .C1(n4902), .C2(n6475), .A(n4887), .B(n4886), .ZN(U3048)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n4897), .B1(n6482), 
        .B2(n4896), .ZN(n4889) );
  AOI22_X1 U6042 ( .A1(n4899), .A2(n6484), .B1(n4898), .B2(n6483), .ZN(n4888)
         );
  OAI211_X1 U6043 ( .C1(n4902), .C2(n6487), .A(n4889), .B(n4888), .ZN(U3050)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4897), .B1(n6476), 
        .B2(n4896), .ZN(n4891) );
  AOI22_X1 U6045 ( .A1(n4899), .A2(n6478), .B1(n4898), .B2(n6477), .ZN(n4890)
         );
  OAI211_X1 U6046 ( .C1(n4902), .C2(n6481), .A(n4891), .B(n4890), .ZN(U3049)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4897), .B1(n6452), 
        .B2(n4896), .ZN(n4893) );
  AOI22_X1 U6048 ( .A1(n4899), .A2(n6454), .B1(n4898), .B2(n6453), .ZN(n4892)
         );
  OAI211_X1 U6049 ( .C1(n4902), .C2(n6457), .A(n4893), .B(n4892), .ZN(U3045)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n4897), .B1(n6464), 
        .B2(n4896), .ZN(n4895) );
  AOI22_X1 U6051 ( .A1(n4899), .A2(n6466), .B1(n4898), .B2(n6465), .ZN(n4894)
         );
  OAI211_X1 U6052 ( .C1(n4902), .C2(n6469), .A(n4895), .B(n4894), .ZN(U3047)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n4897), .B1(n6458), 
        .B2(n4896), .ZN(n4901) );
  AOI22_X1 U6054 ( .A1(n4899), .A2(n6460), .B1(n4898), .B2(n6459), .ZN(n4900)
         );
  OAI211_X1 U6055 ( .C1(n4902), .C2(n6463), .A(n4901), .B(n4900), .ZN(U3046)
         );
  XOR2_X1 U6056 ( .A(n4904), .B(n4903), .Z(n6013) );
  INV_X1 U6057 ( .A(n6013), .ZN(n4910) );
  INV_X1 U6058 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6576) );
  OR2_X1 U6059 ( .A1(n5721), .A2(n6576), .ZN(n6007) );
  INV_X1 U6060 ( .A(n6007), .ZN(n4905) );
  AOI21_X1 U6061 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4905), 
        .ZN(n4906) );
  OAI21_X1 U6062 ( .B1(n5915), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4906), 
        .ZN(n4907) );
  AOI21_X1 U6063 ( .B1(n4908), .B2(n5910), .A(n4907), .ZN(n4909) );
  OAI21_X1 U6064 ( .B1(n4910), .B2(n5918), .A(n4909), .ZN(U2985) );
  OAI21_X1 U6065 ( .B1(n4913), .B2(n4912), .A(n4911), .ZN(n5968) );
  INV_X1 U6066 ( .A(n5921), .ZN(n5416) );
  INV_X1 U6067 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U6068 ( .A1(n5416), .A2(n4915), .B1(n5721), .B2(n4914), .ZN(n4918)
         );
  NOR2_X1 U6069 ( .A1(n4916), .A2(n4644), .ZN(n4917) );
  AOI211_X1 U6070 ( .C1(n5888), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4920)
         );
  OAI21_X1 U6071 ( .B1(n5918), .B2(n5968), .A(n4920), .ZN(U2981) );
  INV_X1 U6072 ( .A(n4921), .ZN(n4927) );
  AOI22_X1 U6073 ( .A1(n5586), .A2(n5819), .B1(n5790), .B2(n6006), .ZN(n4925)
         );
  INV_X1 U6074 ( .A(n4922), .ZN(n4923) );
  AOI22_X1 U6075 ( .A1(n5820), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n4923), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4924) );
  OAI211_X1 U6076 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5813), .A(n4925), 
        .B(n4924), .ZN(n4926) );
  AOI211_X1 U6077 ( .C1(n5818), .C2(EBX_REG_1__SCAN_IN), .A(n4927), .B(n4926), 
        .ZN(n4928) );
  OAI21_X1 U6078 ( .B1(n4929), .B2(n5817), .A(n4928), .ZN(U2826) );
  NOR2_X1 U6079 ( .A1(n4824), .A2(n4931), .ZN(n4932) );
  OR2_X1 U6080 ( .A1(n4930), .A2(n4932), .ZN(n5797) );
  INV_X1 U6081 ( .A(DATAI_9_), .ZN(n6895) );
  INV_X1 U6082 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5866) );
  OAI222_X1 U6083 ( .A1(n5797), .A2(n5653), .B1(n5371), .B2(n6895), .C1(n5369), 
        .C2(n5866), .ZN(U2882) );
  INV_X1 U6084 ( .A(n4933), .ZN(n4935) );
  OAI21_X1 U6085 ( .B1(n5263), .B2(n4935), .A(n4934), .ZN(n4936) );
  INV_X1 U6086 ( .A(n4936), .ZN(n4937) );
  OR2_X1 U6087 ( .A1(n4937), .A2(n4943), .ZN(n5789) );
  INV_X1 U6088 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4938) );
  OAI222_X1 U6089 ( .A1(n5789), .A2(n5336), .B1(n4938), .B2(n5840), .C1(n5343), 
        .C2(n5797), .ZN(U2850) );
  OR2_X1 U6090 ( .A1(n4930), .A2(n4940), .ZN(n4941) );
  AND2_X1 U6091 ( .A1(n4939), .A2(n4941), .ZN(n4988) );
  OR2_X1 U6092 ( .A1(n4943), .A2(n4942), .ZN(n4944) );
  AND2_X1 U6093 ( .A1(n5009), .A2(n4944), .ZN(n5929) );
  AOI22_X1 U6094 ( .A1(n5929), .A2(n5790), .B1(n5818), .B2(EBX_REG_10__SCAN_IN), .ZN(n4946) );
  INV_X1 U6095 ( .A(n5791), .ZN(n5803) );
  AOI21_X1 U6096 ( .B1(n5820), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5803), 
        .ZN(n4945) );
  OAI211_X1 U6097 ( .C1(n4986), .C2(n5813), .A(n4946), .B(n4945), .ZN(n4947)
         );
  AOI21_X1 U6098 ( .B1(n5796), .B2(REIP_REG_10__SCAN_IN), .A(n4947), .ZN(n4950) );
  INV_X1 U6099 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6584) );
  INV_X1 U6100 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6583) );
  AOI21_X1 U6101 ( .B1(n6584), .B2(n6583), .A(n5802), .ZN(n4948) );
  NAND2_X1 U6102 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5781) );
  NAND2_X1 U6103 ( .A1(n4948), .A2(n5781), .ZN(n4949) );
  OAI211_X1 U6104 ( .C1(n4951), .C2(n5646), .A(n4950), .B(n4949), .ZN(U2817)
         );
  INV_X1 U6105 ( .A(DATAI_10_), .ZN(n6775) );
  INV_X1 U6106 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5864) );
  OAI222_X1 U6107 ( .A1(n4951), .A2(n5653), .B1(n5371), .B2(n6775), .C1(n5369), 
        .C2(n5864), .ZN(U2881) );
  INV_X1 U6108 ( .A(n5929), .ZN(n4953) );
  INV_X1 U6109 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4952) );
  OAI222_X1 U6110 ( .A1(n4953), .A2(n5336), .B1(n5840), .B2(n4952), .C1(n5343), 
        .C2(n4951), .ZN(U2849) );
  NAND2_X1 U6111 ( .A1(n4955), .A2(n4954), .ZN(n4956) );
  XNOR2_X1 U6112 ( .A(n4957), .B(n4956), .ZN(n5940) );
  NAND2_X1 U6113 ( .A1(n5940), .A2(n5909), .ZN(n4960) );
  INV_X2 U6114 ( .A(n5721), .ZN(n5990) );
  NAND2_X1 U6115 ( .A1(n5990), .A2(REIP_REG_9__SCAN_IN), .ZN(n5936) );
  OAI21_X1 U6116 ( .B1(n5416), .B2(n5793), .A(n5936), .ZN(n4958) );
  AOI21_X1 U6117 ( .B1(n5888), .B2(n5798), .A(n4958), .ZN(n4959) );
  OAI211_X1 U6118 ( .C1(n4644), .C2(n5797), .A(n4960), .B(n4959), .ZN(U2977)
         );
  OAI21_X1 U6119 ( .B1(n4962), .B2(n4965), .A(n4964), .ZN(n5974) );
  INV_X1 U6120 ( .A(n4966), .ZN(n4968) );
  AOI22_X1 U6121 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4967) );
  OAI21_X1 U6122 ( .B1(n5915), .B2(n4968), .A(n4967), .ZN(n4969) );
  AOI21_X1 U6123 ( .B1(n4970), .B2(n5910), .A(n4969), .ZN(n4971) );
  OAI21_X1 U6124 ( .B1(n5918), .B2(n5974), .A(n4971), .ZN(U2982) );
  OAI21_X1 U6125 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(n5949) );
  NAND2_X1 U6126 ( .A1(n5990), .A2(REIP_REG_8__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U6127 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4975)
         );
  OAI211_X1 U6128 ( .C1(n5915), .C2(n4976), .A(n5946), .B(n4975), .ZN(n4977)
         );
  AOI21_X1 U6129 ( .B1(n4978), .B2(n5910), .A(n4977), .ZN(n4979) );
  OAI21_X1 U6130 ( .B1(n5949), .B2(n5918), .A(n4979), .ZN(U2978) );
  INV_X1 U6131 ( .A(n4980), .ZN(n4981) );
  AOI21_X1 U6132 ( .B1(n4982), .B2(n4939), .A(n4981), .ZN(n5889) );
  INV_X1 U6133 ( .A(n5889), .ZN(n4983) );
  INV_X1 U6134 ( .A(DATAI_11_), .ZN(n6888) );
  INV_X1 U6135 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5862) );
  OAI222_X1 U6136 ( .A1(n4983), .A2(n5653), .B1(n5371), .B2(n6888), .C1(n5369), 
        .C2(n5862), .ZN(U2880) );
  XNOR2_X1 U6137 ( .A(n5065), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4984)
         );
  XNOR2_X1 U6138 ( .A(n3637), .B(n4984), .ZN(n5930) );
  INV_X1 U6139 ( .A(n5930), .ZN(n4990) );
  AOI22_X1 U6140 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n4985) );
  OAI21_X1 U6141 ( .B1(n5915), .B2(n4986), .A(n4985), .ZN(n4987) );
  AOI21_X1 U6142 ( .B1(n4988), .B2(n5910), .A(n4987), .ZN(n4989) );
  OAI21_X1 U6143 ( .B1(n4990), .B2(n5918), .A(n4989), .ZN(U2976) );
  XOR2_X1 U6144 ( .A(n4991), .B(n4980), .Z(n5026) );
  INV_X1 U6145 ( .A(n5026), .ZN(n5002) );
  INV_X1 U6146 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U6147 ( .A1(n5007), .A2(n4992), .ZN(n4993) );
  NAND2_X1 U6148 ( .A1(n5725), .A2(n4993), .ZN(n5036) );
  NAND2_X1 U6149 ( .A1(n4994), .A2(n5138), .ZN(n5774) );
  INV_X1 U6150 ( .A(n5774), .ZN(n5782) );
  NAND2_X1 U6151 ( .A1(n5782), .A2(REIP_REG_12__SCAN_IN), .ZN(n4999) );
  INV_X1 U6152 ( .A(n4995), .ZN(n5024) );
  NAND2_X1 U6153 ( .A1(n5820), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4996)
         );
  OAI211_X1 U6154 ( .C1(n5813), .C2(n5024), .A(n5791), .B(n4996), .ZN(n4997)
         );
  AOI21_X1 U6155 ( .B1(EBX_REG_12__SCAN_IN), .B2(n5818), .A(n4997), .ZN(n4998)
         );
  OAI211_X1 U6156 ( .C1(n5036), .C2(n5825), .A(n4999), .B(n4998), .ZN(n5000)
         );
  AOI21_X1 U6157 ( .B1(n5777), .B2(n6587), .A(n5000), .ZN(n5001) );
  OAI21_X1 U6158 ( .B1(n5002), .B2(n5646), .A(n5001), .ZN(U2815) );
  INV_X1 U6159 ( .A(DATAI_12_), .ZN(n6788) );
  OAI222_X1 U6160 ( .A1(n5653), .A2(n5002), .B1(n5371), .B2(n6788), .C1(n5369), 
        .C2(n3838), .ZN(U2879) );
  INV_X1 U6161 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5003) );
  OAI222_X1 U6162 ( .A1(n5036), .A2(n5336), .B1(n5840), .B2(n5003), .C1(n5343), 
        .C2(n5002), .ZN(U2847) );
  AOI22_X1 U6163 ( .A1(n5004), .A2(n5065), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n3637), .ZN(n5006) );
  XNOR2_X1 U6164 ( .A(n5065), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5005)
         );
  XNOR2_X1 U6165 ( .A(n5006), .B(n5005), .ZN(n5892) );
  INV_X1 U6166 ( .A(n5007), .ZN(n5008) );
  AOI21_X1 U6167 ( .B1(n5010), .B2(n5009), .A(n5008), .ZN(n5835) );
  INV_X1 U6168 ( .A(n5530), .ZN(n5013) );
  INV_X1 U6169 ( .A(n5927), .ZN(n5012) );
  INV_X1 U6170 ( .A(n5011), .ZN(n5924) );
  AOI21_X1 U6171 ( .B1(n5012), .B2(n5014), .A(n5924), .ZN(n5532) );
  OAI21_X1 U6172 ( .B1(n5013), .B2(n5708), .A(n5532), .ZN(n5710) );
  NOR3_X1 U6173 ( .A1(n4308), .A2(n5709), .A3(n5014), .ZN(n5030) );
  AOI21_X1 U6174 ( .B1(n5013), .B2(n5992), .A(n5030), .ZN(n5714) );
  INV_X1 U6175 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U6176 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5710), .B1(n5722), .B2(n5028), .ZN(n5015) );
  OAI21_X1 U6177 ( .B1(n5721), .B2(n6585), .A(n5015), .ZN(n5016) );
  AOI21_X1 U6178 ( .B1(n5835), .B2(n6023), .A(n5016), .ZN(n5017) );
  OAI21_X1 U6179 ( .B1(n5892), .B2(n6018), .A(n5017), .ZN(U3007) );
  INV_X1 U6180 ( .A(n5018), .ZN(n5019) );
  NOR2_X1 U6181 ( .A1(n5020), .A2(n5019), .ZN(n5021) );
  XNOR2_X1 U6182 ( .A(n5022), .B(n5021), .ZN(n5040) );
  NAND2_X1 U6183 ( .A1(n5990), .A2(REIP_REG_12__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6184 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5023)
         );
  OAI211_X1 U6185 ( .C1(n5915), .C2(n5024), .A(n5034), .B(n5023), .ZN(n5025)
         );
  AOI21_X1 U6186 ( .B1(n5026), .B2(n5910), .A(n5025), .ZN(n5027) );
  OAI21_X1 U6187 ( .B1(n5040), .B2(n5918), .A(n5027), .ZN(U2974) );
  NOR2_X1 U6188 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5028), .ZN(n5038)
         );
  INV_X1 U6189 ( .A(n6025), .ZN(n5029) );
  NOR3_X1 U6190 ( .A1(n5030), .A2(n5029), .A3(n5992), .ZN(n5032) );
  INV_X1 U6191 ( .A(n5710), .ZN(n5031) );
  OAI21_X1 U6192 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5032), .A(n5031), 
        .ZN(n5033) );
  NAND2_X1 U6193 ( .A1(n5033), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5035) );
  OAI211_X1 U6194 ( .C1(n6009), .C2(n5036), .A(n5035), .B(n5034), .ZN(n5037)
         );
  AOI21_X1 U6195 ( .B1(n5038), .B2(n5722), .A(n5037), .ZN(n5039) );
  OAI21_X1 U6196 ( .B1(n5040), .B2(n6018), .A(n5039), .ZN(U3006) );
  INV_X1 U6197 ( .A(n5042), .ZN(n5043) );
  NAND2_X1 U6198 ( .A1(n3859), .A2(n5043), .ZN(n5045) );
  INV_X1 U6199 ( .A(n5832), .ZN(n5046) );
  INV_X1 U6200 ( .A(DATAI_13_), .ZN(n6739) );
  INV_X1 U6201 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5859) );
  OAI222_X1 U6202 ( .A1(n5046), .A2(n5653), .B1(n5371), .B2(n6739), .C1(n5369), 
        .C2(n5859), .ZN(U2878) );
  OAI21_X1 U6203 ( .B1(n5049), .B2(n5048), .A(n5047), .ZN(n5450) );
  INV_X1 U6204 ( .A(DATAI_14_), .ZN(n6952) );
  INV_X1 U6205 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5857) );
  OAI222_X1 U6206 ( .A1(n5450), .A2(n5653), .B1(n5371), .B2(n6952), .C1(n5369), 
        .C2(n5857), .ZN(U2877) );
  OAI21_X1 U6207 ( .B1(n5727), .B2(n5050), .A(n5252), .ZN(n5760) );
  INV_X1 U6208 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5762) );
  OAI222_X1 U6209 ( .A1(n5760), .A2(n5336), .B1(n5762), .B2(n5840), .C1(n5450), 
        .C2(n5343), .ZN(U2845) );
  XNOR2_X1 U6210 ( .A(n5448), .B(n5569), .ZN(n5053) );
  XNOR2_X1 U6211 ( .A(n5052), .B(n5053), .ZN(n5570) );
  INV_X1 U6212 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5244) );
  INV_X1 U6213 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5054) );
  OAI22_X1 U6214 ( .A1(n5416), .A2(n5244), .B1(n5721), .B2(n5054), .ZN(n5055)
         );
  AOI21_X1 U6215 ( .B1(n5888), .B2(n5241), .A(n5055), .ZN(n5058) );
  AOI21_X1 U6216 ( .B1(n5056), .B2(n5248), .A(n5223), .ZN(n5849) );
  NAND2_X1 U6217 ( .A1(n5849), .A2(n5910), .ZN(n5057) );
  OAI211_X1 U6218 ( .C1(n5570), .C2(n5918), .A(n5058), .B(n5057), .ZN(U2970)
         );
  NAND3_X1 U6219 ( .A1(n3636), .A2(n5512), .A3(n5540), .ZN(n5066) );
  XNOR2_X1 U6220 ( .A(n5448), .B(n5061), .ZN(n5430) );
  XNOR2_X1 U6221 ( .A(n5448), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5415)
         );
  OAI21_X1 U6222 ( .B1(n5060), .B2(n5066), .A(n5092), .ZN(n5067) );
  XNOR2_X1 U6223 ( .A(n5067), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5083)
         );
  INV_X1 U6224 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U6225 ( .A1(n5721), .A2(n6992), .ZN(n5077) );
  NOR2_X1 U6226 ( .A1(n5068), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5069)
         );
  AOI211_X1 U6227 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5070), .A(n5077), .B(n5069), .ZN(n5074) );
  INV_X1 U6228 ( .A(n5299), .ZN(n5071) );
  AOI21_X1 U6229 ( .B1(n5072), .B2(n5215), .A(n5071), .ZN(n5305) );
  NAND2_X1 U6230 ( .A1(n5305), .A2(n6023), .ZN(n5073) );
  OAI211_X1 U6231 ( .C1(n5083), .C2(n6018), .A(n5074), .B(n5073), .ZN(U2995)
         );
  NOR2_X1 U6232 ( .A1(n5416), .A2(n5075), .ZN(n5076) );
  AOI211_X1 U6233 ( .C1(n5888), .C2(n5205), .A(n5077), .B(n5076), .ZN(n5082)
         );
  OR2_X1 U6234 ( .A1(n5283), .A2(n5213), .ZN(n5211) );
  NAND2_X1 U6235 ( .A1(n5211), .A2(n5079), .ZN(n5080) );
  NAND2_X1 U6236 ( .A1(n5201), .A2(n5910), .ZN(n5081) );
  OAI211_X1 U6237 ( .C1(n5083), .C2(n5918), .A(n5082), .B(n5081), .ZN(U2963)
         );
  AOI21_X1 U6238 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5086), 
        .ZN(n5087) );
  OAI21_X1 U6239 ( .B1(n5915), .B2(n5157), .A(n5087), .ZN(n5088) );
  AOI21_X1 U6240 ( .B1(n5155), .B2(n5910), .A(n5088), .ZN(n5089) );
  OAI21_X1 U6241 ( .B1(n5090), .B2(n5918), .A(n5089), .ZN(U2956) );
  NAND3_X1 U6242 ( .A1(n3636), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5091) );
  XNOR2_X1 U6243 ( .A(n5093), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5108)
         );
  XNOR2_X1 U6244 ( .A(n5299), .B(n5296), .ZN(n5618) );
  AND2_X1 U6245 ( .A1(n5990), .A2(REIP_REG_24__SCAN_IN), .ZN(n5103) );
  NAND3_X1 U6246 ( .A1(n5510), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5512), .ZN(n5095) );
  INV_X1 U6247 ( .A(n5686), .ZN(n5094) );
  AOI21_X1 U6248 ( .B1(n5096), .B2(n5095), .A(n5094), .ZN(n5097) );
  AOI211_X1 U6249 ( .C1(n5618), .C2(n6023), .A(n5103), .B(n5097), .ZN(n5098)
         );
  OAI21_X1 U6250 ( .B1(n5108), .B2(n6018), .A(n5098), .ZN(U2994) );
  AND2_X1 U6251 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  INV_X1 U6252 ( .A(n5616), .ZN(n5105) );
  AOI21_X1 U6253 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5103), 
        .ZN(n5104) );
  OAI21_X1 U6254 ( .B1(n5915), .B2(n5105), .A(n5104), .ZN(n5106) );
  AOI21_X1 U6255 ( .B1(n5662), .B2(n5910), .A(n5106), .ZN(n5107) );
  OAI21_X1 U6256 ( .B1(n5108), .B2(n5918), .A(n5107), .ZN(U2962) );
  INV_X1 U6257 ( .A(n4555), .ZN(n5110) );
  INV_X1 U6258 ( .A(n5737), .ZN(n5115) );
  AOI21_X1 U6259 ( .B1(n5110), .B2(n5590), .A(n5115), .ZN(n5118) );
  INV_X1 U6260 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U6261 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5109), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6015), .ZN(n5592) );
  NOR3_X1 U6262 ( .A1(n5587), .A2(n4308), .A3(n5592), .ZN(n5112) );
  NOR3_X1 U6263 ( .A1(n5110), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6543), 
        .ZN(n5111) );
  AOI211_X1 U6264 ( .C1(n5114), .C2(n5113), .A(n5112), .B(n5111), .ZN(n5116)
         );
  OAI22_X1 U6265 ( .A1(n5118), .A2(n5117), .B1(n5116), .B2(n5115), .ZN(U3459)
         );
  INV_X1 U6266 ( .A(n5345), .ZN(n5154) );
  MUX2_X1 U6267 ( .A(EBX_REG_29__SCAN_IN), .B(n5120), .S(n5119), .Z(n5123) );
  NOR2_X1 U6268 ( .A1(n5121), .A2(EBX_REG_29__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6269 ( .A1(n5123), .A2(n5122), .ZN(n5166) );
  NOR2_X1 U6270 ( .A1(n5179), .A2(n5166), .ZN(n5168) );
  OAI22_X1 U6271 ( .A1(n5127), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5126), .ZN(n5128) );
  XNOR2_X1 U6272 ( .A(n5129), .B(n5128), .ZN(n5468) );
  INV_X1 U6273 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6973) );
  INV_X1 U6274 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6863) );
  NOR2_X1 U6275 ( .A1(n6973), .A2(n6863), .ZN(n5150) );
  INV_X1 U6276 ( .A(n5130), .ZN(n5132) );
  AND3_X1 U6277 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_20__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6278 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U6279 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5214) );
  INV_X1 U6280 ( .A(n5214), .ZN(n5134) );
  NAND2_X1 U6281 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5134), .ZN(n5135) );
  AND2_X1 U6282 ( .A1(n5138), .A2(n5135), .ZN(n5136) );
  NAND3_X1 U6283 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5137) );
  AND2_X1 U6284 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  NOR2_X1 U6285 ( .A1(n5617), .A2(n5139), .ZN(n5601) );
  OAI21_X1 U6286 ( .B1(n5150), .B2(n5140), .A(n5601), .ZN(n5186) );
  NOR2_X1 U6287 ( .A1(n5186), .A2(n6597), .ZN(n5156) );
  AOI211_X1 U6288 ( .C1(n5156), .C2(REIP_REG_30__SCAN_IN), .A(n6786), .B(n5236), .ZN(n5146) );
  NAND3_X1 U6289 ( .A1(n5142), .A2(EBX_REG_31__SCAN_IN), .A3(n5141), .ZN(n5143) );
  OAI21_X1 U6290 ( .B1(n5794), .B2(n5144), .A(n5143), .ZN(n5145) );
  AOI21_X1 U6291 ( .B1(n5468), .B2(n5790), .A(n3206), .ZN(n5153) );
  NAND2_X1 U6292 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5147), .ZN(n5645) );
  NAND2_X1 U6293 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .ZN(
        n5148) );
  NOR2_X2 U6294 ( .A1(n5645), .A2(n5148), .ZN(n5629) );
  NAND3_X1 U6295 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5629), .ZN(n5202) );
  NOR2_X2 U6296 ( .A1(n5202), .A2(n6992), .ZN(n5610) );
  AND2_X1 U6297 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5149) );
  NAND2_X1 U6298 ( .A1(n5608), .A2(n5149), .ZN(n5200) );
  INV_X1 U6299 ( .A(n5150), .ZN(n5151) );
  NOR2_X2 U6300 ( .A1(n5200), .A2(n5151), .ZN(n5175) );
  NAND4_X1 U6301 ( .A1(n5175), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n6786), .ZN(n5152) );
  OAI211_X1 U6302 ( .C1(n5154), .C2(n5646), .A(n5153), .B(n5152), .ZN(U2796)
         );
  INV_X1 U6303 ( .A(n5155), .ZN(n5354) );
  NOR3_X1 U6304 ( .A1(n5156), .A2(n5236), .A3(n6599), .ZN(n5161) );
  INV_X1 U6305 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5278) );
  INV_X1 U6306 ( .A(n5157), .ZN(n5158) );
  AOI22_X1 U6307 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5820), .B1(n5821), 
        .B2(n5158), .ZN(n5159) );
  OAI21_X1 U6308 ( .B1(n5761), .B2(n5278), .A(n5159), .ZN(n5160) );
  AOI211_X1 U6309 ( .C1(n5162), .C2(n5790), .A(n5161), .B(n5160), .ZN(n5164)
         );
  NAND3_X1 U6310 ( .A1(n5175), .A2(REIP_REG_29__SCAN_IN), .A3(n6599), .ZN(
        n5163) );
  OAI211_X1 U6311 ( .C1(n5354), .C2(n5646), .A(n5164), .B(n5163), .ZN(U2797)
         );
  AND2_X1 U6312 ( .A1(n5179), .A2(n5166), .ZN(n5167) );
  NAND2_X1 U6313 ( .A1(n5186), .A2(REIP_REG_29__SCAN_IN), .ZN(n5173) );
  OAI22_X1 U6314 ( .A1(n5170), .A2(n5794), .B1(n5813), .B2(n5169), .ZN(n5171)
         );
  AOI21_X1 U6315 ( .B1(n5818), .B2(EBX_REG_29__SCAN_IN), .A(n5171), .ZN(n5172)
         );
  OAI211_X1 U6316 ( .C1(n5825), .C2(n5472), .A(n5173), .B(n5172), .ZN(n5174)
         );
  AOI21_X1 U6317 ( .B1(n5175), .B2(n6597), .A(n5174), .ZN(n5176) );
  OAI21_X1 U6318 ( .B1(n5165), .B2(n5646), .A(n5176), .ZN(U2798) );
  AOI21_X1 U6319 ( .B1(n5178), .B2(n5177), .A(n4189), .ZN(n5381) );
  INV_X1 U6320 ( .A(n5381), .ZN(n5359) );
  OAI21_X1 U6321 ( .B1(n5193), .B2(n5180), .A(n5179), .ZN(n5486) );
  OAI22_X1 U6322 ( .A1(n5181), .A2(n5794), .B1(n5813), .B2(n5379), .ZN(n5182)
         );
  AOI21_X1 U6323 ( .B1(n5818), .B2(EBX_REG_28__SCAN_IN), .A(n5182), .ZN(n5183)
         );
  OAI21_X1 U6324 ( .B1(n5486), .B2(n5825), .A(n5183), .ZN(n5185) );
  NOR3_X1 U6325 ( .A1(n5200), .A2(REIP_REG_28__SCAN_IN), .A3(n6863), .ZN(n5184) );
  AOI211_X1 U6326 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5186), .A(n5185), .B(n5184), .ZN(n5187) );
  OAI21_X1 U6327 ( .B1(n5359), .B2(n5646), .A(n5187), .ZN(U2799) );
  AND2_X1 U6328 ( .A1(n5189), .A2(n5188), .ZN(n5286) );
  OAI21_X1 U6329 ( .B1(n5286), .B2(n5190), .A(n5177), .ZN(n5362) );
  INV_X1 U6330 ( .A(n5362), .ZN(n5389) );
  NAND2_X1 U6331 ( .A1(n5389), .A2(n5810), .ZN(n5199) );
  INV_X1 U6332 ( .A(n5601), .ZN(n5197) );
  NOR2_X1 U6333 ( .A1(n5287), .A2(n5191), .ZN(n5192) );
  OR2_X1 U6334 ( .A1(n5193), .A2(n5192), .ZN(n5497) );
  AOI22_X1 U6335 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5820), .B1(n5821), 
        .B2(n5385), .ZN(n5195) );
  NAND2_X1 U6336 ( .A1(n5818), .A2(EBX_REG_27__SCAN_IN), .ZN(n5194) );
  OAI211_X1 U6337 ( .C1(n5497), .C2(n5825), .A(n5195), .B(n5194), .ZN(n5196)
         );
  AOI21_X1 U6338 ( .B1(n5197), .B2(REIP_REG_27__SCAN_IN), .A(n5196), .ZN(n5198) );
  OAI211_X1 U6339 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5200), .A(n5199), .B(n5198), .ZN(U2800) );
  NAND2_X1 U6340 ( .A1(n6992), .A2(n5202), .ZN(n5209) );
  INV_X1 U6341 ( .A(n5305), .ZN(n5207) );
  INV_X1 U6342 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5203) );
  OAI22_X1 U6343 ( .A1(n5203), .A2(n5761), .B1(n5075), .B2(n5794), .ZN(n5204)
         );
  AOI21_X1 U6344 ( .B1(n5821), .B2(n5205), .A(n5204), .ZN(n5206) );
  OAI21_X1 U6345 ( .B1(n5207), .B2(n5825), .A(n5206), .ZN(n5208) );
  AOI21_X1 U6346 ( .B1(n5209), .B2(n5617), .A(n5208), .ZN(n5210) );
  OAI21_X1 U6347 ( .B1(n5365), .B2(n5646), .A(n5210), .ZN(U2804) );
  INV_X1 U6348 ( .A(n5211), .ZN(n5212) );
  AOI21_X1 U6349 ( .B1(n5213), .B2(n5283), .A(n5212), .ZN(n5665) );
  INV_X1 U6350 ( .A(n5665), .ZN(n5307) );
  OAI211_X1 U6351 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5629), .B(n5214), .ZN(n5222) );
  OAI21_X1 U6352 ( .B1(n5311), .B2(n5216), .A(n5215), .ZN(n5515) );
  INV_X1 U6353 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5217) );
  OAI22_X1 U6354 ( .A1(n5217), .A2(n5794), .B1(n5813), .B2(n5410), .ZN(n5218)
         );
  AOI21_X1 U6355 ( .B1(n5818), .B2(EBX_REG_22__SCAN_IN), .A(n5218), .ZN(n5219)
         );
  OAI21_X1 U6356 ( .B1(n5515), .B2(n5825), .A(n5219), .ZN(n5220) );
  AOI21_X1 U6357 ( .B1(n5634), .B2(REIP_REG_22__SCAN_IN), .A(n5220), .ZN(n5221) );
  OAI211_X1 U6358 ( .C1(n5307), .C2(n5646), .A(n5222), .B(n5221), .ZN(U2805)
         );
  XOR2_X1 U6359 ( .A(n5224), .B(n5223), .Z(n5844) );
  INV_X1 U6360 ( .A(n5844), .ZN(n5234) );
  NOR2_X1 U6361 ( .A1(n5240), .A2(n5225), .ZN(n5226) );
  OR2_X1 U6362 ( .A1(n5227), .A2(n5226), .ZN(n5557) );
  INV_X1 U6363 ( .A(n5557), .ZN(n5232) );
  AOI22_X1 U6364 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n5820), .B1(n5678), 
        .B2(n5821), .ZN(n5228) );
  OAI211_X1 U6365 ( .C1(n5761), .C2(n5331), .A(n5228), .B(n5791), .ZN(n5231)
         );
  AOI21_X1 U6366 ( .B1(n6969), .B2(n5229), .A(n5652), .ZN(n5230) );
  AOI211_X1 U6367 ( .C1(n5232), .C2(n5790), .A(n5231), .B(n5230), .ZN(n5233)
         );
  OAI21_X1 U6368 ( .B1(n5234), .B2(n5646), .A(n5233), .ZN(U2810) );
  INV_X1 U6369 ( .A(n5849), .ZN(n5334) );
  NOR2_X1 U6370 ( .A1(n5236), .A2(n5235), .ZN(n5758) );
  INV_X1 U6371 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6589) );
  XNOR2_X1 U6372 ( .A(REIP_REG_16__SCAN_IN), .B(n6589), .ZN(n5237) );
  AOI22_X1 U6373 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5758), .B1(n5257), .B2(
        n5237), .ZN(n5247) );
  AND2_X1 U6374 ( .A1(n3203), .A2(n5238), .ZN(n5239) );
  NOR2_X1 U6375 ( .A1(n5240), .A2(n5239), .ZN(n5567) );
  AOI21_X1 U6376 ( .B1(n5241), .B2(n5821), .A(n5803), .ZN(n5243) );
  NAND2_X1 U6377 ( .A1(n5818), .A2(EBX_REG_16__SCAN_IN), .ZN(n5242) );
  OAI211_X1 U6378 ( .C1(n5794), .C2(n5244), .A(n5243), .B(n5242), .ZN(n5245)
         );
  AOI21_X1 U6379 ( .B1(n5567), .B2(n5790), .A(n5245), .ZN(n5246) );
  OAI211_X1 U6380 ( .C1(n5334), .C2(n5646), .A(n5247), .B(n5246), .ZN(U2811)
         );
  INV_X1 U6381 ( .A(n5248), .ZN(n5249) );
  AOI21_X1 U6382 ( .B1(n5250), .B2(n5047), .A(n5249), .ZN(n5443) );
  NAND2_X1 U6383 ( .A1(n5443), .A2(n5810), .ZN(n5259) );
  NAND2_X1 U6384 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  AND2_X1 U6385 ( .A1(n3203), .A2(n5253), .ZN(n5702) );
  AOI22_X1 U6386 ( .A1(n5702), .A2(n5790), .B1(n5818), .B2(EBX_REG_15__SCAN_IN), .ZN(n5254) );
  OAI211_X1 U6387 ( .C1(n5794), .C2(n5255), .A(n5254), .B(n5791), .ZN(n5256)
         );
  AOI221_X1 U6388 ( .B1(n5257), .B2(n6589), .C1(n5758), .C2(
        REIP_REG_15__SCAN_IN), .A(n5256), .ZN(n5258) );
  OAI211_X1 U6389 ( .C1(n5441), .C2(n5813), .A(n5259), .B(n5258), .ZN(U2812)
         );
  OR2_X1 U6390 ( .A1(n4710), .A2(n5260), .ZN(n5261) );
  XOR2_X1 U6391 ( .A(n5262), .B(n5261), .Z(n5461) );
  INV_X1 U6392 ( .A(n5461), .ZN(n5372) );
  INV_X1 U6393 ( .A(n5459), .ZN(n5271) );
  INV_X1 U6394 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5268) );
  INV_X1 U6395 ( .A(n5263), .ZN(n5264) );
  AOI21_X1 U6396 ( .B1(n5266), .B2(n5265), .A(n5264), .ZN(n5956) );
  AOI22_X1 U6397 ( .A1(n5790), .A2(n5956), .B1(n5818), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5267) );
  OAI211_X1 U6398 ( .C1(n5794), .C2(n5268), .A(n5267), .B(n5791), .ZN(n5270)
         );
  INV_X1 U6399 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6580) );
  NOR3_X1 U6400 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5272), .A3(n6580), .ZN(n5269)
         );
  AOI211_X1 U6401 ( .C1(n5821), .C2(n5271), .A(n5270), .B(n5269), .ZN(n5274)
         );
  NOR2_X1 U6402 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5272), .ZN(n5808) );
  OAI21_X1 U6403 ( .B1(n5809), .B2(n5808), .A(REIP_REG_7__SCAN_IN), .ZN(n5273)
         );
  OAI211_X1 U6404 ( .C1(n5372), .C2(n5646), .A(n5274), .B(n5273), .ZN(U2820)
         );
  INV_X1 U6405 ( .A(n5468), .ZN(n5276) );
  OAI22_X1 U6406 ( .A1(n5276), .A2(n5336), .B1(n5275), .B2(n5840), .ZN(U2828)
         );
  OAI222_X1 U6407 ( .A1(n5343), .A2(n5354), .B1(n5840), .B2(n5278), .C1(n5277), 
        .C2(n5336), .ZN(U2829) );
  OAI222_X1 U6408 ( .A1(n5279), .A2(n5840), .B1(n5336), .B2(n5472), .C1(n5165), 
        .C2(n5343), .ZN(U2830) );
  OAI222_X1 U6409 ( .A1(n5280), .A2(n5840), .B1(n5336), .B2(n5486), .C1(n5359), 
        .C2(n5343), .ZN(U2831) );
  INV_X1 U6410 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5281) );
  OAI222_X1 U6411 ( .A1(n5281), .A2(n5840), .B1(n5336), .B2(n5497), .C1(n5362), 
        .C2(n5343), .ZN(U2832) );
  NOR2_X1 U6412 ( .A1(n5283), .A2(n5282), .ZN(n5295) );
  NOR2_X1 U6413 ( .A1(n5295), .A2(n5284), .ZN(n5285) );
  INV_X1 U6414 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5291) );
  INV_X1 U6415 ( .A(n5287), .ZN(n5290) );
  NAND2_X1 U6416 ( .A1(n5300), .A2(n5288), .ZN(n5289) );
  NAND2_X1 U6417 ( .A1(n5290), .A2(n5289), .ZN(n5599) );
  OAI222_X1 U6418 ( .A1(n5343), .A2(n5394), .B1(n5840), .B2(n5291), .C1(n5599), 
        .C2(n5336), .ZN(U2833) );
  NOR2_X1 U6419 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  INV_X1 U6420 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5302) );
  INV_X1 U6421 ( .A(n5296), .ZN(n5298) );
  OAI21_X1 U6422 ( .B1(n5299), .B2(n5298), .A(n5297), .ZN(n5301) );
  NAND2_X1 U6423 ( .A1(n5301), .A2(n5300), .ZN(n5688) );
  OAI222_X1 U6424 ( .A1(n5343), .A2(n5658), .B1(n5840), .B2(n5302), .C1(n5688), 
        .C2(n5336), .ZN(U2834) );
  INV_X1 U6425 ( .A(n5662), .ZN(n5304) );
  AOI22_X1 U6426 ( .A1(n5618), .A2(n5836), .B1(EBX_REG_24__SCAN_IN), .B2(n5341), .ZN(n5303) );
  OAI21_X1 U6427 ( .B1(n5304), .B2(n5343), .A(n5303), .ZN(U2835) );
  AOI22_X1 U6428 ( .A1(n5305), .A2(n5836), .B1(n5341), .B2(EBX_REG_23__SCAN_IN), .ZN(n5306) );
  OAI21_X1 U6429 ( .B1(n5365), .B2(n5343), .A(n5306), .ZN(U2836) );
  INV_X1 U6430 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5308) );
  OAI222_X1 U6431 ( .A1(n5336), .A2(n5515), .B1(n5840), .B2(n5308), .C1(n5307), 
        .C2(n5343), .ZN(U2837) );
  XNOR2_X1 U6432 ( .A(n5309), .B(n5310), .ZN(n5623) );
  INV_X1 U6433 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5313) );
  AOI21_X1 U6434 ( .B1(n3152), .B2(n5312), .A(n5311), .ZN(n5624) );
  INV_X1 U6435 ( .A(n5624), .ZN(n5527) );
  OAI222_X1 U6436 ( .A1(n5343), .A2(n5623), .B1(n5840), .B2(n5313), .C1(n5527), 
        .C2(n5336), .ZN(U2838) );
  INV_X1 U6437 ( .A(n5314), .ZN(n5317) );
  MUX2_X1 U6438 ( .A(n5317), .B(n5316), .S(n5315), .Z(n5319) );
  XNOR2_X1 U6439 ( .A(n5319), .B(n5318), .ZN(n5635) );
  INV_X1 U6440 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5323) );
  NOR2_X1 U6441 ( .A1(n5320), .A2(n5321), .ZN(n5322) );
  OR2_X1 U6442 ( .A1(n5309), .A2(n5322), .ZN(n5632) );
  OAI222_X1 U6443 ( .A1(n5336), .A2(n5635), .B1(n5840), .B2(n5323), .C1(n5343), 
        .C2(n5632), .ZN(U2839) );
  AOI21_X1 U6444 ( .B1(n5324), .B2(n4430), .A(n5320), .ZN(n5435) );
  INV_X1 U6445 ( .A(n5435), .ZN(n5647) );
  XNOR2_X1 U6446 ( .A(n5326), .B(n5325), .ZN(n5695) );
  AOI22_X1 U6447 ( .A1(n5695), .A2(n5836), .B1(n5341), .B2(EBX_REG_19__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U6448 ( .B1(n5647), .B2(n5343), .A(n5327), .ZN(U2840) );
  INV_X1 U6449 ( .A(n5548), .ZN(n5330) );
  OAI222_X1 U6450 ( .A1(n5336), .A2(n5330), .B1(n5840), .B2(n5329), .C1(n5343), 
        .C2(n5328), .ZN(U2841) );
  OAI22_X1 U6451 ( .A1(n5557), .A2(n5336), .B1(n5331), .B2(n5840), .ZN(n5332)
         );
  AOI21_X1 U6452 ( .B1(n5844), .B2(n5837), .A(n5332), .ZN(n5333) );
  INV_X1 U6453 ( .A(n5333), .ZN(U2842) );
  INV_X1 U6454 ( .A(n5567), .ZN(n5337) );
  INV_X1 U6455 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5335) );
  OAI222_X1 U6456 ( .A1(n5337), .A2(n5336), .B1(n5840), .B2(n5335), .C1(n5343), 
        .C2(n5334), .ZN(U2843) );
  INV_X1 U6457 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6458 ( .A1(n5443), .A2(n5837), .ZN(n5339) );
  NAND2_X1 U6459 ( .A1(n5702), .A2(n5836), .ZN(n5338) );
  OAI211_X1 U6460 ( .C1(n5340), .C2(n5840), .A(n5339), .B(n5338), .ZN(U2844)
         );
  AOI22_X1 U6461 ( .A1(n5956), .A2(n5836), .B1(n5341), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5342) );
  OAI21_X1 U6462 ( .B1(n5372), .B2(n5343), .A(n5342), .ZN(U2852) );
  NAND3_X1 U6463 ( .A1(n5345), .A2(n5344), .A3(n5369), .ZN(n5348) );
  AOI22_X1 U6464 ( .A1(n5851), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5850), .ZN(n5347) );
  NAND2_X1 U6465 ( .A1(n5348), .A2(n5347), .ZN(U2860) );
  AND2_X1 U6466 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  AOI22_X1 U6467 ( .A1(n5847), .A2(DATAI_14_), .B1(n5850), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6468 ( .A1(n5851), .A2(DATAI_30_), .ZN(n5352) );
  OAI211_X1 U6469 ( .C1(n5354), .C2(n5653), .A(n5353), .B(n5352), .ZN(U2861)
         );
  AOI22_X1 U6470 ( .A1(n5847), .A2(DATAI_13_), .B1(n5850), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6471 ( .A1(n5851), .A2(DATAI_29_), .ZN(n5355) );
  OAI211_X1 U6472 ( .C1(n5165), .C2(n5653), .A(n5356), .B(n5355), .ZN(U2862)
         );
  AOI22_X1 U6473 ( .A1(n5847), .A2(DATAI_12_), .B1(n5850), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6474 ( .A1(n5851), .A2(DATAI_28_), .ZN(n5357) );
  OAI211_X1 U6475 ( .C1(n5359), .C2(n5653), .A(n5358), .B(n5357), .ZN(U2863)
         );
  AOI22_X1 U6476 ( .A1(n5847), .A2(DATAI_11_), .B1(n5850), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6477 ( .A1(n5851), .A2(DATAI_27_), .ZN(n5360) );
  OAI211_X1 U6478 ( .C1(n5362), .C2(n5653), .A(n5361), .B(n5360), .ZN(U2864)
         );
  AOI22_X1 U6479 ( .A1(n5847), .A2(DATAI_7_), .B1(n5850), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6480 ( .A1(n5851), .A2(DATAI_23_), .ZN(n5363) );
  OAI211_X1 U6481 ( .C1(n5365), .C2(n5653), .A(n5364), .B(n5363), .ZN(U2868)
         );
  AOI22_X1 U6482 ( .A1(n5851), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5850), .ZN(n5367) );
  NAND2_X1 U6483 ( .A1(n5847), .A2(DATAI_3_), .ZN(n5366) );
  OAI211_X1 U6484 ( .C1(n5647), .C2(n5653), .A(n5367), .B(n5366), .ZN(U2872)
         );
  INV_X1 U6485 ( .A(n5443), .ZN(n5368) );
  INV_X1 U6486 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5855) );
  OAI222_X1 U6487 ( .A1(n5368), .A2(n5653), .B1(n5371), .B2(n6927), .C1(n5369), 
        .C2(n5855), .ZN(U2876) );
  OAI222_X1 U6488 ( .A1(n5653), .A2(n5372), .B1(n5371), .B2(n5370), .C1(n5369), 
        .C2(n3764), .ZN(U2884) );
  NAND2_X1 U6489 ( .A1(n5375), .A2(n5391), .ZN(n5501) );
  INV_X1 U6490 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U6491 ( .A(n5377), .B(n5376), .ZN(n5490) );
  NOR2_X1 U6492 ( .A1(n5721), .A2(n6973), .ZN(n5485) );
  AOI21_X1 U6493 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5485), 
        .ZN(n5378) );
  OAI21_X1 U6494 ( .B1(n5915), .B2(n5379), .A(n5378), .ZN(n5380) );
  AOI21_X1 U6495 ( .B1(n5381), .B2(n5910), .A(n5380), .ZN(n5382) );
  OAI21_X1 U6496 ( .B1(n5490), .B2(n5918), .A(n5382), .ZN(U2958) );
  NOR2_X1 U6497 ( .A1(n5383), .A2(n3156), .ZN(n5384) );
  XNOR2_X1 U6498 ( .A(n5384), .B(n5492), .ZN(n5500) );
  INV_X1 U6499 ( .A(n5385), .ZN(n5387) );
  NOR2_X1 U6500 ( .A1(n5721), .A2(n6863), .ZN(n5491) );
  AOI21_X1 U6501 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5491), 
        .ZN(n5386) );
  OAI21_X1 U6502 ( .B1(n5915), .B2(n5387), .A(n5386), .ZN(n5388) );
  AOI21_X1 U6503 ( .B1(n5389), .B2(n5910), .A(n5388), .ZN(n5390) );
  OAI21_X1 U6504 ( .B1(n5500), .B2(n5918), .A(n5390), .ZN(U2959) );
  XNOR2_X1 U6505 ( .A(n5448), .B(n5391), .ZN(n5392) );
  XNOR2_X1 U6506 ( .A(n5393), .B(n5392), .ZN(n5509) );
  INV_X1 U6507 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5395) );
  NOR2_X1 U6508 ( .A1(n5721), .A2(n5395), .ZN(n5505) );
  AOI21_X1 U6509 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5505), 
        .ZN(n5396) );
  OAI21_X1 U6510 ( .B1(n5915), .B2(n5605), .A(n5396), .ZN(n5397) );
  AOI21_X1 U6511 ( .B1(n5654), .B2(n5910), .A(n5397), .ZN(n5398) );
  OAI21_X1 U6512 ( .B1(n5918), .B2(n5509), .A(n5398), .ZN(U2960) );
  AOI21_X1 U6513 ( .B1(n5401), .B2(n5399), .A(n5400), .ZN(n5687) );
  INV_X1 U6514 ( .A(n5658), .ZN(n5609) );
  INV_X1 U6515 ( .A(n5402), .ZN(n5606) );
  AOI22_X1 U6516 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n5403) );
  OAI21_X1 U6517 ( .B1(n5915), .B2(n5606), .A(n5403), .ZN(n5404) );
  AOI21_X1 U6518 ( .B1(n5609), .B2(n5910), .A(n5404), .ZN(n5405) );
  OAI21_X1 U6519 ( .B1(n5687), .B2(n5918), .A(n5405), .ZN(U2961) );
  AOI21_X1 U6520 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5448), .A(n5406), 
        .ZN(n5407) );
  XNOR2_X1 U6521 ( .A(n5408), .B(n5407), .ZN(n5519) );
  INV_X1 U6522 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6887) );
  NOR2_X1 U6523 ( .A1(n5721), .A2(n6887), .ZN(n5514) );
  AOI21_X1 U6524 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5514), 
        .ZN(n5409) );
  OAI21_X1 U6525 ( .B1(n5915), .B2(n5410), .A(n5409), .ZN(n5411) );
  AOI21_X1 U6526 ( .B1(n5665), .B2(n5910), .A(n5411), .ZN(n5412) );
  OAI21_X1 U6527 ( .B1(n5519), .B2(n5918), .A(n5412), .ZN(U2964) );
  OAI21_X1 U6528 ( .B1(n5413), .B2(n5415), .A(n5414), .ZN(n5520) );
  NAND2_X1 U6529 ( .A1(n5520), .A2(n5909), .ZN(n5419) );
  NAND2_X1 U6530 ( .A1(n5990), .A2(REIP_REG_21__SCAN_IN), .ZN(n5521) );
  OAI21_X1 U6531 ( .B1(n5416), .B2(n5627), .A(n5521), .ZN(n5417) );
  AOI21_X1 U6532 ( .B1(n5625), .B2(n5888), .A(n5417), .ZN(n5418) );
  OAI211_X1 U6533 ( .C1(n4644), .C2(n5623), .A(n5419), .B(n5418), .ZN(U2965)
         );
  XNOR2_X1 U6534 ( .A(n5448), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5421)
         );
  XNOR2_X1 U6535 ( .A(n5422), .B(n5421), .ZN(n5528) );
  NAND2_X1 U6536 ( .A1(n5528), .A2(n5909), .ZN(n5426) );
  INV_X1 U6537 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5423) );
  NOR2_X1 U6538 ( .A1(n5721), .A2(n5423), .ZN(n5536) );
  NOR2_X1 U6539 ( .A1(n5915), .A2(n5641), .ZN(n5424) );
  AOI211_X1 U6540 ( .C1(n5921), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5536), 
        .B(n5424), .ZN(n5425) );
  OAI211_X1 U6541 ( .C1(n4644), .C2(n5632), .A(n5426), .B(n5425), .ZN(U2966)
         );
  AOI21_X1 U6542 ( .B1(n5431), .B2(n5430), .A(n5429), .ZN(n5696) );
  INV_X1 U6543 ( .A(n5696), .ZN(n5437) );
  INV_X1 U6544 ( .A(n5642), .ZN(n5433) );
  AOI22_X1 U6545 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5432) );
  OAI21_X1 U6546 ( .B1(n5915), .B2(n5433), .A(n5432), .ZN(n5434) );
  AOI21_X1 U6547 ( .B1(n5435), .B2(n5910), .A(n5434), .ZN(n5436) );
  OAI21_X1 U6548 ( .B1(n5437), .B2(n5918), .A(n5436), .ZN(U2967) );
  XNOR2_X1 U6549 ( .A(n5448), .B(n5706), .ZN(n5438) );
  XNOR2_X1 U6550 ( .A(n5439), .B(n5438), .ZN(n5703) );
  INV_X1 U6551 ( .A(n5703), .ZN(n5445) );
  AOI22_X1 U6552 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5440) );
  OAI21_X1 U6553 ( .B1(n5915), .B2(n5441), .A(n5440), .ZN(n5442) );
  AOI21_X1 U6554 ( .B1(n5443), .B2(n5910), .A(n5442), .ZN(n5444) );
  OAI21_X1 U6555 ( .B1(n5445), .B2(n5918), .A(n5444), .ZN(U2971) );
  XNOR2_X1 U6556 ( .A(n5448), .B(n5447), .ZN(n5449) );
  XNOR2_X1 U6557 ( .A(n5446), .B(n5449), .ZN(n5715) );
  INV_X1 U6558 ( .A(n5450), .ZN(n5765) );
  AOI22_X1 U6559 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n5990), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U6560 ( .B1(n5915), .B2(n5452), .A(n5451), .ZN(n5453) );
  AOI21_X1 U6561 ( .B1(n5765), .B2(n5910), .A(n5453), .ZN(n5454) );
  OAI21_X1 U6562 ( .B1(n5715), .B2(n5918), .A(n5454), .ZN(U2972) );
  OAI21_X1 U6563 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(n5957) );
  NAND2_X1 U6564 ( .A1(n5990), .A2(REIP_REG_7__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U6565 ( .A1(n5921), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5458)
         );
  OAI211_X1 U6566 ( .C1(n5915), .C2(n5459), .A(n5954), .B(n5458), .ZN(n5460)
         );
  AOI21_X1 U6567 ( .B1(n5461), .B2(n5910), .A(n5460), .ZN(n5462) );
  OAI21_X1 U6568 ( .B1(n5957), .B2(n5918), .A(n5462), .ZN(U2979) );
  NOR3_X1 U6569 ( .A1(n5464), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5463), 
        .ZN(n5465) );
  AOI211_X1 U6570 ( .C1(n5467), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5466), .B(n5465), .ZN(n5470) );
  NAND2_X1 U6571 ( .A1(n5468), .A2(n6023), .ZN(n5469) );
  OAI211_X1 U6572 ( .C1(n5471), .C2(n6018), .A(n5470), .B(n5469), .ZN(U2987)
         );
  INV_X1 U6573 ( .A(n5472), .ZN(n5479) );
  AOI21_X1 U6574 ( .B1(n5474), .B2(n5476), .A(n5473), .ZN(n5475) );
  OAI21_X1 U6575 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5478) );
  AOI21_X1 U6576 ( .B1(n5479), .B2(n6023), .A(n5478), .ZN(n5480) );
  OAI21_X1 U6577 ( .B1(n5481), .B2(n6018), .A(n5480), .ZN(U2989) );
  INV_X1 U6578 ( .A(n5493), .ZN(n5483) );
  XNOR2_X1 U6579 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5482) );
  NOR2_X1 U6580 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  AOI211_X1 U6581 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5494), .A(n5485), .B(n5484), .ZN(n5489) );
  INV_X1 U6582 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U6583 ( .A1(n5487), .A2(n6023), .ZN(n5488) );
  OAI211_X1 U6584 ( .C1(n5490), .C2(n6018), .A(n5489), .B(n5488), .ZN(U2990)
         );
  AOI21_X1 U6585 ( .B1(n5493), .B2(n5492), .A(n5491), .ZN(n5496) );
  NAND2_X1 U6586 ( .A1(n5494), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U6587 ( .C1(n5497), .C2(n6009), .A(n5496), .B(n5495), .ZN(n5498)
         );
  INV_X1 U6588 ( .A(n5498), .ZN(n5499) );
  OAI21_X1 U6589 ( .B1(n5500), .B2(n6018), .A(n5499), .ZN(U2991) );
  INV_X1 U6590 ( .A(n5693), .ZN(n5503) );
  AND3_X1 U6591 ( .A1(n5503), .A2(n5502), .A3(n5501), .ZN(n5504) );
  AOI211_X1 U6592 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5686), .A(n5505), .B(n5504), .ZN(n5508) );
  INV_X1 U6593 ( .A(n5599), .ZN(n5506) );
  NAND2_X1 U6594 ( .A1(n5506), .A2(n6023), .ZN(n5507) );
  OAI211_X1 U6595 ( .C1(n5509), .C2(n6018), .A(n5508), .B(n5507), .ZN(U2992)
         );
  INV_X1 U6596 ( .A(n5510), .ZN(n5522) );
  NOR3_X1 U6597 ( .A1(n5522), .A2(n5512), .A3(n5511), .ZN(n5513) );
  AOI211_X1 U6598 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5524), .A(n5514), .B(n5513), .ZN(n5518) );
  INV_X1 U6599 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6600 ( .A1(n5516), .A2(n6023), .ZN(n5517) );
  OAI211_X1 U6601 ( .C1(n5519), .C2(n6018), .A(n5518), .B(n5517), .ZN(U2996)
         );
  NAND2_X1 U6602 ( .A1(n5520), .A2(n6012), .ZN(n5526) );
  OAI21_X1 U6603 ( .B1(n5522), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5521), 
        .ZN(n5523) );
  AOI21_X1 U6604 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5524), .A(n5523), 
        .ZN(n5525) );
  OAI211_X1 U6605 ( .C1(n6009), .C2(n5527), .A(n5526), .B(n5525), .ZN(U2997)
         );
  INV_X1 U6606 ( .A(n5528), .ZN(n5543) );
  NAND2_X1 U6607 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5533), .ZN(n5529) );
  OAI21_X1 U6608 ( .B1(n5530), .B2(n5529), .A(n5992), .ZN(n5531) );
  OAI211_X1 U6609 ( .C1(n5927), .C2(n5533), .A(n5532), .B(n5531), .ZN(n5559)
         );
  NOR2_X1 U6610 ( .A1(n5927), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5534)
         );
  NOR2_X1 U6611 ( .A1(n5559), .A2(n5534), .ZN(n5552) );
  OAI21_X1 U6612 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6005), .A(n5552), 
        .ZN(n5694) );
  NOR2_X1 U6613 ( .A1(n5635), .A2(n6009), .ZN(n5535) );
  AOI211_X1 U6614 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5694), .A(n5536), .B(n5535), .ZN(n5542) );
  INV_X1 U6615 ( .A(n5564), .ZN(n5537) );
  NAND2_X1 U6616 ( .A1(n5537), .A2(n5722), .ZN(n5700) );
  NOR2_X1 U6617 ( .A1(n5573), .A2(n5700), .ZN(n5561) );
  NAND2_X1 U6618 ( .A1(n5561), .A2(n5538), .ZN(n5699) );
  OR3_X1 U6619 ( .A1(n5699), .A2(n5540), .A3(n5539), .ZN(n5541) );
  OAI211_X1 U6620 ( .C1(n5543), .C2(n6018), .A(n5542), .B(n5541), .ZN(U2998)
         );
  NAND3_X1 U6621 ( .A1(n5052), .A2(n5065), .A3(n5569), .ZN(n5553) );
  NOR3_X1 U6622 ( .A1(n5052), .A2(n5065), .A3(n5569), .ZN(n5555) );
  NAND2_X1 U6623 ( .A1(n5555), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5544) );
  OAI21_X1 U6624 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5553), .A(n5544), 
        .ZN(n5545) );
  XNOR2_X1 U6625 ( .A(n5545), .B(n5551), .ZN(n5674) );
  NAND2_X1 U6626 ( .A1(n5674), .A2(n6012), .ZN(n5550) );
  NAND3_X1 U6627 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5561), .A3(n5551), .ZN(n5546) );
  OAI21_X1 U6628 ( .B1(n5721), .B2(n6764), .A(n5546), .ZN(n5547) );
  AOI21_X1 U6629 ( .B1(n5548), .B2(n6023), .A(n5547), .ZN(n5549) );
  OAI211_X1 U6630 ( .C1(n5552), .C2(n5551), .A(n5550), .B(n5549), .ZN(U3000)
         );
  INV_X1 U6631 ( .A(n5553), .ZN(n5554) );
  NOR2_X1 U6632 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  XNOR2_X1 U6633 ( .A(n5556), .B(n5560), .ZN(n5681) );
  OAI22_X1 U6634 ( .A1(n5557), .A2(n6009), .B1(n5721), .B2(n6969), .ZN(n5558)
         );
  AOI21_X1 U6635 ( .B1(n5559), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5558), 
        .ZN(n5563) );
  NAND2_X1 U6636 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  OAI211_X1 U6637 ( .C1(n5681), .C2(n6018), .A(n5563), .B(n5562), .ZN(U3001)
         );
  AOI21_X1 U6638 ( .B1(n5706), .B2(n5569), .A(n5700), .ZN(n5574) );
  AND2_X1 U6639 ( .A1(n5928), .A2(n5564), .ZN(n5565) );
  NOR2_X1 U6640 ( .A1(n5710), .A2(n5565), .ZN(n5707) );
  NOR2_X1 U6641 ( .A1(n5721), .A2(n5054), .ZN(n5566) );
  AOI21_X1 U6642 ( .B1(n5567), .B2(n6023), .A(n5566), .ZN(n5568) );
  OAI21_X1 U6643 ( .B1(n5707), .B2(n5569), .A(n5568), .ZN(n5572) );
  NOR2_X1 U6644 ( .A1(n5570), .A2(n6018), .ZN(n5571) );
  AOI211_X1 U6645 ( .C1(n5574), .C2(n5573), .A(n5572), .B(n5571), .ZN(n5575)
         );
  INV_X1 U6646 ( .A(n5575), .ZN(U3002) );
  OAI211_X1 U6647 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6202), .A(n5578), .B(
        n6612), .ZN(n5576) );
  OAI21_X1 U6648 ( .B1(n5579), .B2(n6029), .A(n5576), .ZN(n5577) );
  MUX2_X1 U6649 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5577), .S(n6610), 
        .Z(U3464) );
  XNOR2_X1 U6650 ( .A(n6027), .B(n5578), .ZN(n5580) );
  OAI22_X1 U6651 ( .A1(n5580), .A2(n6438), .B1(n6030), .B2(n5579), .ZN(n5581)
         );
  MUX2_X1 U6652 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5581), .S(n6610), 
        .Z(U3463) );
  NOR2_X1 U6653 ( .A1(n5583), .A2(n5582), .ZN(n5588) );
  OAI22_X1 U6654 ( .A1(n6507), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n5588), .B2(n3713), .ZN(n5584) );
  AOI21_X1 U6655 ( .B1(n5586), .B2(n5585), .A(n5584), .ZN(n6509) );
  NOR2_X1 U6656 ( .A1(n5587), .A2(n4308), .ZN(n5591) );
  INV_X1 U6657 ( .A(n5588), .ZN(n5589) );
  AOI22_X1 U6658 ( .A1(n5592), .A2(n5591), .B1(n5590), .B2(n5589), .ZN(n5593)
         );
  OAI21_X1 U6659 ( .B1(n6509), .B2(n5732), .A(n5593), .ZN(n5594) );
  MUX2_X1 U6660 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n5594), .S(n5737), 
        .Z(U3460) );
  INV_X1 U6661 ( .A(n5595), .ZN(n5597) );
  OAI22_X1 U6662 ( .A1(n5597), .A2(n5732), .B1(n5596), .B2(n6543), .ZN(n5598)
         );
  MUX2_X1 U6663 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5598), .S(n5737), 
        .Z(U3456) );
  AND2_X1 U6664 ( .A1(n5880), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6665 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5818), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5820), .ZN(n5604) );
  AOI21_X1 U6666 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5608), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5600) );
  OAI22_X1 U6667 ( .A1(n5601), .A2(n5600), .B1(n5599), .B2(n5825), .ZN(n5602)
         );
  AOI21_X1 U6668 ( .B1(n5654), .B2(n5810), .A(n5602), .ZN(n5603) );
  OAI211_X1 U6669 ( .C1(n5605), .C2(n5813), .A(n5604), .B(n5603), .ZN(U2801)
         );
  AOI22_X1 U6670 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5818), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5820), .ZN(n5615) );
  OAI22_X1 U6671 ( .A1(n5688), .A2(n5825), .B1(n5606), .B2(n5813), .ZN(n5607)
         );
  INV_X1 U6672 ( .A(n5607), .ZN(n5614) );
  INV_X1 U6673 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6594) );
  AOI22_X1 U6674 ( .A1(n5609), .A2(n5810), .B1(n5608), .B2(n6594), .ZN(n5613)
         );
  INV_X1 U6675 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U6676 ( .A1(n6747), .A2(n5610), .ZN(n5619) );
  INV_X1 U6677 ( .A(n5619), .ZN(n5611) );
  OAI21_X1 U6678 ( .B1(n5611), .B2(n5617), .A(REIP_REG_25__SCAN_IN), .ZN(n5612) );
  NAND4_X1 U6679 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(U2802)
         );
  AOI22_X1 U6680 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5818), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5820), .ZN(n5622) );
  AOI22_X1 U6681 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5617), .B1(n5616), .B2(
        n5821), .ZN(n5621) );
  AOI22_X1 U6682 ( .A1(n5662), .A2(n5810), .B1(n5790), .B2(n5618), .ZN(n5620)
         );
  NAND4_X1 U6683 ( .A1(n5622), .A2(n5621), .A3(n5620), .A4(n5619), .ZN(U2803)
         );
  INV_X1 U6684 ( .A(n5623), .ZN(n5668) );
  AOI22_X1 U6685 ( .A1(n5668), .A2(n5810), .B1(n5624), .B2(n5790), .ZN(n5631)
         );
  INV_X1 U6686 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6897) );
  AOI22_X1 U6687 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5818), .B1(n5625), .B2(n5821), .ZN(n5626) );
  OAI21_X1 U6688 ( .B1(n5627), .B2(n5794), .A(n5626), .ZN(n5628) );
  AOI221_X1 U6689 ( .B1(n5634), .B2(REIP_REG_21__SCAN_IN), .C1(n5629), .C2(
        n6897), .A(n5628), .ZN(n5630) );
  NAND2_X1 U6690 ( .A1(n5631), .A2(n5630), .ZN(U2806) );
  AOI22_X1 U6691 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5818), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5820), .ZN(n5640) );
  INV_X1 U6692 ( .A(n5632), .ZN(n5671) );
  INV_X1 U6693 ( .A(n5645), .ZN(n5633) );
  AOI21_X1 U6694 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5633), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5637) );
  INV_X1 U6695 ( .A(n5634), .ZN(n5636) );
  OAI22_X1 U6696 ( .A1(n5637), .A2(n5636), .B1(n5635), .B2(n5825), .ZN(n5638)
         );
  AOI21_X1 U6697 ( .B1(n5671), .B2(n5810), .A(n5638), .ZN(n5639) );
  OAI211_X1 U6698 ( .C1(n5641), .C2(n5813), .A(n5640), .B(n5639), .ZN(U2807)
         );
  INV_X1 U6699 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6727) );
  INV_X1 U6700 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5644) );
  AOI22_X1 U6701 ( .A1(n5695), .A2(n5790), .B1(n5821), .B2(n5642), .ZN(n5643)
         );
  OAI211_X1 U6702 ( .C1(n5794), .C2(n5644), .A(n5643), .B(n5791), .ZN(n5649)
         );
  OAI22_X1 U6703 ( .A1(n5647), .A2(n5646), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5645), .ZN(n5648) );
  AOI211_X1 U6704 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5818), .A(n5649), .B(n5648), 
        .ZN(n5650) );
  OAI221_X1 U6705 ( .B1(n6727), .B2(n5652), .C1(n6727), .C2(n5651), .A(n5650), 
        .ZN(U2808) );
  AOI22_X1 U6706 ( .A1(n5654), .A2(n5848), .B1(n5847), .B2(DATAI_10_), .ZN(
        n5656) );
  AOI22_X1 U6707 ( .A1(n5851), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5850), .ZN(n5655) );
  NAND2_X1 U6708 ( .A1(n5656), .A2(n5655), .ZN(U2865) );
  INV_X1 U6709 ( .A(n5847), .ZN(n5657) );
  OAI22_X1 U6710 ( .A1(n5658), .A2(n5653), .B1(n5657), .B2(n6895), .ZN(n5659)
         );
  INV_X1 U6711 ( .A(n5659), .ZN(n5661) );
  AOI22_X1 U6712 ( .A1(n5851), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5850), .ZN(n5660) );
  NAND2_X1 U6713 ( .A1(n5661), .A2(n5660), .ZN(U2866) );
  AOI22_X1 U6714 ( .A1(n5662), .A2(n5848), .B1(n5847), .B2(DATAI_8_), .ZN(
        n5664) );
  AOI22_X1 U6715 ( .A1(n5851), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5850), .ZN(n5663) );
  NAND2_X1 U6716 ( .A1(n5664), .A2(n5663), .ZN(U2867) );
  AOI22_X1 U6717 ( .A1(n5665), .A2(n5848), .B1(n5847), .B2(DATAI_6_), .ZN(
        n5667) );
  AOI22_X1 U6718 ( .A1(n5851), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5850), .ZN(n5666) );
  NAND2_X1 U6719 ( .A1(n5667), .A2(n5666), .ZN(U2869) );
  AOI22_X1 U6720 ( .A1(n5668), .A2(n5848), .B1(n5847), .B2(DATAI_5_), .ZN(
        n5670) );
  AOI22_X1 U6721 ( .A1(n5851), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5850), .ZN(n5669) );
  NAND2_X1 U6722 ( .A1(n5670), .A2(n5669), .ZN(U2870) );
  AOI22_X1 U6723 ( .A1(n5671), .A2(n5848), .B1(n5847), .B2(DATAI_4_), .ZN(
        n5673) );
  AOI22_X1 U6724 ( .A1(n5851), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5850), .ZN(n5672) );
  NAND2_X1 U6725 ( .A1(n5673), .A2(n5672), .ZN(U2871) );
  AOI22_X1 U6726 ( .A1(n5990), .A2(REIP_REG_18__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5676) );
  AOI22_X1 U6727 ( .A1(n5674), .A2(n5909), .B1(n5910), .B2(n5841), .ZN(n5675)
         );
  OAI211_X1 U6728 ( .C1(n5915), .C2(n5677), .A(n5676), .B(n5675), .ZN(U2968)
         );
  AOI22_X1 U6729 ( .A1(n5990), .A2(REIP_REG_17__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5680) );
  AOI22_X1 U6730 ( .A1(n5844), .A2(n5910), .B1(n5888), .B2(n5678), .ZN(n5679)
         );
  OAI211_X1 U6731 ( .C1(n5681), .C2(n5918), .A(n5680), .B(n5679), .ZN(U2969)
         );
  AOI22_X1 U6732 ( .A1(n5990), .A2(REIP_REG_13__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U6733 ( .A(n5682), .B(n5683), .ZN(n5728) );
  AOI22_X1 U6734 ( .A1(n5728), .A2(n5909), .B1(n5910), .B2(n5832), .ZN(n5684)
         );
  OAI211_X1 U6735 ( .C1(n5915), .C2(n5780), .A(n5685), .B(n5684), .ZN(U2973)
         );
  AOI22_X1 U6736 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5686), .B1(n5990), .B2(REIP_REG_25__SCAN_IN), .ZN(n5692) );
  INV_X1 U6737 ( .A(n5687), .ZN(n5690) );
  INV_X1 U6738 ( .A(n5688), .ZN(n5689) );
  AOI22_X1 U6739 ( .A1(n5690), .A2(n6012), .B1(n6023), .B2(n5689), .ZN(n5691)
         );
  OAI211_X1 U6740 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5693), .A(n5692), .B(n5691), .ZN(U2993) );
  AOI22_X1 U6741 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5694), .B1(n5990), .B2(REIP_REG_19__SCAN_IN), .ZN(n5698) );
  AOI22_X1 U6742 ( .A1(n5696), .A2(n6012), .B1(n6023), .B2(n5695), .ZN(n5697)
         );
  OAI211_X1 U6743 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5699), .A(n5698), .B(n5697), .ZN(U2999) );
  INV_X1 U6744 ( .A(n5700), .ZN(n5701) );
  AOI22_X1 U6745 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5990), .B1(n5701), .B2(
        n5706), .ZN(n5705) );
  AOI22_X1 U6746 ( .A1(n5703), .A2(n6012), .B1(n6023), .B2(n5702), .ZN(n5704)
         );
  OAI211_X1 U6747 ( .C1(n5707), .C2(n5706), .A(n5705), .B(n5704), .ZN(U3003)
         );
  NOR2_X1 U6748 ( .A1(n5712), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5723)
         );
  INV_X1 U6749 ( .A(n5723), .ZN(n5713) );
  NAND2_X1 U6750 ( .A1(n5709), .A2(n5708), .ZN(n6003) );
  NOR2_X1 U6751 ( .A1(n5718), .A2(n6025), .ZN(n5711) );
  AOI211_X1 U6752 ( .C1(n5712), .C2(n6003), .A(n5711), .B(n5710), .ZN(n5731)
         );
  OAI21_X1 U6753 ( .B1(n5714), .B2(n5713), .A(n5731), .ZN(n5717) );
  OAI22_X1 U6754 ( .A1(n5715), .A2(n6018), .B1(n6009), .B2(n5760), .ZN(n5716)
         );
  AOI21_X1 U6755 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5717), .A(n5716), 
        .ZN(n5720) );
  NAND3_X1 U6756 ( .A1(n5718), .A2(n5447), .A3(n5722), .ZN(n5719) );
  OAI211_X1 U6757 ( .C1(n6588), .C2(n5721), .A(n5720), .B(n5719), .ZN(U3004)
         );
  AOI22_X1 U6758 ( .A1(n5990), .A2(REIP_REG_13__SCAN_IN), .B1(n5723), .B2(
        n5722), .ZN(n5730) );
  AND2_X1 U6759 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  NOR2_X1 U6760 ( .A1(n5727), .A2(n5726), .ZN(n5831) );
  AOI22_X1 U6761 ( .A1(n5728), .A2(n6012), .B1(n6023), .B2(n5831), .ZN(n5729)
         );
  OAI211_X1 U6762 ( .C1(n5731), .C2(n3641), .A(n5730), .B(n5729), .ZN(U3005)
         );
  OR3_X1 U6763 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n5735) );
  OAI21_X1 U6764 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(U3455) );
  INV_X1 U6765 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6965) );
  INV_X1 U6766 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6872) );
  NAND2_X1 U6767 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6575), .ZN(n5738) );
  AOI21_X2 U6768 ( .B1(STATE_REG_0__SCAN_IN), .B2(n5738), .A(n7027), .ZN(n6605) );
  INV_X1 U6769 ( .A(n6605), .ZN(n6603) );
  OAI21_X1 U6770 ( .B1(n7027), .B2(n6872), .A(n6603), .ZN(U2789) );
  INV_X1 U6771 ( .A(n6549), .ZN(n5741) );
  INV_X1 U6772 ( .A(n6548), .ZN(n6546) );
  OAI21_X1 U6773 ( .B1(n5739), .B2(n6546), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5740) );
  OAI21_X1 U6774 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5741), .A(n5740), .ZN(
        U2790) );
  NOR2_X1 U6775 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5743) );
  OAI21_X1 U6776 ( .B1(n5743), .B2(D_C_N_REG_SCAN_IN), .A(n7026), .ZN(n5742)
         );
  OAI21_X1 U6777 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7026), .A(n5742), .ZN(
        U2791) );
  OAI21_X1 U6778 ( .B1(BS16_N), .B2(n5743), .A(n6605), .ZN(n6604) );
  OAI21_X1 U6779 ( .B1(n6605), .B2(n6793), .A(n6604), .ZN(U2792) );
  OAI21_X1 U6780 ( .B1(n5744), .B2(n6721), .A(n5918), .ZN(U2793) );
  NOR4_X1 U6781 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(n5748) );
  NOR4_X1 U6782 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5747)
         );
  NOR4_X1 U6783 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5746) );
  NOR4_X1 U6784 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5745) );
  NAND4_X1 U6785 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(n5754)
         );
  NOR4_X1 U6786 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n5752) );
  AOI211_X1 U6787 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_8__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n5751) );
  NOR4_X1 U6788 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5750) );
  NOR4_X1 U6789 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(n5749) );
  NAND4_X1 U6790 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n5753)
         );
  NOR2_X1 U6791 ( .A1(n5754), .A2(n5753), .ZN(n6624) );
  INV_X1 U6792 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6736) );
  NOR3_X1 U6793 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5756) );
  OAI21_X1 U6794 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5756), .A(n6624), .ZN(n5755)
         );
  OAI21_X1 U6795 ( .B1(n6624), .B2(n6736), .A(n5755), .ZN(U2794) );
  INV_X1 U6796 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6883) );
  AOI21_X1 U6797 ( .B1(n6576), .B2(n6883), .A(n5756), .ZN(n5757) );
  INV_X1 U6798 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6741) );
  INV_X1 U6799 ( .A(n6624), .ZN(n6622) );
  AOI22_X1 U6800 ( .A1(n6624), .A2(n5757), .B1(n6741), .B2(n6622), .ZN(U2795)
         );
  INV_X1 U6801 ( .A(n5758), .ZN(n5759) );
  OAI222_X1 U6802 ( .A1(n5762), .A2(n5761), .B1(n5760), .B2(n5825), .C1(n6588), 
        .C2(n5759), .ZN(n5763) );
  AOI211_X1 U6803 ( .C1(n5820), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5803), 
        .B(n5763), .ZN(n5767) );
  AOI22_X1 U6804 ( .A1(n5765), .A2(n5810), .B1(n5821), .B2(n5764), .ZN(n5766)
         );
  OAI211_X1 U6805 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5768), .A(n5767), .B(n5766), .ZN(U2813) );
  INV_X1 U6806 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U6807 ( .A1(n5818), .A2(EBX_REG_13__SCAN_IN), .ZN(n5770) );
  AOI21_X1 U6808 ( .B1(n5820), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5803), 
        .ZN(n5769) );
  NAND2_X1 U6809 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  AOI21_X1 U6810 ( .B1(n5831), .B2(n5790), .A(n5771), .ZN(n5772) );
  OAI21_X1 U6811 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  AOI21_X1 U6812 ( .B1(n5832), .B2(n5810), .A(n5775), .ZN(n5779) );
  OAI211_X1 U6813 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n5777), .B(n5776), .ZN(n5778) );
  OAI211_X1 U6814 ( .C1(n5813), .C2(n5780), .A(n5779), .B(n5778), .ZN(U2814)
         );
  AOI22_X1 U6815 ( .A1(n5889), .A2(n5810), .B1(n5821), .B2(n5887), .ZN(n5788)
         );
  NOR3_X1 U6816 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5802), .A3(n5781), .ZN(n5786) );
  AOI22_X1 U6817 ( .A1(n5782), .A2(REIP_REG_11__SCAN_IN), .B1(n5790), .B2(
        n5835), .ZN(n5783) );
  OAI211_X1 U6818 ( .C1(n5794), .C2(n5784), .A(n5783), .B(n5791), .ZN(n5785)
         );
  AOI211_X1 U6819 ( .C1(n5818), .C2(EBX_REG_11__SCAN_IN), .A(n5786), .B(n5785), 
        .ZN(n5787) );
  NAND2_X1 U6820 ( .A1(n5788), .A2(n5787), .ZN(U2816) );
  INV_X1 U6821 ( .A(n5789), .ZN(n5938) );
  AOI22_X1 U6822 ( .A1(n5938), .A2(n5790), .B1(n5818), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5792) );
  OAI211_X1 U6823 ( .C1(n5794), .C2(n5793), .A(n5792), .B(n5791), .ZN(n5795)
         );
  AOI21_X1 U6824 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5796), .A(n5795), .ZN(n5801)
         );
  INV_X1 U6825 ( .A(n5797), .ZN(n5799) );
  AOI22_X1 U6826 ( .A1(n5799), .A2(n5810), .B1(n5821), .B2(n5798), .ZN(n5800)
         );
  OAI211_X1 U6827 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5802), .A(n5801), .B(n5800), 
        .ZN(U2818) );
  AOI21_X1 U6828 ( .B1(n5820), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5803), 
        .ZN(n5805) );
  NAND2_X1 U6829 ( .A1(n5818), .A2(EBX_REG_6__SCAN_IN), .ZN(n5804) );
  OAI211_X1 U6830 ( .C1(n5825), .C2(n5806), .A(n5805), .B(n5804), .ZN(n5807)
         );
  AOI211_X1 U6831 ( .C1(n5809), .C2(REIP_REG_6__SCAN_IN), .A(n5808), .B(n5807), 
        .ZN(n5812) );
  NAND2_X1 U6832 ( .A1(n5893), .A2(n5810), .ZN(n5811) );
  OAI211_X1 U6833 ( .C1(n5813), .C2(n5897), .A(n5812), .B(n5811), .ZN(U2821)
         );
  INV_X1 U6834 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6578) );
  INV_X1 U6835 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U6836 ( .A1(n5815), .A2(REIP_REG_2__SCAN_IN), .ZN(n5829) );
  INV_X1 U6837 ( .A(n5816), .ZN(n5902) );
  INV_X1 U6838 ( .A(n5817), .ZN(n5827) );
  AOI22_X1 U6839 ( .A1(n5819), .A2(n6392), .B1(n5818), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5824) );
  INV_X1 U6840 ( .A(n5905), .ZN(n5822) );
  AOI22_X1 U6841 ( .A1(n5822), .A2(n5821), .B1(n5820), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U6842 ( .C1(n5825), .C2(n5982), .A(n5824), .B(n5823), .ZN(n5826)
         );
  AOI21_X1 U6843 ( .B1(n5902), .B2(n5827), .A(n5826), .ZN(n5828) );
  OAI221_X1 U6844 ( .B1(n5830), .B2(n6578), .C1(n5830), .C2(n5829), .A(n5828), 
        .ZN(U2824) );
  INV_X1 U6845 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5834) );
  AOI22_X1 U6846 ( .A1(n5832), .A2(n5837), .B1(n5836), .B2(n5831), .ZN(n5833)
         );
  OAI21_X1 U6847 ( .B1(n5840), .B2(n5834), .A(n5833), .ZN(U2846) );
  INV_X1 U6848 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5839) );
  AOI22_X1 U6849 ( .A1(n5889), .A2(n5837), .B1(n5836), .B2(n5835), .ZN(n5838)
         );
  OAI21_X1 U6850 ( .B1(n5840), .B2(n5839), .A(n5838), .ZN(U2848) );
  AOI22_X1 U6851 ( .A1(n5841), .A2(n5848), .B1(n5847), .B2(DATAI_2_), .ZN(
        n5843) );
  AOI22_X1 U6852 ( .A1(n5851), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5850), .ZN(n5842) );
  NAND2_X1 U6853 ( .A1(n5843), .A2(n5842), .ZN(U2873) );
  AOI22_X1 U6854 ( .A1(n5844), .A2(n5848), .B1(n5847), .B2(DATAI_1_), .ZN(
        n5846) );
  AOI22_X1 U6855 ( .A1(n5851), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5850), .ZN(n5845) );
  NAND2_X1 U6856 ( .A1(n5846), .A2(n5845), .ZN(U2874) );
  AOI22_X1 U6857 ( .A1(n5849), .A2(n5848), .B1(n5847), .B2(DATAI_0_), .ZN(
        n5853) );
  AOI22_X1 U6858 ( .A1(n5851), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5850), .ZN(n5852) );
  NAND2_X1 U6859 ( .A1(n5853), .A2(n5852), .ZN(U2875) );
  AOI22_X1 U6860 ( .A1(n6534), .A2(LWORD_REG_15__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5854) );
  OAI21_X1 U6861 ( .B1(n5855), .B2(n5885), .A(n5854), .ZN(U2908) );
  AOI22_X1 U6862 ( .A1(n6534), .A2(LWORD_REG_14__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U6863 ( .B1(n5857), .B2(n5885), .A(n5856), .ZN(U2909) );
  AOI22_X1 U6864 ( .A1(n6534), .A2(LWORD_REG_13__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5858) );
  OAI21_X1 U6865 ( .B1(n5859), .B2(n5885), .A(n5858), .ZN(U2910) );
  AOI22_X1 U6866 ( .A1(n6534), .A2(LWORD_REG_12__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U6867 ( .B1(n3838), .B2(n5885), .A(n5860), .ZN(U2911) );
  AOI22_X1 U6868 ( .A1(n6534), .A2(LWORD_REG_11__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5861) );
  OAI21_X1 U6869 ( .B1(n5862), .B2(n5885), .A(n5861), .ZN(U2912) );
  AOI22_X1 U6870 ( .A1(n6534), .A2(LWORD_REG_10__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5863) );
  OAI21_X1 U6871 ( .B1(n5864), .B2(n5885), .A(n5863), .ZN(U2913) );
  AOI22_X1 U6872 ( .A1(n6534), .A2(LWORD_REG_9__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5865) );
  OAI21_X1 U6873 ( .B1(n5866), .B2(n5885), .A(n5865), .ZN(U2914) );
  AOI22_X1 U6874 ( .A1(n6534), .A2(LWORD_REG_8__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5867) );
  OAI21_X1 U6875 ( .B1(n5868), .B2(n5885), .A(n5867), .ZN(U2915) );
  AOI22_X1 U6876 ( .A1(n6534), .A2(LWORD_REG_7__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U6877 ( .B1(n3764), .B2(n5885), .A(n5869), .ZN(U2916) );
  AOI22_X1 U6878 ( .A1(n6534), .A2(LWORD_REG_6__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U6879 ( .B1(n5871), .B2(n5885), .A(n5870), .ZN(U2917) );
  AOI22_X1 U6880 ( .A1(n6534), .A2(LWORD_REG_5__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5872) );
  OAI21_X1 U6881 ( .B1(n5873), .B2(n5885), .A(n5872), .ZN(U2918) );
  AOI22_X1 U6882 ( .A1(n6534), .A2(LWORD_REG_4__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5874) );
  OAI21_X1 U6883 ( .B1(n5875), .B2(n5885), .A(n5874), .ZN(U2919) );
  AOI22_X1 U6884 ( .A1(n6534), .A2(LWORD_REG_3__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5876) );
  OAI21_X1 U6885 ( .B1(n5877), .B2(n5885), .A(n5876), .ZN(U2920) );
  AOI22_X1 U6886 ( .A1(n6534), .A2(LWORD_REG_2__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6887 ( .B1(n5879), .B2(n5885), .A(n5878), .ZN(U2921) );
  AOI22_X1 U6888 ( .A1(n6534), .A2(LWORD_REG_1__SCAN_IN), .B1(n5880), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5881) );
  OAI21_X1 U6889 ( .B1(n5882), .B2(n5885), .A(n5881), .ZN(U2922) );
  AOI22_X1 U6890 ( .A1(n6534), .A2(LWORD_REG_0__SCAN_IN), .B1(n5883), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U6891 ( .B1(n5886), .B2(n5885), .A(n5884), .ZN(U2923) );
  AOI22_X1 U6892 ( .A1(n5990), .A2(REIP_REG_11__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5891) );
  AOI22_X1 U6893 ( .A1(n5889), .A2(n5910), .B1(n5888), .B2(n5887), .ZN(n5890)
         );
  OAI211_X1 U6894 ( .C1(n5892), .C2(n5918), .A(n5891), .B(n5890), .ZN(U2975)
         );
  AOI22_X1 U6895 ( .A1(n5990), .A2(REIP_REG_6__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5896) );
  AOI22_X1 U6896 ( .A1(n5894), .A2(n5909), .B1(n5893), .B2(n5910), .ZN(n5895)
         );
  OAI211_X1 U6897 ( .C1(n5915), .C2(n5897), .A(n5896), .B(n5895), .ZN(U2980)
         );
  AOI22_X1 U6898 ( .A1(n5990), .A2(REIP_REG_3__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U6899 ( .B1(n5900), .B2(n5898), .A(n5899), .ZN(n5901) );
  INV_X1 U6900 ( .A(n5901), .ZN(n5984) );
  AOI22_X1 U6901 ( .A1(n5909), .A2(n5984), .B1(n5902), .B2(n5910), .ZN(n5903)
         );
  OAI211_X1 U6902 ( .C1(n5915), .C2(n5905), .A(n5904), .B(n5903), .ZN(U2983)
         );
  AOI22_X1 U6903 ( .A1(n5990), .A2(REIP_REG_2__SCAN_IN), .B1(n5921), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5913) );
  XNOR2_X1 U6904 ( .A(n5906), .B(n5997), .ZN(n5907) );
  XNOR2_X1 U6905 ( .A(n5908), .B(n5907), .ZN(n5995) );
  AOI22_X1 U6906 ( .A1(n5911), .A2(n5910), .B1(n5909), .B2(n5995), .ZN(n5912)
         );
  OAI211_X1 U6907 ( .C1(n5915), .C2(n5914), .A(n5913), .B(n5912), .ZN(U2984)
         );
  XNOR2_X1 U6908 ( .A(n5916), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6017)
         );
  OAI22_X1 U6909 ( .A1(n5918), .A2(n6017), .B1(n4644), .B2(n5917), .ZN(n5919)
         );
  AOI221_X1 U6910 ( .B1(n5921), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n5920), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5919), .ZN(n5922) );
  NAND2_X1 U6911 ( .A1(n5990), .A2(REIP_REG_0__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U6912 ( .A1(n5922), .A2(n6016), .ZN(U2986) );
  INV_X1 U6913 ( .A(n5923), .ZN(n5931) );
  AOI21_X1 U6914 ( .B1(n5992), .B2(n5931), .A(n5924), .ZN(n5925) );
  OAI21_X1 U6915 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5958) );
  AOI21_X1 U6916 ( .B1(n5945), .B2(n5928), .A(n5958), .ZN(n5944) );
  INV_X1 U6917 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5935) );
  AOI222_X1 U6918 ( .A1(n5930), .A2(n6012), .B1(n6023), .B2(n5929), .C1(
        REIP_REG_10__SCAN_IN), .C2(n5990), .ZN(n5934) );
  NOR2_X1 U6919 ( .A1(n5945), .A2(n5962), .ZN(n5939) );
  OAI211_X1 U6920 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5939), .B(n5932), .ZN(n5933) );
  OAI211_X1 U6921 ( .C1(n5944), .C2(n5935), .A(n5934), .B(n5933), .ZN(U3008)
         );
  INV_X1 U6922 ( .A(n5936), .ZN(n5937) );
  AOI21_X1 U6923 ( .B1(n5938), .B2(n6023), .A(n5937), .ZN(n5942) );
  AOI22_X1 U6924 ( .A1(n5940), .A2(n6012), .B1(n5939), .B2(n5943), .ZN(n5941)
         );
  OAI211_X1 U6925 ( .C1(n5944), .C2(n5943), .A(n5942), .B(n5941), .ZN(U3009)
         );
  OAI21_X1 U6926 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5945), .ZN(n5953) );
  INV_X1 U6927 ( .A(n5946), .ZN(n5947) );
  AOI21_X1 U6928 ( .B1(n6023), .B2(n5948), .A(n5947), .ZN(n5952) );
  INV_X1 U6929 ( .A(n5949), .ZN(n5950) );
  AOI22_X1 U6930 ( .A1(n5950), .A2(n6012), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n5958), .ZN(n5951) );
  OAI211_X1 U6931 ( .C1(n5962), .C2(n5953), .A(n5952), .B(n5951), .ZN(U3010)
         );
  INV_X1 U6932 ( .A(n5954), .ZN(n5955) );
  AOI21_X1 U6933 ( .B1(n5956), .B2(n6023), .A(n5955), .ZN(n5961) );
  INV_X1 U6934 ( .A(n5957), .ZN(n5959) );
  AOI22_X1 U6935 ( .A1(n5959), .A2(n6012), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n5958), .ZN(n5960) );
  OAI211_X1 U6936 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n5962), .A(n5961), 
        .B(n5960), .ZN(U3011) );
  OAI21_X1 U6937 ( .B1(n5965), .B2(n5964), .A(n5963), .ZN(n5966) );
  AOI21_X1 U6938 ( .B1(n5992), .B2(n5967), .A(n5966), .ZN(n5972) );
  INV_X1 U6939 ( .A(n5968), .ZN(n5969) );
  AOI22_X1 U6940 ( .A1(n5969), .A2(n6012), .B1(n6023), .B2(n3201), .ZN(n5971)
         );
  NAND2_X1 U6941 ( .A1(n5990), .A2(REIP_REG_5__SCAN_IN), .ZN(n5970) );
  OAI211_X1 U6942 ( .C1(n5973), .C2(n5972), .A(n5971), .B(n5970), .ZN(U3013)
         );
  AOI21_X1 U6943 ( .B1(n5992), .B2(n5994), .A(n5996), .ZN(n5989) );
  INV_X1 U6944 ( .A(n5974), .ZN(n5975) );
  AOI222_X1 U6945 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5990), .B1(n6023), .B2(
        n5976), .C1(n6012), .C2(n5975), .ZN(n5980) );
  NOR2_X1 U6946 ( .A1(n5994), .A2(n5977), .ZN(n5985) );
  OAI211_X1 U6947 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5985), .B(n5978), .ZN(n5979) );
  OAI211_X1 U6948 ( .C1(n5989), .C2(n5981), .A(n5980), .B(n5979), .ZN(U3014)
         );
  INV_X1 U6949 ( .A(n5982), .ZN(n5983) );
  AOI22_X1 U6950 ( .A1(n6023), .A2(n5983), .B1(n5990), .B2(REIP_REG_3__SCAN_IN), .ZN(n5987) );
  AOI22_X1 U6951 ( .A1(n5985), .A2(n5988), .B1(n5984), .B2(n6012), .ZN(n5986)
         );
  OAI211_X1 U6952 ( .C1(n5989), .C2(n5988), .A(n5987), .B(n5986), .ZN(U3015)
         );
  AOI22_X1 U6953 ( .A1(n6023), .A2(n5991), .B1(n5990), .B2(REIP_REG_2__SCAN_IN), .ZN(n6002) );
  OAI221_X1 U6954 ( .B1(n5994), .B2(n5993), .C1(n5994), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5992), .ZN(n6001) );
  AOI22_X1 U6955 ( .A1(n5996), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6012), 
        .B2(n5995), .ZN(n6000) );
  NAND3_X1 U6956 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5998), .A3(n5997), 
        .ZN(n5999) );
  NAND4_X1 U6957 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(U3016)
         );
  NAND2_X1 U6958 ( .A1(n4308), .A2(n6003), .ZN(n6019) );
  NOR3_X1 U6959 ( .A1(n6005), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6004), 
        .ZN(n6011) );
  INV_X1 U6960 ( .A(n6006), .ZN(n6008) );
  OAI21_X1 U6961 ( .B1(n6009), .B2(n6008), .A(n6007), .ZN(n6010) );
  AOI211_X1 U6962 ( .C1(n6013), .C2(n6012), .A(n6011), .B(n6010), .ZN(n6014)
         );
  OAI221_X1 U6963 ( .B1(n6015), .B2(n6026), .C1(n6015), .C2(n6019), .A(n6014), 
        .ZN(U3017) );
  OAI21_X1 U6964 ( .B1(n6018), .B2(n6017), .A(n6016), .ZN(n6021) );
  INV_X1 U6965 ( .A(n6019), .ZN(n6020) );
  AOI211_X1 U6966 ( .C1(n6023), .C2(n6022), .A(n6021), .B(n6020), .ZN(n6024)
         );
  OAI221_X1 U6967 ( .B1(n4308), .B2(n6026), .C1(n4308), .C2(n6025), .A(n6024), 
        .ZN(U3018) );
  INV_X1 U6968 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6523) );
  NOR2_X1 U6969 ( .A1(n6523), .A2(n6610), .ZN(U3019) );
  NAND2_X1 U6970 ( .A1(n6027), .A2(n6238), .ZN(n6028) );
  NAND3_X1 U6971 ( .A1(n6525), .A2(n6517), .A3(n6512), .ZN(n6066) );
  NOR2_X1 U6972 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6066), .ZN(n6055)
         );
  NAND2_X1 U6973 ( .A1(n6030), .A2(n6029), .ZN(n6206) );
  INV_X1 U6974 ( .A(n6206), .ZN(n6237) );
  NAND2_X1 U6975 ( .A1(n6207), .A2(n6237), .ZN(n6060) );
  INV_X1 U6976 ( .A(n6287), .ZN(n6330) );
  INV_X1 U6977 ( .A(n6031), .ZN(n6032) );
  OAI22_X1 U6978 ( .A1(n6060), .A2(n6438), .B1(n6330), .B2(n6032), .ZN(n6054)
         );
  AOI22_X1 U6979 ( .A1(n6440), .A2(n6055), .B1(n6439), .B2(n6054), .ZN(n6041)
         );
  INV_X1 U6980 ( .A(n6090), .ZN(n6034) );
  AND2_X1 U6981 ( .A1(n6383), .A2(n6611), .ZN(n6033) );
  OAI21_X1 U6982 ( .B1(n6034), .B2(n6492), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6035) );
  NAND3_X1 U6983 ( .A1(n6035), .A2(n6612), .A3(n6060), .ZN(n6039) );
  INV_X1 U6984 ( .A(n6055), .ZN(n6037) );
  AOI211_X1 U6985 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6037), .A(n6386), .B(
        n6036), .ZN(n6038) );
  NAND2_X1 U6986 ( .A1(n6039), .A2(n6038), .ZN(n6056) );
  AOI22_X1 U6987 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n6056), .B1(n6397), 
        .B2(n6492), .ZN(n6040) );
  OAI211_X1 U6988 ( .C1(n6400), .C2(n6090), .A(n6041), .B(n6040), .ZN(U3020)
         );
  AOI22_X1 U6989 ( .A1(n6453), .A2(n6055), .B1(n6452), .B2(n6054), .ZN(n6043)
         );
  AOI22_X1 U6990 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n6056), .B1(n6401), 
        .B2(n6492), .ZN(n6042) );
  OAI211_X1 U6991 ( .C1(n6404), .C2(n6090), .A(n6043), .B(n6042), .ZN(U3021)
         );
  AOI22_X1 U6992 ( .A1(n6459), .A2(n6055), .B1(n6458), .B2(n6054), .ZN(n6045)
         );
  AOI22_X1 U6993 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n6056), .B1(n6405), 
        .B2(n6492), .ZN(n6044) );
  OAI211_X1 U6994 ( .C1(n6408), .C2(n6090), .A(n6045), .B(n6044), .ZN(U3022)
         );
  AOI22_X1 U6995 ( .A1(n6465), .A2(n6055), .B1(n6464), .B2(n6054), .ZN(n6047)
         );
  AOI22_X1 U6996 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n6056), .B1(n6409), 
        .B2(n6492), .ZN(n6046) );
  OAI211_X1 U6997 ( .C1(n6412), .C2(n6090), .A(n6047), .B(n6046), .ZN(U3023)
         );
  AOI22_X1 U6998 ( .A1(n6471), .A2(n6055), .B1(n6470), .B2(n6054), .ZN(n6049)
         );
  AOI22_X1 U6999 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n6056), .B1(n6413), 
        .B2(n6492), .ZN(n6048) );
  OAI211_X1 U7000 ( .C1(n6416), .C2(n6090), .A(n6049), .B(n6048), .ZN(U3024)
         );
  AOI22_X1 U7001 ( .A1(n6477), .A2(n6055), .B1(n6476), .B2(n6054), .ZN(n6051)
         );
  AOI22_X1 U7002 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n6056), .B1(n6417), 
        .B2(n6492), .ZN(n6050) );
  OAI211_X1 U7003 ( .C1(n6420), .C2(n6090), .A(n6051), .B(n6050), .ZN(U3025)
         );
  AOI22_X1 U7004 ( .A1(n6483), .A2(n6055), .B1(n6482), .B2(n6054), .ZN(n6053)
         );
  AOI22_X1 U7005 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n6056), .B1(n6421), 
        .B2(n6492), .ZN(n6052) );
  OAI211_X1 U7006 ( .C1(n6424), .C2(n6090), .A(n6053), .B(n6052), .ZN(U3026)
         );
  AOI22_X1 U7007 ( .A1(n6491), .A2(n6055), .B1(n6489), .B2(n6054), .ZN(n6058)
         );
  AOI22_X1 U7008 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n6056), .B1(n6428), 
        .B2(n6492), .ZN(n6057) );
  OAI211_X1 U7009 ( .C1(n6432), .C2(n6090), .A(n6058), .B(n6057), .ZN(U3027)
         );
  NOR2_X1 U7010 ( .A1(n6619), .A2(n6066), .ZN(n6061) );
  INV_X1 U7011 ( .A(n6061), .ZN(n6089) );
  OAI22_X1 U7012 ( .A1(n6123), .A2(n6400), .B1(n6234), .B2(n6089), .ZN(n6059)
         );
  INV_X1 U7013 ( .A(n6059), .ZN(n6070) );
  INV_X1 U7014 ( .A(n6060), .ZN(n6062) );
  AOI21_X1 U7015 ( .B1(n6062), .B2(n6614), .A(n6061), .ZN(n6067) );
  AOI21_X1 U7016 ( .B1(n6063), .B2(STATEBS16_REG_SCAN_IN), .A(n6438), .ZN(
        n6065) );
  AOI22_X1 U7017 ( .A1(n6067), .A2(n6065), .B1(n6438), .B2(n6066), .ZN(n6064)
         );
  NAND2_X1 U7018 ( .A1(n6446), .A2(n6064), .ZN(n6093) );
  INV_X1 U7019 ( .A(n6065), .ZN(n6068) );
  OAI22_X1 U7020 ( .A1(n6068), .A2(n6067), .B1(n6436), .B2(n6066), .ZN(n6092)
         );
  AOI22_X1 U7021 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6093), .B1(n6439), 
        .B2(n6092), .ZN(n6069) );
  OAI211_X1 U7022 ( .C1(n6451), .C2(n6090), .A(n6070), .B(n6069), .ZN(U3028)
         );
  INV_X1 U7023 ( .A(n6453), .ZN(n6249) );
  OAI22_X1 U7024 ( .A1(n6090), .A2(n6457), .B1(n6249), .B2(n6089), .ZN(n6071)
         );
  INV_X1 U7025 ( .A(n6071), .ZN(n6073) );
  AOI22_X1 U7026 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6093), .B1(n6452), 
        .B2(n6092), .ZN(n6072) );
  OAI211_X1 U7027 ( .C1(n6123), .C2(n6404), .A(n6073), .B(n6072), .ZN(U3029)
         );
  OAI22_X1 U7028 ( .A1(n6123), .A2(n6408), .B1(n6253), .B2(n6089), .ZN(n6074)
         );
  INV_X1 U7029 ( .A(n6074), .ZN(n6076) );
  AOI22_X1 U7030 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6093), .B1(n6458), 
        .B2(n6092), .ZN(n6075) );
  OAI211_X1 U7031 ( .C1(n6463), .C2(n6090), .A(n6076), .B(n6075), .ZN(U3030)
         );
  INV_X1 U7032 ( .A(n6465), .ZN(n6257) );
  OAI22_X1 U7033 ( .A1(n6123), .A2(n6412), .B1(n6257), .B2(n6089), .ZN(n6077)
         );
  INV_X1 U7034 ( .A(n6077), .ZN(n6079) );
  AOI22_X1 U7035 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6093), .B1(n6464), 
        .B2(n6092), .ZN(n6078) );
  OAI211_X1 U7036 ( .C1(n6469), .C2(n6090), .A(n6079), .B(n6078), .ZN(U3031)
         );
  INV_X1 U7037 ( .A(n6471), .ZN(n6261) );
  OAI22_X1 U7038 ( .A1(n6123), .A2(n6416), .B1(n6261), .B2(n6089), .ZN(n6080)
         );
  INV_X1 U7039 ( .A(n6080), .ZN(n6082) );
  AOI22_X1 U7040 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6093), .B1(n6470), 
        .B2(n6092), .ZN(n6081) );
  OAI211_X1 U7041 ( .C1(n6475), .C2(n6090), .A(n6082), .B(n6081), .ZN(U3032)
         );
  INV_X1 U7042 ( .A(n6477), .ZN(n6265) );
  OAI22_X1 U7043 ( .A1(n6090), .A2(n6481), .B1(n6265), .B2(n6089), .ZN(n6083)
         );
  INV_X1 U7044 ( .A(n6083), .ZN(n6085) );
  AOI22_X1 U7045 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6093), .B1(n6476), 
        .B2(n6092), .ZN(n6084) );
  OAI211_X1 U7046 ( .C1(n6123), .C2(n6420), .A(n6085), .B(n6084), .ZN(U3033)
         );
  INV_X1 U7047 ( .A(n6483), .ZN(n6269) );
  OAI22_X1 U7048 ( .A1(n6123), .A2(n6424), .B1(n6269), .B2(n6089), .ZN(n6086)
         );
  INV_X1 U7049 ( .A(n6086), .ZN(n6088) );
  AOI22_X1 U7050 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6093), .B1(n6482), 
        .B2(n6092), .ZN(n6087) );
  OAI211_X1 U7051 ( .C1(n6487), .C2(n6090), .A(n6088), .B(n6087), .ZN(U3034)
         );
  OAI22_X1 U7052 ( .A1(n6090), .A2(n6498), .B1(n6274), .B2(n6089), .ZN(n6091)
         );
  INV_X1 U7053 ( .A(n6091), .ZN(n6095) );
  AOI22_X1 U7054 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6093), .B1(n6489), 
        .B2(n6092), .ZN(n6094) );
  OAI211_X1 U7055 ( .C1(n6123), .C2(n6432), .A(n6095), .B(n6094), .ZN(U3035)
         );
  NOR2_X1 U7056 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6096), .ZN(n6118)
         );
  NAND3_X1 U7057 ( .A1(n6287), .A2(n6385), .A3(n6525), .ZN(n6097) );
  OAI21_X1 U7058 ( .B1(n6099), .B2(n6438), .A(n6097), .ZN(n6117) );
  AOI22_X1 U7059 ( .A1(n6440), .A2(n6118), .B1(n6439), .B2(n6117), .ZN(n6104)
         );
  INV_X1 U7060 ( .A(n6123), .ZN(n6098) );
  OAI21_X1 U7061 ( .B1(n6119), .B2(n6098), .A(n6162), .ZN(n6100) );
  NAND2_X1 U7062 ( .A1(n6100), .A2(n6099), .ZN(n6102) );
  OAI21_X1 U7063 ( .B1(n6385), .B2(n6436), .A(n6101), .ZN(n6165) );
  NOR2_X1 U7064 ( .A1(n6386), .A2(n6165), .ZN(n6285) );
  AOI22_X1 U7065 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n6120), .B1(n6448), 
        .B2(n6119), .ZN(n6103) );
  OAI211_X1 U7066 ( .C1(n6451), .C2(n6123), .A(n6104), .B(n6103), .ZN(U3036)
         );
  AOI22_X1 U7067 ( .A1(n6453), .A2(n6118), .B1(n6452), .B2(n6117), .ZN(n6106)
         );
  AOI22_X1 U7068 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6454), .ZN(n6105) );
  OAI211_X1 U7069 ( .C1(n6123), .C2(n6457), .A(n6106), .B(n6105), .ZN(U3037)
         );
  AOI22_X1 U7070 ( .A1(n6459), .A2(n6118), .B1(n6458), .B2(n6117), .ZN(n6108)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6460), .ZN(n6107) );
  OAI211_X1 U7072 ( .C1(n6123), .C2(n6463), .A(n6108), .B(n6107), .ZN(U3038)
         );
  AOI22_X1 U7073 ( .A1(n6465), .A2(n6118), .B1(n6464), .B2(n6117), .ZN(n6110)
         );
  AOI22_X1 U7074 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6466), .ZN(n6109) );
  OAI211_X1 U7075 ( .C1(n6123), .C2(n6469), .A(n6110), .B(n6109), .ZN(U3039)
         );
  AOI22_X1 U7076 ( .A1(n6471), .A2(n6118), .B1(n6470), .B2(n6117), .ZN(n6112)
         );
  AOI22_X1 U7077 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6472), .ZN(n6111) );
  OAI211_X1 U7078 ( .C1(n6123), .C2(n6475), .A(n6112), .B(n6111), .ZN(U3040)
         );
  AOI22_X1 U7079 ( .A1(n6477), .A2(n6118), .B1(n6476), .B2(n6117), .ZN(n6114)
         );
  AOI22_X1 U7080 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6478), .ZN(n6113) );
  OAI211_X1 U7081 ( .C1(n6123), .C2(n6481), .A(n6114), .B(n6113), .ZN(U3041)
         );
  AOI22_X1 U7082 ( .A1(n6483), .A2(n6118), .B1(n6482), .B2(n6117), .ZN(n6116)
         );
  AOI22_X1 U7083 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6484), .ZN(n6115) );
  OAI211_X1 U7084 ( .C1(n6123), .C2(n6487), .A(n6116), .B(n6115), .ZN(U3042)
         );
  AOI22_X1 U7085 ( .A1(n6491), .A2(n6118), .B1(n6489), .B2(n6117), .ZN(n6122)
         );
  AOI22_X1 U7086 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n6120), .B1(n6119), 
        .B2(n6493), .ZN(n6121) );
  OAI211_X1 U7087 ( .C1(n6123), .C2(n6498), .A(n6122), .B(n6121), .ZN(U3043)
         );
  NOR2_X2 U7088 ( .A1(n6124), .A2(n6361), .ZN(n6183) );
  NOR2_X1 U7089 ( .A1(n6619), .A2(n6132), .ZN(n6149) );
  AOI22_X1 U7090 ( .A1(n6183), .A2(n6448), .B1(n6440), .B2(n6149), .ZN(n6136)
         );
  OR2_X1 U7091 ( .A1(n6126), .A2(n6125), .ZN(n6128) );
  INV_X1 U7092 ( .A(n6149), .ZN(n6127) );
  AND2_X1 U7093 ( .A1(n6128), .A2(n6127), .ZN(n6134) );
  INV_X1 U7094 ( .A(n6134), .ZN(n6131) );
  AOI21_X1 U7095 ( .B1(n6438), .B2(n6132), .A(n6129), .ZN(n6130) );
  OAI21_X1 U7096 ( .B1(n6133), .B2(n6131), .A(n6130), .ZN(n6151) );
  OAI22_X1 U7097 ( .A1(n6134), .A2(n6133), .B1(n6436), .B2(n6132), .ZN(n6150)
         );
  AOI22_X1 U7098 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6151), .B1(n6439), 
        .B2(n6150), .ZN(n6135) );
  OAI211_X1 U7099 ( .C1(n6451), .C2(n6154), .A(n6136), .B(n6135), .ZN(U3060)
         );
  AOI22_X1 U7100 ( .A1(n6183), .A2(n6454), .B1(n6453), .B2(n6149), .ZN(n6138)
         );
  AOI22_X1 U7101 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6151), .B1(n6452), 
        .B2(n6150), .ZN(n6137) );
  OAI211_X1 U7102 ( .C1(n6457), .C2(n6154), .A(n6138), .B(n6137), .ZN(U3061)
         );
  AOI22_X1 U7103 ( .A1(n6183), .A2(n6460), .B1(n6459), .B2(n6149), .ZN(n6140)
         );
  AOI22_X1 U7104 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6151), .B1(n6458), 
        .B2(n6150), .ZN(n6139) );
  OAI211_X1 U7105 ( .C1(n6463), .C2(n6154), .A(n6140), .B(n6139), .ZN(U3062)
         );
  AOI22_X1 U7106 ( .A1(n6183), .A2(n6466), .B1(n6465), .B2(n6149), .ZN(n6142)
         );
  AOI22_X1 U7107 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6151), .B1(n6464), 
        .B2(n6150), .ZN(n6141) );
  OAI211_X1 U7108 ( .C1(n6469), .C2(n6154), .A(n6142), .B(n6141), .ZN(U3063)
         );
  AOI22_X1 U7109 ( .A1(n6183), .A2(n6472), .B1(n6471), .B2(n6149), .ZN(n6144)
         );
  AOI22_X1 U7110 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6151), .B1(n6470), 
        .B2(n6150), .ZN(n6143) );
  OAI211_X1 U7111 ( .C1(n6475), .C2(n6154), .A(n6144), .B(n6143), .ZN(U3064)
         );
  AOI22_X1 U7112 ( .A1(n6183), .A2(n6478), .B1(n6477), .B2(n6149), .ZN(n6146)
         );
  AOI22_X1 U7113 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6151), .B1(n6476), 
        .B2(n6150), .ZN(n6145) );
  OAI211_X1 U7114 ( .C1(n6481), .C2(n6154), .A(n6146), .B(n6145), .ZN(U3065)
         );
  AOI22_X1 U7115 ( .A1(n6183), .A2(n6484), .B1(n6483), .B2(n6149), .ZN(n6148)
         );
  AOI22_X1 U7116 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6151), .B1(n6482), 
        .B2(n6150), .ZN(n6147) );
  OAI211_X1 U7117 ( .C1(n6487), .C2(n6154), .A(n6148), .B(n6147), .ZN(U3066)
         );
  AOI22_X1 U7118 ( .A1(n6183), .A2(n6493), .B1(n6491), .B2(n6149), .ZN(n6153)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6151), .B1(n6489), 
        .B2(n6150), .ZN(n6152) );
  OAI211_X1 U7120 ( .C1(n6498), .C2(n6154), .A(n6153), .B(n6152), .ZN(U3067)
         );
  INV_X1 U7121 ( .A(n6434), .ZN(n6389) );
  INV_X1 U7122 ( .A(n6385), .ZN(n6158) );
  NOR2_X1 U7123 ( .A1(n6436), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6393)
         );
  INV_X1 U7124 ( .A(n6393), .ZN(n6157) );
  INV_X1 U7125 ( .A(n6155), .ZN(n6156) );
  OAI33_X1 U7126 ( .A1(n6392), .A2(n6389), .A3(n6438), .B1(n6158), .B2(n6157), 
        .B3(n6156), .ZN(n6182) );
  NOR2_X1 U7127 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6159), .ZN(n6181)
         );
  AOI22_X1 U7128 ( .A1(n3165), .A2(n6439), .B1(n6440), .B2(n6181), .ZN(n6168)
         );
  INV_X1 U7129 ( .A(n6181), .ZN(n6164) );
  INV_X1 U7130 ( .A(n6183), .ZN(n6160) );
  NAND3_X1 U7131 ( .A1(n6160), .A2(n6612), .A3(n6201), .ZN(n6161) );
  AOI21_X1 U7132 ( .B1(n6162), .B2(n6161), .A(n6434), .ZN(n6163) );
  AOI21_X1 U7133 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6164), .A(n6163), .ZN(
        n6166) );
  NOR2_X1 U7134 ( .A1(n6287), .A2(n6165), .ZN(n6396) );
  NAND3_X1 U7135 ( .A1(n6525), .A2(n6166), .A3(n6396), .ZN(n6184) );
  AOI22_X1 U7136 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n6184), .B1(n6397), 
        .B2(n6183), .ZN(n6167) );
  OAI211_X1 U7137 ( .C1(n6400), .C2(n6201), .A(n6168), .B(n6167), .ZN(U3068)
         );
  AOI22_X1 U7138 ( .A1(n3165), .A2(n6452), .B1(n6453), .B2(n6181), .ZN(n6170)
         );
  AOI22_X1 U7139 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6184), .B1(n6401), 
        .B2(n6183), .ZN(n6169) );
  OAI211_X1 U7140 ( .C1(n6404), .C2(n6201), .A(n6170), .B(n6169), .ZN(U3069)
         );
  AOI22_X1 U7141 ( .A1(n3165), .A2(n6458), .B1(n6459), .B2(n6181), .ZN(n6172)
         );
  AOI22_X1 U7142 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n6184), .B1(n6405), 
        .B2(n6183), .ZN(n6171) );
  OAI211_X1 U7143 ( .C1(n6408), .C2(n6201), .A(n6172), .B(n6171), .ZN(U3070)
         );
  AOI22_X1 U7144 ( .A1(n3165), .A2(n6464), .B1(n6465), .B2(n6181), .ZN(n6174)
         );
  AOI22_X1 U7145 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n6184), .B1(n6409), 
        .B2(n6183), .ZN(n6173) );
  OAI211_X1 U7146 ( .C1(n6412), .C2(n6201), .A(n6174), .B(n6173), .ZN(U3071)
         );
  AOI22_X1 U7147 ( .A1(n3165), .A2(n6470), .B1(n6471), .B2(n6181), .ZN(n6176)
         );
  AOI22_X1 U7148 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n6184), .B1(n6413), 
        .B2(n6183), .ZN(n6175) );
  OAI211_X1 U7149 ( .C1(n6416), .C2(n6201), .A(n6176), .B(n6175), .ZN(U3072)
         );
  AOI22_X1 U7150 ( .A1(n3165), .A2(n6476), .B1(n6477), .B2(n6181), .ZN(n6178)
         );
  AOI22_X1 U7151 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n6184), .B1(n6417), 
        .B2(n6183), .ZN(n6177) );
  OAI211_X1 U7152 ( .C1(n6420), .C2(n6201), .A(n6178), .B(n6177), .ZN(U3073)
         );
  AOI22_X1 U7153 ( .A1(n3165), .A2(n6482), .B1(n6483), .B2(n6181), .ZN(n6180)
         );
  AOI22_X1 U7154 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6184), .B1(n6421), 
        .B2(n6183), .ZN(n6179) );
  OAI211_X1 U7155 ( .C1(n6424), .C2(n6201), .A(n6180), .B(n6179), .ZN(U3074)
         );
  AOI22_X1 U7156 ( .A1(n3165), .A2(n6489), .B1(n6491), .B2(n6181), .ZN(n6186)
         );
  AOI22_X1 U7157 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n6184), .B1(n6428), 
        .B2(n6183), .ZN(n6185) );
  OAI211_X1 U7158 ( .C1(n6432), .C2(n6201), .A(n6186), .B(n6185), .ZN(U3075)
         );
  INV_X1 U7159 ( .A(n6187), .ZN(n6196) );
  AOI22_X1 U7160 ( .A1(n6229), .A2(n6454), .B1(n6196), .B2(n6453), .ZN(n6189)
         );
  AOI22_X1 U7161 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6198), .B1(n6452), 
        .B2(n6197), .ZN(n6188) );
  OAI211_X1 U7162 ( .C1(n6457), .C2(n6201), .A(n6189), .B(n6188), .ZN(U3077)
         );
  AOI22_X1 U7163 ( .A1(n6229), .A2(n6466), .B1(n6196), .B2(n6465), .ZN(n6191)
         );
  AOI22_X1 U7164 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6198), .B1(n6464), 
        .B2(n6197), .ZN(n6190) );
  OAI211_X1 U7165 ( .C1(n6469), .C2(n6201), .A(n6191), .B(n6190), .ZN(U3079)
         );
  AOI22_X1 U7166 ( .A1(n6229), .A2(n6472), .B1(n6196), .B2(n6471), .ZN(n6193)
         );
  AOI22_X1 U7167 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6198), .B1(n6470), 
        .B2(n6197), .ZN(n6192) );
  OAI211_X1 U7168 ( .C1(n6475), .C2(n6201), .A(n6193), .B(n6192), .ZN(U3080)
         );
  AOI22_X1 U7169 ( .A1(n6229), .A2(n6478), .B1(n6196), .B2(n6477), .ZN(n6195)
         );
  AOI22_X1 U7170 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6198), .B1(n6476), 
        .B2(n6197), .ZN(n6194) );
  OAI211_X1 U7171 ( .C1(n6481), .C2(n6201), .A(n6195), .B(n6194), .ZN(U3081)
         );
  AOI22_X1 U7172 ( .A1(n6229), .A2(n6484), .B1(n6196), .B2(n6483), .ZN(n6200)
         );
  AOI22_X1 U7173 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6198), .B1(n6482), 
        .B2(n6197), .ZN(n6199) );
  OAI211_X1 U7174 ( .C1(n6487), .C2(n6201), .A(n6200), .B(n6199), .ZN(U3082)
         );
  NAND3_X1 U7175 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6517), .A3(n6512), .ZN(n6244) );
  NOR2_X1 U7176 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6244), .ZN(n6228)
         );
  NAND2_X1 U7177 ( .A1(n6392), .A2(n6612), .ZN(n6388) );
  INV_X1 U7178 ( .A(n6203), .ZN(n6204) );
  OR2_X1 U7179 ( .A1(n6204), .A2(n6385), .ZN(n6322) );
  OAI22_X1 U7180 ( .A1(n6388), .A2(n6206), .B1(n6330), .B2(n6322), .ZN(n6227)
         );
  AOI22_X1 U7181 ( .A1(n6440), .A2(n6228), .B1(n6439), .B2(n6227), .ZN(n6214)
         );
  AOI21_X1 U7182 ( .B1(n6280), .B2(n6205), .A(n6793), .ZN(n6212) );
  OAI21_X1 U7183 ( .B1(n6207), .B2(n6206), .A(n6612), .ZN(n6211) );
  AOI21_X1 U7184 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6322), .A(n6208), .ZN(
        n6331) );
  INV_X1 U7185 ( .A(n6228), .ZN(n6209) );
  AOI21_X1 U7186 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6209), .A(n6386), .ZN(
        n6210) );
  OAI211_X1 U7187 ( .C1(n6212), .C2(n6211), .A(n6331), .B(n6210), .ZN(n6230)
         );
  AOI22_X1 U7188 ( .A1(n6230), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6397), 
        .B2(n6229), .ZN(n6213) );
  OAI211_X1 U7189 ( .C1(n6400), .C2(n6280), .A(n6214), .B(n6213), .ZN(U3084)
         );
  AOI22_X1 U7190 ( .A1(n6453), .A2(n6228), .B1(n6452), .B2(n6227), .ZN(n6216)
         );
  AOI22_X1 U7191 ( .A1(n6230), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6401), 
        .B2(n6229), .ZN(n6215) );
  OAI211_X1 U7192 ( .C1(n6404), .C2(n6280), .A(n6216), .B(n6215), .ZN(U3085)
         );
  AOI22_X1 U7193 ( .A1(n6459), .A2(n6228), .B1(n6458), .B2(n6227), .ZN(n6218)
         );
  AOI22_X1 U7194 ( .A1(n6230), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6405), 
        .B2(n6229), .ZN(n6217) );
  OAI211_X1 U7195 ( .C1(n6408), .C2(n6280), .A(n6218), .B(n6217), .ZN(U3086)
         );
  AOI22_X1 U7196 ( .A1(n6465), .A2(n6228), .B1(n6464), .B2(n6227), .ZN(n6220)
         );
  AOI22_X1 U7197 ( .A1(n6230), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6409), 
        .B2(n6229), .ZN(n6219) );
  OAI211_X1 U7198 ( .C1(n6412), .C2(n6280), .A(n6220), .B(n6219), .ZN(U3087)
         );
  AOI22_X1 U7199 ( .A1(n6471), .A2(n6228), .B1(n6470), .B2(n6227), .ZN(n6222)
         );
  AOI22_X1 U7200 ( .A1(n6230), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6413), 
        .B2(n6229), .ZN(n6221) );
  OAI211_X1 U7201 ( .C1(n6416), .C2(n6280), .A(n6222), .B(n6221), .ZN(U3088)
         );
  AOI22_X1 U7202 ( .A1(n6477), .A2(n6228), .B1(n6476), .B2(n6227), .ZN(n6224)
         );
  AOI22_X1 U7203 ( .A1(n6230), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6417), 
        .B2(n6229), .ZN(n6223) );
  OAI211_X1 U7204 ( .C1(n6420), .C2(n6280), .A(n6224), .B(n6223), .ZN(U3089)
         );
  AOI22_X1 U7205 ( .A1(n6483), .A2(n6228), .B1(n6482), .B2(n6227), .ZN(n6226)
         );
  AOI22_X1 U7206 ( .A1(n6230), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6421), 
        .B2(n6229), .ZN(n6225) );
  OAI211_X1 U7207 ( .C1(n6424), .C2(n6280), .A(n6226), .B(n6225), .ZN(U3090)
         );
  AOI22_X1 U7208 ( .A1(n6491), .A2(n6228), .B1(n6489), .B2(n6227), .ZN(n6232)
         );
  AOI22_X1 U7209 ( .A1(n6230), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6428), 
        .B2(n6229), .ZN(n6231) );
  OAI211_X1 U7210 ( .C1(n6432), .C2(n6280), .A(n6232), .B(n6231), .ZN(U3091)
         );
  NOR2_X1 U7211 ( .A1(n6619), .A2(n6244), .ZN(n6236) );
  INV_X1 U7212 ( .A(n6236), .ZN(n6273) );
  OAI22_X1 U7213 ( .A1(n6280), .A2(n6451), .B1(n6234), .B2(n6273), .ZN(n6235)
         );
  INV_X1 U7214 ( .A(n6235), .ZN(n6248) );
  AND2_X1 U7215 ( .A1(n6392), .A2(n6614), .ZN(n6435) );
  AOI21_X1 U7216 ( .B1(n6435), .B2(n6237), .A(n6236), .ZN(n6246) );
  NAND2_X1 U7217 ( .A1(n6238), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6239) );
  OR2_X1 U7218 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  AND2_X1 U7219 ( .A1(n6241), .A2(n6612), .ZN(n6243) );
  AOI22_X1 U7220 ( .A1(n6246), .A2(n6243), .B1(n6438), .B2(n6244), .ZN(n6242)
         );
  NAND2_X1 U7221 ( .A1(n6446), .A2(n6242), .ZN(n6277) );
  INV_X1 U7222 ( .A(n6243), .ZN(n6245) );
  OAI22_X1 U7223 ( .A1(n6246), .A2(n6245), .B1(n6436), .B2(n6244), .ZN(n6276)
         );
  AOI22_X1 U7224 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6277), .B1(n6439), 
        .B2(n6276), .ZN(n6247) );
  OAI211_X1 U7225 ( .C1(n6400), .C2(n6311), .A(n6248), .B(n6247), .ZN(U3092)
         );
  OAI22_X1 U7226 ( .A1(n6311), .A2(n6404), .B1(n6249), .B2(n6273), .ZN(n6250)
         );
  INV_X1 U7227 ( .A(n6250), .ZN(n6252) );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6277), .B1(n6452), 
        .B2(n6276), .ZN(n6251) );
  OAI211_X1 U7229 ( .C1(n6457), .C2(n6280), .A(n6252), .B(n6251), .ZN(U3093)
         );
  OAI22_X1 U7230 ( .A1(n6311), .A2(n6408), .B1(n6253), .B2(n6273), .ZN(n6254)
         );
  INV_X1 U7231 ( .A(n6254), .ZN(n6256) );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6277), .B1(n6458), 
        .B2(n6276), .ZN(n6255) );
  OAI211_X1 U7233 ( .C1(n6463), .C2(n6280), .A(n6256), .B(n6255), .ZN(U3094)
         );
  OAI22_X1 U7234 ( .A1(n6311), .A2(n6412), .B1(n6257), .B2(n6273), .ZN(n6258)
         );
  INV_X1 U7235 ( .A(n6258), .ZN(n6260) );
  AOI22_X1 U7236 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6277), .B1(n6464), 
        .B2(n6276), .ZN(n6259) );
  OAI211_X1 U7237 ( .C1(n6469), .C2(n6280), .A(n6260), .B(n6259), .ZN(U3095)
         );
  OAI22_X1 U7238 ( .A1(n6280), .A2(n6475), .B1(n6261), .B2(n6273), .ZN(n6262)
         );
  INV_X1 U7239 ( .A(n6262), .ZN(n6264) );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6277), .B1(n6470), 
        .B2(n6276), .ZN(n6263) );
  OAI211_X1 U7241 ( .C1(n6416), .C2(n6311), .A(n6264), .B(n6263), .ZN(U3096)
         );
  OAI22_X1 U7242 ( .A1(n6311), .A2(n6420), .B1(n6265), .B2(n6273), .ZN(n6266)
         );
  INV_X1 U7243 ( .A(n6266), .ZN(n6268) );
  AOI22_X1 U7244 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6277), .B1(n6476), 
        .B2(n6276), .ZN(n6267) );
  OAI211_X1 U7245 ( .C1(n6481), .C2(n6280), .A(n6268), .B(n6267), .ZN(U3097)
         );
  OAI22_X1 U7246 ( .A1(n6311), .A2(n6424), .B1(n6269), .B2(n6273), .ZN(n6270)
         );
  INV_X1 U7247 ( .A(n6270), .ZN(n6272) );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6277), .B1(n6482), 
        .B2(n6276), .ZN(n6271) );
  OAI211_X1 U7249 ( .C1(n6487), .C2(n6280), .A(n6272), .B(n6271), .ZN(U3098)
         );
  OAI22_X1 U7250 ( .A1(n6311), .A2(n6432), .B1(n6274), .B2(n6273), .ZN(n6275)
         );
  INV_X1 U7251 ( .A(n6275), .ZN(n6279) );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6277), .B1(n6489), 
        .B2(n6276), .ZN(n6278) );
  OAI211_X1 U7253 ( .C1(n6498), .C2(n6280), .A(n6279), .B(n6278), .ZN(U3099)
         );
  NOR2_X1 U7254 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6281), .ZN(n6305)
         );
  AOI22_X1 U7255 ( .A1(n6306), .A2(n6448), .B1(n6440), .B2(n6305), .ZN(n6292)
         );
  NAND2_X1 U7256 ( .A1(n6311), .A2(n6321), .ZN(n6282) );
  AOI21_X1 U7257 ( .B1(n6282), .B2(STATEBS16_REG_SCAN_IN), .A(n6438), .ZN(
        n6286) );
  NOR2_X1 U7258 ( .A1(n6305), .A2(n6609), .ZN(n6283) );
  AOI21_X1 U7259 ( .B1(n6286), .B2(n6289), .A(n6283), .ZN(n6284) );
  OAI211_X1 U7260 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6436), .A(n6285), .B(n6284), .ZN(n6308) );
  INV_X1 U7261 ( .A(n6286), .ZN(n6290) );
  NAND3_X1 U7262 ( .A1(n6287), .A2(n6385), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6288) );
  AOI22_X1 U7263 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6308), .B1(n6439), 
        .B2(n6307), .ZN(n6291) );
  OAI211_X1 U7264 ( .C1(n6451), .C2(n6311), .A(n6292), .B(n6291), .ZN(U3100)
         );
  AOI22_X1 U7265 ( .A1(n6306), .A2(n6454), .B1(n6453), .B2(n6305), .ZN(n6294)
         );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6308), .B1(n6452), 
        .B2(n6307), .ZN(n6293) );
  OAI211_X1 U7267 ( .C1(n6457), .C2(n6311), .A(n6294), .B(n6293), .ZN(U3101)
         );
  AOI22_X1 U7268 ( .A1(n6306), .A2(n6460), .B1(n6459), .B2(n6305), .ZN(n6296)
         );
  AOI22_X1 U7269 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6308), .B1(n6458), 
        .B2(n6307), .ZN(n6295) );
  OAI211_X1 U7270 ( .C1(n6463), .C2(n6311), .A(n6296), .B(n6295), .ZN(U3102)
         );
  AOI22_X1 U7271 ( .A1(n6306), .A2(n6466), .B1(n6465), .B2(n6305), .ZN(n6298)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6308), .B1(n6464), 
        .B2(n6307), .ZN(n6297) );
  OAI211_X1 U7273 ( .C1(n6469), .C2(n6311), .A(n6298), .B(n6297), .ZN(U3103)
         );
  AOI22_X1 U7274 ( .A1(n6306), .A2(n6472), .B1(n6471), .B2(n6305), .ZN(n6300)
         );
  AOI22_X1 U7275 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6308), .B1(n6470), 
        .B2(n6307), .ZN(n6299) );
  OAI211_X1 U7276 ( .C1(n6475), .C2(n6311), .A(n6300), .B(n6299), .ZN(U3104)
         );
  AOI22_X1 U7277 ( .A1(n6306), .A2(n6478), .B1(n6477), .B2(n6305), .ZN(n6302)
         );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6308), .B1(n6476), 
        .B2(n6307), .ZN(n6301) );
  OAI211_X1 U7279 ( .C1(n6481), .C2(n6311), .A(n6302), .B(n6301), .ZN(U3105)
         );
  AOI22_X1 U7280 ( .A1(n6306), .A2(n6484), .B1(n6483), .B2(n6305), .ZN(n6304)
         );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6308), .B1(n6482), 
        .B2(n6307), .ZN(n6303) );
  OAI211_X1 U7282 ( .C1(n6487), .C2(n6311), .A(n6304), .B(n6303), .ZN(U3106)
         );
  AOI22_X1 U7283 ( .A1(n6306), .A2(n6493), .B1(n6491), .B2(n6305), .ZN(n6310)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6308), .B1(n6489), 
        .B2(n6307), .ZN(n6309) );
  OAI211_X1 U7285 ( .C1(n6498), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3107)
         );
  AOI22_X1 U7286 ( .A1(n6349), .A2(n6472), .B1(n6471), .B2(n6316), .ZN(n6313)
         );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6318), .B1(n6470), 
        .B2(n6317), .ZN(n6312) );
  OAI211_X1 U7288 ( .C1(n6475), .C2(n6321), .A(n6313), .B(n6312), .ZN(U3112)
         );
  AOI22_X1 U7289 ( .A1(n6349), .A2(n6478), .B1(n6477), .B2(n6316), .ZN(n6315)
         );
  AOI22_X1 U7290 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6318), .B1(n6476), 
        .B2(n6317), .ZN(n6314) );
  OAI211_X1 U7291 ( .C1(n6481), .C2(n6321), .A(n6315), .B(n6314), .ZN(U3113)
         );
  AOI22_X1 U7292 ( .A1(n6349), .A2(n6484), .B1(n6483), .B2(n6316), .ZN(n6320)
         );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6318), .B1(n6482), 
        .B2(n6317), .ZN(n6319) );
  OAI211_X1 U7294 ( .C1(n6487), .C2(n6321), .A(n6320), .B(n6319), .ZN(U3114)
         );
  NOR2_X1 U7295 ( .A1(n6525), .A2(n6354), .ZN(n6359) );
  NAND2_X1 U7296 ( .A1(n6619), .A2(n6359), .ZN(n6328) );
  INV_X1 U7297 ( .A(n6328), .ZN(n6348) );
  INV_X1 U7298 ( .A(n6353), .ZN(n6326) );
  INV_X1 U7299 ( .A(n6386), .ZN(n6323) );
  OAI22_X1 U7300 ( .A1(n6326), .A2(n6388), .B1(n6323), .B2(n6322), .ZN(n6347)
         );
  AOI22_X1 U7301 ( .A1(n6440), .A2(n6348), .B1(n6439), .B2(n6347), .ZN(n6334)
         );
  INV_X1 U7302 ( .A(n6382), .ZN(n6324) );
  OAI21_X1 U7303 ( .B1(n6324), .B2(n6349), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6325) );
  OAI211_X1 U7304 ( .C1(n6327), .C2(n6326), .A(n6325), .B(n6612), .ZN(n6332)
         );
  NAND2_X1 U7305 ( .A1(n6328), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6329) );
  NAND4_X1 U7306 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n6350)
         );
  AOI22_X1 U7307 ( .A1(n6350), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6397), 
        .B2(n6349), .ZN(n6333) );
  OAI211_X1 U7308 ( .C1(n6400), .C2(n6382), .A(n6334), .B(n6333), .ZN(U3116)
         );
  AOI22_X1 U7309 ( .A1(n6453), .A2(n6348), .B1(n6452), .B2(n6347), .ZN(n6336)
         );
  AOI22_X1 U7310 ( .A1(n6350), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6401), 
        .B2(n6349), .ZN(n6335) );
  OAI211_X1 U7311 ( .C1(n6404), .C2(n6382), .A(n6336), .B(n6335), .ZN(U3117)
         );
  AOI22_X1 U7312 ( .A1(n6459), .A2(n6348), .B1(n6458), .B2(n6347), .ZN(n6338)
         );
  AOI22_X1 U7313 ( .A1(n6350), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6405), 
        .B2(n6349), .ZN(n6337) );
  OAI211_X1 U7314 ( .C1(n6408), .C2(n6382), .A(n6338), .B(n6337), .ZN(U3118)
         );
  AOI22_X1 U7315 ( .A1(n6465), .A2(n6348), .B1(n6464), .B2(n6347), .ZN(n6340)
         );
  AOI22_X1 U7316 ( .A1(n6350), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6409), 
        .B2(n6349), .ZN(n6339) );
  OAI211_X1 U7317 ( .C1(n6412), .C2(n6382), .A(n6340), .B(n6339), .ZN(U3119)
         );
  AOI22_X1 U7318 ( .A1(n6471), .A2(n6348), .B1(n6470), .B2(n6347), .ZN(n6342)
         );
  AOI22_X1 U7319 ( .A1(n6350), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6413), 
        .B2(n6349), .ZN(n6341) );
  OAI211_X1 U7320 ( .C1(n6416), .C2(n6382), .A(n6342), .B(n6341), .ZN(U3120)
         );
  AOI22_X1 U7321 ( .A1(n6477), .A2(n6348), .B1(n6476), .B2(n6347), .ZN(n6344)
         );
  AOI22_X1 U7322 ( .A1(n6350), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6417), 
        .B2(n6349), .ZN(n6343) );
  OAI211_X1 U7323 ( .C1(n6420), .C2(n6382), .A(n6344), .B(n6343), .ZN(U3121)
         );
  AOI22_X1 U7324 ( .A1(n6483), .A2(n6348), .B1(n6482), .B2(n6347), .ZN(n6346)
         );
  AOI22_X1 U7325 ( .A1(n6350), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6421), 
        .B2(n6349), .ZN(n6345) );
  OAI211_X1 U7326 ( .C1(n6424), .C2(n6382), .A(n6346), .B(n6345), .ZN(U3122)
         );
  AOI22_X1 U7327 ( .A1(n6491), .A2(n6348), .B1(n6489), .B2(n6347), .ZN(n6352)
         );
  AOI22_X1 U7328 ( .A1(n6350), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6428), 
        .B2(n6349), .ZN(n6351) );
  OAI211_X1 U7329 ( .C1(n6432), .C2(n6382), .A(n6352), .B(n6351), .ZN(U3123)
         );
  AND2_X1 U7330 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6359), .ZN(n6378)
         );
  AOI21_X1 U7331 ( .B1(n6435), .B2(n6353), .A(n6378), .ZN(n6357) );
  NAND2_X1 U7332 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6355) );
  OAI22_X1 U7333 ( .A1(n6357), .A2(n6438), .B1(n6355), .B2(n6354), .ZN(n6377)
         );
  AOI22_X1 U7334 ( .A1(n6440), .A2(n6378), .B1(n6439), .B2(n6377), .ZN(n6364)
         );
  NAND2_X1 U7335 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  OAI221_X1 U7336 ( .B1(n6612), .B2(n6359), .C1(n6438), .C2(n6358), .A(n6446), 
        .ZN(n6379) );
  INV_X1 U7337 ( .A(n6360), .ZN(n6362) );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6379), .B1(n6448), 
        .B2(n6427), .ZN(n6363) );
  OAI211_X1 U7339 ( .C1(n6451), .C2(n6382), .A(n6364), .B(n6363), .ZN(U3124)
         );
  AOI22_X1 U7340 ( .A1(n6453), .A2(n6378), .B1(n6452), .B2(n6377), .ZN(n6366)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6379), .B1(n6454), 
        .B2(n6427), .ZN(n6365) );
  OAI211_X1 U7342 ( .C1(n6457), .C2(n6382), .A(n6366), .B(n6365), .ZN(U3125)
         );
  AOI22_X1 U7343 ( .A1(n6459), .A2(n6378), .B1(n6458), .B2(n6377), .ZN(n6368)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6379), .B1(n6460), 
        .B2(n6427), .ZN(n6367) );
  OAI211_X1 U7345 ( .C1(n6463), .C2(n6382), .A(n6368), .B(n6367), .ZN(U3126)
         );
  AOI22_X1 U7346 ( .A1(n6465), .A2(n6378), .B1(n6464), .B2(n6377), .ZN(n6370)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6379), .B1(n6466), 
        .B2(n6427), .ZN(n6369) );
  OAI211_X1 U7348 ( .C1(n6469), .C2(n6382), .A(n6370), .B(n6369), .ZN(U3127)
         );
  AOI22_X1 U7349 ( .A1(n6471), .A2(n6378), .B1(n6470), .B2(n6377), .ZN(n6372)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6379), .B1(n6472), 
        .B2(n6427), .ZN(n6371) );
  OAI211_X1 U7351 ( .C1(n6475), .C2(n6382), .A(n6372), .B(n6371), .ZN(U3128)
         );
  AOI22_X1 U7352 ( .A1(n6477), .A2(n6378), .B1(n6476), .B2(n6377), .ZN(n6374)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6379), .B1(n6478), 
        .B2(n6427), .ZN(n6373) );
  OAI211_X1 U7354 ( .C1(n6481), .C2(n6382), .A(n6374), .B(n6373), .ZN(U3129)
         );
  AOI22_X1 U7355 ( .A1(n6483), .A2(n6378), .B1(n6482), .B2(n6377), .ZN(n6376)
         );
  AOI22_X1 U7356 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6379), .B1(n6484), 
        .B2(n6427), .ZN(n6375) );
  OAI211_X1 U7357 ( .C1(n6487), .C2(n6382), .A(n6376), .B(n6375), .ZN(U3130)
         );
  AOI22_X1 U7358 ( .A1(n6491), .A2(n6378), .B1(n6489), .B2(n6377), .ZN(n6381)
         );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6379), .B1(n6493), 
        .B2(n6427), .ZN(n6380) );
  OAI211_X1 U7360 ( .C1(n6498), .C2(n6382), .A(n6381), .B(n6380), .ZN(U3131)
         );
  NAND2_X1 U7361 ( .A1(n6384), .A2(n6383), .ZN(n6441) );
  NOR2_X1 U7362 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6437), .ZN(n6426)
         );
  NAND3_X1 U7363 ( .A1(n6386), .A2(n6385), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U7364 ( .B1(n6389), .B2(n6388), .A(n6387), .ZN(n6425) );
  AOI22_X1 U7365 ( .A1(n6440), .A2(n6426), .B1(n6439), .B2(n6425), .ZN(n6399)
         );
  INV_X1 U7366 ( .A(n6427), .ZN(n6390) );
  AOI21_X1 U7367 ( .B1(n6390), .B2(n6497), .A(n6793), .ZN(n6391) );
  AOI211_X1 U7368 ( .C1(n6434), .C2(n6392), .A(n6438), .B(n6391), .ZN(n6394)
         );
  NOR2_X1 U7369 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6429), .B1(n6397), 
        .B2(n6427), .ZN(n6398) );
  OAI211_X1 U7371 ( .C1(n6400), .C2(n6497), .A(n6399), .B(n6398), .ZN(U3132)
         );
  AOI22_X1 U7372 ( .A1(n6453), .A2(n6426), .B1(n6452), .B2(n6425), .ZN(n6403)
         );
  AOI22_X1 U7373 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6429), .B1(n6401), 
        .B2(n6427), .ZN(n6402) );
  OAI211_X1 U7374 ( .C1(n6404), .C2(n6497), .A(n6403), .B(n6402), .ZN(U3133)
         );
  AOI22_X1 U7375 ( .A1(n6459), .A2(n6426), .B1(n6458), .B2(n6425), .ZN(n6407)
         );
  AOI22_X1 U7376 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6429), .B1(n6405), 
        .B2(n6427), .ZN(n6406) );
  OAI211_X1 U7377 ( .C1(n6408), .C2(n6497), .A(n6407), .B(n6406), .ZN(U3134)
         );
  AOI22_X1 U7378 ( .A1(n6465), .A2(n6426), .B1(n6464), .B2(n6425), .ZN(n6411)
         );
  AOI22_X1 U7379 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6429), .B1(n6409), 
        .B2(n6427), .ZN(n6410) );
  OAI211_X1 U7380 ( .C1(n6412), .C2(n6497), .A(n6411), .B(n6410), .ZN(U3135)
         );
  AOI22_X1 U7381 ( .A1(n6471), .A2(n6426), .B1(n6470), .B2(n6425), .ZN(n6415)
         );
  AOI22_X1 U7382 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6429), .B1(n6413), 
        .B2(n6427), .ZN(n6414) );
  OAI211_X1 U7383 ( .C1(n6416), .C2(n6497), .A(n6415), .B(n6414), .ZN(U3136)
         );
  AOI22_X1 U7384 ( .A1(n6477), .A2(n6426), .B1(n6476), .B2(n6425), .ZN(n6419)
         );
  AOI22_X1 U7385 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6429), .B1(n6417), 
        .B2(n6427), .ZN(n6418) );
  OAI211_X1 U7386 ( .C1(n6420), .C2(n6497), .A(n6419), .B(n6418), .ZN(U3137)
         );
  AOI22_X1 U7387 ( .A1(n6483), .A2(n6426), .B1(n6482), .B2(n6425), .ZN(n6423)
         );
  AOI22_X1 U7388 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6429), .B1(n6421), 
        .B2(n6427), .ZN(n6422) );
  OAI211_X1 U7389 ( .C1(n6424), .C2(n6497), .A(n6423), .B(n6422), .ZN(U3138)
         );
  AOI22_X1 U7390 ( .A1(n6491), .A2(n6426), .B1(n6489), .B2(n6425), .ZN(n6431)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6427), .ZN(n6430) );
  OAI211_X1 U7392 ( .C1(n6432), .C2(n6497), .A(n6431), .B(n6430), .ZN(U3139)
         );
  INV_X1 U7393 ( .A(n6433), .ZN(n6490) );
  AOI21_X1 U7394 ( .B1(n6435), .B2(n6434), .A(n6490), .ZN(n6442) );
  OAI22_X1 U7395 ( .A1(n6442), .A2(n6438), .B1(n6437), .B2(n6436), .ZN(n6488)
         );
  AOI22_X1 U7396 ( .A1(n6440), .A2(n6490), .B1(n6439), .B2(n6488), .ZN(n6450)
         );
  AND2_X1 U7397 ( .A1(n6441), .A2(n5910), .ZN(n6444) );
  OAI21_X1 U7398 ( .B1(n6444), .B2(n6443), .A(n6442), .ZN(n6445) );
  OAI211_X1 U7399 ( .C1(n6447), .C2(n6612), .A(n6446), .B(n6445), .ZN(n6494)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6494), .B1(n6448), 
        .B2(n6492), .ZN(n6449) );
  OAI211_X1 U7401 ( .C1(n6451), .C2(n6497), .A(n6450), .B(n6449), .ZN(U3140)
         );
  AOI22_X1 U7402 ( .A1(n6453), .A2(n6490), .B1(n6452), .B2(n6488), .ZN(n6456)
         );
  AOI22_X1 U7403 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6494), .B1(n6454), 
        .B2(n6492), .ZN(n6455) );
  OAI211_X1 U7404 ( .C1(n6457), .C2(n6497), .A(n6456), .B(n6455), .ZN(U3141)
         );
  AOI22_X1 U7405 ( .A1(n6459), .A2(n6490), .B1(n6458), .B2(n6488), .ZN(n6462)
         );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6494), .B1(n6460), 
        .B2(n6492), .ZN(n6461) );
  OAI211_X1 U7407 ( .C1(n6463), .C2(n6497), .A(n6462), .B(n6461), .ZN(U3142)
         );
  AOI22_X1 U7408 ( .A1(n6465), .A2(n6490), .B1(n6464), .B2(n6488), .ZN(n6468)
         );
  AOI22_X1 U7409 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6494), .B1(n6466), 
        .B2(n6492), .ZN(n6467) );
  OAI211_X1 U7410 ( .C1(n6469), .C2(n6497), .A(n6468), .B(n6467), .ZN(U3143)
         );
  AOI22_X1 U7411 ( .A1(n6471), .A2(n6490), .B1(n6470), .B2(n6488), .ZN(n6474)
         );
  AOI22_X1 U7412 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6494), .B1(n6472), 
        .B2(n6492), .ZN(n6473) );
  OAI211_X1 U7413 ( .C1(n6475), .C2(n6497), .A(n6474), .B(n6473), .ZN(U3144)
         );
  AOI22_X1 U7414 ( .A1(n6477), .A2(n6490), .B1(n6476), .B2(n6488), .ZN(n6480)
         );
  AOI22_X1 U7415 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6494), .B1(n6478), 
        .B2(n6492), .ZN(n6479) );
  OAI211_X1 U7416 ( .C1(n6481), .C2(n6497), .A(n6480), .B(n6479), .ZN(U3145)
         );
  AOI22_X1 U7417 ( .A1(n6483), .A2(n6490), .B1(n6482), .B2(n6488), .ZN(n6486)
         );
  AOI22_X1 U7418 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6494), .B1(n6484), 
        .B2(n6492), .ZN(n6485) );
  OAI211_X1 U7419 ( .C1(n6487), .C2(n6497), .A(n6486), .B(n6485), .ZN(U3146)
         );
  AOI22_X1 U7420 ( .A1(n6491), .A2(n6490), .B1(n6489), .B2(n6488), .ZN(n6496)
         );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6494), .B1(n6493), 
        .B2(n6492), .ZN(n6495) );
  OAI211_X1 U7422 ( .C1(n6498), .C2(n6497), .A(n6496), .B(n6495), .ZN(U3147)
         );
  INV_X1 U7423 ( .A(n6499), .ZN(n6529) );
  NOR2_X1 U7424 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6504) );
  NOR2_X1 U7425 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  OAI211_X1 U7426 ( .C1(n6504), .C2(n6503), .A(n6532), .B(n6502), .ZN(n6505)
         );
  INV_X1 U7427 ( .A(n6505), .ZN(n6528) );
  NAND2_X1 U7428 ( .A1(n6526), .A2(n6525), .ZN(n6522) );
  OAI211_X1 U7429 ( .C1(n6508), .C2(n6507), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6506), .ZN(n6511) );
  INV_X1 U7430 ( .A(n6509), .ZN(n6510) );
  OAI21_X1 U7431 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6514) );
  NAND2_X1 U7432 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  OAI21_X1 U7433 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6518) );
  INV_X1 U7434 ( .A(n6518), .ZN(n6516) );
  NOR2_X1 U7435 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6516), .ZN(n6519)
         );
  OAI22_X1 U7436 ( .A1(n6520), .A2(n6519), .B1(n6518), .B2(n6517), .ZN(n6521)
         );
  NAND2_X1 U7437 ( .A1(n6522), .A2(n6521), .ZN(n6524) );
  OAI211_X1 U7438 ( .C1(n6526), .C2(n6525), .A(n6524), .B(n6523), .ZN(n6527)
         );
  INV_X1 U7439 ( .A(n6530), .ZN(n6531) );
  AND3_X1 U7440 ( .A1(n6533), .A2(n6532), .A3(n6531), .ZN(n6615) );
  NAND2_X1 U7441 ( .A1(n6547), .A2(n6548), .ZN(n6536) );
  NAND2_X1 U7442 ( .A1(READY_N), .A2(n6534), .ZN(n6535) );
  NAND2_X1 U7443 ( .A1(n6536), .A2(n6535), .ZN(n6540) );
  OR2_X1 U7444 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  OAI21_X1 U7445 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6627), .A(n6608), .ZN(
        n6550) );
  AOI221_X1 U7446 ( .B1(n6615), .B2(STATE2_REG_0__SCAN_IN), .C1(n6550), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6541), .ZN(n6545) );
  OAI211_X1 U7447 ( .C1(n6555), .C2(n6543), .A(n6542), .B(n6608), .ZN(n6544)
         );
  OAI211_X1 U7448 ( .C1(n6547), .C2(n6546), .A(n6545), .B(n6544), .ZN(U3148)
         );
  AOI21_X1 U7449 ( .B1(n6549), .B2(n6627), .A(n6548), .ZN(n6553) );
  OAI211_X1 U7450 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6550), .ZN(n6551) );
  OAI211_X1 U7451 ( .C1(n6554), .C2(n6553), .A(n6552), .B(n6551), .ZN(U3149)
         );
  INV_X1 U7452 ( .A(n6555), .ZN(n6631) );
  OAI221_X1 U7453 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6627), .A(n6606), .ZN(n6557) );
  OAI21_X1 U7454 ( .B1(n6631), .B2(n6557), .A(n6556), .ZN(U3150) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6603), .ZN(U3151) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6603), .ZN(U3152) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6603), .ZN(U3153) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6603), .ZN(U3154) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6603), .ZN(U3155) );
  AND2_X1 U7460 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6603), .ZN(U3156) );
  AND2_X1 U7461 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6603), .ZN(U3157) );
  AND2_X1 U7462 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6603), .ZN(U3158) );
  AND2_X1 U7463 ( .A1(n6603), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7464 ( .A1(n6603), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  INV_X1 U7465 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U7466 ( .A1(n6605), .A2(n6733), .ZN(U3161) );
  AND2_X1 U7467 ( .A1(n6603), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7468 ( .A1(n6603), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7469 ( .A1(n6603), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  INV_X1 U7470 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U7471 ( .A1(n6605), .A2(n6800), .ZN(U3165) );
  AND2_X1 U7472 ( .A1(n6603), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  INV_X1 U7473 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6805) );
  NOR2_X1 U7474 ( .A1(n6605), .A2(n6805), .ZN(U3167) );
  AND2_X1 U7475 ( .A1(n6603), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  INV_X1 U7476 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U7477 ( .A1(n6605), .A2(n6751), .ZN(U3169) );
  INV_X1 U7478 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U7479 ( .A1(n6605), .A2(n6738), .ZN(U3170) );
  INV_X1 U7480 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7021) );
  NOR2_X1 U7481 ( .A1(n6605), .A2(n7021), .ZN(U3171) );
  AND2_X1 U7482 ( .A1(n6603), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  INV_X1 U7483 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6806) );
  NOR2_X1 U7484 ( .A1(n6605), .A2(n6806), .ZN(U3173) );
  INV_X1 U7485 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U7486 ( .A1(n6605), .A2(n6709), .ZN(U3174) );
  INV_X1 U7487 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6794) );
  NOR2_X1 U7488 ( .A1(n6605), .A2(n6794), .ZN(U3175) );
  INV_X1 U7489 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U7490 ( .A1(n6605), .A2(n6964), .ZN(U3176) );
  AND2_X1 U7491 ( .A1(n6603), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  INV_X1 U7492 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U7493 ( .A1(n6605), .A2(n6687), .ZN(U3178) );
  INV_X1 U7494 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U7495 ( .A1(n6605), .A2(n6980), .ZN(U3179) );
  INV_X1 U7496 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U7497 ( .A1(n6605), .A2(n6791), .ZN(U3180) );
  NAND2_X1 U7498 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6573) );
  INV_X1 U7499 ( .A(n6573), .ZN(n6559) );
  NOR2_X1 U7500 ( .A1(n6627), .A2(n6965), .ZN(n6570) );
  AOI21_X1 U7501 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6570), .ZN(n6574)
         );
  OAI221_X1 U7502 ( .B1(n6575), .B2(NA_N), .C1(n6575), .C2(n6965), .A(n4260), 
        .ZN(n6567) );
  INV_X1 U7503 ( .A(HOLD), .ZN(n6565) );
  NOR2_X1 U7504 ( .A1(n6965), .A2(n6565), .ZN(n6560) );
  INV_X1 U7505 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6866) );
  OAI21_X1 U7506 ( .B1(n6560), .B2(n6866), .A(n7026), .ZN(n6558) );
  OAI211_X1 U7507 ( .C1(n6559), .C2(n6574), .A(n6567), .B(n6558), .ZN(U3181)
         );
  INV_X1 U7508 ( .A(n6570), .ZN(n6563) );
  NOR2_X1 U7509 ( .A1(n4260), .A2(n6866), .ZN(n6561) );
  OAI22_X1 U7510 ( .A1(n6561), .A2(n6560), .B1(n6575), .B2(n6565), .ZN(n6562)
         );
  NAND3_X1 U7511 ( .A1(n6564), .A2(n6563), .A3(n6562), .ZN(U3182) );
  INV_X1 U7512 ( .A(NA_N), .ZN(n6569) );
  AOI21_X1 U7513 ( .B1(n6569), .B2(READY_N), .A(n6965), .ZN(n6566) );
  AOI211_X1 U7514 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6575), .A(n6566), 
        .B(n6565), .ZN(n6568) );
  OAI21_X1 U7515 ( .B1(n6568), .B2(n4260), .A(n6567), .ZN(n6572) );
  NAND4_X1 U7516 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6570), .A4(n6569), .ZN(n6571) );
  OAI211_X1 U7517 ( .C1(n6574), .C2(n6573), .A(n6572), .B(n6571), .ZN(U3183)
         );
  NAND2_X1 U7518 ( .A1(n7027), .A2(n6575), .ZN(n6600) );
  INV_X1 U7519 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6577) );
  INV_X2 U7520 ( .A(n7026), .ZN(n7027) );
  OAI222_X1 U7521 ( .A1(n6600), .A2(n4832), .B1(n6577), .B2(n7027), .C1(n6576), 
        .C2(n6598), .ZN(U3184) );
  INV_X1 U7522 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6767) );
  OAI222_X1 U7523 ( .A1(n6598), .A2(n4832), .B1(n6767), .B2(n7027), .C1(n6578), 
        .C2(n6596), .ZN(U3185) );
  INV_X1 U7524 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6803) );
  OAI222_X1 U7525 ( .A1(n6598), .A2(n6578), .B1(n6803), .B2(n7027), .C1(n6579), 
        .C2(n6596), .ZN(U3186) );
  INV_X1 U7526 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6723) );
  OAI222_X1 U7527 ( .A1(n6598), .A2(n6579), .B1(n6723), .B2(n7027), .C1(n4914), 
        .C2(n6596), .ZN(U3187) );
  INV_X1 U7528 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6875) );
  OAI222_X1 U7529 ( .A1(n6600), .A2(n6580), .B1(n6875), .B2(n7027), .C1(n4914), 
        .C2(n6598), .ZN(U3188) );
  INV_X1 U7530 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6949) );
  INV_X1 U7531 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6581) );
  OAI222_X1 U7532 ( .A1(n6598), .A2(n6580), .B1(n6949), .B2(n7027), .C1(n6581), 
        .C2(n6596), .ZN(U3189) );
  INV_X1 U7533 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7000) );
  OAI222_X1 U7534 ( .A1(n6598), .A2(n6581), .B1(n7000), .B2(n7027), .C1(n6582), 
        .C2(n6600), .ZN(U3190) );
  INV_X1 U7535 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6982) );
  OAI222_X1 U7536 ( .A1(n6596), .A2(n6583), .B1(n6982), .B2(n7027), .C1(n6582), 
        .C2(n6598), .ZN(U3191) );
  INV_X1 U7537 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6753) );
  OAI222_X1 U7538 ( .A1(n6598), .A2(n6583), .B1(n6753), .B2(n7027), .C1(n6584), 
        .C2(n6600), .ZN(U3192) );
  INV_X1 U7539 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6970) );
  INV_X1 U7540 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6585) );
  OAI222_X1 U7541 ( .A1(n6598), .A2(n6584), .B1(n6970), .B2(n7027), .C1(n6585), 
        .C2(n6600), .ZN(U3193) );
  INV_X1 U7542 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6860) );
  OAI222_X1 U7543 ( .A1(n6600), .A2(n6587), .B1(n6860), .B2(n7027), .C1(n6585), 
        .C2(n6598), .ZN(U3194) );
  INV_X1 U7544 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6586) );
  OAI222_X1 U7545 ( .A1(n6598), .A2(n6587), .B1(n6586), .B2(n7027), .C1(n5773), 
        .C2(n6600), .ZN(U3195) );
  INV_X1 U7546 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6876) );
  OAI222_X1 U7547 ( .A1(n6598), .A2(n5773), .B1(n6876), .B2(n7027), .C1(n6588), 
        .C2(n6600), .ZN(U3196) );
  INV_X1 U7548 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6967) );
  OAI222_X1 U7549 ( .A1(n6600), .A2(n6589), .B1(n6967), .B2(n7027), .C1(n6588), 
        .C2(n6598), .ZN(U3197) );
  INV_X1 U7550 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6856) );
  OAI222_X1 U7551 ( .A1(n6598), .A2(n6589), .B1(n6856), .B2(n7027), .C1(n5054), 
        .C2(n6596), .ZN(U3198) );
  INV_X1 U7552 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6985) );
  OAI222_X1 U7553 ( .A1(n6598), .A2(n5054), .B1(n6985), .B2(n7027), .C1(n6969), 
        .C2(n6596), .ZN(U3199) );
  INV_X1 U7554 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6998) );
  OAI222_X1 U7555 ( .A1(n6598), .A2(n6969), .B1(n6998), .B2(n7027), .C1(n6764), 
        .C2(n6596), .ZN(U3200) );
  INV_X1 U7556 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6590) );
  OAI222_X1 U7557 ( .A1(n6596), .A2(n6727), .B1(n6590), .B2(n7027), .C1(n6764), 
        .C2(n6598), .ZN(U3201) );
  INV_X1 U7558 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6780) );
  OAI222_X1 U7559 ( .A1(n6600), .A2(n5423), .B1(n6780), .B2(n7027), .C1(n6727), 
        .C2(n6598), .ZN(U3202) );
  INV_X1 U7560 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U7561 ( .A1(n6598), .A2(n5423), .B1(n6591), .B2(n7027), .C1(n6897), 
        .C2(n6596), .ZN(U3203) );
  INV_X1 U7562 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6592) );
  OAI222_X1 U7563 ( .A1(n6598), .A2(n6897), .B1(n6592), .B2(n7027), .C1(n6887), 
        .C2(n6596), .ZN(U3204) );
  INV_X1 U7564 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6862) );
  OAI222_X1 U7565 ( .A1(n6598), .A2(n6887), .B1(n6862), .B2(n7027), .C1(n6992), 
        .C2(n6596), .ZN(U3205) );
  INV_X1 U7566 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U7567 ( .A1(n6598), .A2(n6992), .B1(n6593), .B2(n7027), .C1(n6747), 
        .C2(n6596), .ZN(U3206) );
  INV_X1 U7568 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7001) );
  OAI222_X1 U7569 ( .A1(n6596), .A2(n6594), .B1(n7001), .B2(n7027), .C1(n6747), 
        .C2(n6598), .ZN(U3207) );
  INV_X1 U7570 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6857) );
  OAI222_X1 U7571 ( .A1(n6598), .A2(n6594), .B1(n6857), .B2(n7027), .C1(n5395), 
        .C2(n6596), .ZN(U3208) );
  INV_X1 U7572 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6595) );
  OAI222_X1 U7573 ( .A1(n6598), .A2(n5395), .B1(n6595), .B2(n7027), .C1(n6863), 
        .C2(n6596), .ZN(U3209) );
  INV_X1 U7574 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6754) );
  OAI222_X1 U7575 ( .A1(n6598), .A2(n6863), .B1(n6754), .B2(n7027), .C1(n6973), 
        .C2(n6596), .ZN(U3210) );
  INV_X1 U7576 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6900) );
  OAI222_X1 U7577 ( .A1(n6598), .A2(n6973), .B1(n6900), .B2(n7027), .C1(n6597), 
        .C2(n6596), .ZN(U3211) );
  INV_X1 U7578 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U7579 ( .A1(n6598), .A2(n6597), .B1(n6766), .B2(n7027), .C1(n6599), 
        .C2(n6596), .ZN(U3212) );
  INV_X1 U7580 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6865) );
  OAI222_X1 U7581 ( .A1(n6600), .A2(n6786), .B1(n6865), .B2(n7027), .C1(n6599), 
        .C2(n6598), .ZN(U3213) );
  INV_X1 U7582 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6991) );
  INV_X1 U7583 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7584 ( .A1(n7027), .A2(n6991), .B1(n6777), .B2(n7026), .ZN(U3446)
         );
  INV_X1 U7585 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7586 ( .A1(n7027), .A2(n6736), .B1(n6950), .B2(n7026), .ZN(U3447)
         );
  INV_X1 U7587 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6984) );
  INV_X1 U7588 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7589 ( .A1(n7027), .A2(n6984), .B1(n6601), .B2(n7026), .ZN(U3448)
         );
  INV_X1 U7590 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6994) );
  INV_X1 U7591 ( .A(n6604), .ZN(n6602) );
  AOI21_X1 U7592 ( .B1(n6994), .B2(n6603), .A(n6602), .ZN(U3451) );
  OAI21_X1 U7593 ( .B1(n6605), .B2(n6883), .A(n6604), .ZN(U3452) );
  OAI211_X1 U7594 ( .C1(n6609), .C2(n6608), .A(n6607), .B(n6606), .ZN(U3453)
         );
  INV_X1 U7595 ( .A(n6610), .ZN(n6618) );
  AOI22_X1 U7596 ( .A1(n6614), .A2(n6613), .B1(n6612), .B2(n6611), .ZN(n6617)
         );
  NOR2_X1 U7597 ( .A1(n6618), .A2(n6615), .ZN(n6616) );
  AOI22_X1 U7598 ( .A1(n6619), .A2(n6618), .B1(n6617), .B2(n6616), .ZN(U3465)
         );
  AOI211_X1 U7599 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6620) );
  AOI21_X1 U7600 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6620), .ZN(n6621) );
  AOI22_X1 U7601 ( .A1(n6624), .A2(n6621), .B1(n6991), .B2(n6622), .ZN(U3468)
         );
  NOR2_X1 U7602 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6623) );
  AOI22_X1 U7603 ( .A1(n6624), .A2(n6623), .B1(n6984), .B2(n6622), .ZN(U3469)
         );
  INV_X1 U7604 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6879) );
  AOI22_X1 U7605 ( .A1(n7027), .A2(READREQUEST_REG_SCAN_IN), .B1(n6879), .B2(
        n7026), .ZN(U3470) );
  AOI211_X1 U7606 ( .C1(n6628), .C2(n6627), .A(n6626), .B(n6625), .ZN(n6635)
         );
  OAI211_X1 U7607 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6630), .A(n6629), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6632) );
  AOI21_X1 U7608 ( .B1(n6632), .B2(STATE2_REG_0__SCAN_IN), .A(n6631), .ZN(
        n6634) );
  NAND2_X1 U7609 ( .A1(n6635), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6633) );
  OAI21_X1 U7610 ( .B1(n6635), .B2(n6634), .A(n6633), .ZN(U3472) );
  INV_X1 U7611 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6749) );
  AOI22_X1 U7612 ( .A1(n7027), .A2(n6636), .B1(n6749), .B2(n7026), .ZN(U3473)
         );
  OAI22_X1 U7613 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g86), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n6637) );
  AOI221_X1 U7614 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_g101), .C1(
        ADDRESS_REG_14__SCAN_IN), .C2(keyinput_g86), .A(n6637), .ZN(n6644) );
  OAI22_X1 U7615 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(keyinput_g81), .ZN(n6638) );
  AOI221_X1 U7616 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(keyinput_g81), .C2(
        ADDRESS_REG_19__SCAN_IN), .A(n6638), .ZN(n6643) );
  OAI22_X1 U7617 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput_g124), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput_g70), .ZN(n6639) );
  AOI221_X1 U7618 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g70), .C2(BE_N_REG_0__SCAN_IN), .A(n6639), .ZN(n6642) );
  OAI22_X1 U7619 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .ZN(n6640) );
  AOI221_X1 U7620 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(keyinput_g85), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6640), .ZN(n6641) );
  NAND4_X1 U7621 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6672)
         );
  OAI22_X1 U7622 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .ZN(n6645) );
  AOI221_X1 U7623 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(keyinput_g37), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6645), .ZN(n6652) );
  OAI22_X1 U7624 ( .A1(DATAI_30_), .A2(keyinput_g1), .B1(keyinput_g93), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n6646) );
  AOI221_X1 U7625 ( .B1(DATAI_30_), .B2(keyinput_g1), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput_g93), .A(n6646), .ZN(n6651) );
  OAI22_X1 U7626 ( .A1(NA_N), .A2(keyinput_g33), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(keyinput_g96), .ZN(n6647) );
  AOI221_X1 U7627 ( .B1(NA_N), .B2(keyinput_g33), .C1(keyinput_g96), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6647), .ZN(n6650) );
  OAI22_X1 U7628 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(keyinput_g120), .B2(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6648) );
  AOI221_X1 U7629 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput_g120), .A(n6648), .ZN(n6649)
         );
  NAND4_X1 U7630 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6671)
         );
  OAI22_X1 U7631 ( .A1(ADDRESS_REG_20__SCAN_IN), .A2(keyinput_g80), .B1(
        keyinput_g91), .B2(ADDRESS_REG_9__SCAN_IN), .ZN(n6653) );
  AOI221_X1 U7632 ( .B1(ADDRESS_REG_20__SCAN_IN), .B2(keyinput_g80), .C1(
        ADDRESS_REG_9__SCAN_IN), .C2(keyinput_g91), .A(n6653), .ZN(n6660) );
  OAI22_X1 U7633 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_g52), .B1(DATAI_14_), .B2(keyinput_g17), .ZN(n6654) );
  AOI221_X1 U7634 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g17), .C2(DATAI_14_), .A(n6654), .ZN(n6659) );
  OAI22_X1 U7635 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_g57), .B1(
        DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput_g126), .ZN(n6655) );
  AOI221_X1 U7636 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g126), .C2(DATAWIDTH_REG_22__SCAN_IN), .A(n6655), .ZN(n6658)
         );
  OAI22_X1 U7637 ( .A1(ADDRESS_REG_22__SCAN_IN), .A2(keyinput_g78), .B1(
        BE_N_REG_3__SCAN_IN), .B2(keyinput_g67), .ZN(n6656) );
  AOI221_X1 U7638 ( .B1(ADDRESS_REG_22__SCAN_IN), .B2(keyinput_g78), .C1(
        keyinput_g67), .C2(BE_N_REG_3__SCAN_IN), .A(n6656), .ZN(n6657) );
  NAND4_X1 U7639 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6670)
         );
  OAI22_X1 U7640 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(keyinput_g79), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n6661) );
  AOI221_X1 U7641 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(
        ADDRESS_REG_21__SCAN_IN), .C2(keyinput_g79), .A(n6661), .ZN(n6668) );
  OAI22_X1 U7642 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(keyinput_g42), .B2(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6662) );
  AOI221_X1 U7643 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g42), .A(n6662), .ZN(n6667)
         );
  OAI22_X1 U7644 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(
        DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_g118), .ZN(n6663) );
  AOI221_X1 U7645 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(keyinput_g118), 
        .C2(DATAWIDTH_REG_14__SCAN_IN), .A(n6663), .ZN(n6666) );
  OAI22_X1 U7646 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_19_), .B2(
        keyinput_g12), .ZN(n6664) );
  AOI221_X1 U7647 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(keyinput_g12), .C2(
        DATAI_19_), .A(n6664), .ZN(n6665) );
  NAND4_X1 U7648 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6669)
         );
  NOR4_X1 U7649 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n7025)
         );
  OAI22_X1 U7650 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput_g83), .B1(
        keyinput_g123), .B2(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6673) );
  AOI221_X1 U7651 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput_g83), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput_g123), .A(n6673), .ZN(n6680)
         );
  OAI22_X1 U7652 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .ZN(n6674) );
  AOI221_X1 U7653 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        keyinput_g88), .C2(ADDRESS_REG_12__SCAN_IN), .A(n6674), .ZN(n6679) );
  OAI22_X1 U7654 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(keyinput_g107), .B2(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6675) );
  AOI221_X1 U7655 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(
        DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput_g107), .A(n6675), .ZN(n6678)
         );
  OAI22_X1 U7656 ( .A1(DATAI_0_), .A2(keyinput_g31), .B1(
        DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .ZN(n6676) );
  AOI221_X1 U7657 ( .B1(DATAI_0_), .B2(keyinput_g31), .C1(keyinput_g110), .C2(
        DATAWIDTH_REG_6__SCAN_IN), .A(n6676), .ZN(n6677) );
  NAND4_X1 U7658 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n6818)
         );
  OAI22_X1 U7659 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        HOLD), .B2(keyinput_g36), .ZN(n6681) );
  AOI221_X1 U7660 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g36), .C2(HOLD), .A(n6681), .ZN(n6707) );
  OAI22_X1 U7661 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g114), .B2(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6682) );
  AOI221_X1 U7662 ( .B1(ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .C1(
        DATAWIDTH_REG_10__SCAN_IN), .C2(keyinput_g114), .A(n6682), .ZN(n6685)
         );
  OAI22_X1 U7663 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput_g122), .B1(
        DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput_g105), .ZN(n6683) );
  AOI221_X1 U7664 ( .B1(DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g105), .C2(DATAWIDTH_REG_1__SCAN_IN), .A(n6683), .ZN(n6684)
         );
  OAI211_X1 U7665 ( .C1(n6687), .C2(keyinput_g108), .A(n6685), .B(n6684), .ZN(
        n6686) );
  AOI21_X1 U7666 ( .B1(n6687), .B2(keyinput_g108), .A(n6686), .ZN(n6706) );
  AOI22_X1 U7667 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(DATAI_17_), 
        .B2(keyinput_g14), .ZN(n6688) );
  OAI221_X1 U7668 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(DATAI_17_), 
        .C2(keyinput_g14), .A(n6688), .ZN(n6695) );
  AOI22_X1 U7669 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_g90), .B1(
        DATAI_1_), .B2(keyinput_g30), .ZN(n6689) );
  OAI221_X1 U7670 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_g90), .C1(
        DATAI_1_), .C2(keyinput_g30), .A(n6689), .ZN(n6694) );
  AOI22_X1 U7671 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6690) );
  OAI221_X1 U7672 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6690), .ZN(n6693) );
  AOI22_X1 U7673 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(DATAI_28_), 
        .B2(keyinput_g3), .ZN(n6691) );
  OAI221_X1 U7674 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(DATAI_28_), 
        .C2(keyinput_g3), .A(n6691), .ZN(n6692) );
  NOR4_X1 U7675 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6705)
         );
  AOI22_X1 U7676 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput_g94), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(keyinput_g100), .ZN(n6696) );
  OAI221_X1 U7677 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .C1(
        ADDRESS_REG_0__SCAN_IN), .C2(keyinput_g100), .A(n6696), .ZN(n6703) );
  AOI22_X1 U7678 ( .A1(DATAI_25_), .A2(keyinput_g6), .B1(READY_N), .B2(
        keyinput_g35), .ZN(n6697) );
  OAI221_X1 U7679 ( .B1(DATAI_25_), .B2(keyinput_g6), .C1(READY_N), .C2(
        keyinput_g35), .A(n6697), .ZN(n6702) );
  AOI22_X1 U7680 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput_g109), .B1(
        D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .ZN(n6698) );
  OAI221_X1 U7681 ( .B1(DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput_g109), .C1(
        D_C_N_REG_SCAN_IN), .C2(keyinput_g41), .A(n6698), .ZN(n6701) );
  AOI22_X1 U7682 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput_g89), .B1(
        REIP_REG_29__SCAN_IN), .B2(keyinput_g53), .ZN(n6699) );
  OAI221_X1 U7683 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput_g89), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_g53), .A(n6699), .ZN(n6700) );
  NOR4_X1 U7684 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6704)
         );
  NAND4_X1 U7685 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6817)
         );
  AOI22_X1 U7686 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_g66), .B1(n6709), 
        .B2(keyinput_g112), .ZN(n6708) );
  OAI221_X1 U7687 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_g66), .C1(n6709), 
        .C2(keyinput_g112), .A(n6708), .ZN(n6719) );
  AOI22_X1 U7688 ( .A1(n6873), .A2(keyinput_g29), .B1(keyinput_g38), .B2(n6872), .ZN(n6710) );
  OAI221_X1 U7689 ( .B1(n6873), .B2(keyinput_g29), .C1(n6872), .C2(
        keyinput_g38), .A(n6710), .ZN(n6718) );
  INV_X1 U7690 ( .A(BS16_N), .ZN(n6712) );
  AOI22_X1 U7691 ( .A1(n6712), .A2(keyinput_g34), .B1(keyinput_g76), .B2(n6857), .ZN(n6711) );
  OAI221_X1 U7692 ( .B1(n6712), .B2(keyinput_g34), .C1(n6857), .C2(
        keyinput_g76), .A(n6711), .ZN(n6717) );
  AOI22_X1 U7693 ( .A1(n6715), .A2(keyinput_g9), .B1(n6714), .B2(keyinput_g23), 
        .ZN(n6713) );
  OAI221_X1 U7694 ( .B1(n6715), .B2(keyinput_g9), .C1(n6714), .C2(keyinput_g23), .A(n6713), .ZN(n6716) );
  NOR4_X1 U7695 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6762)
         );
  AOI22_X1 U7696 ( .A1(n6950), .A2(keyinput_g69), .B1(n6721), .B2(keyinput_g45), .ZN(n6720) );
  OAI221_X1 U7697 ( .B1(n6950), .B2(keyinput_g69), .C1(n6721), .C2(
        keyinput_g45), .A(n6720), .ZN(n6731) );
  AOI22_X1 U7698 ( .A1(n4260), .A2(keyinput_g103), .B1(keyinput_g97), .B2(
        n6723), .ZN(n6722) );
  OAI221_X1 U7699 ( .B1(n4260), .B2(keyinput_g103), .C1(n6723), .C2(
        keyinput_g97), .A(n6722), .ZN(n6730) );
  AOI22_X1 U7700 ( .A1(n6725), .A2(keyinput_g15), .B1(n4763), .B2(keyinput_g2), 
        .ZN(n6724) );
  OAI221_X1 U7701 ( .B1(n6725), .B2(keyinput_g15), .C1(n4763), .C2(keyinput_g2), .A(n6724), .ZN(n6729) );
  AOI22_X1 U7702 ( .A1(n6969), .A2(keyinput_g65), .B1(keyinput_g63), .B2(n6727), .ZN(n6726) );
  OAI221_X1 U7703 ( .B1(n6969), .B2(keyinput_g65), .C1(n6727), .C2(
        keyinput_g63), .A(n6726), .ZN(n6728) );
  NOR4_X1 U7704 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6761)
         );
  AOI22_X1 U7705 ( .A1(n6992), .A2(keyinput_g59), .B1(keyinput_g125), .B2(
        n6733), .ZN(n6732) );
  OAI221_X1 U7706 ( .B1(n6992), .B2(keyinput_g59), .C1(n6733), .C2(
        keyinput_g125), .A(n6732), .ZN(n6745) );
  AOI22_X1 U7707 ( .A1(n6736), .A2(keyinput_g48), .B1(n6735), .B2(keyinput_g26), .ZN(n6734) );
  OAI221_X1 U7708 ( .B1(n6736), .B2(keyinput_g48), .C1(n6735), .C2(
        keyinput_g26), .A(n6734), .ZN(n6744) );
  AOI22_X1 U7709 ( .A1(n6739), .A2(keyinput_g18), .B1(keyinput_g116), .B2(
        n6738), .ZN(n6737) );
  OAI221_X1 U7710 ( .B1(n6739), .B2(keyinput_g18), .C1(n6738), .C2(
        keyinput_g116), .A(n6737), .ZN(n6743) );
  AOI22_X1 U7711 ( .A1(n6741), .A2(keyinput_g50), .B1(n6863), .B2(keyinput_g55), .ZN(n6740) );
  OAI221_X1 U7712 ( .B1(n6741), .B2(keyinput_g50), .C1(n6863), .C2(
        keyinput_g55), .A(n6740), .ZN(n6742) );
  NOR4_X1 U7713 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6760)
         );
  AOI22_X1 U7714 ( .A1(n6984), .A2(keyinput_g47), .B1(n6747), .B2(keyinput_g58), .ZN(n6746) );
  OAI221_X1 U7715 ( .B1(n6984), .B2(keyinput_g47), .C1(n6747), .C2(
        keyinput_g58), .A(n6746), .ZN(n6758) );
  AOI22_X1 U7716 ( .A1(n6749), .A2(keyinput_g40), .B1(n4736), .B2(keyinput_g4), 
        .ZN(n6748) );
  OAI221_X1 U7717 ( .B1(n6749), .B2(keyinput_g40), .C1(n4736), .C2(keyinput_g4), .A(n6748), .ZN(n6757) );
  AOI22_X1 U7718 ( .A1(n6995), .A2(keyinput_g8), .B1(keyinput_g117), .B2(n6751), .ZN(n6750) );
  OAI221_X1 U7719 ( .B1(n6995), .B2(keyinput_g8), .C1(n6751), .C2(
        keyinput_g117), .A(n6750), .ZN(n6756) );
  AOI22_X1 U7720 ( .A1(n6754), .A2(keyinput_g74), .B1(n6753), .B2(keyinput_g92), .ZN(n6752) );
  OAI221_X1 U7721 ( .B1(n6754), .B2(keyinput_g74), .C1(n6753), .C2(
        keyinput_g92), .A(n6752), .ZN(n6755) );
  NOR4_X1 U7722 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6759)
         );
  NAND4_X1 U7723 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6816)
         );
  AOI22_X1 U7724 ( .A1(n5423), .A2(keyinput_g62), .B1(n6764), .B2(keyinput_g64), .ZN(n6763) );
  OAI221_X1 U7725 ( .B1(n5423), .B2(keyinput_g62), .C1(n6764), .C2(
        keyinput_g64), .A(n6763), .ZN(n6773) );
  AOI22_X1 U7726 ( .A1(n6767), .A2(keyinput_g99), .B1(keyinput_g72), .B2(n6766), .ZN(n6765) );
  OAI221_X1 U7727 ( .B1(n6767), .B2(keyinput_g99), .C1(n6766), .C2(
        keyinput_g72), .A(n6765), .ZN(n6772) );
  AOI22_X1 U7728 ( .A1(n6887), .A2(keyinput_g60), .B1(n6965), .B2(
        keyinput_g102), .ZN(n6768) );
  OAI221_X1 U7729 ( .B1(n6887), .B2(keyinput_g60), .C1(n6965), .C2(
        keyinput_g102), .A(n6768), .ZN(n6771) );
  INV_X1 U7730 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7731 ( .A1(n6967), .A2(keyinput_g87), .B1(n6899), .B2(keyinput_g39), .ZN(n6769) );
  OAI221_X1 U7732 ( .B1(n6967), .B2(keyinput_g87), .C1(n6899), .C2(
        keyinput_g39), .A(n6769), .ZN(n6770) );
  NOR4_X1 U7733 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6814)
         );
  AOI22_X1 U7734 ( .A1(n6775), .A2(keyinput_g21), .B1(keyinput_g28), .B2(n6997), .ZN(n6774) );
  OAI221_X1 U7735 ( .B1(n6775), .B2(keyinput_g21), .C1(n6997), .C2(
        keyinput_g28), .A(n6774), .ZN(n6784) );
  AOI22_X1 U7736 ( .A1(n6777), .A2(keyinput_g68), .B1(keyinput_g73), .B2(n6900), .ZN(n6776) );
  OAI221_X1 U7737 ( .B1(n6777), .B2(keyinput_g68), .C1(n6900), .C2(
        keyinput_g73), .A(n6776), .ZN(n6783) );
  AOI22_X1 U7738 ( .A1(n6949), .A2(keyinput_g95), .B1(n4645), .B2(keyinput_g0), 
        .ZN(n6778) );
  OAI221_X1 U7739 ( .B1(n6949), .B2(keyinput_g95), .C1(n4645), .C2(keyinput_g0), .A(n6778), .ZN(n6782) );
  AOI22_X1 U7740 ( .A1(n6958), .A2(keyinput_g13), .B1(keyinput_g82), .B2(n6780), .ZN(n6779) );
  OAI221_X1 U7741 ( .B1(n6958), .B2(keyinput_g13), .C1(n6780), .C2(
        keyinput_g82), .A(n6779), .ZN(n6781) );
  NOR4_X1 U7742 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(n6813)
         );
  AOI22_X1 U7743 ( .A1(n6998), .A2(keyinput_g84), .B1(n6786), .B2(keyinput_g51), .ZN(n6785) );
  OAI221_X1 U7744 ( .B1(n6998), .B2(keyinput_g84), .C1(n6786), .C2(
        keyinput_g51), .A(n6785), .ZN(n6798) );
  AOI22_X1 U7745 ( .A1(n6788), .A2(keyinput_g19), .B1(keyinput_g49), .B2(n6991), .ZN(n6787) );
  OAI221_X1 U7746 ( .B1(n6788), .B2(keyinput_g19), .C1(n6991), .C2(
        keyinput_g49), .A(n6787), .ZN(n6797) );
  AOI22_X1 U7747 ( .A1(n6791), .A2(keyinput_g106), .B1(n6790), .B2(
        keyinput_g27), .ZN(n6789) );
  OAI221_X1 U7748 ( .B1(n6791), .B2(keyinput_g106), .C1(n6790), .C2(
        keyinput_g27), .A(n6789), .ZN(n6796) );
  AOI22_X1 U7749 ( .A1(n6794), .A2(keyinput_g111), .B1(n6793), .B2(
        keyinput_g43), .ZN(n6792) );
  OAI221_X1 U7750 ( .B1(n6794), .B2(keyinput_g111), .C1(n6793), .C2(
        keyinput_g43), .A(n6792), .ZN(n6795) );
  NOR4_X1 U7751 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n6812)
         );
  AOI22_X1 U7752 ( .A1(n6800), .A2(keyinput_g121), .B1(n6865), .B2(
        keyinput_g71), .ZN(n6799) );
  OAI221_X1 U7753 ( .B1(n6800), .B2(keyinput_g121), .C1(n6865), .C2(
        keyinput_g71), .A(n6799), .ZN(n6810) );
  AOI22_X1 U7754 ( .A1(n7001), .A2(keyinput_g77), .B1(n6897), .B2(keyinput_g61), .ZN(n6801) );
  OAI221_X1 U7755 ( .B1(n7001), .B2(keyinput_g77), .C1(n6897), .C2(
        keyinput_g61), .A(n6801), .ZN(n6809) );
  AOI22_X1 U7756 ( .A1(n5395), .A2(keyinput_g56), .B1(keyinput_g98), .B2(n6803), .ZN(n6802) );
  OAI221_X1 U7757 ( .B1(n5395), .B2(keyinput_g56), .C1(n6803), .C2(
        keyinput_g98), .A(n6802), .ZN(n6808) );
  AOI22_X1 U7758 ( .A1(n6806), .A2(keyinput_g113), .B1(keyinput_g119), .B2(
        n6805), .ZN(n6804) );
  OAI221_X1 U7759 ( .B1(n6806), .B2(keyinput_g113), .C1(n6805), .C2(
        keyinput_g119), .A(n6804), .ZN(n6807) );
  NOR4_X1 U7760 ( .A1(n6810), .A2(n6809), .A3(n6808), .A4(n6807), .ZN(n6811)
         );
  NAND4_X1 U7761 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6815)
         );
  NOR4_X1 U7762 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n7024)
         );
  OAI22_X1 U7763 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_f101), .B1(
        DATAI_27_), .B2(keyinput_f4), .ZN(n6819) );
  AOI221_X1 U7764 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f4), .C2(DATAI_27_), .A(n6819), .ZN(n6826) );
  OAI22_X1 U7765 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(keyinput_f83), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n6820) );
  AOI221_X1 U7766 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput_f83), .A(n6820), .ZN(n6825) );
  OAI22_X1 U7767 ( .A1(keyinput_f92), .A2(ADDRESS_REG_8__SCAN_IN), .B1(
        keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .ZN(n6821) );
  AOI221_X1 U7768 ( .B1(keyinput_f92), .B2(ADDRESS_REG_8__SCAN_IN), .C1(
        ADDRESS_REG_25__SCAN_IN), .C2(keyinput_f75), .A(n6821), .ZN(n6824) );
  OAI22_X1 U7769 ( .A1(keyinput_f81), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        keyinput_f108), .B2(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6822) );
  AOI221_X1 U7770 ( .B1(keyinput_f81), .B2(ADDRESS_REG_19__SCAN_IN), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput_f108), .A(n6822), .ZN(n6823)
         );
  NAND4_X1 U7771 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6854)
         );
  OAI22_X1 U7772 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_f123), .ZN(n6827) );
  AOI221_X1 U7773 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f123), .C2(DATAWIDTH_REG_19__SCAN_IN), .A(n6827), .ZN(n6834)
         );
  OAI22_X1 U7774 ( .A1(keyinput_f106), .A2(DATAWIDTH_REG_2__SCAN_IN), .B1(
        keyinput_f114), .B2(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6828) );
  AOI221_X1 U7775 ( .B1(keyinput_f106), .B2(DATAWIDTH_REG_2__SCAN_IN), .C1(
        DATAWIDTH_REG_10__SCAN_IN), .C2(keyinput_f114), .A(n6828), .ZN(n6833)
         );
  OAI22_X1 U7776 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_24_), .B2(
        keyinput_f7), .ZN(n6829) );
  AOI221_X1 U7777 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(keyinput_f7), .C2(
        DATAI_24_), .A(n6829), .ZN(n6832) );
  OAI22_X1 U7778 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(DATAI_22_), .B2(keyinput_f9), .ZN(n6830) );
  AOI221_X1 U7779 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f9), .C2(DATAI_22_), .A(n6830), .ZN(n6831) );
  NAND4_X1 U7780 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n6853)
         );
  OAI22_X1 U7781 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_19_), .B2(
        keyinput_f12), .ZN(n6835) );
  AOI221_X1 U7782 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(keyinput_f12), .C2(
        DATAI_19_), .A(n6835), .ZN(n6842) );
  OAI22_X1 U7783 ( .A1(keyinput_f111), .A2(DATAWIDTH_REG_7__SCAN_IN), .B1(
        keyinput_f127), .B2(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6836) );
  AOI221_X1 U7784 ( .B1(keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .C1(
        DATAWIDTH_REG_23__SCAN_IN), .C2(keyinput_f127), .A(n6836), .ZN(n6841)
         );
  OAI22_X1 U7785 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f124), .B2(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6837) );
  AOI221_X1 U7786 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput_f124), .A(n6837), .ZN(n6840)
         );
  OAI22_X1 U7787 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        keyinput_f97), .B2(ADDRESS_REG_3__SCAN_IN), .ZN(n6838) );
  AOI221_X1 U7788 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        ADDRESS_REG_3__SCAN_IN), .C2(keyinput_f97), .A(n6838), .ZN(n6839) );
  NAND4_X1 U7789 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6852)
         );
  OAI22_X1 U7790 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f32), .B2(MEMORYFETCH_REG_SCAN_IN), .ZN(n6843) );
  AOI221_X1 U7791 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_f32), .A(n6843), .ZN(n6850) );
  OAI22_X1 U7792 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_f103), .B1(
        DATAI_17_), .B2(keyinput_f14), .ZN(n6844) );
  AOI221_X1 U7793 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f14), .C2(DATAI_17_), .A(n6844), .ZN(n6849) );
  OAI22_X1 U7794 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_f64), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n6845) );
  AOI221_X1 U7795 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .C1(
        keyinput_f44), .C2(MORE_REG_SCAN_IN), .A(n6845), .ZN(n6848) );
  OAI22_X1 U7796 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(keyinput_f98), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n6846) );
  AOI221_X1 U7797 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(
        ADDRESS_REG_2__SCAN_IN), .C2(keyinput_f98), .A(n6846), .ZN(n6847) );
  NAND4_X1 U7798 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6851)
         );
  NOR4_X1 U7799 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n7017)
         );
  AOI22_X1 U7800 ( .A1(n6857), .A2(keyinput_f76), .B1(keyinput_f86), .B2(n6856), .ZN(n6855) );
  OAI221_X1 U7801 ( .B1(n6857), .B2(keyinput_f76), .C1(n6856), .C2(
        keyinput_f86), .A(n6855), .ZN(n6870) );
  AOI22_X1 U7802 ( .A1(n6860), .A2(keyinput_f90), .B1(n6859), .B2(keyinput_f30), .ZN(n6858) );
  OAI221_X1 U7803 ( .B1(n6860), .B2(keyinput_f90), .C1(n6859), .C2(
        keyinput_f30), .A(n6858), .ZN(n6869) );
  AOI22_X1 U7804 ( .A1(n6863), .A2(keyinput_f55), .B1(keyinput_f79), .B2(n6862), .ZN(n6861) );
  OAI221_X1 U7805 ( .B1(n6863), .B2(keyinput_f55), .C1(n6862), .C2(
        keyinput_f79), .A(n6861), .ZN(n6868) );
  AOI22_X1 U7806 ( .A1(n6866), .A2(keyinput_f42), .B1(keyinput_f71), .B2(n6865), .ZN(n6864) );
  OAI221_X1 U7807 ( .B1(n6866), .B2(keyinput_f42), .C1(n6865), .C2(
        keyinput_f71), .A(n6864), .ZN(n6867) );
  NOR4_X1 U7808 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n7016)
         );
  AOI22_X1 U7809 ( .A1(n6873), .A2(keyinput_f29), .B1(keyinput_f38), .B2(n6872), .ZN(n6871) );
  OAI221_X1 U7810 ( .B1(n6873), .B2(keyinput_f29), .C1(n6872), .C2(
        keyinput_f38), .A(n6871), .ZN(n6912) );
  AOI22_X1 U7811 ( .A1(n6876), .A2(keyinput_f88), .B1(keyinput_f96), .B2(n6875), .ZN(n6874) );
  OAI221_X1 U7812 ( .B1(n6876), .B2(keyinput_f88), .C1(n6875), .C2(
        keyinput_f96), .A(n6874), .ZN(n6911) );
  XOR2_X1 U7813 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_f82), .Z(n6881) );
  INV_X1 U7814 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7815 ( .A1(n6879), .A2(keyinput_f46), .B1(n6878), .B2(keyinput_f37), .ZN(n6877) );
  OAI221_X1 U7816 ( .B1(n6879), .B2(keyinput_f46), .C1(n6878), .C2(
        keyinput_f37), .A(n6877), .ZN(n6880) );
  AOI211_X1 U7817 ( .C1(n6883), .C2(keyinput_f105), .A(n6881), .B(n6880), .ZN(
        n6882) );
  OAI21_X1 U7818 ( .B1(n6883), .B2(keyinput_f105), .A(n6882), .ZN(n6910) );
  OAI22_X1 U7819 ( .A1(keyinput_f119), .A2(DATAWIDTH_REG_15__SCAN_IN), .B1(
        keyinput_f34), .B2(BS16_N), .ZN(n6884) );
  AOI221_X1 U7820 ( .B1(keyinput_f119), .B2(DATAWIDTH_REG_15__SCAN_IN), .C1(
        BS16_N), .C2(keyinput_f34), .A(n6884), .ZN(n6908) );
  XOR2_X1 U7821 ( .A(keyinput_f125), .B(DATAWIDTH_REG_21__SCAN_IN), .Z(n6892)
         );
  XOR2_X1 U7822 ( .A(ADDRESS_REG_28__SCAN_IN), .B(keyinput_f72), .Z(n6891) );
  AOI22_X1 U7823 ( .A1(keyinput_f100), .A2(ADDRESS_REG_0__SCAN_IN), .B1(
        keyinput_f122), .B2(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6885) );
  OAI221_X1 U7824 ( .B1(keyinput_f100), .B2(ADDRESS_REG_0__SCAN_IN), .C1(
        keyinput_f122), .C2(DATAWIDTH_REG_18__SCAN_IN), .A(n6885), .ZN(n6890)
         );
  AOI22_X1 U7825 ( .A1(n6888), .A2(keyinput_f20), .B1(n6887), .B2(keyinput_f60), .ZN(n6886) );
  OAI221_X1 U7826 ( .B1(n6888), .B2(keyinput_f20), .C1(n6887), .C2(
        keyinput_f60), .A(n6886), .ZN(n6889) );
  NOR4_X1 U7827 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6907)
         );
  INV_X1 U7828 ( .A(keyinput_f67), .ZN(n6894) );
  OAI22_X1 U7829 ( .A1(n6895), .A2(keyinput_f22), .B1(n6894), .B2(
        BE_N_REG_3__SCAN_IN), .ZN(n6893) );
  AOI221_X1 U7830 ( .B1(n6895), .B2(keyinput_f22), .C1(BE_N_REG_3__SCAN_IN), 
        .C2(n6894), .A(n6893), .ZN(n6906) );
  XOR2_X1 U7831 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_f70), .Z(n6904) );
  XOR2_X1 U7832 ( .A(keyinput_f36), .B(HOLD), .Z(n6903) );
  AOI22_X1 U7833 ( .A1(n4645), .A2(keyinput_f0), .B1(n6897), .B2(keyinput_f61), 
        .ZN(n6896) );
  OAI221_X1 U7834 ( .B1(n4645), .B2(keyinput_f0), .C1(n6897), .C2(keyinput_f61), .A(n6896), .ZN(n6902) );
  AOI22_X1 U7835 ( .A1(n6900), .A2(keyinput_f73), .B1(n6899), .B2(keyinput_f39), .ZN(n6898) );
  OAI221_X1 U7836 ( .B1(n6900), .B2(keyinput_f73), .C1(n6899), .C2(
        keyinput_f39), .A(n6898), .ZN(n6901) );
  NOR4_X1 U7837 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6905)
         );
  NAND4_X1 U7838 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), .ZN(n6909)
         );
  NOR4_X1 U7839 ( .A1(n6912), .A2(n6911), .A3(n6910), .A4(n6909), .ZN(n7015)
         );
  OAI22_X1 U7840 ( .A1(keyinput_f126), .A2(DATAWIDTH_REG_22__SCAN_IN), .B1(
        keyinput_f78), .B2(ADDRESS_REG_22__SCAN_IN), .ZN(n6913) );
  AOI221_X1 U7841 ( .B1(keyinput_f126), .B2(DATAWIDTH_REG_22__SCAN_IN), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_f78), .A(n6913), .ZN(n6920) );
  OAI22_X1 U7842 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(
        BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_f50), .ZN(n6914) );
  AOI221_X1 U7843 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(keyinput_f50), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n6914), .ZN(n6919) );
  OAI22_X1 U7844 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f118), .B2(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6915) );
  AOI221_X1 U7845 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(
        DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput_f118), .A(n6915), .ZN(n6918)
         );
  OAI22_X1 U7846 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(FLUSH_REG_SCAN_IN), 
        .B2(keyinput_f45), .ZN(n6916) );
  AOI221_X1 U7847 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(keyinput_f45), .C2(
        FLUSH_REG_SCAN_IN), .A(n6916), .ZN(n6917) );
  NAND4_X1 U7848 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n7013)
         );
  OAI22_X1 U7849 ( .A1(keyinput_f68), .A2(BE_N_REG_2__SCAN_IN), .B1(
        keyinput_f112), .B2(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6921) );
  AOI221_X1 U7850 ( .B1(keyinput_f68), .B2(BE_N_REG_2__SCAN_IN), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput_f112), .A(n6921), .ZN(n6947)
         );
  OAI22_X1 U7851 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(keyinput_f89), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n6922) );
  AOI221_X1 U7852 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(
        ADDRESS_REG_11__SCAN_IN), .C2(keyinput_f89), .A(n6922), .ZN(n6925) );
  OAI22_X1 U7853 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f113), .B2(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6923) );
  AOI221_X1 U7854 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_f113), .A(n6923), .ZN(n6924)
         );
  OAI211_X1 U7855 ( .C1(n6927), .C2(keyinput_f16), .A(n6925), .B(n6924), .ZN(
        n6926) );
  AOI21_X1 U7856 ( .B1(n6927), .B2(keyinput_f16), .A(n6926), .ZN(n6946) );
  AOI22_X1 U7857 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(READY_N), .B2(
        keyinput_f35), .ZN(n6928) );
  OAI221_X1 U7858 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(READY_N), .C2(
        keyinput_f35), .A(n6928), .ZN(n6935) );
  AOI22_X1 U7859 ( .A1(keyinput_f33), .A2(NA_N), .B1(keyinput_f41), .B2(
        D_C_N_REG_SCAN_IN), .ZN(n6929) );
  OAI221_X1 U7860 ( .B1(keyinput_f33), .B2(NA_N), .C1(keyinput_f41), .C2(
        D_C_N_REG_SCAN_IN), .A(n6929), .ZN(n6934) );
  AOI22_X1 U7861 ( .A1(keyinput_f99), .A2(ADDRESS_REG_1__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .ZN(n6930) );
  OAI221_X1 U7862 ( .B1(keyinput_f99), .B2(ADDRESS_REG_1__SCAN_IN), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n6930), .ZN(n6933) );
  AOI22_X1 U7863 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(DATAI_20_), .B2(
        keyinput_f11), .ZN(n6931) );
  OAI221_X1 U7864 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(DATAI_20_), .C2(
        keyinput_f11), .A(n6931), .ZN(n6932) );
  NOR4_X1 U7865 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(n6945)
         );
  AOI22_X1 U7866 ( .A1(keyinput_f80), .A2(ADDRESS_REG_20__SCAN_IN), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .ZN(n6936) );
  OAI221_X1 U7867 ( .B1(keyinput_f80), .B2(ADDRESS_REG_20__SCAN_IN), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6936), .ZN(n6943) );
  AOI22_X1 U7868 ( .A1(keyinput_f117), .A2(DATAWIDTH_REG_13__SCAN_IN), .B1(
        keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6937) );
  OAI221_X1 U7869 ( .B1(keyinput_f117), .B2(DATAWIDTH_REG_13__SCAN_IN), .C1(
        keyinput_f48), .C2(BYTEENABLE_REG_1__SCAN_IN), .A(n6937), .ZN(n6942)
         );
  AOI22_X1 U7870 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(DATAI_26_), .B2(
        keyinput_f5), .ZN(n6938) );
  OAI221_X1 U7871 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n6938), .ZN(n6941) );
  AOI22_X1 U7872 ( .A1(keyinput_f40), .A2(M_IO_N_REG_SCAN_IN), .B1(DATAI_10_), 
        .B2(keyinput_f21), .ZN(n6939) );
  OAI221_X1 U7873 ( .B1(keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .C1(DATAI_10_), 
        .C2(keyinput_f21), .A(n6939), .ZN(n6940) );
  NOR4_X1 U7874 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n6944)
         );
  NAND4_X1 U7875 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n7012)
         );
  OAI22_X1 U7876 ( .A1(n6950), .A2(keyinput_f69), .B1(n6949), .B2(keyinput_f95), .ZN(n6948) );
  AOI221_X1 U7877 ( .B1(n6950), .B2(keyinput_f69), .C1(keyinput_f95), .C2(
        n6949), .A(n6948), .ZN(n6962) );
  OAI22_X1 U7878 ( .A1(n5423), .A2(keyinput_f62), .B1(n6952), .B2(keyinput_f17), .ZN(n6951) );
  AOI221_X1 U7879 ( .B1(n5423), .B2(keyinput_f62), .C1(keyinput_f17), .C2(
        n6952), .A(n6951), .ZN(n6961) );
  INV_X1 U7880 ( .A(keyinput_f120), .ZN(n6954) );
  OAI22_X1 U7881 ( .A1(n6955), .A2(keyinput_f25), .B1(n6954), .B2(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6953) );
  AOI221_X1 U7882 ( .B1(n6955), .B2(keyinput_f25), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(n6954), .A(n6953), .ZN(n6960) );
  INV_X1 U7883 ( .A(keyinput_f116), .ZN(n6957) );
  OAI22_X1 U7884 ( .A1(n6958), .A2(keyinput_f13), .B1(n6957), .B2(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n6956) );
  AOI221_X1 U7885 ( .B1(n6958), .B2(keyinput_f13), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(n6957), .A(n6956), .ZN(n6959) );
  NAND4_X1 U7886 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n7011)
         );
  AOI22_X1 U7887 ( .A1(n6965), .A2(keyinput_f102), .B1(keyinput_f110), .B2(
        n6964), .ZN(n6963) );
  OAI221_X1 U7888 ( .B1(n6965), .B2(keyinput_f102), .C1(n6964), .C2(
        keyinput_f110), .A(n6963), .ZN(n6977) );
  AOI22_X1 U7889 ( .A1(n4781), .A2(keyinput_f3), .B1(keyinput_f87), .B2(n6967), 
        .ZN(n6966) );
  OAI221_X1 U7890 ( .B1(n4781), .B2(keyinput_f3), .C1(n6967), .C2(keyinput_f87), .A(n6966), .ZN(n6976) );
  AOI22_X1 U7891 ( .A1(n6970), .A2(keyinput_f91), .B1(n6969), .B2(keyinput_f65), .ZN(n6968) );
  OAI221_X1 U7892 ( .B1(n6970), .B2(keyinput_f91), .C1(n6969), .C2(
        keyinput_f65), .A(n6968), .ZN(n6975) );
  AOI22_X1 U7893 ( .A1(n6973), .A2(keyinput_f54), .B1(keyinput_f31), .B2(n6972), .ZN(n6971) );
  OAI221_X1 U7894 ( .B1(n6973), .B2(keyinput_f54), .C1(n6972), .C2(
        keyinput_f31), .A(n6971), .ZN(n6974) );
  NOR4_X1 U7895 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n7009)
         );
  INV_X1 U7896 ( .A(keyinput_f109), .ZN(n6979) );
  OAI22_X1 U7897 ( .A1(keyinput_f107), .A2(n6980), .B1(n6979), .B2(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6978) );
  AOI221_X1 U7898 ( .B1(n6980), .B2(keyinput_f107), .C1(n6979), .C2(
        DATAWIDTH_REG_5__SCAN_IN), .A(n6978), .ZN(n7008) );
  XOR2_X1 U7899 ( .A(keyinput_f121), .B(DATAWIDTH_REG_17__SCAN_IN), .Z(n6989)
         );
  XOR2_X1 U7900 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_f74), .Z(n6988) );
  AOI22_X1 U7901 ( .A1(n5395), .A2(keyinput_f56), .B1(keyinput_f93), .B2(n6982), .ZN(n6981) );
  OAI221_X1 U7902 ( .B1(n5395), .B2(keyinput_f56), .C1(n6982), .C2(
        keyinput_f93), .A(n6981), .ZN(n6987) );
  AOI22_X1 U7903 ( .A1(n6985), .A2(keyinput_f85), .B1(keyinput_f47), .B2(n6984), .ZN(n6983) );
  OAI221_X1 U7904 ( .B1(n6985), .B2(keyinput_f85), .C1(n6984), .C2(
        keyinput_f47), .A(n6983), .ZN(n6986) );
  NOR4_X1 U7905 ( .A1(n6989), .A2(n6988), .A3(n6987), .A4(n6986), .ZN(n7007)
         );
  AOI22_X1 U7906 ( .A1(n6992), .A2(keyinput_f59), .B1(keyinput_f49), .B2(n6991), .ZN(n6990) );
  OAI221_X1 U7907 ( .B1(n6992), .B2(keyinput_f59), .C1(n6991), .C2(
        keyinput_f49), .A(n6990), .ZN(n7005) );
  AOI22_X1 U7908 ( .A1(n6995), .A2(keyinput_f8), .B1(keyinput_f104), .B2(n6994), .ZN(n6993) );
  OAI221_X1 U7909 ( .B1(n6995), .B2(keyinput_f8), .C1(n6994), .C2(
        keyinput_f104), .A(n6993), .ZN(n7004) );
  AOI22_X1 U7910 ( .A1(n6998), .A2(keyinput_f84), .B1(n6997), .B2(keyinput_f28), .ZN(n6996) );
  OAI221_X1 U7911 ( .B1(n6998), .B2(keyinput_f84), .C1(n6997), .C2(
        keyinput_f28), .A(n6996), .ZN(n7003) );
  AOI22_X1 U7912 ( .A1(n7001), .A2(keyinput_f77), .B1(keyinput_f94), .B2(n7000), .ZN(n6999) );
  OAI221_X1 U7913 ( .B1(n7001), .B2(keyinput_f77), .C1(n7000), .C2(
        keyinput_f94), .A(n6999), .ZN(n7002) );
  NOR4_X1 U7914 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n7006)
         );
  NAND4_X1 U7915 ( .A1(n7009), .A2(n7008), .A3(n7007), .A4(n7006), .ZN(n7010)
         );
  NOR4_X1 U7916 ( .A1(n7013), .A2(n7012), .A3(n7011), .A4(n7010), .ZN(n7014)
         );
  NAND4_X1 U7917 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(n7019)
         );
  AOI21_X1 U7918 ( .B1(keyinput_f115), .B2(n7019), .A(n7021), .ZN(n7022) );
  INV_X1 U7919 ( .A(keyinput_f115), .ZN(n7018) );
  AOI21_X1 U7920 ( .B1(n7019), .B2(n7018), .A(keyinput_g115), .ZN(n7020) );
  AOI22_X1 U7921 ( .A1(keyinput_g115), .A2(n7022), .B1(n7021), .B2(n7020), 
        .ZN(n7023) );
  AOI21_X1 U7922 ( .B1(n7025), .B2(n7024), .A(n7023), .ZN(n7029) );
  AOI22_X1 U7923 ( .A1(n7027), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7026), .ZN(n7028) );
  XNOR2_X1 U7924 ( .A(n7029), .B(n7028), .ZN(U3445) );
  INV_X1 U3618 ( .A(n4053), .ZN(n7030) );
  INV_X2 U3640 ( .A(n7030), .ZN(n7031) );
  CLKBUF_X1 U3676 ( .A(n3150), .Z(n4053) );
  CLKBUF_X1 U3934 ( .A(n3380), .Z(n4608) );
  INV_X1 U4031 ( .A(n4524), .ZN(n5126) );
  CLKBUF_X1 U4746 ( .A(n4665), .Z(n4706) );
  CLKBUF_X1 U7925 ( .A(n5883), .Z(n5880) );
endmodule

