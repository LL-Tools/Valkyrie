

module b15_C_AntiSAT_k_256_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3187, n3189, n3190, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212;

  INV_X1 U3635 ( .A(n5599), .ZN(n4298) );
  NAND2_X1 U3636 ( .A1(n4473), .A2(n3448), .ZN(n4215) );
  INV_X4 U3637 ( .A(n4301), .ZN(n4861) );
  AND2_X1 U3638 ( .A1(n3494), .A2(n3472), .ZN(n3526) );
  INV_X1 U3639 ( .A(n3207), .ZN(n3208) );
  CLKBUF_X2 U3640 ( .A(n3361), .Z(n4596) );
  INV_X2 U3641 ( .A(n3452), .ZN(n4488) );
  CLKBUF_X2 U3642 ( .A(n3206), .Z(n3192) );
  AND2_X1 U3643 ( .A1(n4519), .A2(n4593), .ZN(n3527) );
  AND2_X1 U3644 ( .A1(n3321), .A2(n4591), .ZN(n3561) );
  CLKBUF_X1 U3645 ( .A(n3514), .Z(n3189) );
  CLKBUF_X2 U3646 ( .A(n3507), .Z(n3193) );
  AND2_X2 U3647 ( .A1(n4519), .A2(n4592), .ZN(n3205) );
  INV_X1 U3648 ( .A(n3207), .ZN(n3210) );
  NAND2_X1 U3649 ( .A1(n3502), .A2(n3501), .ZN(n3611) );
  NOR2_X1 U3650 ( .A1(n5526), .A2(n5525), .ZN(n3274) );
  NOR2_X2 U3651 ( .A1(n4883), .A2(n4884), .ZN(n6206) );
  NAND4_X2 U3652 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3452)
         );
  INV_X1 U3653 ( .A(n6198), .ZN(n6210) );
  INV_X1 U3654 ( .A(n3491), .ZN(n3463) );
  OR2_X1 U3655 ( .A1(n4877), .A2(n4791), .ZN(n4883) );
  INV_X1 U3656 ( .A(n3658), .ZN(n4145) );
  INV_X1 U3657 ( .A(n6212), .ZN(n6257) );
  XNOR2_X1 U3658 ( .A(n4300), .B(n4299), .ZN(n5785) );
  AND2_X1 U3659 ( .A1(n5727), .A2(n5728), .ZN(n3187) );
  INV_X1 U3660 ( .A(n3393), .ZN(n3475) );
  INV_X1 U3662 ( .A(n3207), .ZN(n3209) );
  INV_X1 U3663 ( .A(n3207), .ZN(n3211) );
  INV_X1 U3664 ( .A(n3540), .ZN(n3207) );
  XNOR2_X2 U3665 ( .A(n3524), .B(n3523), .ZN(n3642) );
  OAI22_X2 U3666 ( .A1(n4604), .A2(STATE2_REG_0__SCAN_IN), .B1(n4345), .B2(
        n3618), .ZN(n3524) );
  INV_X2 U3667 ( .A(n3448), .ZN(n4472) );
  NOR2_X2 U3668 ( .A1(n4471), .A2(n4543), .ZN(n4552) );
  OAI21_X2 U3670 ( .B1(n5575), .B2(n3296), .A(n5574), .ZN(n6012) );
  NAND2_X2 U3671 ( .A1(n3594), .A2(n3593), .ZN(n5108) );
  BUF_X8 U3673 ( .A(n3514), .Z(n3190) );
  AND2_X2 U3674 ( .A1(n4523), .A2(n4592), .ZN(n3514) );
  AND2_X1 U3675 ( .A1(n4519), .A2(n4592), .ZN(n3206) );
  OAI22_X1 U3676 ( .A1(n5711), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5719), .B2(n5702), .ZN(n5703) );
  AOI21_X1 U3677 ( .B1(n3247), .B2(n3244), .A(n3213), .ZN(n3243) );
  AND2_X1 U3678 ( .A1(n4686), .A2(n3710), .ZN(n4786) );
  AND2_X2 U3679 ( .A1(n4654), .A2(n3666), .ZN(n4686) );
  INV_X4 U3680 ( .A(n4396), .ZN(n3194) );
  AND2_X1 U3681 ( .A1(n4340), .A2(n4339), .ZN(n6396) );
  OR2_X1 U3682 ( .A1(n3642), .A2(n3640), .ZN(n3580) );
  NAND2_X1 U3684 ( .A1(n6285), .A2(n4651), .ZN(n6054) );
  NAND2_X1 U3685 ( .A1(n4199), .A2(n4198), .ZN(n4540) );
  AND2_X1 U3686 ( .A1(n4641), .A2(n3585), .ZN(n3420) );
  AND2_X1 U3687 ( .A1(n3573), .A2(n4691), .ZN(n4420) );
  INV_X1 U3688 ( .A(n3419), .ZN(n3573) );
  NAND2_X2 U3689 ( .A1(n3340), .A2(n3339), .ZN(n3393) );
  CLKBUF_X2 U3690 ( .A(n3433), .Z(n4123) );
  CLKBUF_X2 U3691 ( .A(n3560), .Z(n4121) );
  CLKBUF_X2 U3692 ( .A(n3527), .Z(n4128) );
  BUF_X2 U3693 ( .A(n3366), .Z(n3506) );
  CLKBUF_X2 U3694 ( .A(n3566), .Z(n4130) );
  CLKBUF_X2 U3695 ( .A(n3561), .Z(n3539) );
  CLKBUF_X2 U3696 ( .A(n3382), .Z(n4129) );
  CLKBUF_X2 U3697 ( .A(n3434), .Z(n4122) );
  INV_X1 U3698 ( .A(n3508), .ZN(n3195) );
  INV_X2 U3699 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3307) );
  INV_X2 U3700 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3604) );
  AND2_X1 U3701 ( .A1(n3306), .A2(n4430), .ZN(n3231) );
  NOR2_X1 U3702 ( .A1(n5677), .A2(n5801), .ZN(n5658) );
  AOI21_X1 U3703 ( .B1(n5656), .B2(n6400), .A(n5655), .ZN(n5657) );
  AND2_X1 U3704 ( .A1(n5566), .A2(n3217), .ZN(n5996) );
  XNOR2_X1 U3705 ( .A(n3216), .B(n4149), .ZN(n5656) );
  NAND2_X1 U3706 ( .A1(n5647), .A2(n4412), .ZN(n4413) );
  OR2_X1 U3707 ( .A1(n5680), .A2(n5564), .ZN(n6050) );
  CLKBUF_X1 U3708 ( .A(n5506), .Z(n5507) );
  OR2_X2 U3709 ( .A1(n5755), .A2(n5754), .ZN(n5740) );
  AND2_X1 U3710 ( .A1(n3285), .A2(n3286), .ZN(n5434) );
  INV_X1 U3711 ( .A(n3820), .ZN(n5376) );
  OR2_X1 U3712 ( .A1(n5468), .A2(n5467), .ZN(n5817) );
  AND2_X1 U3713 ( .A1(n5320), .A2(n3253), .ZN(n3252) );
  AND2_X1 U3714 ( .A1(n3248), .A2(n5768), .ZN(n3247) );
  NOR2_X1 U3715 ( .A1(n5569), .A2(n3269), .ZN(n5468) );
  OR2_X1 U3716 ( .A1(n3194), .A2(n6108), .ZN(n4400) );
  OR2_X1 U3717 ( .A1(n3194), .A2(n5386), .ZN(n5405) );
  NAND2_X1 U3718 ( .A1(n6388), .A2(n4352), .ZN(n4775) );
  INV_X1 U3719 ( .A(n4408), .ZN(n4396) );
  XNOR2_X1 U3720 ( .A(n4367), .B(n4873), .ZN(n4864) );
  NAND2_X1 U3721 ( .A1(n4366), .A2(n4365), .ZN(n4367) );
  NAND2_X1 U3722 ( .A1(n5497), .A2(n3228), .ZN(n5587) );
  AND2_X1 U3723 ( .A1(n4688), .A2(n4687), .ZN(n3666) );
  NOR2_X2 U3724 ( .A1(n5030), .A2(n5196), .ZN(n5986) );
  NAND2_X1 U3725 ( .A1(n4333), .A2(n4332), .ZN(n6398) );
  NAND2_X1 U3726 ( .A1(n3639), .A2(n3638), .ZN(n4688) );
  NAND2_X1 U3727 ( .A1(n4446), .A2(n4445), .ZN(n6224) );
  AND2_X1 U3728 ( .A1(n5441), .A2(n5440), .ZN(n5439) );
  CLKBUF_X1 U3729 ( .A(n4675), .Z(n4676) );
  OAI21_X1 U3730 ( .B1(n3582), .B2(n3581), .A(n3583), .ZN(n3579) );
  XNOR2_X1 U3731 ( .A(n3584), .B(n3583), .ZN(n4675) );
  OR3_X2 U3732 ( .A1(n6793), .A2(n4211), .A3(n4210), .ZN(n5548) );
  NAND2_X2 U3733 ( .A1(n4661), .A2(n4660), .ZN(n6272) );
  OAI21_X1 U3734 ( .B1(n3595), .B2(STATE2_REG_0__SCAN_IN), .A(n3591), .ZN(
        n3576) );
  NAND2_X1 U3735 ( .A1(n3559), .A2(n3558), .ZN(n3595) );
  NAND2_X1 U3736 ( .A1(n5391), .A2(n4250), .ZN(n5394) );
  AND2_X2 U3737 ( .A1(n6206), .A2(n4242), .ZN(n5391) );
  NAND2_X1 U3738 ( .A1(n3493), .A2(n4470), .ZN(n3555) );
  AND4_X1 U3739 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3493)
         );
  AND2_X1 U3740 ( .A1(n4667), .A2(n4663), .ZN(n3273) );
  NOR2_X1 U3741 ( .A1(n4462), .A2(n3461), .ZN(n4491) );
  AND2_X1 U3742 ( .A1(n4230), .A2(n4229), .ZN(n4791) );
  INV_X1 U3743 ( .A(n4477), .ZN(n6651) );
  NAND2_X1 U3744 ( .A1(n4488), .A2(n4472), .ZN(n3491) );
  NAND2_X1 U3745 ( .A1(n3618), .A2(n3617), .ZN(n4196) );
  NAND2_X1 U3746 ( .A1(n3460), .A2(n3393), .ZN(n4641) );
  INV_X1 U3747 ( .A(n3460), .ZN(n3372) );
  INV_X1 U3748 ( .A(n3460), .ZN(n4691) );
  AND4_X2 U3749 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3460)
         );
  NAND2_X1 U3750 ( .A1(n3299), .A2(n3371), .ZN(n4700) );
  NAND2_X2 U3751 ( .A1(n3218), .A2(n3381), .ZN(n3483) );
  OR2_X2 U3752 ( .A1(n3392), .A2(n3391), .ZN(n3585) );
  AND4_X1 U3753 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3418)
         );
  AND4_X1 U3754 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3446)
         );
  AND4_X1 U3755 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3447)
         );
  AND4_X1 U3756 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3416)
         );
  AND4_X1 U3757 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3330)
         );
  AND4_X1 U3758 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3359)
         );
  AND4_X1 U3759 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3340)
         );
  AND4_X1 U3760 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3360)
         );
  AND4_X1 U3761 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3444)
         );
  AND4_X1 U3762 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3445)
         );
  AND4_X1 U3763 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3327)
         );
  AND4_X1 U3764 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3328)
         );
  AND4_X1 U3765 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3329)
         );
  AND4_X1 U3766 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3381)
         );
  AND4_X1 U3767 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3371)
         );
  AND4_X1 U3768 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  AND4_X1 U3769 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3358)
         );
  AND4_X1 U3770 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3339)
         );
  AND4_X1 U3771 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3415)
         );
  AND4_X1 U3772 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3417)
         );
  OAI221_X1 U3774 ( .B1(n7009), .B2(keyinput240), .C1(n7107), .C2(keyinput217), 
        .A(n7008), .ZN(n7017) );
  NAND2_X1 U3775 ( .A1(n4523), .A2(n4593), .ZN(n3201) );
  NAND2_X1 U3776 ( .A1(n4523), .A2(n4593), .ZN(n3508) );
  AND2_X1 U3777 ( .A1(n3604), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3321)
         );
  AND2_X2 U3778 ( .A1(n3307), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4523)
         );
  NOR2_X2 U3779 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4592) );
  AND2_X2 U3780 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4593) );
  NOR2_X2 U3781 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4621) );
  CLKBUF_X1 U3782 ( .A(n6376), .Z(n3196) );
  CLKBUF_X1 U3783 ( .A(n4886), .Z(n3197) );
  INV_X1 U3784 ( .A(n4624), .ZN(n3198) );
  NAND2_X1 U3785 ( .A1(n5727), .A2(n5728), .ZN(n3199) );
  NAND2_X1 U3786 ( .A1(n4207), .A2(n4488), .ZN(n4499) );
  AOI21_X2 U3787 ( .B1(n5734), .B2(n5701), .A(n5700), .ZN(n5727) );
  OR2_X2 U3788 ( .A1(n5574), .A2(n3290), .ZN(n3217) );
  NAND2_X2 U3789 ( .A1(n5476), .A2(n3296), .ZN(n5574) );
  NAND2_X2 U3790 ( .A1(n3580), .A2(n3631), .ZN(n4673) );
  OR2_X2 U3791 ( .A1(n5667), .A2(n5692), .ZN(n5647) );
  XNOR2_X2 U3792 ( .A(n3631), .B(n3641), .ZN(n4715) );
  NAND2_X1 U3793 ( .A1(n3594), .A2(n3577), .ZN(n3583) );
  NAND2_X1 U3794 ( .A1(n3579), .A2(n3578), .ZN(n3640) );
  NAND2_X2 U3795 ( .A1(n4775), .A2(n4774), .ZN(n4773) );
  NAND2_X2 U3796 ( .A1(n5381), .A2(n5382), .ZN(n5406) );
  NAND2_X2 U3797 ( .A1(n3249), .A2(n3250), .ZN(n5381) );
  NAND2_X2 U3798 ( .A1(n3475), .A2(n3372), .ZN(n3450) );
  XNOR2_X1 U3799 ( .A(n3582), .B(n3581), .ZN(n3584) );
  AND2_X2 U3800 ( .A1(n5491), .A2(n3292), .ZN(n5476) );
  NOR2_X4 U3801 ( .A1(n5506), .A2(n5508), .ZN(n5491) );
  NOR2_X2 U3802 ( .A1(n3490), .A2(n3459), .ZN(n4207) );
  NAND2_X1 U3803 ( .A1(n3554), .A2(n3555), .ZN(n3559) );
  OAI21_X4 U3804 ( .B1(n5406), .B2(n4399), .A(n4398), .ZN(n5775) );
  AND2_X4 U3805 ( .A1(n3452), .A2(n3483), .ZN(n5599) );
  OAI211_X2 U3806 ( .C1(n3424), .C2(n3462), .A(n3398), .B(n3397), .ZN(n3490)
         );
  AND2_X2 U3807 ( .A1(n3480), .A2(n3585), .ZN(n3398) );
  AOI21_X2 U3808 ( .B1(n3490), .B2(n4472), .A(n3422), .ZN(n4419) );
  XNOR2_X1 U3809 ( .A(n3611), .B(n5099), .ZN(n4589) );
  INV_X1 U3810 ( .A(n3508), .ZN(n3202) );
  INV_X1 U3811 ( .A(n3201), .ZN(n3203) );
  INV_X1 U3812 ( .A(n3201), .ZN(n3204) );
  AND2_X1 U3813 ( .A1(n4519), .A2(n4592), .ZN(n3507) );
  XNOR2_X2 U3814 ( .A(n3526), .B(n3525), .ZN(n4512) );
  NAND2_X1 U3815 ( .A1(n4540), .A2(n6673), .ZN(n4639) );
  NAND2_X1 U3816 ( .A1(n3424), .A2(n3585), .ZN(n4462) );
  AND2_X1 U3817 ( .A1(n3293), .A2(n3294), .ZN(n3292) );
  INV_X1 U3818 ( .A(n5478), .ZN(n3293) );
  AND2_X1 U3819 ( .A1(n3259), .A2(n3258), .ZN(n3257) );
  INV_X1 U3820 ( .A(n4404), .ZN(n3258) );
  AND2_X1 U3821 ( .A1(n4298), .A2(n4215), .ZN(n4464) );
  NAND2_X1 U3822 ( .A1(n3393), .A2(n3585), .ZN(n4543) );
  INV_X1 U3823 ( .A(n3618), .ZN(n4644) );
  NAND2_X1 U3824 ( .A1(n3275), .A2(n3494), .ZN(n3504) );
  NAND4_X1 U3825 ( .A1(n3475), .A2(n3462), .A3(n3585), .A4(n3419), .ZN(n4477)
         );
  NAND2_X1 U3826 ( .A1(n3242), .A2(n3240), .ZN(n5755) );
  AND2_X1 U3827 ( .A1(n3241), .A2(n4400), .ZN(n3240) );
  INV_X1 U3828 ( .A(n6690), .ZN(n6673) );
  INV_X1 U3829 ( .A(n5108), .ZN(n5196) );
  NAND2_X1 U3830 ( .A1(n6125), .A2(n4424), .ZN(n5780) );
  NOR2_X1 U3831 ( .A1(n4188), .A2(n4187), .ZN(n4186) );
  AND2_X1 U3832 ( .A1(n3701), .A2(n3700), .ZN(n3712) );
  INV_X1 U3833 ( .A(n3667), .ZN(n3689) );
  NAND3_X1 U3834 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(n3667) );
  NAND2_X1 U3835 ( .A1(n3654), .A2(n3653), .ZN(n3688) );
  AOI21_X1 U3836 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6669), .A(n4186), 
        .ZN(n4184) );
  NAND2_X1 U3837 ( .A1(n5565), .A2(n3291), .ZN(n3290) );
  INV_X1 U3838 ( .A(n5679), .ZN(n3291) );
  AND2_X1 U3839 ( .A1(n3295), .A2(n5584), .ZN(n3294) );
  AND2_X1 U3840 ( .A1(n5588), .A2(n3974), .ZN(n3295) );
  NOR2_X1 U3841 ( .A1(n3222), .A2(n3277), .ZN(n3276) );
  INV_X1 U3842 ( .A(n5603), .ZN(n3277) );
  OR2_X1 U3843 ( .A1(n4477), .A2(n6685), .ZN(n4116) );
  NAND2_X1 U3844 ( .A1(n3804), .A2(n3803), .ZN(n3820) );
  NAND2_X1 U3845 ( .A1(n3738), .A2(n3282), .ZN(n3281) );
  INV_X1 U3846 ( .A(n5074), .ZN(n3282) );
  NOR2_X1 U3847 ( .A1(n3393), .A2(n6680), .ZN(n3845) );
  INV_X1 U3848 ( .A(n3603), .ZN(n3657) );
  AND2_X1 U3849 ( .A1(n5456), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3603) );
  INV_X1 U3850 ( .A(n5496), .ZN(n3264) );
  AND2_X1 U3851 ( .A1(n3194), .A2(n5912), .ZN(n4404) );
  AND2_X1 U3852 ( .A1(n3301), .A2(n4401), .ZN(n3259) );
  NAND2_X1 U3853 ( .A1(n5777), .A2(n5776), .ZN(n3248) );
  INV_X1 U3854 ( .A(n5321), .ZN(n3251) );
  NAND2_X1 U3855 ( .A1(n3254), .A2(n4395), .ZN(n3253) );
  INV_X1 U3856 ( .A(n5241), .ZN(n3254) );
  AND3_X1 U3857 ( .A1(n4473), .A2(n3462), .A3(n3460), .ZN(n3464) );
  NAND2_X1 U3858 ( .A1(n3562), .A2(n3261), .ZN(n4334) );
  NOR2_X1 U3859 ( .A1(n3571), .A2(n3262), .ZN(n3261) );
  OR2_X1 U3860 ( .A1(n3419), .A2(n6685), .ZN(n3618) );
  INV_X1 U3861 ( .A(n3483), .ZN(n4473) );
  INV_X1 U3862 ( .A(n4423), .ZN(n3614) );
  AND2_X1 U3863 ( .A1(n3613), .A2(n4781), .ZN(n5010) );
  AND2_X1 U3864 ( .A1(n5027), .A2(n3498), .ZN(n4720) );
  INV_X1 U3865 ( .A(n3504), .ZN(n3502) );
  OR2_X1 U3866 ( .A1(n6782), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U3867 ( .A1(n3274), .A2(n3223), .ZN(n5512) );
  AND2_X1 U3868 ( .A1(n4254), .A2(n4253), .ZN(n5262) );
  INV_X1 U3869 ( .A(n4017), .ZN(n4146) );
  NAND2_X1 U3870 ( .A1(n3289), .A2(n4421), .ZN(n3287) );
  NAND2_X1 U3871 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4060)
         );
  AND2_X1 U3872 ( .A1(n3884), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3885)
         );
  NAND2_X1 U3873 ( .A1(n4773), .A2(n3237), .ZN(n3236) );
  NAND2_X1 U3874 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3633) );
  NOR2_X2 U3875 ( .A1(n5587), .A2(n5480), .ZN(n5578) );
  INV_X1 U3876 ( .A(n3247), .ZN(n3245) );
  OAI21_X1 U3877 ( .B1(n5407), .B2(n3194), .A(n5405), .ZN(n4397) );
  CLKBUF_X1 U3878 ( .A(n4491), .Z(n4492) );
  NAND2_X1 U3879 ( .A1(n4548), .A2(n4547), .ZN(n4561) );
  OR2_X1 U3880 ( .A1(n4639), .A2(n4546), .ZN(n4547) );
  INV_X1 U3881 ( .A(n5008), .ZN(n5101) );
  NAND2_X1 U3882 ( .A1(n6685), .A2(n4677), .ZN(n5283) );
  INV_X1 U3883 ( .A(n4958), .ZN(n4953) );
  AOI22_X1 U3884 ( .A1(n3361), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3388) );
  NOR2_X1 U3885 ( .A1(n4820), .A2(n4913), .ZN(n4679) );
  NAND2_X1 U3886 ( .A1(n4444), .A2(n4302), .ZN(n6234) );
  NAND2_X1 U3887 ( .A1(n6328), .A2(n4650), .ZN(n6285) );
  AND2_X1 U3888 ( .A1(n4649), .A2(n4648), .ZN(n4650) );
  NAND2_X1 U3889 ( .A1(n5780), .A2(n4427), .ZN(n6406) );
  OR2_X1 U3890 ( .A1(n4639), .A2(n6646), .ZN(n6125) );
  NAND2_X1 U3891 ( .A1(n4438), .A2(n3271), .ZN(n4300) );
  NAND2_X1 U3892 ( .A1(n5468), .A2(n4440), .ZN(n3271) );
  OR2_X1 U3893 ( .A1(n5647), .A2(n5649), .ZN(n5650) );
  CLKBUF_X1 U3894 ( .A(n4604), .Z(n4605) );
  AND2_X1 U3895 ( .A1(n3491), .A2(n4164), .ZN(n4178) );
  AOI21_X1 U3896 ( .B1(n4161), .B2(n4158), .A(n4157), .ZN(n4188) );
  OR2_X1 U3897 ( .A1(n3699), .A2(n3698), .ZN(n4382) );
  OR2_X1 U3898 ( .A1(n3652), .A2(n3651), .ZN(n4371) );
  OR2_X1 U3899 ( .A1(n3677), .A2(n3676), .ZN(n4370) );
  NAND2_X1 U3900 ( .A1(n3449), .A2(n4513), .ZN(n3479) );
  OR2_X1 U3901 ( .A1(n3537), .A2(n3536), .ZN(n4335) );
  NAND2_X1 U3902 ( .A1(n4420), .A2(n5599), .ZN(n4513) );
  AND2_X1 U3903 ( .A1(n3632), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3322)
         );
  NOR2_X1 U3904 ( .A1(n4163), .A2(n4162), .ZN(n4183) );
  OR2_X1 U3905 ( .A1(n3448), .A2(n6685), .ZN(n3617) );
  AND2_X1 U3906 ( .A1(n3908), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3926)
         );
  INV_X1 U3907 ( .A(n3230), .ZN(n3278) );
  NOR2_X1 U3908 ( .A1(n5436), .A2(n3284), .ZN(n3283) );
  INV_X1 U3909 ( .A(n5625), .ZN(n3284) );
  INV_X1 U3910 ( .A(n5237), .ZN(n3279) );
  NAND2_X1 U3911 ( .A1(n6680), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4017) );
  XNOR2_X1 U3912 ( .A(n3680), .B(n3687), .ZN(n4361) );
  XNOR2_X1 U3913 ( .A(n3667), .B(n3688), .ZN(n4353) );
  NAND2_X1 U3914 ( .A1(n4635), .A2(n4634), .ZN(n3608) );
  INV_X1 U3915 ( .A(n3845), .ZN(n3799) );
  NAND3_X1 U3916 ( .A1(n3419), .A2(n3448), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4179) );
  OR2_X1 U3917 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  INV_X1 U3918 ( .A(n3522), .ZN(n4345) );
  AOI21_X1 U3919 ( .B1(n3612), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3500), 
        .ZN(n3503) );
  OR2_X1 U3920 ( .A1(n3628), .A2(n3627), .ZN(n4354) );
  AND2_X1 U3921 ( .A1(n4509), .A2(n4508), .ZN(n4615) );
  INV_X1 U3922 ( .A(n3495), .ZN(n3612) );
  NOR2_X1 U3923 ( .A1(n6500), .A2(n4676), .ZN(n4922) );
  INV_X1 U3924 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6658) );
  AOI22_X1 U3925 ( .A1(n3560), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U3926 ( .A1(n3189), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U3927 ( .A1(n3566), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U3928 ( .A1(n3560), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3385) );
  OAI21_X1 U3929 ( .B1(n6799), .B2(n4628), .A(n6771), .ZN(n4677) );
  OR2_X1 U3930 ( .A1(n4673), .A2(n4674), .ZN(n4820) );
  INV_X1 U3931 ( .A(n4676), .ZN(n4913) );
  NOR2_X1 U3932 ( .A1(n4179), .A2(n4379), .ZN(n4191) );
  AOI221_X1 U3933 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4184), .C1(
        n6115), .C2(n4184), .A(n4159), .ZN(n4203) );
  NAND2_X1 U3934 ( .A1(n3421), .A2(n3212), .ZN(n3422) );
  INV_X1 U3935 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6662) );
  OR2_X1 U3936 ( .A1(n4639), .A2(n4460), .ZN(n4489) );
  INV_X1 U3937 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5553) );
  OAI21_X1 U3938 ( .B1(n6002), .B2(n3658), .A(n4079), .ZN(n5679) );
  AND2_X1 U3939 ( .A1(n4003), .A2(n4002), .ZN(n5588) );
  AND2_X1 U3940 ( .A1(n4261), .A2(n4260), .ZN(n5440) );
  AND2_X1 U3941 ( .A1(n4549), .A2(n4535), .ZN(n4656) );
  INV_X1 U3942 ( .A(n3608), .ZN(n4637) );
  AOI21_X1 U3943 ( .B1(n4449), .B2(n4145), .A(n4144), .ZN(n4421) );
  AOI21_X1 U3944 ( .B1(n5993), .B2(n4145), .A(n4097), .ZN(n5565) );
  OR2_X1 U3945 ( .A1(n4060), .A2(n6018), .ZN(n4061) );
  NOR2_X1 U3946 ( .A1(n4023), .A2(n5704), .ZN(n4024) );
  OR2_X1 U3947 ( .A1(n5694), .A2(n3658), .ZN(n4042) );
  INV_X1 U3948 ( .A(n5476), .ZN(n5573) );
  OR2_X1 U3949 ( .A1(n6019), .A2(n3658), .ZN(n4022) );
  NAND2_X1 U3950 ( .A1(n3975), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3976)
         );
  OR2_X1 U3951 ( .A1(n3976), .A2(n3998), .ZN(n4023) );
  NOR2_X1 U3952 ( .A1(n3941), .A2(n3953), .ZN(n3975) );
  NAND2_X1 U3953 ( .A1(n3926), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3941)
         );
  NAND2_X1 U3954 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3907)
         );
  NOR2_X1 U3955 ( .A1(n3854), .A2(n3853), .ZN(n3884) );
  CLKBUF_X1 U3956 ( .A(n5607), .Z(n5608) );
  NAND2_X1 U3957 ( .A1(n3836), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3854)
         );
  NOR2_X1 U3958 ( .A1(n3832), .A2(n5424), .ZN(n3836) );
  NAND2_X1 U3959 ( .A1(n5376), .A2(n3821), .ZN(n5435) );
  NAND2_X1 U3960 ( .A1(n3805), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3832)
         );
  CLKBUF_X1 U3961 ( .A(n5417), .Z(n5418) );
  NOR2_X1 U3962 ( .A1(n3786), .A2(n5313), .ZN(n3805) );
  NAND2_X1 U3963 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3786)
         );
  NAND2_X1 U3964 ( .A1(n3740), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3741)
         );
  INV_X1 U3965 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7009) );
  NOR2_X1 U3966 ( .A1(n7009), .A2(n3741), .ZN(n3781) );
  AOI21_X1 U3967 ( .B1(n4145), .B2(n5324), .A(n3757), .ZN(n5074) );
  INV_X1 U3968 ( .A(n4980), .ZN(n3280) );
  NAND2_X1 U3969 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3717), .ZN(n3739)
         );
  INV_X1 U3970 ( .A(n4360), .ZN(n3238) );
  NOR2_X1 U3971 ( .A1(n5251), .A2(n3703), .ZN(n3717) );
  CLKBUF_X1 U3972 ( .A(n4786), .Z(n4787) );
  NOR2_X1 U3973 ( .A1(n3659), .A2(n5553), .ZN(n3681) );
  INV_X1 U3974 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U3975 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3634), .ZN(n3659)
         );
  OAI211_X1 U3976 ( .C1(n3657), .C2(n3604), .A(n3606), .B(n3605), .ZN(n4655)
         );
  AND2_X1 U3977 ( .A1(n3270), .A2(n5464), .ZN(n3269) );
  OR2_X1 U3978 ( .A1(n5465), .A2(n5599), .ZN(n3270) );
  NAND2_X1 U3979 ( .A1(n5647), .A2(n3224), .ZN(n5677) );
  OR2_X1 U3980 ( .A1(n3194), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5684)
         );
  INV_X1 U3981 ( .A(n5585), .ZN(n3263) );
  NAND2_X1 U3982 ( .A1(n5497), .A2(n3227), .ZN(n5592) );
  INV_X1 U3983 ( .A(n3274), .ZN(n5598) );
  NAND2_X1 U3984 ( .A1(n5740), .A2(n3257), .ZN(n3256) );
  OR2_X1 U3985 ( .A1(n3194), .A2(n4403), .ZN(n4405) );
  NAND2_X1 U3986 ( .A1(n5439), .A2(n5621), .ZN(n5623) );
  AND2_X1 U3987 ( .A1(n4259), .A2(n4258), .ZN(n5421) );
  NOR2_X1 U3988 ( .A1(n5956), .A2(n5421), .ZN(n5441) );
  INV_X1 U3989 ( .A(n5262), .ZN(n3267) );
  INV_X1 U3990 ( .A(n5394), .ZN(n3268) );
  NAND2_X1 U3991 ( .A1(n3266), .A2(n3265), .ZN(n5956) );
  INV_X1 U3992 ( .A(n5959), .ZN(n3265) );
  AND2_X1 U3993 ( .A1(n6484), .A2(n5792), .ZN(n5937) );
  AOI21_X1 U3994 ( .B1(n3252), .B2(n3255), .A(n3251), .ZN(n3250) );
  INV_X1 U3995 ( .A(n4395), .ZN(n3255) );
  NAND2_X1 U3996 ( .A1(n5242), .A2(n5241), .ZN(n5240) );
  INV_X1 U3997 ( .A(n6493), .ZN(n5906) );
  NAND2_X1 U3998 ( .A1(n4886), .A2(n4378), .ZN(n6376) );
  NAND2_X1 U3999 ( .A1(n3273), .A2(n4664), .ZN(n4879) );
  NAND2_X1 U4000 ( .A1(n4342), .A2(n7097), .ZN(n4343) );
  INV_X1 U4001 ( .A(n6398), .ZN(n4342) );
  NAND2_X1 U4002 ( .A1(n4561), .A2(n4656), .ZN(n5792) );
  AND2_X1 U4003 ( .A1(n5945), .A2(n4868), .ZN(n5935) );
  INV_X1 U4004 ( .A(n4464), .ZN(n4558) );
  OAI21_X1 U4005 ( .B1(n3495), .B2(n3308), .A(n3474), .ZN(n3554) );
  XNOR2_X1 U4006 ( .A(n4334), .B(n3260), .ZN(n3572) );
  OAI211_X1 U4007 ( .C1(n3495), .C2(n3307), .A(n3469), .B(n3468), .ZN(n3494)
         );
  AND2_X2 U4008 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4519)
         );
  OR3_X1 U4009 ( .A1(n4715), .A2(n4913), .A3(n5024), .ZN(n5030) );
  INV_X1 U4010 ( .A(n4922), .ZN(n5109) );
  OR2_X1 U4011 ( .A1(n5022), .A2(n4676), .ZN(n4899) );
  AND2_X1 U4012 ( .A1(n4894), .A2(n6567), .ZN(n4896) );
  AND3_X1 U4013 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6685), .A3(n4677), .ZN(
        n4754) );
  AOI21_X1 U4014 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6504), .A(n5283), .ZN(
        n6565) );
  INV_X1 U4015 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6669) );
  INV_X1 U4016 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6680) );
  INV_X1 U4017 ( .A(n6224), .ZN(n6251) );
  AND2_X1 U4018 ( .A1(n5654), .A2(n4448), .ZN(n6212) );
  AND2_X1 U4019 ( .A1(n5548), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6244) );
  INV_X1 U4020 ( .A(n5996), .ZN(n5636) );
  INV_X1 U4021 ( .A(n6054), .ZN(n6277) );
  AND2_X1 U4022 ( .A1(n6285), .A2(n5456), .ZN(n6276) );
  AND2_X1 U4023 ( .A1(n6285), .A2(n5457), .ZN(n6280) );
  INV_X1 U4024 ( .A(n6285), .ZN(n6279) );
  NAND2_X1 U4025 ( .A1(n6285), .A2(n4652), .ZN(n6284) );
  AND2_X1 U4026 ( .A1(n4534), .A2(n4533), .ZN(n6298) );
  CLKBUF_X1 U4027 ( .A(n4587), .Z(n6796) );
  INV_X2 U4028 ( .A(n6302), .ZN(n6308) );
  XNOR2_X1 U4029 ( .A(n5461), .B(n4421), .ZN(n5455) );
  INV_X2 U4030 ( .A(n5766), .ZN(n6400) );
  INV_X1 U4031 ( .A(n6125), .ZN(n6402) );
  NAND2_X1 U4032 ( .A1(n5740), .A2(n4401), .ZN(n5749) );
  OR2_X1 U4033 ( .A1(n5775), .A2(n3245), .ZN(n3239) );
  OR2_X1 U4034 ( .A1(n5775), .A2(n5777), .ZN(n3246) );
  INV_X1 U4035 ( .A(n6463), .ZN(n6487) );
  AND2_X1 U4036 ( .A1(n4561), .A2(n4555), .ZN(n6477) );
  INV_X1 U4037 ( .A(n6567), .ZN(n6559) );
  NAND2_X1 U4038 ( .A1(n6776), .A2(n6769), .ZN(n6782) );
  OR2_X1 U4039 ( .A1(n6500), .A2(n5138), .ZN(n6605) );
  AOI22_X1 U4040 ( .A1(n5345), .A2(n5342), .B1(n5339), .B2(n5338), .ZN(n5375)
         );
  AND2_X1 U4041 ( .A1(n5016), .A2(n5015), .ZN(n7201) );
  INV_X1 U4042 ( .A(n7210), .ZN(n5019) );
  NOR2_X1 U4043 ( .A1(n6283), .A2(n5283), .ZN(n6629) );
  OR2_X1 U4044 ( .A1(n4824), .A2(n4823), .ZN(n4852) );
  INV_X1 U4045 ( .A(n4978), .ZN(n4856) );
  INV_X1 U4046 ( .A(n6520), .ZN(n6579) );
  INV_X1 U4047 ( .A(n6526), .ZN(n6586) );
  INV_X1 U4048 ( .A(n6534), .ZN(n7200) );
  INV_X1 U4049 ( .A(n6538), .ZN(n6603) );
  INV_X1 U4050 ( .A(n6542), .ZN(n6612) );
  AND2_X1 U4051 ( .A1(n4672), .A2(n4671), .ZN(n4780) );
  NAND2_X1 U4052 ( .A1(n4679), .A2(n5196), .ZN(n4769) );
  INV_X1 U4053 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U4054 ( .A1(n6776), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6682) );
  INV_X1 U4055 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6776) );
  OR2_X1 U4056 ( .A1(n6682), .A2(n6685), .ZN(n6690) );
  AND2_X1 U4057 ( .A1(n6679), .A2(n6678), .ZN(n6766) );
  OR2_X1 U4058 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  OAI21_X1 U4059 ( .B1(n5654), .B2(n6406), .A(n5653), .ZN(n5655) );
  AND2_X2 U4060 ( .A1(n4488), .A2(n3448), .ZN(n3481) );
  AND2_X1 U4061 ( .A1(n3462), .A2(n3483), .ZN(n3212) );
  INV_X1 U4062 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3632) );
  NOR2_X1 U4063 ( .A1(n5537), .A2(n3222), .ZN(n5520) );
  NAND2_X1 U4064 ( .A1(n3280), .A2(n3738), .ZN(n4979) );
  NAND2_X1 U4065 ( .A1(n5491), .A2(n3294), .ZN(n5477) );
  AND2_X1 U4066 ( .A1(n3322), .A2(n4519), .ZN(n3560) );
  NAND2_X1 U4067 ( .A1(n5538), .A2(n3230), .ZN(n5521) );
  AND2_X1 U4068 ( .A1(n3194), .A2(n5949), .ZN(n3213) );
  AND2_X2 U4069 ( .A1(n4621), .A2(n4592), .ZN(n3439) );
  OR2_X1 U4070 ( .A1(n3585), .A2(n6680), .ZN(n3214) );
  AND3_X1 U4071 ( .A1(n3835), .A2(n3834), .A3(n3833), .ZN(n5436) );
  NAND2_X1 U4072 ( .A1(n5740), .A2(n3259), .ZN(n5708) );
  AND2_X1 U4073 ( .A1(n4367), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3215)
         );
  OR2_X1 U4074 ( .A1(n5574), .A2(n3287), .ZN(n3216) );
  AND2_X1 U4075 ( .A1(n3322), .A2(n4591), .ZN(n3361) );
  AND2_X1 U4076 ( .A1(n4592), .A2(n4591), .ZN(n3434) );
  AND2_X1 U4077 ( .A1(n5491), .A2(n3974), .ZN(n5493) );
  NOR2_X1 U4078 ( .A1(n5574), .A2(n5679), .ZN(n5564) );
  AND2_X1 U4079 ( .A1(n5491), .A2(n3295), .ZN(n5583) );
  AND4_X1 U4080 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3218)
         );
  AND2_X1 U4081 ( .A1(n3322), .A2(n4523), .ZN(n3366) );
  NAND2_X1 U4082 ( .A1(n4641), .A2(n3573), .ZN(n3423) );
  AND2_X1 U4083 ( .A1(n3322), .A2(n4621), .ZN(n3433) );
  OR2_X1 U4084 ( .A1(n5569), .A2(n5465), .ZN(n3219) );
  NAND2_X1 U4085 ( .A1(n3457), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3495) );
  OR2_X1 U4086 ( .A1(n3550), .A2(n3549), .ZN(n4389) );
  INV_X1 U4087 ( .A(n4389), .ZN(n3260) );
  AND2_X1 U4089 ( .A1(n3321), .A2(n4621), .ZN(n3566) );
  NAND2_X1 U4090 ( .A1(n3450), .A2(n3483), .ZN(n3480) );
  OAI21_X1 U4091 ( .B1(n4673), .B2(n3799), .A(n4017), .ZN(n3607) );
  NAND2_X1 U4092 ( .A1(n3194), .A2(n6108), .ZN(n3220) );
  OR2_X1 U4093 ( .A1(n5463), .A2(n4434), .ZN(n3221) );
  AND2_X1 U4094 ( .A1(n5578), .A2(n5577), .ZN(n5576) );
  NAND2_X1 U4095 ( .A1(n5611), .A2(n5612), .ZN(n5525) );
  NOR2_X1 U4096 ( .A1(n4980), .A2(n3281), .ZN(n5073) );
  AND2_X1 U4097 ( .A1(n3285), .A2(n3283), .ZN(n5616) );
  NAND2_X1 U4098 ( .A1(n5497), .A2(n5496), .ZN(n5495) );
  OR2_X1 U4099 ( .A1(n5522), .A2(n3278), .ZN(n3222) );
  AND2_X1 U4100 ( .A1(n4491), .A2(n3448), .ZN(n4200) );
  NAND2_X1 U4101 ( .A1(n5240), .A2(n4395), .ZN(n5319) );
  NAND2_X1 U4102 ( .A1(n3239), .A2(n3243), .ZN(n5761) );
  NAND2_X1 U4103 ( .A1(n3246), .A2(n5776), .ZN(n5767) );
  INV_X1 U4104 ( .A(n5776), .ZN(n3244) );
  NAND2_X1 U4105 ( .A1(n3236), .A2(n3234), .ZN(n4886) );
  XNOR2_X1 U4106 ( .A(n3820), .B(n3821), .ZN(n5416) );
  AND2_X1 U4107 ( .A1(n4273), .A2(n4272), .ZN(n3223) );
  AND2_X1 U4108 ( .A1(n4412), .A2(n5686), .ZN(n3224) );
  OR2_X1 U4109 ( .A1(n4404), .A2(n4405), .ZN(n3225) );
  INV_X1 U4110 ( .A(n3289), .ZN(n3288) );
  NOR2_X1 U4111 ( .A1(n5462), .A2(n3290), .ZN(n3289) );
  NOR2_X1 U4112 ( .A1(n5623), .A2(n5618), .ZN(n5611) );
  OR2_X1 U4113 ( .A1(n3281), .A2(n3279), .ZN(n3226) );
  OR2_X1 U4114 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3658) );
  NAND2_X1 U4115 ( .A1(n3610), .A2(n3609), .ZN(n4654) );
  NOR2_X1 U4116 ( .A1(n5590), .A2(n3264), .ZN(n3227) );
  NAND2_X1 U4117 ( .A1(n3602), .A2(n3608), .ZN(n4653) );
  NAND2_X1 U4118 ( .A1(n3268), .A2(n3267), .ZN(n5958) );
  INV_X1 U4119 ( .A(n5958), .ZN(n3266) );
  AND2_X1 U4120 ( .A1(n3227), .A2(n3263), .ZN(n3228) );
  AND2_X1 U4121 ( .A1(n3283), .A2(n5617), .ZN(n3229) );
  AND2_X2 U4122 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4591) );
  INV_X1 U4123 ( .A(n3272), .ZN(n4662) );
  NAND2_X1 U4124 ( .A1(n4664), .A2(n4663), .ZN(n3272) );
  AND2_X1 U4125 ( .A1(n3905), .A2(n3904), .ZN(n3230) );
  INV_X1 U4126 ( .A(n5436), .ZN(n3286) );
  OAI21_X1 U4127 ( .B1(n5816), .B2(n6125), .A(n3231), .ZN(U2956) );
  OAI21_X1 U4128 ( .B1(n4773), .B2(n3233), .A(n3232), .ZN(n4888) );
  AOI21_X1 U4129 ( .B1(n4864), .B2(n3238), .A(n3215), .ZN(n3232) );
  INV_X1 U4130 ( .A(n4864), .ZN(n3233) );
  INV_X1 U4131 ( .A(n3235), .ZN(n3234) );
  OAI21_X1 U4132 ( .B1(n4864), .B2(n3215), .A(n4887), .ZN(n3235) );
  NOR2_X1 U4133 ( .A1(n3215), .A2(n3238), .ZN(n3237) );
  NAND2_X1 U4134 ( .A1(n4865), .A2(n4864), .ZN(n4867) );
  NAND2_X1 U4135 ( .A1(n4773), .A2(n4360), .ZN(n4865) );
  NAND3_X1 U4136 ( .A1(n3243), .A2(n3245), .A3(n3220), .ZN(n3241) );
  NAND3_X1 U4137 ( .A1(n5775), .A2(n3243), .A3(n3220), .ZN(n3242) );
  NAND2_X1 U4138 ( .A1(n5242), .A2(n3252), .ZN(n3249) );
  NAND2_X2 U4139 ( .A1(n3256), .A2(n3225), .ZN(n5910) );
  NAND3_X1 U4140 ( .A1(n3563), .A2(n3564), .A3(n3565), .ZN(n3262) );
  NAND3_X1 U4141 ( .A1(n4664), .A2(n3273), .A3(n4228), .ZN(n4877) );
  NAND2_X1 U4142 ( .A1(n3559), .A2(n3472), .ZN(n3275) );
  NAND2_X1 U4143 ( .A1(n5538), .A2(n3276), .ZN(n5506) );
  NOR2_X1 U4144 ( .A1(n4980), .A2(n3226), .ZN(n5236) );
  NAND2_X1 U4145 ( .A1(n5417), .A2(n5435), .ZN(n3285) );
  NAND2_X1 U4146 ( .A1(n3285), .A2(n3229), .ZN(n5607) );
  INV_X1 U4147 ( .A(n5607), .ZN(n3889) );
  NOR2_X2 U4148 ( .A1(n5574), .A2(n3288), .ZN(n5461) );
  NOR2_X1 U4149 ( .A1(n5910), .A2(n5697), .ZN(n5698) );
  INV_X1 U4150 ( .A(n3423), .ZN(n3424) );
  AND2_X1 U4151 ( .A1(n4059), .A2(n4058), .ZN(n3296) );
  OR2_X1 U4152 ( .A1(n4432), .A2(n4431), .ZN(n3297) );
  NAND2_X1 U4153 ( .A1(n4327), .A2(n4326), .ZN(n4762) );
  NAND2_X1 U4154 ( .A1(n4350), .A2(n4349), .ZN(n4351) );
  OR2_X1 U4155 ( .A1(n3470), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3298)
         );
  AND4_X1 U4156 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3299)
         );
  AND2_X1 U4157 ( .A1(n3194), .A2(n5913), .ZN(n3300) );
  NAND2_X1 U4158 ( .A1(n3194), .A2(n6098), .ZN(n3301) );
  AND2_X1 U4159 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3302) );
  INV_X1 U4160 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4414) );
  AND2_X1 U4161 ( .A1(n3688), .A2(n3687), .ZN(n3303) );
  INV_X1 U4162 ( .A(n5647), .ZN(n5691) );
  INV_X1 U4163 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5313) );
  NOR2_X1 U4164 ( .A1(n5010), .A2(n5277), .ZN(n3304) );
  OR2_X1 U4165 ( .A1(n5455), .A2(n6198), .ZN(n3305) );
  OR2_X1 U4166 ( .A1(n5455), .A2(n5766), .ZN(n3306) );
  INV_X1 U4167 ( .A(n3712), .ZN(n3713) );
  INV_X1 U4168 ( .A(n4179), .ZN(n4189) );
  NAND2_X1 U4169 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6504), .ZN(n4166) );
  OAI21_X1 U4170 ( .B1(n4165), .B2(n4166), .A(n4154), .ZN(n4161) );
  NAND2_X1 U4171 ( .A1(n3212), .A2(n3460), .ZN(n3461) );
  INV_X1 U4172 ( .A(n5609), .ZN(n3888) );
  XNOR2_X1 U4173 ( .A(n4368), .B(n3715), .ZN(n4380) );
  NAND2_X1 U4174 ( .A1(n3630), .A2(n3629), .ZN(n3641) );
  AOI22_X1 U4175 ( .A1(n3189), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3369) );
  INV_X1 U4176 ( .A(n5492), .ZN(n3974) );
  INV_X1 U4177 ( .A(n4981), .ZN(n3738) );
  AND2_X1 U4178 ( .A1(n4767), .A2(n4788), .ZN(n3710) );
  INV_X1 U4179 ( .A(n4397), .ZN(n4398) );
  NAND2_X1 U4180 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  INV_X1 U4181 ( .A(n3739), .ZN(n3740) );
  OR2_X1 U4182 ( .A1(n6029), .A2(n3658), .ZN(n4003) );
  INV_X1 U4183 ( .A(n4880), .ZN(n4228) );
  NAND2_X1 U4184 ( .A1(n4368), .A2(n4391), .ZN(n4408) );
  NAND2_X1 U4185 ( .A1(n3616), .A2(n3615), .ZN(n5099) );
  OR2_X1 U4186 ( .A1(n4061), .A2(n4075), .ZN(n4098) );
  INV_X1 U4187 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5424) );
  INV_X1 U4188 ( .A(n6247), .ZN(n6217) );
  NAND2_X1 U4189 ( .A1(n5548), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5267) );
  AND3_X1 U4190 ( .A1(n3737), .A2(n3736), .A3(n3735), .ZN(n4981) );
  OR2_X1 U4191 ( .A1(n4100), .A2(n7126), .ZN(n4150) );
  NOR2_X1 U4192 ( .A1(n3907), .A2(n3906), .ZN(n3908) );
  INV_X1 U4193 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5251) );
  OR2_X1 U4194 ( .A1(n5835), .A2(n5834), .ZN(n6049) );
  AND2_X1 U4195 ( .A1(n4249), .A2(n4248), .ZN(n5389) );
  NAND2_X1 U4196 ( .A1(n4561), .A2(n4560), .ZN(n6463) );
  OR3_X1 U4197 ( .A1(n4715), .A2(n5024), .A3(n4676), .ZN(n4719) );
  INV_X1 U4198 ( .A(n4949), .ZN(n5180) );
  OR2_X1 U4199 ( .A1(n4899), .A2(n5108), .ZN(n5340) );
  OR2_X1 U4200 ( .A1(n4820), .A2(n4676), .ZN(n4958) );
  NAND2_X1 U4201 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  NAND2_X1 U4202 ( .A1(n4489), .A2(n4454), .ZN(n6793) );
  NOR2_X1 U4203 ( .A1(n5735), .A2(n6047), .ZN(n6028) );
  NOR2_X1 U4204 ( .A1(n6732), .A2(n6172), .ZN(n6163) );
  INV_X1 U4205 ( .A(n6234), .ZN(n6249) );
  XNOR2_X1 U4206 ( .A(n4153), .B(n4152), .ZN(n5654) );
  OR2_X1 U4207 ( .A1(n5267), .A2(n4308), .ZN(n6247) );
  INV_X1 U4208 ( .A(n5627), .ZN(n6259) );
  INV_X1 U4209 ( .A(n6301), .ZN(n4587) );
  INV_X1 U4210 ( .A(n6313), .ZN(n6353) );
  OR3_X1 U4211 ( .A1(n4489), .A2(n4488), .A3(READY_N), .ZN(n6328) );
  INV_X1 U4212 ( .A(n6328), .ZN(n6371) );
  INV_X1 U4213 ( .A(n6406), .ZN(n5782) );
  NAND2_X1 U4214 ( .A1(n3681), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3703)
         );
  INV_X1 U4215 ( .A(n5780), .ZN(n6395) );
  AND2_X1 U4216 ( .A1(n6455), .A2(n5385), .ZN(n6435) );
  OR2_X1 U4217 ( .A1(n5893), .A2(n6495), .ZN(n6479) );
  INV_X1 U4218 ( .A(n6461), .ZN(n6471) );
  INV_X1 U4219 ( .A(n4615), .ZN(n6655) );
  INV_X1 U4220 ( .A(n4719), .ZN(n5197) );
  OAI211_X1 U4221 ( .C1(n5035), .C2(n5034), .A(n6565), .B(n5033), .ZN(n5059)
         );
  NOR2_X1 U4222 ( .A1(n5109), .A2(n5196), .ZN(n4949) );
  OAI211_X1 U4223 ( .C1(n4918), .C2(n4917), .A(n4916), .B(n6507), .ZN(n4945)
         );
  INV_X1 U4224 ( .A(n6605), .ZN(n6618) );
  INV_X1 U4225 ( .A(n5177), .ZN(n5139) );
  INV_X1 U4226 ( .A(n5340), .ZN(n5373) );
  NAND2_X1 U4227 ( .A1(n4715), .A2(n4673), .ZN(n5022) );
  NOR2_X2 U4228 ( .A1(n4958), .A2(n5196), .ZN(n7205) );
  INV_X1 U4229 ( .A(n6623), .ZN(n6549) );
  INV_X1 U4230 ( .A(n6616), .ZN(n6547) );
  INV_X1 U4231 ( .A(n4769), .ZN(n4783) );
  NAND2_X1 U4232 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4540), .ZN(n6771) );
  OR2_X1 U4233 ( .A1(n6782), .A2(n6685), .ZN(n6689) );
  NOR2_X1 U4234 ( .A1(n4321), .A2(n4320), .ZN(n4322) );
  INV_X1 U4235 ( .A(n6244), .ZN(n6227) );
  OR2_X1 U4236 ( .A1(n5654), .A2(n4447), .ZN(n6198) );
  NAND2_X1 U4237 ( .A1(n6298), .A2(n3448), .ZN(n6287) );
  OR2_X1 U4238 ( .A1(n6298), .A2(n6796), .ZN(n6302) );
  INV_X1 U4239 ( .A(n6298), .ZN(n6310) );
  INV_X1 U4240 ( .A(n6366), .ZN(n6313) );
  OR2_X2 U4241 ( .A1(n4639), .A2(n6677), .ZN(n6373) );
  OR2_X1 U4242 ( .A1(n6695), .A2(n6559), .ZN(n5766) );
  INV_X1 U4243 ( .A(n6477), .ZN(n6489) );
  OR2_X1 U4244 ( .A1(n6782), .A2(n4208), .ZN(n6461) );
  INV_X1 U4245 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6504) );
  INV_X1 U4246 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7080) );
  INV_X1 U4247 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6115) );
  AND3_X1 U4248 ( .A1(n4718), .A2(n4717), .A3(n6503), .ZN(n4761) );
  NAND2_X1 U4249 ( .A1(n5197), .A2(n5196), .ZN(n5989) );
  NAND2_X1 U4250 ( .A1(n4914), .A2(n5196), .ZN(n5057) );
  AOI21_X1 U4251 ( .B1(n5104), .B2(n5106), .A(n5103), .ZN(n5185) );
  OR2_X1 U4252 ( .A1(n6500), .A2(n6499), .ZN(n6614) );
  OR2_X1 U4253 ( .A1(n4899), .A2(n5196), .ZN(n5177) );
  INV_X1 U4254 ( .A(n6638), .ZN(n6591) );
  OR2_X1 U4255 ( .A1(n5022), .A2(n6499), .ZN(n6642) );
  OR2_X1 U4256 ( .A1(n5022), .A2(n5138), .ZN(n7210) );
  NAND2_X1 U4257 ( .A1(n4953), .A2(n5196), .ZN(n4978) );
  INV_X1 U4258 ( .A(n6629), .ZN(n6572) );
  NAND2_X1 U4259 ( .A1(n4679), .A2(n5108), .ZN(n4859) );
  INV_X1 U4260 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6769) );
  INV_X1 U4261 ( .A(n6765), .ZN(n6762) );
  NAND2_X1 U4262 ( .A1(n3203), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3312)
         );
  INV_X1 U4263 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4264 ( .A1(n3540), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4265 ( .A1(n3193), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3310) );
  AND2_X4 U4266 ( .A1(n4621), .A2(n4593), .ZN(n3509) );
  NAND2_X1 U4267 ( .A1(n3509), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3309)
         );
  NAND2_X1 U4268 ( .A1(n3560), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4269 ( .A1(n3189), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4270 ( .A1(n3433), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4271 ( .A1(n3434), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4272 ( .A1(n3566), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4273 ( .A1(n3561), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3319)
         );
  NAND2_X1 U4274 ( .A1(n3439), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3318) );
  AND2_X4 U4275 ( .A1(n4593), .A2(n4591), .ZN(n3515) );
  NAND2_X1 U4276 ( .A1(n3515), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3317)
         );
  NAND2_X1 U4277 ( .A1(n3527), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4278 ( .A1(n3366), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4279 ( .A1(n3382), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4280 ( .A1(n3361), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4281 ( .A1(n3366), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3527), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4282 ( .A1(n3560), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4283 ( .A1(n3540), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4284 ( .A1(n3202), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4285 ( .A1(n3361), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4286 ( .A1(n3439), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3335) );
  NAND2_X1 U4287 ( .A1(n3366), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4288 ( .A1(n3527), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3343)
         );
  NAND2_X1 U4289 ( .A1(n3204), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4290 ( .A1(n3509), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4291 ( .A1(n3382), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4292 ( .A1(n3540), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3347)
         );
  NAND2_X1 U4293 ( .A1(n3560), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4294 ( .A1(n3193), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4295 ( .A1(n3361), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4296 ( .A1(n3189), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4297 ( .A1(n3433), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4298 ( .A1(n3434), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4299 ( .A1(n3566), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4300 ( .A1(n3561), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3355)
         );
  NAND2_X1 U4301 ( .A1(n3439), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4302 ( .A1(n3515), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3353)
         );
  NAND4_X2 U4303 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3419)
         );
  AOI22_X1 U4304 ( .A1(n3540), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4305 ( .A1(n3204), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3527), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4306 ( .A1(n3361), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4307 ( .A1(n3566), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4308 ( .A1(n3366), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4309 ( .A1(n3561), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4310 ( .A1(n3560), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3367) );
  INV_X2 U4311 ( .A(n4700), .ZN(n3462) );
  AOI22_X1 U4312 ( .A1(n3366), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3527), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4313 ( .A1(n3540), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4314 ( .A1(n3203), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4315 ( .A1(n3190), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4316 ( .A1(n3566), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4317 ( .A1(n3361), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4318 ( .A1(n3439), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4319 ( .A1(n3366), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3527), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4320 ( .A1(n3540), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4321 ( .A1(n3204), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3383) );
  NAND4_X1 U4322 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3392)
         );
  AOI22_X1 U4323 ( .A1(n3190), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4324 ( .A1(n3566), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4325 ( .A1(n3439), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4326 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3391)
         );
  NAND2_X1 U4327 ( .A1(n3423), .A2(n3475), .ZN(n3396) );
  NAND2_X1 U4328 ( .A1(n3462), .A2(n4641), .ZN(n3394) );
  NAND2_X1 U4329 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  NAND2_X1 U4330 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  NAND2_X1 U4331 ( .A1(n3366), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4332 ( .A1(n3560), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3401) );
  NAND2_X1 U4333 ( .A1(n3540), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3400)
         );
  NAND2_X1 U4334 ( .A1(n3205), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4335 ( .A1(n3433), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3406) );
  NAND2_X1 U4336 ( .A1(n3361), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3405) );
  NAND2_X1 U4337 ( .A1(n3566), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4338 ( .A1(n3439), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4339 ( .A1(n3527), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3410)
         );
  NAND2_X1 U4340 ( .A1(n3382), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4341 ( .A1(n3202), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3408)
         );
  NAND2_X1 U4342 ( .A1(n3509), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3407)
         );
  NAND2_X1 U4343 ( .A1(n3189), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4344 ( .A1(n3561), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3413)
         );
  NAND2_X1 U4345 ( .A1(n3434), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3412) );
  NAND2_X1 U4346 ( .A1(n3515), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3411)
         );
  NAND4_X4 U4347 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3448)
         );
  OAI21_X1 U4348 ( .B1(n3419), .B2(n3450), .A(n3420), .ZN(n3482) );
  INV_X1 U4349 ( .A(n3482), .ZN(n3421) );
  NAND2_X1 U4350 ( .A1(n3527), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3428)
         );
  NAND2_X1 U4351 ( .A1(n3366), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U4352 ( .A1(n3202), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3426)
         );
  NAND2_X1 U4353 ( .A1(n3509), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3425)
         );
  NAND2_X1 U4354 ( .A1(n3540), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3432)
         );
  NAND2_X1 U4355 ( .A1(n3382), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3431) );
  NAND2_X1 U4356 ( .A1(n3560), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4357 ( .A1(n3192), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3429) );
  NAND2_X1 U4358 ( .A1(n3361), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U4359 ( .A1(n3190), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3437) );
  NAND2_X1 U4360 ( .A1(n3433), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4361 ( .A1(n3434), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4362 ( .A1(n3566), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4363 ( .A1(n3561), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3442)
         );
  NAND2_X1 U4364 ( .A1(n3439), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U4365 ( .A1(n3515), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3440)
         );
  NAND2_X1 U4366 ( .A1(n4462), .A2(n3481), .ZN(n3449) );
  INV_X1 U4367 ( .A(n4420), .ZN(n3451) );
  NAND2_X1 U4368 ( .A1(n3451), .A2(n3450), .ZN(n3454) );
  NAND2_X1 U4369 ( .A1(n4472), .A2(n3452), .ZN(n5266) );
  XNOR2_X1 U4370 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4303) );
  NAND2_X1 U4371 ( .A1(n4488), .A2(n4303), .ZN(n3465) );
  INV_X1 U4372 ( .A(n3465), .ZN(n3453) );
  AOI21_X1 U4373 ( .B1(n3454), .B2(n5266), .A(n3453), .ZN(n3455) );
  NOR2_X1 U4374 ( .A1(n3479), .A2(n3455), .ZN(n3456) );
  NAND2_X1 U4375 ( .A1(n4419), .A2(n3456), .ZN(n3457) );
  XNOR2_X1 U4376 ( .A(n6504), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5277)
         );
  AND2_X1 U4377 ( .A1(n6682), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3458)
         );
  AOI21_X1 U4378 ( .B1(n3614), .B2(n5277), .A(n3458), .ZN(n3469) );
  NAND2_X1 U4379 ( .A1(n4420), .A2(n4472), .ZN(n3459) );
  AOI21_X1 U4380 ( .B1(n4200), .B2(n3465), .A(n4552), .ZN(n3466) );
  NAND2_X1 U4381 ( .A1(n4499), .A2(n3466), .ZN(n3467) );
  NAND2_X1 U4382 ( .A1(n3467), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3468) );
  INV_X1 U4383 ( .A(n3468), .ZN(n3471) );
  INV_X1 U4384 ( .A(n3469), .ZN(n3470) );
  NAND2_X1 U4385 ( .A1(n3471), .A2(n3298), .ZN(n3472) );
  MUX2_X1 U4386 ( .A(n6682), .B(n3614), .S(n6504), .Z(n3473) );
  INV_X1 U4387 ( .A(n3473), .ZN(n3474) );
  NAND2_X1 U4388 ( .A1(n6651), .A2(n4473), .ZN(n3476) );
  NAND2_X1 U4389 ( .A1(n3476), .A2(n4472), .ZN(n3478) );
  NAND2_X1 U4390 ( .A1(n3448), .A2(n3462), .ZN(n3477) );
  NAND2_X1 U4391 ( .A1(n3478), .A2(n3477), .ZN(n3489) );
  INV_X1 U4392 ( .A(n3479), .ZN(n3488) );
  AOI21_X1 U4393 ( .B1(n3480), .B2(n3481), .A(n6689), .ZN(n3487) );
  NAND2_X1 U4394 ( .A1(n3450), .A2(n3419), .ZN(n3484) );
  NAND2_X1 U4395 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  OAI21_X1 U4396 ( .B1(n3482), .B2(n3485), .A(n3452), .ZN(n3486) );
  NOR2_X1 U4397 ( .A1(n4420), .A2(n5266), .ZN(n3492) );
  AOI21_X1 U4398 ( .B1(n3490), .B2(n3463), .A(n3492), .ZN(n4470) );
  AND2_X1 U4399 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4400 ( .A1(n3496), .A2(n6662), .ZN(n5027) );
  INV_X1 U4401 ( .A(n3496), .ZN(n3497) );
  NAND2_X1 U4402 ( .A1(n3497), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3498) );
  INV_X1 U4403 ( .A(n6682), .ZN(n3499) );
  OAI22_X1 U4404 ( .A1(n4720), .A2(n4423), .B1(n3499), .B2(n6662), .ZN(n3500)
         );
  INV_X1 U4405 ( .A(n3503), .ZN(n3501) );
  NAND2_X1 U4406 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND2_X1 U4407 ( .A1(n3611), .A2(n3505), .ZN(n4604) );
  AOI22_X1 U4408 ( .A1(n3506), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4409 ( .A1(n4121), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4410 ( .A1(n3208), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4411 ( .A1(n3195), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4412 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3521)
         );
  AOI22_X1 U4413 ( .A1(n3190), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4414 ( .A1(n4130), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4415 ( .A1(n4596), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4416 ( .A1(n3439), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4417 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3520)
         );
  INV_X1 U4418 ( .A(n3617), .ZN(n3551) );
  AOI22_X1 U4419 ( .A1(n4189), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3551), 
        .B2(n3522), .ZN(n3523) );
  INV_X1 U4420 ( .A(n3559), .ZN(n3525) );
  AOI22_X1 U4421 ( .A1(n3506), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4422 ( .A1(n4121), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4423 ( .A1(n3210), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4424 ( .A1(n3195), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3528) );
  NAND4_X1 U4425 ( .A1(n3531), .A2(n3530), .A3(n3529), .A4(n3528), .ZN(n3537)
         );
  AOI22_X1 U4426 ( .A1(n3190), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4427 ( .A1(n4130), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4428 ( .A1(n4596), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4429 ( .A1(n3439), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4430 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  NAND2_X1 U4431 ( .A1(n4644), .A2(n4335), .ZN(n3538) );
  OAI21_X2 U4432 ( .B1(n4512), .B2(STATE2_REG_0__SCAN_IN), .A(n3538), .ZN(
        n3582) );
  INV_X1 U4433 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U4434 ( .A1(n3506), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4435 ( .A1(n4121), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4436 ( .A1(n4123), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4437 ( .A1(n3209), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4438 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3550)
         );
  AOI22_X1 U4439 ( .A1(n3195), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4440 ( .A1(n3190), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4441 ( .A1(n4596), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4442 ( .A1(n3439), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3545) );
  NAND4_X1 U4443 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3549)
         );
  NAND2_X1 U4444 ( .A1(n4644), .A2(n3260), .ZN(n3553) );
  NAND2_X1 U4445 ( .A1(n3551), .A2(n4335), .ZN(n3552) );
  OAI211_X1 U4446 ( .C1(n4179), .C2(n4739), .A(n3553), .B(n3552), .ZN(n3581)
         );
  INV_X1 U4447 ( .A(n3554), .ZN(n3557) );
  INV_X1 U4448 ( .A(n3555), .ZN(n3556) );
  AOI22_X1 U4449 ( .A1(n3211), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4450 ( .A1(n3382), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4451 ( .A1(n3506), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4452 ( .A1(n3539), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4453 ( .A1(n3204), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4454 ( .A1(n4123), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4455 ( .A1(n3205), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4456 ( .A1(n3566), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4457 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  NAND2_X1 U4458 ( .A1(n3572), .A2(n4644), .ZN(n3591) );
  INV_X1 U4459 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4752) );
  AOI21_X1 U4460 ( .B1(n3573), .B2(n4389), .A(n6685), .ZN(n3575) );
  NAND2_X1 U4461 ( .A1(n4472), .A2(n4334), .ZN(n3574) );
  OAI211_X1 U4462 ( .C1(n4179), .C2(n4752), .A(n3575), .B(n3574), .ZN(n3590)
         );
  NAND2_X1 U4463 ( .A1(n3576), .A2(n3590), .ZN(n3594) );
  NAND2_X1 U4464 ( .A1(n4644), .A2(n4389), .ZN(n3577) );
  NAND2_X1 U4465 ( .A1(n3582), .A2(n3581), .ZN(n3578) );
  NAND2_X2 U4466 ( .A1(n3642), .A2(n3640), .ZN(n3631) );
  INV_X1 U4467 ( .A(n3607), .ZN(n3602) );
  NAND2_X1 U4468 ( .A1(n4675), .A2(n3845), .ZN(n3589) );
  INV_X2 U4469 ( .A(n3214), .ZN(n4147) );
  AOI22_X1 U4470 ( .A1(n4147), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6680), .ZN(n3587) );
  INV_X1 U4471 ( .A(n4543), .ZN(n5456) );
  NAND2_X1 U4472 ( .A1(n3603), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3586) );
  AND2_X1 U4473 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  NAND2_X1 U4474 ( .A1(n3589), .A2(n3588), .ZN(n4635) );
  INV_X1 U4475 ( .A(n3590), .ZN(n3592) );
  AOI21_X1 U4476 ( .B1(n5108), .B2(n3475), .A(n6680), .ZN(n4567) );
  OR2_X1 U4477 ( .A1(n3595), .A2(n3799), .ZN(n3599) );
  AOI22_X1 U4478 ( .A1(n4147), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6680), .ZN(n3597) );
  NAND2_X1 U4479 ( .A1(n3603), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3596) );
  AND2_X1 U4480 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  NAND2_X1 U4481 ( .A1(n3599), .A2(n3598), .ZN(n4566) );
  NAND2_X1 U4482 ( .A1(n4567), .A2(n4566), .ZN(n4565) );
  INV_X1 U4483 ( .A(n4566), .ZN(n3600) );
  NAND2_X1 U4484 ( .A1(n3600), .A2(n4145), .ZN(n3601) );
  NAND2_X1 U4485 ( .A1(n4565), .A2(n3601), .ZN(n4634) );
  OAI21_X1 U4486 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3633), .ZN(n6405) );
  AOI22_X1 U4487 ( .A1(n4145), .A2(n6405), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4488 ( .A1(n4147), .A2(EAX_REG_2__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4489 ( .A1(n4653), .A2(n4655), .ZN(n3610) );
  NAND2_X1 U4490 ( .A1(n3607), .A2(n4637), .ZN(n3609) );
  NAND2_X1 U4491 ( .A1(n3612), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3616) );
  NOR3_X1 U4492 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6662), .A3(n6658), 
        .ZN(n6568) );
  NAND2_X1 U4493 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6568), .ZN(n6615) );
  NAND2_X1 U4494 ( .A1(n6669), .A2(n6615), .ZN(n3613) );
  NAND3_X1 U4495 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4822) );
  INV_X1 U4496 ( .A(n4822), .ZN(n4683) );
  NAND2_X1 U4497 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4683), .ZN(n4781) );
  AOI22_X1 U4498 ( .A1(n3614), .A2(n5010), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6682), .ZN(n3615) );
  NAND2_X1 U4499 ( .A1(n4589), .A2(n6685), .ZN(n3630) );
  AOI22_X1 U4500 ( .A1(n3506), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4501 ( .A1(n4121), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4502 ( .A1(n3208), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4503 ( .A1(n3195), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4504 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3628)
         );
  AOI22_X1 U4505 ( .A1(n3190), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4506 ( .A1(n4130), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4507 ( .A1(n4596), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4508 ( .A1(n3727), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4509 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  AOI22_X1 U4510 ( .A1(n4189), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4196), 
        .B2(n4354), .ZN(n3629) );
  NAND2_X1 U4511 ( .A1(n4715), .A2(n3845), .ZN(n3639) );
  OAI21_X1 U4512 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3634), .A(n3659), 
        .ZN(n6394) );
  AOI22_X1 U4513 ( .A1(n4145), .A2(n6394), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4514 ( .A1(n4147), .A2(EAX_REG_3__SCAN_IN), .ZN(n3635) );
  OAI211_X1 U4515 ( .C1(n3657), .C2(n3632), .A(n3636), .B(n3635), .ZN(n3637)
         );
  INV_X1 U4516 ( .A(n3637), .ZN(n3638) );
  AOI22_X1 U4517 ( .A1(n3506), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4518 ( .A1(n4121), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4519 ( .A1(n3208), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4520 ( .A1(n3195), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4521 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3652)
         );
  AOI22_X1 U4522 ( .A1(n3190), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4523 ( .A1(n4130), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4524 ( .A1(n4596), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4525 ( .A1(n3727), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4526 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3651)
         );
  NAND2_X1 U4527 ( .A1(n4196), .A2(n4371), .ZN(n3654) );
  INV_X1 U4528 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4743) );
  OR2_X1 U4529 ( .A1(n4179), .A2(n4743), .ZN(n3653) );
  NAND2_X1 U4530 ( .A1(n4353), .A2(n3845), .ZN(n3665) );
  NAND2_X1 U4531 ( .A1(n6680), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3656)
         );
  NAND2_X1 U4532 ( .A1(n4147), .A2(EAX_REG_4__SCAN_IN), .ZN(n3655) );
  OAI211_X1 U4533 ( .C1(n3657), .C2(n6115), .A(n3656), .B(n3655), .ZN(n3663)
         );
  INV_X1 U4534 ( .A(n3659), .ZN(n3661) );
  INV_X1 U4535 ( .A(n3681), .ZN(n3660) );
  OAI21_X1 U4536 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3661), .A(n3660), 
        .ZN(n5555) );
  AND2_X1 U4537 ( .A1(n4145), .A2(n5555), .ZN(n3662) );
  AOI21_X1 U4538 ( .B1(n3663), .B2(n3658), .A(n3662), .ZN(n3664) );
  NAND2_X1 U4539 ( .A1(n3665), .A2(n3664), .ZN(n4687) );
  NAND2_X1 U4540 ( .A1(n3689), .A2(n3688), .ZN(n3680) );
  AOI22_X1 U4541 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n3506), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4542 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4129), .B1(n4121), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3670) );
  INV_X1 U4543 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n7028) );
  AOI22_X1 U4544 ( .A1(n3208), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4545 ( .A1(n3195), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4546 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3677)
         );
  AOI22_X1 U4547 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n3190), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4548 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3539), .B1(n4130), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4549 ( .A1(n4596), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4550 ( .A1(n3439), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3672) );
  NAND4_X1 U4551 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3676)
         );
  NAND2_X1 U4552 ( .A1(n4196), .A2(n4370), .ZN(n3679) );
  INV_X1 U4553 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4748) );
  OR2_X1 U4554 ( .A1(n4179), .A2(n4748), .ZN(n3678) );
  NAND2_X1 U4555 ( .A1(n3679), .A2(n3678), .ZN(n3687) );
  NAND2_X1 U4556 ( .A1(n4361), .A2(n3845), .ZN(n3686) );
  INV_X1 U4557 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3683) );
  OAI21_X1 U4558 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3681), .A(n3703), 
        .ZN(n6386) );
  NAND2_X1 U4559 ( .A1(n6386), .A2(n4145), .ZN(n3682) );
  OAI21_X1 U4560 ( .B1(n3683), .B2(n4017), .A(n3682), .ZN(n3684) );
  AOI21_X1 U4561 ( .B1(n4147), .B2(EAX_REG_5__SCAN_IN), .A(n3684), .ZN(n3685)
         );
  NAND2_X1 U4562 ( .A1(n3686), .A2(n3685), .ZN(n4767) );
  NAND2_X1 U4563 ( .A1(n3689), .A2(n3303), .ZN(n3711) );
  NAND2_X1 U4564 ( .A1(n4189), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4565 ( .A1(n3506), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4566 ( .A1(n4121), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4567 ( .A1(n3208), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4568 ( .A1(n3195), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3690) );
  NAND4_X1 U4569 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3699)
         );
  AOI22_X1 U4570 ( .A1(n3190), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4571 ( .A1(n4130), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4572 ( .A1(n4596), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4573 ( .A1(n3727), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4574 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3698)
         );
  NAND2_X1 U4575 ( .A1(n4196), .A2(n4382), .ZN(n3700) );
  NAND2_X1 U4576 ( .A1(n3711), .A2(n3712), .ZN(n4369) );
  NAND2_X1 U4577 ( .A1(n4369), .A2(n3845), .ZN(n3709) );
  INV_X1 U4578 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3702) );
  OAI22_X1 U4579 ( .A1(n3214), .A2(n3702), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5251), .ZN(n3707) );
  INV_X1 U4580 ( .A(n3703), .ZN(n3705) );
  INV_X1 U4581 ( .A(n3717), .ZN(n3704) );
  OAI21_X1 U4582 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3705), .A(n3704), 
        .ZN(n5255) );
  AND2_X1 U4583 ( .A1(n4145), .A2(n5255), .ZN(n3706) );
  AOI21_X1 U4584 ( .B1(n3707), .B2(n3658), .A(n3706), .ZN(n3708) );
  NAND2_X1 U4585 ( .A1(n3709), .A2(n3708), .ZN(n4788) );
  INV_X1 U4586 ( .A(n3711), .ZN(n3714) );
  NAND2_X1 U4587 ( .A1(n3714), .A2(n3713), .ZN(n4368) );
  AOI22_X1 U4588 ( .A1(n4189), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4196), 
        .B2(n4389), .ZN(n3715) );
  INV_X1 U4589 ( .A(n4380), .ZN(n3716) );
  NAND2_X1 U4590 ( .A1(n3716), .A2(n3845), .ZN(n3722) );
  INV_X1 U4591 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3719) );
  OAI21_X1 U4592 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3717), .A(n3739), 
        .ZN(n6381) );
  NAND2_X1 U4593 ( .A1(n6381), .A2(n4145), .ZN(n3718) );
  OAI21_X1 U4594 ( .B1(n4017), .B2(n3719), .A(n3718), .ZN(n3720) );
  AOI21_X1 U4595 ( .B1(n4147), .B2(EAX_REG_7__SCAN_IN), .A(n3720), .ZN(n3721)
         );
  NAND2_X1 U4596 ( .A1(n3722), .A2(n3721), .ZN(n5003) );
  NAND2_X1 U4597 ( .A1(n4786), .A2(n5003), .ZN(n4980) );
  AOI22_X1 U4598 ( .A1(n3203), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4599 ( .A1(n3208), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4600 ( .A1(n3190), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4601 ( .A1(n4596), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4602 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3733)
         );
  AOI22_X1 U4603 ( .A1(n4129), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4604 ( .A1(n4123), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4605 ( .A1(n3506), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4606 ( .A1(n3727), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3728) );
  NAND4_X1 U4607 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3732)
         );
  OAI21_X1 U4608 ( .B1(n3733), .B2(n3732), .A(n3845), .ZN(n3737) );
  XNOR2_X1 U4609 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3739), .ZN(n5247) );
  INV_X1 U4610 ( .A(n5247), .ZN(n3734) );
  AOI22_X1 U4611 ( .A1(n4146), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4145), 
        .B2(n3734), .ZN(n3736) );
  NAND2_X1 U4612 ( .A1(n4147), .A2(EAX_REG_8__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4613 ( .A1(n3741), .A2(n7009), .ZN(n3743) );
  INV_X1 U4614 ( .A(n3781), .ZN(n3742) );
  NAND2_X1 U4615 ( .A1(n3743), .A2(n3742), .ZN(n5324) );
  AOI22_X1 U4616 ( .A1(n3202), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4617 ( .A1(n3208), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4618 ( .A1(n4596), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4619 ( .A1(n4130), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4620 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4621 ( .A1(n4121), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4622 ( .A1(n3506), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4623 ( .A1(n3190), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4624 ( .A1(n4123), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4625 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OAI21_X1 U4626 ( .B1(n3753), .B2(n3752), .A(n3845), .ZN(n3756) );
  NAND2_X1 U4627 ( .A1(n4147), .A2(EAX_REG_9__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4628 ( .A1(n4146), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3754)
         );
  NAND3_X1 U4629 ( .A1(n3756), .A2(n3755), .A3(n3754), .ZN(n3757) );
  AOI22_X1 U4630 ( .A1(n3205), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4631 ( .A1(n3208), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4632 ( .A1(n3190), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4633 ( .A1(n4596), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4634 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3767)
         );
  AOI22_X1 U4635 ( .A1(n4121), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4636 ( .A1(n4123), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4637 ( .A1(n3506), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4638 ( .A1(n3727), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3762) );
  NAND4_X1 U4639 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3766)
         );
  NOR2_X1 U4640 ( .A1(n3767), .A2(n3766), .ZN(n3770) );
  XOR2_X1 U4641 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3781), .Z(n6192) );
  INV_X1 U4642 ( .A(n6192), .ZN(n5400) );
  AOI22_X1 U4643 ( .A1(n4146), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n4145), 
        .B2(n5400), .ZN(n3769) );
  NAND2_X1 U4644 ( .A1(n4147), .A2(EAX_REG_10__SCAN_IN), .ZN(n3768) );
  OAI211_X1 U4645 ( .C1(n3799), .C2(n3770), .A(n3769), .B(n3768), .ZN(n5237)
         );
  AOI22_X1 U4646 ( .A1(n3208), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4647 ( .A1(n3204), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4648 ( .A1(n3190), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4649 ( .A1(n4130), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4650 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3780)
         );
  AOI22_X1 U4651 ( .A1(n4121), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4652 ( .A1(n4123), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4653 ( .A1(n3506), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4654 ( .A1(n3539), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4655 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4656 ( .A1(n3780), .A2(n3779), .ZN(n3785) );
  INV_X1 U4657 ( .A(n3786), .ZN(n3782) );
  XNOR2_X1 U4658 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3782), .ZN(n5410)
         );
  AOI22_X1 U4659 ( .A1(n4145), .A2(n5410), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4660 ( .A1(n4147), .A2(EAX_REG_11__SCAN_IN), .ZN(n3783) );
  OAI211_X1 U4661 ( .C1(n3799), .C2(n3785), .A(n3784), .B(n3783), .ZN(n5259)
         );
  NAND2_X1 U4662 ( .A1(n5236), .A2(n5259), .ZN(n5258) );
  INV_X1 U4663 ( .A(n5258), .ZN(n3804) );
  XOR2_X1 U4664 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3805), .Z(n6187) );
  NAND2_X1 U4665 ( .A1(n6187), .A2(n4145), .ZN(n3802) );
  INV_X1 U4666 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5379) );
  INV_X1 U4667 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6124) );
  OAI21_X1 U4668 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6124), .A(n6680), 
        .ZN(n3787) );
  OAI21_X1 U4669 ( .B1(n3214), .B2(n5379), .A(n3787), .ZN(n3801) );
  AOI22_X1 U4670 ( .A1(n3208), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4671 ( .A1(n3190), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4672 ( .A1(n4129), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4673 ( .A1(n3539), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4674 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4675 ( .A1(n3203), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4676 ( .A1(n4121), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4677 ( .A1(n4128), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4678 ( .A1(n4130), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4679 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  NOR2_X1 U4680 ( .A1(n3797), .A2(n3796), .ZN(n3798) );
  NOR2_X1 U4681 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  AOI21_X1 U4682 ( .B1(n3802), .B2(n3801), .A(n3800), .ZN(n5377) );
  INV_X1 U4683 ( .A(n5377), .ZN(n3803) );
  XNOR2_X1 U4684 ( .A(n3832), .B(n5424), .ZN(n5771) );
  NAND2_X1 U4685 ( .A1(n5771), .A2(n4145), .ZN(n3808) );
  NOR2_X1 U4686 ( .A1(n4017), .A2(n5424), .ZN(n3806) );
  AOI21_X1 U4687 ( .B1(n4147), .B2(EAX_REG_13__SCAN_IN), .A(n3806), .ZN(n3807)
         );
  NAND2_X1 U4688 ( .A1(n3808), .A2(n3807), .ZN(n3821) );
  AOI22_X1 U4689 ( .A1(n4121), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4690 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3208), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4691 ( .A1(n3195), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4692 ( .A1(n3192), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4693 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3818)
         );
  AOI22_X1 U4694 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n4123), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4695 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n3190), .B1(n4596), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4696 ( .A1(n4129), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4697 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4130), .B1(n3727), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4698 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3817)
         );
  OR2_X1 U4699 ( .A1(n3818), .A2(n3817), .ZN(n3819) );
  AND2_X1 U4700 ( .A1(n3845), .A2(n3819), .ZN(n5419) );
  NAND2_X1 U4701 ( .A1(n5416), .A2(n5419), .ZN(n5417) );
  AOI22_X1 U4702 ( .A1(n3190), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4703 ( .A1(n3210), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4704 ( .A1(n4129), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4705 ( .A1(n3727), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3822) );
  NAND4_X1 U4706 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3831)
         );
  AOI22_X1 U4707 ( .A1(n3506), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4708 ( .A1(n3195), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4709 ( .A1(n4121), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4710 ( .A1(n4130), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4711 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3830)
         );
  OAI21_X1 U4712 ( .B1(n3831), .B2(n3830), .A(n3845), .ZN(n3835) );
  XNOR2_X1 U4713 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3836), .ZN(n6179)
         );
  AOI22_X1 U4714 ( .A1(n4145), .A2(n6179), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4715 ( .A1(n4147), .A2(EAX_REG_14__SCAN_IN), .ZN(n3833) );
  XOR2_X1 U4716 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3854), .Z(n6166) );
  NAND2_X1 U4717 ( .A1(n6166), .A2(n4145), .ZN(n3852) );
  AOI22_X1 U4718 ( .A1(n3506), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4719 ( .A1(n3208), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4720 ( .A1(n4129), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4721 ( .A1(n4123), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4722 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3847)
         );
  AOI22_X1 U4723 ( .A1(n4121), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4724 ( .A1(n3190), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4725 ( .A1(n3205), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4726 ( .A1(n4130), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4727 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3846)
         );
  OAI21_X1 U4728 ( .B1(n3847), .B2(n3846), .A(n3845), .ZN(n3850) );
  NAND2_X1 U4729 ( .A1(n4147), .A2(EAX_REG_15__SCAN_IN), .ZN(n3849) );
  NAND2_X1 U4730 ( .A1(n4146), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3848)
         );
  AND3_X1 U4731 ( .A1(n3850), .A2(n3849), .A3(n3848), .ZN(n3851) );
  NAND2_X1 U4732 ( .A1(n3852), .A2(n3851), .ZN(n5625) );
  INV_X1 U4733 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3853) );
  XNOR2_X1 U4734 ( .A(n3884), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6151)
         );
  NAND2_X1 U4735 ( .A1(n6151), .A2(n4145), .ZN(n3869) );
  AOI22_X1 U4736 ( .A1(n3195), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4737 ( .A1(n4121), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4738 ( .A1(n3190), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4739 ( .A1(n3506), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4740 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3864)
         );
  AOI22_X1 U4741 ( .A1(n3210), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4742 ( .A1(n4596), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4743 ( .A1(n4129), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4744 ( .A1(n3727), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4745 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  NOR2_X1 U4746 ( .A1(n3864), .A2(n3863), .ZN(n3866) );
  AOI22_X1 U4747 ( .A1(n4147), .A2(EAX_REG_16__SCAN_IN), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3865) );
  OAI21_X1 U4748 ( .B1(n4116), .B2(n3866), .A(n3865), .ZN(n3867) );
  INV_X1 U4749 ( .A(n3867), .ZN(n3868) );
  NAND2_X1 U4750 ( .A1(n3869), .A2(n3868), .ZN(n5617) );
  AOI22_X1 U4751 ( .A1(n3208), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4752 ( .A1(n4121), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4753 ( .A1(n3190), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4754 ( .A1(n4130), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4755 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4756 ( .A1(n3506), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4757 ( .A1(n3205), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4758 ( .A1(n4129), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4759 ( .A1(n4123), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4760 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  NOR2_X1 U4761 ( .A1(n3879), .A2(n3878), .ZN(n3883) );
  OAI21_X1 U4762 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6124), .A(n6680), 
        .ZN(n3880) );
  INV_X1 U4763 ( .A(n3880), .ZN(n3881) );
  AOI21_X1 U4764 ( .B1(n4147), .B2(EAX_REG_17__SCAN_IN), .A(n3881), .ZN(n3882)
         );
  OAI21_X1 U4765 ( .B1(n4116), .B2(n3883), .A(n3882), .ZN(n3887) );
  OAI21_X1 U4766 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3885), .A(n3907), 
        .ZN(n6142) );
  OR2_X1 U4767 ( .A1(n3658), .A2(n6142), .ZN(n3886) );
  NAND2_X1 U4768 ( .A1(n3887), .A2(n3886), .ZN(n5609) );
  NAND2_X1 U4769 ( .A1(n3889), .A2(n3888), .ZN(n5537) );
  AOI22_X1 U4770 ( .A1(n3506), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4771 ( .A1(n4121), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4772 ( .A1(n3195), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4773 ( .A1(n4130), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4774 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3899)
         );
  AOI22_X1 U4775 ( .A1(n3208), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4776 ( .A1(n3190), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4777 ( .A1(n4596), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4778 ( .A1(n3539), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4779 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  NOR2_X1 U4780 ( .A1(n3899), .A2(n3898), .ZN(n3903) );
  NAND2_X1 U4781 ( .A1(n6680), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U4782 ( .A1(n3658), .A2(n3900), .ZN(n3901) );
  AOI21_X1 U4783 ( .B1(n4147), .B2(EAX_REG_18__SCAN_IN), .A(n3901), .ZN(n3902)
         );
  OAI21_X1 U4784 ( .B1(n4116), .B2(n3903), .A(n3902), .ZN(n3905) );
  XNOR2_X1 U4785 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3907), .ZN(n5743)
         );
  NAND2_X1 U4786 ( .A1(n4145), .A2(n5743), .ZN(n3904) );
  INV_X1 U4787 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3906) );
  INV_X1 U4788 ( .A(n3926), .ZN(n3925) );
  OR2_X1 U4789 ( .A1(n3908), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3909)
         );
  NAND2_X1 U4790 ( .A1(n3925), .A2(n3909), .ZN(n6077) );
  AOI22_X1 U4791 ( .A1(n3506), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4792 ( .A1(n3208), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4793 ( .A1(n3190), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4794 ( .A1(n4130), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4795 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4796 ( .A1(n4129), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4797 ( .A1(n4128), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4798 ( .A1(n3539), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3727), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4799 ( .A1(n4123), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4800 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NOR2_X1 U4801 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  NOR2_X1 U4802 ( .A1(n4116), .A2(n3920), .ZN(n3924) );
  INV_X1 U4803 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4804 ( .A1(n6680), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3921)
         );
  OAI211_X1 U4805 ( .C1(n3214), .C2(n3922), .A(n3658), .B(n3921), .ZN(n3923)
         );
  OAI22_X1 U4806 ( .A1(n6077), .A2(n3658), .B1(n3924), .B2(n3923), .ZN(n5522)
         );
  INV_X1 U4807 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U4808 ( .A1(n3925), .A2(n6039), .ZN(n3927) );
  AND2_X1 U4809 ( .A1(n3927), .A2(n3941), .ZN(n6045) );
  AOI21_X1 U4810 ( .B1(n6039), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3928) );
  AOI21_X1 U4811 ( .B1(n4147), .B2(EAX_REG_20__SCAN_IN), .A(n3928), .ZN(n3940)
         );
  AOI22_X1 U4812 ( .A1(n3506), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4813 ( .A1(n4121), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4814 ( .A1(n3210), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4815 ( .A1(n3195), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4816 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3938)
         );
  AOI22_X1 U4817 ( .A1(n3190), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4818 ( .A1(n4130), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4819 ( .A1(n4596), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4820 ( .A1(n3727), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3933) );
  NAND4_X1 U4821 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3937)
         );
  INV_X1 U4822 ( .A(n4116), .ZN(n4142) );
  OAI21_X1 U4823 ( .B1(n3938), .B2(n3937), .A(n4142), .ZN(n3939) );
  AOI22_X1 U4824 ( .A1(n6045), .A2(n4145), .B1(n3940), .B2(n3939), .ZN(n5603)
         );
  INV_X1 U4825 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3953) );
  AND2_X1 U4826 ( .A1(n3941), .A2(n3953), .ZN(n3942) );
  OR2_X1 U4827 ( .A1(n3942), .A2(n3975), .ZN(n5729) );
  AOI22_X1 U4828 ( .A1(n3506), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4829 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n3210), .B1(n3192), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4830 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4596), .B1(n3190), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4831 ( .A1(n4129), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4832 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3952)
         );
  AOI22_X1 U4833 ( .A1(n4121), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4834 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n3539), .B1(n4130), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4835 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4128), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4836 ( .A1(n3727), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4837 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  NOR2_X1 U4838 ( .A1(n3952), .A2(n3951), .ZN(n3956) );
  OAI21_X1 U4839 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3953), .A(n3658), .ZN(
        n3954) );
  AOI21_X1 U4840 ( .B1(n4147), .B2(EAX_REG_21__SCAN_IN), .A(n3954), .ZN(n3955)
         );
  OAI21_X1 U4841 ( .B1(n4116), .B2(n3956), .A(n3955), .ZN(n3957) );
  OAI21_X1 U4842 ( .B1(n5729), .B2(n3658), .A(n3957), .ZN(n5508) );
  INV_X1 U4843 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5720) );
  XNOR2_X1 U4844 ( .A(n3975), .B(n5720), .ZN(n5724) );
  NAND2_X1 U4845 ( .A1(n5724), .A2(n4145), .ZN(n3973) );
  AOI22_X1 U4846 ( .A1(n4121), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4847 ( .A1(n3506), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4848 ( .A1(n3539), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4849 ( .A1(n4130), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4850 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3967)
         );
  AOI22_X1 U4851 ( .A1(n3210), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4852 ( .A1(n4123), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4853 ( .A1(n4128), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4854 ( .A1(n3190), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4855 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3966)
         );
  NOR2_X1 U4856 ( .A1(n3967), .A2(n3966), .ZN(n3971) );
  NAND2_X1 U4857 ( .A1(n6680), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3968)
         );
  NAND2_X1 U4858 ( .A1(n3658), .A2(n3968), .ZN(n3969) );
  AOI21_X1 U4859 ( .B1(n4147), .B2(EAX_REG_22__SCAN_IN), .A(n3969), .ZN(n3970)
         );
  OAI21_X1 U4860 ( .B1(n4116), .B2(n3971), .A(n3970), .ZN(n3972) );
  NAND2_X1 U4861 ( .A1(n3973), .A2(n3972), .ZN(n5492) );
  INV_X1 U4862 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4863 ( .A1(n3976), .A2(n3998), .ZN(n3977) );
  NAND2_X1 U4864 ( .A1(n4023), .A2(n3977), .ZN(n6029) );
  AOI22_X1 U4865 ( .A1(n3506), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4866 ( .A1(n3204), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4867 ( .A1(n3208), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4868 ( .A1(n4596), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4869 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4870 ( .A1(n3190), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4871 ( .A1(n4121), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4872 ( .A1(n4123), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4873 ( .A1(n3727), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4874 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  NOR2_X1 U4875 ( .A1(n3987), .A2(n3986), .ZN(n4004) );
  AOI22_X1 U4876 ( .A1(n3208), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4877 ( .A1(n4123), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4878 ( .A1(n4121), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4879 ( .A1(n3727), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4880 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3997)
         );
  AOI22_X1 U4881 ( .A1(n3506), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4882 ( .A1(n4129), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4883 ( .A1(n3190), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4884 ( .A1(n3204), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U4885 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n3996)
         );
  NOR2_X1 U4886 ( .A1(n3997), .A2(n3996), .ZN(n4005) );
  XNOR2_X1 U4887 ( .A(n4004), .B(n4005), .ZN(n4001) );
  OAI21_X1 U4888 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3998), .A(n3658), .ZN(
        n3999) );
  AOI21_X1 U4889 ( .B1(n4147), .B2(EAX_REG_23__SCAN_IN), .A(n3999), .ZN(n4000)
         );
  OAI21_X1 U4890 ( .B1(n4001), .B2(n4116), .A(n4000), .ZN(n4002) );
  XNOR2_X1 U4891 ( .A(n4023), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6019)
         );
  NOR2_X1 U4892 ( .A1(n4005), .A2(n4004), .ZN(n4037) );
  AOI22_X1 U4893 ( .A1(n3506), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4894 ( .A1(n4121), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4895 ( .A1(n3210), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4896 ( .A1(n3204), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4897 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4015)
         );
  AOI22_X1 U4898 ( .A1(n3190), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4899 ( .A1(n4130), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4900 ( .A1(n4596), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4901 ( .A1(n3727), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4902 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4014)
         );
  OR2_X1 U4903 ( .A1(n4015), .A2(n4014), .ZN(n4036) );
  INV_X1 U4904 ( .A(n4036), .ZN(n4016) );
  XNOR2_X1 U4905 ( .A(n4037), .B(n4016), .ZN(n4020) );
  INV_X1 U4906 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4018) );
  INV_X1 U4907 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5704) );
  OAI22_X1 U4908 ( .A1(n3214), .A2(n4018), .B1(n5704), .B2(n4017), .ZN(n4019)
         );
  AOI21_X1 U4909 ( .B1(n4020), .B2(n4142), .A(n4019), .ZN(n4021) );
  NAND2_X1 U4910 ( .A1(n4022), .A2(n4021), .ZN(n5584) );
  OR2_X1 U4911 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4025)
         );
  NAND2_X1 U4912 ( .A1(n4060), .A2(n4025), .ZN(n5694) );
  AOI22_X1 U4913 ( .A1(n3506), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4914 ( .A1(n4121), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4915 ( .A1(n4123), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4916 ( .A1(n3727), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4917 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4035)
         );
  AOI22_X1 U4918 ( .A1(n3208), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4919 ( .A1(n4130), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4920 ( .A1(n4128), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4921 ( .A1(n3190), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4922 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4034)
         );
  NOR2_X1 U4923 ( .A1(n4035), .A2(n4034), .ZN(n4044) );
  NAND2_X1 U4924 ( .A1(n4037), .A2(n4036), .ZN(n4043) );
  XNOR2_X1 U4925 ( .A(n4044), .B(n4043), .ZN(n4040) );
  INV_X1 U4926 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5483) );
  AOI21_X1 U4927 ( .B1(n5483), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4038) );
  AOI21_X1 U4928 ( .B1(n4147), .B2(EAX_REG_25__SCAN_IN), .A(n4038), .ZN(n4039)
         );
  OAI21_X1 U4929 ( .B1(n4040), .B2(n4116), .A(n4039), .ZN(n4041) );
  NAND2_X1 U4930 ( .A1(n4042), .A2(n4041), .ZN(n5478) );
  XNOR2_X1 U4931 ( .A(n4060), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6008)
         );
  NAND2_X1 U4932 ( .A1(n6008), .A2(n4145), .ZN(n4059) );
  NOR2_X1 U4933 ( .A1(n4044), .A2(n4043), .ZN(n4074) );
  AOI22_X1 U4934 ( .A1(n3506), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4935 ( .A1(n4121), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4129), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4936 ( .A1(n3210), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4937 ( .A1(n3202), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U4938 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4054)
         );
  AOI22_X1 U4939 ( .A1(n3190), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4940 ( .A1(n4130), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4941 ( .A1(n4596), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4942 ( .A1(n3727), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U4943 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4053)
         );
  OR2_X1 U4944 ( .A1(n4054), .A2(n4053), .ZN(n4073) );
  XNOR2_X1 U4945 ( .A(n4074), .B(n4073), .ZN(n4057) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U4947 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6018), .A(n3658), .ZN(
        n4055) );
  AOI21_X1 U4948 ( .B1(n4147), .B2(EAX_REG_26__SCAN_IN), .A(n4055), .ZN(n4056)
         );
  OAI21_X1 U4949 ( .B1(n4057), .B2(n4116), .A(n4056), .ZN(n4058) );
  INV_X1 U4950 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U4951 ( .A1(n4061), .A2(n4075), .ZN(n4062) );
  NAND2_X1 U4952 ( .A1(n4098), .A2(n4062), .ZN(n6002) );
  AOI22_X1 U4953 ( .A1(n3506), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4954 ( .A1(n3210), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4955 ( .A1(n4130), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4956 ( .A1(n3193), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U4957 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4072)
         );
  AOI22_X1 U4958 ( .A1(n4129), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4959 ( .A1(n3190), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4960 ( .A1(n4596), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4961 ( .A1(n3439), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U4962 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4071)
         );
  NOR2_X1 U4963 ( .A1(n4072), .A2(n4071), .ZN(n4081) );
  NAND2_X1 U4964 ( .A1(n4074), .A2(n4073), .ZN(n4080) );
  XNOR2_X1 U4965 ( .A(n4081), .B(n4080), .ZN(n4078) );
  OAI21_X1 U4966 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4075), .A(n3658), .ZN(
        n4076) );
  AOI21_X1 U4967 ( .B1(n4147), .B2(EAX_REG_27__SCAN_IN), .A(n4076), .ZN(n4077)
         );
  OAI21_X1 U4968 ( .B1(n4078), .B2(n4116), .A(n4077), .ZN(n4079) );
  XNOR2_X1 U4969 ( .A(n4098), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5993)
         );
  NOR2_X1 U4970 ( .A1(n4081), .A2(n4080), .ZN(n4113) );
  AOI22_X1 U4971 ( .A1(n3506), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4972 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4129), .B1(n4121), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4973 ( .A1(n3210), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4974 ( .A1(n3204), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U4975 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4091)
         );
  AOI22_X1 U4976 ( .A1(n3190), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4977 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4130), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4978 ( .A1(n4596), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4979 ( .A1(n3727), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U4980 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  OR2_X1 U4981 ( .A1(n4091), .A2(n4090), .ZN(n4112) );
  INV_X1 U4982 ( .A(n4112), .ZN(n4092) );
  XNOR2_X1 U4983 ( .A(n4113), .B(n4092), .ZN(n4096) );
  INV_X1 U4984 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4094) );
  NAND2_X1 U4985 ( .A1(n6680), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4093)
         );
  OAI211_X1 U4986 ( .C1(n3214), .C2(n4094), .A(n3658), .B(n4093), .ZN(n4095)
         );
  AOI21_X1 U4987 ( .B1(n4096), .B2(n4142), .A(n4095), .ZN(n4097) );
  INV_X1 U4988 ( .A(n4098), .ZN(n4099) );
  NAND2_X1 U4989 ( .A1(n4099), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4100)
         );
  INV_X1 U4990 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n7126) );
  NAND2_X1 U4991 ( .A1(n4100), .A2(n7126), .ZN(n4101) );
  NAND2_X1 U4992 ( .A1(n4150), .A2(n4101), .ZN(n5663) );
  AOI22_X1 U4993 ( .A1(n4129), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U4994 ( .A1(n3506), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U4995 ( .A1(n4123), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U4996 ( .A1(n3439), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U4997 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4111)
         );
  AOI22_X1 U4998 ( .A1(n3193), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4999 ( .A1(n3208), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5000 ( .A1(n3190), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4596), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5001 ( .A1(n4130), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5002 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  NOR2_X1 U5003 ( .A1(n4111), .A2(n4110), .ZN(n4120) );
  NAND2_X1 U5004 ( .A1(n4113), .A2(n4112), .ZN(n4119) );
  XNOR2_X1 U5005 ( .A(n4120), .B(n4119), .ZN(n4117) );
  NOR2_X1 U5006 ( .A1(n7126), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4114) );
  AOI211_X1 U5007 ( .C1(n4147), .C2(EAX_REG_29__SCAN_IN), .A(n4145), .B(n4114), 
        .ZN(n4115) );
  OAI21_X1 U5008 ( .B1(n4117), .B2(n4116), .A(n4115), .ZN(n4118) );
  OAI21_X1 U5009 ( .B1(n5663), .B2(n3658), .A(n4118), .ZN(n5462) );
  XNOR2_X1 U5010 ( .A(n4150), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4449)
         );
  NOR2_X1 U5011 ( .A1(n4120), .A2(n4119), .ZN(n4138) );
  AOI22_X1 U5012 ( .A1(n3210), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5013 ( .A1(n3190), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3539), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5014 ( .A1(n4123), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5015 ( .A1(n3727), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3515), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5016 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4136)
         );
  AOI22_X1 U5017 ( .A1(n3506), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5018 ( .A1(n4129), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5019 ( .A1(n4596), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4130), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5020 ( .A1(n3204), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4131) );
  NAND4_X1 U5021 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4135)
         );
  NOR2_X1 U5022 ( .A1(n4136), .A2(n4135), .ZN(n4137) );
  XNOR2_X1 U5023 ( .A(n4138), .B(n4137), .ZN(n4143) );
  INV_X1 U5024 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4140) );
  OAI21_X1 U5025 ( .B1(n6124), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6680), 
        .ZN(n4139) );
  OAI21_X1 U5026 ( .B1(n3214), .B2(n4140), .A(n4139), .ZN(n4141) );
  AOI21_X1 U5027 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4144) );
  AOI22_X1 U5028 ( .A1(n4147), .A2(EAX_REG_31__SCAN_IN), .B1(n4146), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4148) );
  INV_X1 U5029 ( .A(n4148), .ZN(n4149) );
  INV_X1 U5030 ( .A(n5656), .ZN(n4323) );
  INV_X1 U5031 ( .A(n4150), .ZN(n4151) );
  NAND2_X1 U5032 ( .A1(n4151), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4153)
         );
  INV_X1 U5033 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4152) );
  NAND2_X1 U5034 ( .A1(n6658), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4154) );
  OAI21_X1 U5035 ( .B1(n6658), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4154), 
        .ZN(n4165) );
  NAND2_X1 U5036 ( .A1(n6662), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5037 ( .A1(n3604), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5038 ( .A1(n4156), .A2(n4155), .ZN(n4160) );
  INV_X1 U5039 ( .A(n4160), .ZN(n4158) );
  INV_X1 U5040 ( .A(n4156), .ZN(n4157) );
  XNOR2_X1 U5041 ( .A(n3632), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4187)
         );
  NOR2_X1 U5042 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n7080), .ZN(n4159)
         );
  NAND2_X1 U5043 ( .A1(n4691), .A2(n3452), .ZN(n4379) );
  NAND2_X1 U5044 ( .A1(n4203), .A2(n4191), .ZN(n4199) );
  INV_X1 U5045 ( .A(n4196), .ZN(n4163) );
  XNOR2_X1 U5046 ( .A(n4161), .B(n4160), .ZN(n4202) );
  INV_X1 U5047 ( .A(n4202), .ZN(n4162) );
  NAND2_X1 U5048 ( .A1(n4488), .A2(n4691), .ZN(n4164) );
  INV_X1 U5049 ( .A(n4178), .ZN(n4182) );
  AOI21_X1 U5050 ( .B1(n3452), .B2(n4196), .A(n3460), .ZN(n4176) );
  XOR2_X1 U5051 ( .A(n4166), .B(n4165), .Z(n4201) );
  NAND2_X1 U5052 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4201), .ZN(n4175) );
  INV_X1 U5053 ( .A(n4166), .ZN(n4167) );
  AOI21_X1 U5054 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n3308), .A(n4167), 
        .ZN(n4170) );
  INV_X1 U5055 ( .A(n4170), .ZN(n4168) );
  OAI21_X1 U5056 ( .B1(n4420), .B2(n4168), .A(n3448), .ZN(n4169) );
  AOI22_X1 U5057 ( .A1(n4178), .A2(n4169), .B1(n4176), .B2(n4175), .ZN(n4171)
         );
  NAND3_X1 U5058 ( .A1(n4170), .A2(n4171), .A3(n4196), .ZN(n4174) );
  INV_X1 U5059 ( .A(n4201), .ZN(n4172) );
  OAI21_X1 U5060 ( .B1(n4172), .B2(n4171), .A(n4191), .ZN(n4173) );
  OAI211_X1 U5061 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4173), .ZN(n4181)
         );
  INV_X1 U5062 ( .A(n4183), .ZN(n4177) );
  OAI211_X1 U5063 ( .C1(n4179), .C2(n4202), .A(n4178), .B(n4177), .ZN(n4180)
         );
  AOI22_X1 U5064 ( .A1(n4183), .A2(n4182), .B1(n4181), .B2(n4180), .ZN(n4194)
         );
  AND3_X1 U5065 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4184), .A3(n6115), 
        .ZN(n4185) );
  AOI211_X1 U5066 ( .C1(n4188), .C2(n4187), .A(n4186), .B(n4185), .ZN(n4190)
         );
  NOR2_X1 U5067 ( .A1(n4189), .A2(n4190), .ZN(n4193) );
  INV_X1 U5068 ( .A(n4190), .ZN(n4206) );
  AOI22_X1 U5069 ( .A1(n4191), .A2(n4206), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6685), .ZN(n4192) );
  OAI21_X1 U5070 ( .B1(n4194), .B2(n4193), .A(n4192), .ZN(n4195) );
  AOI21_X1 U5071 ( .B1(n4196), .B2(n4203), .A(n4195), .ZN(n4197) );
  INV_X1 U5072 ( .A(n4197), .ZN(n4198) );
  INV_X1 U5073 ( .A(n4200), .ZN(n4460) );
  NAND2_X1 U5074 ( .A1(n4202), .A2(n4201), .ZN(n4205) );
  INV_X1 U5075 ( .A(n4203), .ZN(n4204) );
  OAI21_X1 U5076 ( .B1(n4206), .B2(n4205), .A(n4204), .ZN(n4500) );
  INV_X1 U5077 ( .A(n4207), .ZN(n4503) );
  NOR2_X1 U5078 ( .A1(n4500), .A2(n4503), .ZN(n4456) );
  NAND2_X1 U5079 ( .A1(n4456), .A2(n6673), .ZN(n4454) );
  NAND2_X1 U5080 ( .A1(n6776), .A2(n6680), .ZN(n6694) );
  NOR3_X1 U5081 ( .A1(n6685), .A2(n6769), .A3(n6694), .ZN(n4211) );
  AND2_X1 U5082 ( .A1(n6685), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4422) );
  AND2_X1 U5083 ( .A1(n4422), .A2(n4145), .ZN(n6693) );
  INV_X1 U5084 ( .A(n6693), .ZN(n4209) );
  NOR2_X1 U5085 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6697) );
  INV_X1 U5086 ( .A(n6697), .ZN(n4208) );
  NAND2_X1 U5087 ( .A1(n4209), .A2(n6461), .ZN(n4210) );
  NAND2_X1 U5088 ( .A1(n5548), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4447) );
  NAND2_X2 U5089 ( .A1(n3452), .A2(n3448), .ZN(n4301) );
  NOR2_X2 U5090 ( .A1(n5599), .A2(n4301), .ZN(n4287) );
  INV_X1 U5091 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U5092 ( .A1(n4287), .A2(n6252), .ZN(n4214) );
  INV_X1 U5093 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U5094 ( .A1(n4861), .A2(n6252), .ZN(n4212) );
  OAI211_X1 U5095 ( .C1(n5599), .C2(n6494), .A(n4212), .B(n4215), .ZN(n4213)
         );
  NAND2_X1 U5096 ( .A1(n4214), .A2(n4213), .ZN(n4218) );
  INV_X1 U5097 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5270) );
  OR2_X1 U5098 ( .A1(n4215), .A2(n5270), .ZN(n4217) );
  NAND2_X1 U5099 ( .A1(n5599), .A2(n5270), .ZN(n4216) );
  NAND2_X1 U5100 ( .A1(n4217), .A2(n4216), .ZN(n4556) );
  XNOR2_X1 U5101 ( .A(n4218), .B(n4556), .ZN(n4860) );
  AOI21_X2 U5102 ( .B1(n4860), .B2(n4861), .A(n4218), .ZN(n4664) );
  INV_X1 U5103 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5104 ( .A1(n4287), .A2(n4665), .ZN(n4221) );
  INV_X1 U5105 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U5106 ( .A1(n4861), .A2(n4665), .ZN(n4219) );
  OAI211_X1 U5107 ( .C1(n5599), .C2(n7097), .A(n4219), .B(n4215), .ZN(n4220)
         );
  AND2_X1 U5108 ( .A1(n4221), .A2(n4220), .ZN(n4663) );
  MUX2_X1 U5109 ( .A(n4298), .B(n4215), .S(EBX_REG_3__SCAN_IN), .Z(n4223) );
  NAND2_X1 U5110 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4222)
         );
  NAND2_X1 U5111 ( .A1(n4223), .A2(n4222), .ZN(n4667) );
  INV_X1 U5112 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4224) );
  NAND2_X1 U5113 ( .A1(n4287), .A2(n4224), .ZN(n4227) );
  INV_X1 U5114 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U5115 ( .A1(n4861), .A2(n4224), .ZN(n4225) );
  OAI211_X1 U5116 ( .C1(n5599), .C2(n7065), .A(n4225), .B(n4215), .ZN(n4226)
         );
  NAND2_X1 U5117 ( .A1(n4227), .A2(n4226), .ZN(n4880) );
  MUX2_X1 U5118 ( .A(n4298), .B(n4215), .S(EBX_REG_5__SCAN_IN), .Z(n4230) );
  NAND2_X1 U5119 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4229)
         );
  INV_X1 U5120 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U5121 ( .A1(n4287), .A2(n4231), .ZN(n4234) );
  INV_X1 U5122 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U5123 ( .A1(n4861), .A2(n4231), .ZN(n4232) );
  OAI211_X1 U5124 ( .C1(n5599), .C2(n6450), .A(n4232), .B(n4215), .ZN(n4233)
         );
  NAND2_X1 U5125 ( .A1(n4234), .A2(n4233), .ZN(n4884) );
  INV_X1 U5126 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U5127 ( .A1(n4287), .A2(n5065), .ZN(n4237) );
  INV_X1 U5128 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U5129 ( .A1(n4861), .A2(n5065), .ZN(n4235) );
  OAI211_X1 U5130 ( .C1(n5599), .C2(n6432), .A(n4235), .B(n4215), .ZN(n4236)
         );
  NAND2_X1 U5131 ( .A1(n4237), .A2(n4236), .ZN(n4985) );
  INV_X1 U5132 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U5133 ( .A1(n4215), .A2(n6439), .ZN(n4239) );
  INV_X1 U5134 ( .A(EBX_REG_7__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U5135 ( .A1(n4861), .A2(n7076), .ZN(n4238) );
  NAND3_X1 U5136 ( .A1(n4239), .A2(n4298), .A3(n4238), .ZN(n4241) );
  NAND2_X1 U5137 ( .A1(n5599), .A2(n7076), .ZN(n4240) );
  AND2_X1 U5138 ( .A1(n4241), .A2(n4240), .ZN(n4983) );
  NOR2_X1 U5139 ( .A1(n4985), .A2(n4983), .ZN(n4242) );
  INV_X1 U5140 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U5141 ( .A1(n4287), .A2(n6268), .ZN(n4245) );
  INV_X1 U5142 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U5143 ( .A1(n4861), .A2(n6268), .ZN(n4243) );
  OAI211_X1 U5144 ( .C1(n5599), .C2(n5386), .A(n4243), .B(n4215), .ZN(n4244)
         );
  NAND2_X1 U5145 ( .A1(n4245), .A2(n4244), .ZN(n5392) );
  INV_X1 U5146 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U5147 ( .A1(n4215), .A2(n5387), .ZN(n4247) );
  INV_X1 U5148 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5149 ( .A1(n4861), .A2(n5230), .ZN(n4246) );
  NAND3_X1 U5150 ( .A1(n4247), .A2(n4298), .A3(n4246), .ZN(n4249) );
  NAND2_X1 U5151 ( .A1(n5599), .A2(n5230), .ZN(n4248) );
  NOR2_X1 U5152 ( .A1(n5392), .A2(n5389), .ZN(n4250) );
  INV_X1 U5153 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U5154 ( .A1(n4215), .A2(n5407), .ZN(n4252) );
  INV_X1 U5155 ( .A(EBX_REG_11__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U5156 ( .A1(n4861), .A2(n7115), .ZN(n4251) );
  NAND3_X1 U5157 ( .A1(n4252), .A2(n4298), .A3(n4251), .ZN(n4254) );
  NAND2_X1 U5158 ( .A1(n5599), .A2(n7115), .ZN(n4253) );
  INV_X1 U5159 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U5160 ( .A1(n4287), .A2(n6262), .ZN(n4257) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U5162 ( .A1(n4861), .A2(n6262), .ZN(n4255) );
  OAI211_X1 U5163 ( .C1(n5599), .C2(n6974), .A(n4255), .B(n4215), .ZN(n4256)
         );
  NAND2_X1 U5164 ( .A1(n4257), .A2(n4256), .ZN(n5959) );
  MUX2_X1 U5165 ( .A(n4298), .B(n4215), .S(EBX_REG_13__SCAN_IN), .Z(n4259) );
  NAND2_X1 U5166 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4258) );
  INV_X1 U5167 ( .A(n4287), .ZN(n4283) );
  MUX2_X1 U5168 ( .A(n4283), .B(n4298), .S(EBX_REG_14__SCAN_IN), .Z(n4261) );
  INV_X1 U5169 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U5170 ( .A1(n4464), .A2(n6108), .ZN(n4260) );
  MUX2_X1 U5171 ( .A(n4298), .B(n4215), .S(EBX_REG_15__SCAN_IN), .Z(n4263) );
  NAND2_X1 U5172 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U5173 ( .A1(n4263), .A2(n4262), .ZN(n5621) );
  MUX2_X1 U5174 ( .A(n4283), .B(n4298), .S(EBX_REG_16__SCAN_IN), .Z(n4265) );
  INV_X1 U5175 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U5176 ( .A1(n4464), .A2(n6098), .ZN(n4264) );
  NAND2_X1 U5177 ( .A1(n4265), .A2(n4264), .ZN(n5618) );
  MUX2_X1 U5178 ( .A(n4298), .B(n4215), .S(EBX_REG_17__SCAN_IN), .Z(n4267) );
  NAND2_X1 U5179 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U5180 ( .A1(n4267), .A2(n4266), .ZN(n5612) );
  MUX2_X1 U5181 ( .A(n4283), .B(n4298), .S(EBX_REG_19__SCAN_IN), .Z(n4268) );
  OAI21_X1 U5182 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4558), .A(n4268), 
        .ZN(n5526) );
  OAI22_X1 U5183 ( .A1(n4558), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4301), .ZN(n5601) );
  OR2_X1 U5184 ( .A1(n4558), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4270)
         );
  INV_X1 U5185 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U5186 ( .A1(n4861), .A2(n5605), .ZN(n4269) );
  NAND2_X1 U5187 ( .A1(n4270), .A2(n4269), .ZN(n5524) );
  INV_X1 U5188 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U5189 ( .A1(n5524), .A2(n6040), .ZN(n4271) );
  OAI21_X1 U5190 ( .B1(n5601), .B2(n5599), .A(n4271), .ZN(n4273) );
  NAND2_X1 U5191 ( .A1(n5524), .A2(n4298), .ZN(n4272) );
  MUX2_X1 U5192 ( .A(n4283), .B(n4298), .S(EBX_REG_21__SCAN_IN), .Z(n4274) );
  OAI21_X1 U5193 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4558), .A(n4274), 
        .ZN(n5511) );
  NOR2_X2 U5194 ( .A1(n5512), .A2(n5511), .ZN(n5497) );
  INV_X1 U5195 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U5196 ( .A1(n4215), .A2(n4275), .ZN(n4277) );
  INV_X1 U5197 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U5198 ( .A1(n4861), .A2(n5594), .ZN(n4276) );
  NAND3_X1 U5199 ( .A1(n4277), .A2(n4298), .A3(n4276), .ZN(n4279) );
  NAND2_X1 U5200 ( .A1(n5599), .A2(n5594), .ZN(n4278) );
  NAND2_X1 U5201 ( .A1(n4279), .A2(n4278), .ZN(n5496) );
  MUX2_X1 U5202 ( .A(n4283), .B(n4298), .S(EBX_REG_23__SCAN_IN), .Z(n4280) );
  OAI21_X1 U5203 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4558), .A(n4280), 
        .ZN(n5590) );
  MUX2_X1 U5204 ( .A(n4298), .B(n4215), .S(EBX_REG_24__SCAN_IN), .Z(n4282) );
  NAND2_X1 U5205 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4281) );
  AND2_X1 U5206 ( .A1(n4282), .A2(n4281), .ZN(n5585) );
  MUX2_X1 U5207 ( .A(n4283), .B(n4298), .S(EBX_REG_25__SCAN_IN), .Z(n4284) );
  OAI21_X1 U5208 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4558), .A(n4284), 
        .ZN(n5480) );
  MUX2_X1 U5209 ( .A(n4298), .B(n4215), .S(EBX_REG_26__SCAN_IN), .Z(n4286) );
  NAND2_X1 U5210 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U5211 ( .A1(n4286), .A2(n4285), .ZN(n5577) );
  INV_X1 U5212 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U5213 ( .A1(n4287), .A2(n6053), .ZN(n4290) );
  INV_X1 U5214 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U5215 ( .A1(n4861), .A2(n6053), .ZN(n4288) );
  OAI211_X1 U5216 ( .C1(n5599), .C2(n7106), .A(n4288), .B(n4215), .ZN(n4289)
         );
  AND2_X1 U5217 ( .A1(n4290), .A2(n4289), .ZN(n5833) );
  AND2_X2 U5218 ( .A1(n5576), .A2(n5833), .ZN(n5835) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U5220 ( .A1(n4215), .A2(n7066), .ZN(n4292) );
  INV_X1 U5221 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5222 ( .A1(n4861), .A2(n5570), .ZN(n4291) );
  NAND3_X1 U5223 ( .A1(n4292), .A2(n4298), .A3(n4291), .ZN(n4294) );
  NAND2_X1 U5224 ( .A1(n5599), .A2(n5570), .ZN(n4293) );
  NAND2_X1 U5225 ( .A1(n4294), .A2(n4293), .ZN(n5567) );
  NAND2_X2 U5226 ( .A1(n5835), .A2(n5567), .ZN(n5569) );
  OR2_X1 U5227 ( .A1(n4558), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4296)
         );
  INV_X1 U5228 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5229 ( .A1(n4861), .A2(n5563), .ZN(n4295) );
  NAND2_X1 U5230 ( .A1(n4296), .A2(n4295), .ZN(n5465) );
  NAND2_X1 U5231 ( .A1(n5599), .A2(n5563), .ZN(n5464) );
  AND2_X1 U5232 ( .A1(n4301), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4297)
         );
  AOI21_X1 U5233 ( .B1(n4558), .B2(EBX_REG_30__SCAN_IN), .A(n4297), .ZN(n4440)
         );
  NAND2_X1 U5234 ( .A1(n3219), .A2(n4298), .ZN(n4438) );
  OAI22_X1 U5235 ( .A1(n4558), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4301), .ZN(n4299) );
  NOR2_X1 U5236 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4307) );
  NOR2_X1 U5237 ( .A1(n5267), .A2(n4307), .ZN(n4444) );
  INV_X1 U5238 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5562) );
  NOR2_X1 U5239 ( .A1(n4301), .A2(n5562), .ZN(n4302) );
  INV_X1 U5240 ( .A(n4303), .ZN(n4304) );
  INV_X1 U5241 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U5242 ( .A1(n4304), .A2(n6707), .ZN(n6702) );
  OR3_X1 U5243 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6702), .ZN(
        n6676) );
  NAND2_X1 U5244 ( .A1(n3481), .A2(n6676), .ZN(n4305) );
  NOR2_X1 U5245 ( .A1(n5267), .A2(n4305), .ZN(n4443) );
  AOI22_X1 U5246 ( .A1(n4443), .A2(EBX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n6244), .ZN(n4306) );
  OAI21_X1 U5247 ( .B1(n5785), .B2(n6234), .A(n4306), .ZN(n4321) );
  INV_X1 U5248 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6738) );
  INV_X1 U5249 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U5250 ( .A1(n4488), .A2(n6702), .ZN(n4542) );
  NAND3_X1 U5251 ( .A1(n4542), .A2(n4307), .A3(n3448), .ZN(n4308) );
  INV_X1 U5252 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6906) );
  INV_X1 U5253 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6728) );
  INV_X1 U5254 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6722) );
  INV_X1 U5255 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6720) );
  INV_X1 U5256 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6718) );
  NAND3_X1 U5257 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5557) );
  NOR2_X1 U5258 ( .A1(n6718), .A2(n5557), .ZN(n6216) );
  NAND2_X1 U5259 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6216), .ZN(n5249) );
  NOR3_X1 U5260 ( .A1(n6722), .A2(n6720), .A3(n5249), .ZN(n5069) );
  NAND2_X1 U5261 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5069), .ZN(n5067) );
  NAND2_X1 U5262 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5311) );
  NOR3_X1 U5263 ( .A1(n6728), .A2(n5067), .A3(n5311), .ZN(n5425) );
  NAND2_X1 U5264 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5425), .ZN(n5420) );
  NOR2_X1 U5265 ( .A1(n6906), .A2(n5420), .ZN(n4311) );
  NAND2_X1 U5266 ( .A1(n6217), .A2(n4311), .ZN(n6172) );
  NAND4_X1 U5267 ( .A1(n6163), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U5268 ( .A1(n6738), .A2(n5540), .ZN(n5531) );
  NAND2_X1 U5269 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5531), .ZN(n6047) );
  NAND4_X1 U5270 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n6028), .ZN(n6026) );
  NAND3_X1 U5271 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4315) );
  NOR2_X1 U5272 ( .A1(n6026), .A2(n4315), .ZN(n6004) );
  AND2_X1 U5273 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4309) );
  NAND2_X1 U5274 ( .A1(n6004), .A2(n4309), .ZN(n5463) );
  INV_X1 U5275 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6759) );
  NAND3_X1 U5276 ( .A1(n6759), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n4310) );
  NOR2_X1 U5277 ( .A1(n5463), .A2(n4310), .ZN(n4319) );
  NAND3_X1 U5278 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U5279 ( .A1(n6247), .A2(n5548), .ZN(n5273) );
  INV_X1 U5280 ( .A(n5273), .ZN(n5991) );
  INV_X1 U5281 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6736) );
  NOR3_X1 U5282 ( .A1(n5735), .A2(n6736), .A3(n6738), .ZN(n4313) );
  NAND3_X1 U5283 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4312) );
  OAI221_X1 U5284 ( .B1(n6247), .B2(n4311), .C1(n6247), .C2(
        REIP_REG_14__SCAN_IN), .A(n5548), .ZN(n6174) );
  AOI21_X1 U5285 ( .B1(n4312), .B2(n5273), .A(n6174), .ZN(n6150) );
  OAI21_X1 U5286 ( .B1(n5991), .B2(n4313), .A(n6150), .ZN(n6038) );
  AOI21_X1 U5287 ( .B1(n4314), .B2(n5273), .A(n6038), .ZN(n6037) );
  NAND2_X1 U5288 ( .A1(n5273), .A2(n4315), .ZN(n4316) );
  NAND2_X1 U5289 ( .A1(n6037), .A2(n4316), .ZN(n6015) );
  NAND2_X1 U5290 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4317) );
  NOR2_X1 U5291 ( .A1(n6015), .A2(n4317), .ZN(n5990) );
  AND2_X1 U5292 ( .A1(n5990), .A2(REIP_REG_29__SCAN_IN), .ZN(n4432) );
  AOI211_X1 U5293 ( .C1(n4432), .C2(REIP_REG_30__SCAN_IN), .A(n5991), .B(n6759), .ZN(n4318) );
  OAI21_X1 U5294 ( .B1(n4323), .B2(n6198), .A(n4322), .ZN(U2796) );
  INV_X1 U5295 ( .A(n4379), .ZN(n4390) );
  NAND2_X1 U5296 ( .A1(n4675), .A2(n4390), .ZN(n4327) );
  XNOR2_X1 U5297 ( .A(n4335), .B(n4334), .ZN(n4324) );
  INV_X1 U5298 ( .A(n3481), .ZN(n6798) );
  OAI211_X1 U5299 ( .C1(n4324), .C2(n6798), .A(n3212), .B(n4691), .ZN(n4325)
         );
  INV_X1 U5300 ( .A(n4325), .ZN(n4326) );
  NAND2_X1 U5301 ( .A1(n4472), .A2(n3483), .ZN(n4336) );
  OAI21_X1 U5302 ( .B1(n6798), .B2(n4334), .A(n4336), .ZN(n4328) );
  INV_X1 U5303 ( .A(n4328), .ZN(n4329) );
  OAI21_X2 U5304 ( .B1(n5108), .B2(n4379), .A(n4329), .ZN(n4551) );
  NAND2_X1 U5305 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4330)
         );
  NAND2_X1 U5306 ( .A1(n4330), .A2(n6494), .ZN(n4331) );
  AND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U5308 ( .A1(n4551), .A2(n6474), .ZN(n4332) );
  AND2_X1 U5309 ( .A1(n4331), .A2(n4332), .ZN(n4763) );
  NAND2_X1 U5310 ( .A1(n4762), .A2(n4763), .ZN(n4333) );
  NAND2_X1 U5311 ( .A1(n6398), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4341)
         );
  OR2_X1 U5312 ( .A1(n4673), .A2(n4379), .ZN(n4340) );
  NAND2_X1 U5313 ( .A1(n4335), .A2(n4334), .ZN(n4346) );
  XNOR2_X1 U5314 ( .A(n4346), .B(n4345), .ZN(n4338) );
  INV_X1 U5315 ( .A(n4336), .ZN(n4337) );
  AOI21_X1 U5316 ( .B1(n4338), .B2(n3481), .A(n4337), .ZN(n4339) );
  NAND2_X1 U5317 ( .A1(n4341), .A2(n6396), .ZN(n4344) );
  AND2_X1 U5318 ( .A1(n4344), .A2(n4343), .ZN(n6387) );
  NAND2_X1 U5319 ( .A1(n4715), .A2(n4390), .ZN(n4350) );
  NAND2_X1 U5320 ( .A1(n4346), .A2(n4345), .ZN(n4355) );
  INV_X1 U5321 ( .A(n4354), .ZN(n4347) );
  XNOR2_X1 U5322 ( .A(n4355), .B(n4347), .ZN(n4348) );
  NAND2_X1 U5323 ( .A1(n4348), .A2(n3481), .ZN(n4349) );
  INV_X1 U5324 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6468) );
  XNOR2_X1 U5325 ( .A(n4351), .B(n6468), .ZN(n6389) );
  NAND2_X1 U5326 ( .A1(n6387), .A2(n6389), .ZN(n6388) );
  NAND2_X1 U5327 ( .A1(n4351), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4352)
         );
  NAND2_X1 U5328 ( .A1(n4353), .A2(n4390), .ZN(n4358) );
  NAND2_X1 U5329 ( .A1(n4355), .A2(n4354), .ZN(n4373) );
  XNOR2_X1 U5330 ( .A(n4373), .B(n4371), .ZN(n4356) );
  NAND2_X1 U5331 ( .A1(n4356), .A2(n3481), .ZN(n4357) );
  NAND2_X1 U5332 ( .A1(n4358), .A2(n4357), .ZN(n4359) );
  XNOR2_X1 U5333 ( .A(n4359), .B(n7065), .ZN(n4774) );
  NAND2_X1 U5334 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4360)
         );
  NAND2_X1 U5335 ( .A1(n4361), .A2(n4390), .ZN(n4366) );
  INV_X1 U5336 ( .A(n4371), .ZN(n4362) );
  OR2_X1 U5337 ( .A1(n4373), .A2(n4362), .ZN(n4363) );
  XNOR2_X1 U5338 ( .A(n4363), .B(n4370), .ZN(n4364) );
  NAND2_X1 U5339 ( .A1(n4364), .A2(n3481), .ZN(n4365) );
  INV_X1 U5340 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4873) );
  NAND3_X1 U5341 ( .A1(n4368), .A2(n4390), .A3(n4369), .ZN(n4376) );
  NAND2_X1 U5342 ( .A1(n4371), .A2(n4370), .ZN(n4372) );
  OR2_X1 U5343 ( .A1(n4373), .A2(n4372), .ZN(n4381) );
  XNOR2_X1 U5344 ( .A(n4381), .B(n4382), .ZN(n4374) );
  NAND2_X1 U5345 ( .A1(n4374), .A2(n3481), .ZN(n4375) );
  NAND2_X1 U5346 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  XNOR2_X1 U5347 ( .A(n4377), .B(n6450), .ZN(n4887) );
  NAND2_X1 U5348 ( .A1(n4377), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4378)
         );
  OR2_X1 U5349 ( .A1(n4380), .A2(n4379), .ZN(n4386) );
  INV_X1 U5350 ( .A(n4381), .ZN(n4383) );
  NAND2_X1 U5351 ( .A1(n4383), .A2(n4382), .ZN(n4392) );
  XNOR2_X1 U5352 ( .A(n4392), .B(n4389), .ZN(n4384) );
  NAND2_X1 U5353 ( .A1(n4384), .A2(n3481), .ZN(n4385) );
  NAND2_X1 U5354 ( .A1(n4386), .A2(n4385), .ZN(n4387) );
  XNOR2_X1 U5355 ( .A(n4387), .B(n6439), .ZN(n6375) );
  NAND2_X1 U5356 ( .A1(n6376), .A2(n6375), .ZN(n6374) );
  NAND2_X1 U5357 ( .A1(n4387), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4388)
         );
  NAND2_X2 U5358 ( .A1(n6374), .A2(n4388), .ZN(n5242) );
  AND3_X1 U5359 ( .A1(n4390), .A2(n4644), .A3(n4389), .ZN(n4391) );
  OR3_X1 U5360 ( .A1(n4392), .A2(n3260), .A3(n6798), .ZN(n4393) );
  NAND2_X1 U5361 ( .A1(n4408), .A2(n4393), .ZN(n4394) );
  XNOR2_X1 U5362 ( .A(n4394), .B(n6432), .ZN(n5241) );
  NAND2_X1 U5363 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4395)
         );
  NAND2_X1 U5364 ( .A1(n3194), .A2(n5387), .ZN(n5320) );
  OR2_X1 U5365 ( .A1(n3194), .A2(n5387), .ZN(n5321) );
  NAND2_X1 U5366 ( .A1(n3194), .A2(n5386), .ZN(n5382) );
  AND2_X1 U5367 ( .A1(n3194), .A2(n5407), .ZN(n4399) );
  NOR2_X1 U5368 ( .A1(n3194), .A2(n6974), .ZN(n5777) );
  NAND2_X1 U5369 ( .A1(n3194), .A2(n6974), .ZN(n5776) );
  XNOR2_X1 U5370 ( .A(n3194), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5768)
         );
  INV_X1 U5371 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5949) );
  INV_X1 U5372 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6092) );
  XNOR2_X1 U5373 ( .A(n3194), .B(n6092), .ZN(n5754) );
  NAND2_X1 U5374 ( .A1(n3194), .A2(n6092), .ZN(n4401) );
  INV_X1 U5375 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4402) );
  INV_X1 U5376 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6082) );
  AND3_X1 U5377 ( .A1(n6098), .A2(n4402), .A3(n6082), .ZN(n4403) );
  NAND2_X1 U5378 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5912) );
  AND2_X1 U5379 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5873) );
  AND2_X1 U5380 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5896) );
  AND2_X1 U5381 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5798) );
  NAND3_X1 U5382 ( .A1(n5873), .A2(n5896), .A3(n5798), .ZN(n4406) );
  NAND2_X1 U5383 ( .A1(n3194), .A2(n4406), .ZN(n4407) );
  NAND2_X1 U5384 ( .A1(n5910), .A2(n4407), .ZN(n4411) );
  NOR2_X1 U5385 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5897) );
  NOR2_X1 U5386 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5874) );
  INV_X1 U5387 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5859) );
  INV_X1 U5388 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5858) );
  NAND4_X1 U5389 ( .A1(n5897), .A2(n5874), .A3(n5859), .A4(n5858), .ZN(n4409)
         );
  NAND2_X1 U5390 ( .A1(n4396), .A2(n4409), .ZN(n4410) );
  NAND2_X1 U5391 ( .A1(n4411), .A2(n4410), .ZN(n5667) );
  XOR2_X1 U5392 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n3194), .Z(n5692) );
  INV_X1 U5393 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U5394 ( .A1(n3194), .A2(n5850), .ZN(n4412) );
  INV_X1 U5395 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n7109) );
  NOR2_X1 U5396 ( .A1(n4396), .A2(n7109), .ZN(n5686) );
  NAND2_X1 U5397 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5398 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4417) );
  NOR3_X1 U5399 ( .A1(n5684), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U5400 ( .A1(n4413), .A2(n5648), .ZN(n5659) );
  INV_X1 U5401 ( .A(n5659), .ZN(n4415) );
  NAND2_X1 U5402 ( .A1(n4415), .A2(n4414), .ZN(n4416) );
  NAND2_X1 U5403 ( .A1(n4417), .A2(n4416), .ZN(n4418) );
  XNOR2_X1 U5404 ( .A(n4418), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5816)
         );
  NAND2_X1 U5405 ( .A1(n4419), .A2(n4420), .ZN(n6646) );
  NAND2_X1 U5406 ( .A1(n4422), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6695) );
  NOR2_X2 U5407 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6567) );
  NAND2_X1 U5408 ( .A1(n6559), .A2(n4423), .ZN(n6794) );
  NAND2_X1 U5409 ( .A1(n6794), .A2(n6685), .ZN(n4424) );
  NAND2_X1 U5410 ( .A1(n6685), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U5411 ( .A1(n6124), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4425) );
  AND2_X1 U5412 ( .A1(n4426), .A2(n4425), .ZN(n4569) );
  INV_X1 U5413 ( .A(n4569), .ZN(n4427) );
  INV_X1 U5414 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U5415 ( .A1(n6471), .A2(REIP_REG_30__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U5416 ( .B1(n5780), .B2(n4428), .A(n5810), .ZN(n4429) );
  AOI21_X1 U5417 ( .B1(n4449), .B2(n5782), .A(n4429), .ZN(n4430) );
  NAND2_X1 U5418 ( .A1(n5273), .A2(REIP_REG_30__SCAN_IN), .ZN(n4431) );
  INV_X1 U5419 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U5420 ( .A1(n4433), .A2(REIP_REG_29__SCAN_IN), .ZN(n4434) );
  INV_X1 U5421 ( .A(n4440), .ZN(n4437) );
  INV_X1 U5422 ( .A(n5569), .ZN(n4435) );
  NAND2_X1 U5423 ( .A1(n3219), .A2(n4435), .ZN(n4436) );
  NAND3_X1 U5424 ( .A1(n4438), .A2(n4437), .A3(n4436), .ZN(n4442) );
  NAND2_X1 U5425 ( .A1(n5569), .A2(n5599), .ZN(n4439) );
  NAND3_X1 U5426 ( .A1(n3219), .A2(n4440), .A3(n4439), .ZN(n4441) );
  NAND2_X1 U5427 ( .A1(n4442), .A2(n4441), .ZN(n5812) );
  INV_X1 U5428 ( .A(n4443), .ZN(n4446) );
  NAND3_X1 U5429 ( .A1(n4444), .A2(n3448), .A3(n5562), .ZN(n4445) );
  AOI22_X1 U5430 ( .A1(n6224), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6244), .ZN(n4451) );
  INV_X1 U5431 ( .A(n4447), .ZN(n4448) );
  NAND2_X1 U5432 ( .A1(n6212), .A2(n4449), .ZN(n4450) );
  OAI211_X1 U5433 ( .C1(n5812), .C2(n6234), .A(n4451), .B(n4450), .ZN(n4452)
         );
  INV_X1 U5434 ( .A(n4452), .ZN(n4453) );
  NAND4_X1 U5435 ( .A1(n3305), .A2(n3297), .A3(n3221), .A4(n4453), .ZN(U2797)
         );
  AND2_X1 U5436 ( .A1(n6567), .A2(n6776), .ZN(n5063) );
  INV_X1 U5437 ( .A(n4489), .ZN(n4487) );
  AOI211_X1 U5438 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4454), .A(n5063), .B(
        n4487), .ZN(n4455) );
  INV_X1 U5439 ( .A(n4455), .ZN(U2788) );
  OR2_X1 U5440 ( .A1(n4540), .A2(n3463), .ZN(n4458) );
  OR2_X1 U5441 ( .A1(n4456), .A2(n4200), .ZN(n4457) );
  NAND2_X1 U5442 ( .A1(n4458), .A2(n4457), .ZN(n6119) );
  INV_X1 U5443 ( .A(n5266), .ZN(n4459) );
  OR2_X1 U5444 ( .A1(n3481), .A2(n4459), .ZN(n4485) );
  AOI21_X1 U5445 ( .B1(n4485), .B2(n6702), .A(READY_N), .ZN(n6797) );
  NOR2_X1 U5446 ( .A1(n6119), .A2(n6797), .ZN(n6644) );
  OR2_X1 U5447 ( .A1(n6644), .A2(n6690), .ZN(n4481) );
  INV_X1 U5448 ( .A(n4481), .ZN(n6126) );
  INV_X1 U5449 ( .A(MORE_REG_SCAN_IN), .ZN(n4483) );
  INV_X1 U5450 ( .A(n4540), .ZN(n4657) );
  NAND2_X1 U5451 ( .A1(n4419), .A2(n3463), .ZN(n4638) );
  AND2_X1 U5452 ( .A1(n4638), .A2(n6646), .ZN(n4554) );
  NAND2_X1 U5453 ( .A1(n4554), .A2(n4460), .ZN(n4461) );
  NAND2_X1 U5454 ( .A1(n4657), .A2(n4461), .ZN(n4480) );
  NAND2_X1 U5455 ( .A1(n4462), .A2(n3448), .ZN(n4463) );
  MUX2_X1 U5456 ( .A(n6798), .B(n4463), .S(n3450), .Z(n4501) );
  OR2_X1 U5457 ( .A1(n5266), .A2(n4700), .ZN(n4504) );
  AOI21_X1 U5458 ( .B1(n4464), .B2(n4504), .A(n3212), .ZN(n4468) );
  NAND2_X1 U5459 ( .A1(n3482), .A2(n5599), .ZN(n4466) );
  OAI21_X1 U5460 ( .B1(n4543), .B2(n3448), .A(n4700), .ZN(n4465) );
  NAND2_X1 U5461 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  NOR2_X1 U5462 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  NAND3_X1 U5463 ( .A1(n4470), .A2(n4501), .A3(n4469), .ZN(n4516) );
  NAND3_X1 U5464 ( .A1(n4473), .A2(n4472), .A3(n4691), .ZN(n4474) );
  OR2_X1 U5465 ( .A1(n4477), .A2(n4474), .ZN(n4609) );
  OR2_X1 U5466 ( .A1(n4513), .A2(n3448), .ZN(n4475) );
  OAI211_X1 U5467 ( .C1(n4471), .C2(n3393), .A(n4609), .B(n4475), .ZN(n4476)
         );
  NOR2_X1 U5468 ( .A1(n4516), .A2(n4476), .ZN(n4549) );
  NOR2_X1 U5469 ( .A1(n4477), .A2(n4488), .ZN(n4535) );
  NAND2_X1 U5470 ( .A1(n4656), .A2(n4540), .ZN(n4479) );
  NAND2_X1 U5471 ( .A1(n4500), .A2(n4207), .ZN(n4478) );
  AND3_X1 U5472 ( .A1(n4480), .A2(n4479), .A3(n4478), .ZN(n6647) );
  OR2_X1 U5473 ( .A1(n4481), .A2(n6647), .ZN(n4482) );
  OAI21_X1 U5474 ( .B1(n6126), .B2(n4483), .A(n4482), .ZN(U3471) );
  INV_X1 U5475 ( .A(n6793), .ZN(n4486) );
  OAI21_X1 U5476 ( .B1(n5063), .B2(READREQUEST_REG_SCAN_IN), .A(n4486), .ZN(
        n4484) );
  OAI21_X1 U5477 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(U3474) );
  INV_X1 U5478 ( .A(READY_N), .ZN(n6795) );
  OAI21_X1 U5479 ( .B1(n3481), .B2(n6795), .A(n4487), .ZN(n6366) );
  INV_X1 U5480 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n7029) );
  INV_X1 U5481 ( .A(DATAI_9_), .ZN(n4490) );
  NOR2_X1 U5482 ( .A1(n6328), .A2(n4490), .ZN(n6325) );
  INV_X1 U5483 ( .A(n6325), .ZN(n4494) );
  NAND2_X1 U5484 ( .A1(n4492), .A2(n3481), .ZN(n6677) );
  INV_X1 U5485 ( .A(n6373), .ZN(n6368) );
  NAND2_X1 U5486 ( .A1(n6368), .A2(EAX_REG_9__SCAN_IN), .ZN(n4493) );
  OAI211_X1 U5487 ( .C1(n6313), .C2(n7029), .A(n4494), .B(n4493), .ZN(U2948)
         );
  AND2_X1 U5488 ( .A1(n4207), .A2(n3452), .ZN(n6654) );
  INV_X1 U5489 ( .A(n6702), .ZN(n4533) );
  NAND2_X1 U5490 ( .A1(n6654), .A2(n4533), .ZN(n4496) );
  OAI21_X1 U5491 ( .B1(n4533), .B2(n4861), .A(n4492), .ZN(n4495) );
  NAND2_X1 U5492 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  NAND2_X1 U5493 ( .A1(n4497), .A2(n6795), .ZN(n4498) );
  NAND2_X1 U5494 ( .A1(n4498), .A2(n4638), .ZN(n4507) );
  NOR2_X1 U5495 ( .A1(READY_N), .A2(n4500), .ZN(n4640) );
  INV_X1 U5496 ( .A(n4640), .ZN(n4505) );
  NAND2_X1 U5497 ( .A1(n4419), .A2(n4501), .ZN(n4502) );
  NAND2_X1 U5498 ( .A1(n4503), .A2(n4502), .ZN(n4538) );
  OAI211_X1 U5499 ( .C1(n4499), .C2(n4505), .A(n4538), .B(n4504), .ZN(n4506)
         );
  AOI21_X1 U5500 ( .B1(n4507), .B2(n4540), .A(n4506), .ZN(n4509) );
  NAND2_X1 U5501 ( .A1(n4657), .A2(n4656), .ZN(n4508) );
  INV_X1 U5502 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7090) );
  NOR2_X1 U5503 ( .A1(n6776), .A2(n6680), .ZN(n4628) );
  NAND2_X1 U5504 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4628), .ZN(n6767) );
  NOR2_X1 U5505 ( .A1(n7090), .A2(n6767), .ZN(n4510) );
  AOI21_X1 U5506 ( .B1(n6673), .B2(n6655), .A(n4510), .ZN(n6117) );
  OAI21_X1 U5507 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6769), .A(n6117), .ZN(
        n6780) );
  OAI21_X1 U5508 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6771), .A(n6780), 
        .ZN(n6778) );
  INV_X1 U5509 ( .A(n6778), .ZN(n4525) );
  INV_X1 U5510 ( .A(n6780), .ZN(n6774) );
  INV_X1 U5511 ( .A(n6771), .ZN(n5451) );
  INV_X1 U5512 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5513 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4511), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6494), .ZN(n5447) );
  NAND2_X1 U5514 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5446) );
  INV_X1 U5515 ( .A(n5446), .ZN(n4522) );
  NAND2_X1 U5516 ( .A1(n4513), .A2(n4471), .ZN(n4514) );
  NOR2_X1 U5517 ( .A1(n4492), .A2(n4514), .ZN(n4515) );
  AND2_X1 U5518 ( .A1(n4499), .A2(n4515), .ZN(n4518) );
  INV_X1 U5519 ( .A(n4516), .ZN(n4517) );
  NAND2_X1 U5520 ( .A1(n4518), .A2(n4517), .ZN(n6652) );
  INV_X1 U5521 ( .A(n6652), .ZN(n4606) );
  NAND2_X1 U5522 ( .A1(n6654), .A2(n3307), .ZN(n4521) );
  OAI21_X1 U5523 ( .B1(n4523), .B2(n4519), .A(n6651), .ZN(n4520) );
  OAI211_X1 U5524 ( .C1(n4512), .C2(n4606), .A(n4521), .B(n4520), .ZN(n6656)
         );
  INV_X1 U5525 ( .A(n6782), .ZN(n6113) );
  AOI222_X1 U5526 ( .A1(n5451), .A2(n4523), .B1(n5447), .B2(n4522), .C1(n6656), 
        .C2(n6113), .ZN(n4524) );
  OAI22_X1 U5527 ( .A1(n4525), .A2(n3307), .B1(n6774), .B2(n4524), .ZN(U3460)
         );
  INV_X1 U5528 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n7145) );
  INV_X1 U5529 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5005) );
  OAI22_X1 U5530 ( .A1(n6313), .A2(n7145), .B1(n5005), .B2(n6373), .ZN(n4526)
         );
  INV_X1 U5531 ( .A(DATAI_7_), .ZN(n5007) );
  NOR2_X1 U5532 ( .A1(n6328), .A2(n5007), .ZN(n6322) );
  OR2_X1 U5533 ( .A1(n4526), .A2(n6322), .ZN(U2946) );
  INV_X1 U5534 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n7138) );
  AND2_X1 U5535 ( .A1(n6371), .A2(DATAI_13_), .ZN(n6365) );
  INV_X1 U5536 ( .A(n6365), .ZN(n4528) );
  NAND2_X1 U5537 ( .A1(n6368), .A2(EAX_REG_29__SCAN_IN), .ZN(n4527) );
  OAI211_X1 U5538 ( .C1(n6313), .C2(n7138), .A(n4528), .B(n4527), .ZN(U2937)
         );
  INV_X1 U5539 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n7001) );
  AND2_X1 U5540 ( .A1(n6371), .A2(DATAI_11_), .ZN(n6331) );
  INV_X1 U5541 ( .A(n6331), .ZN(n4530) );
  NAND2_X1 U5542 ( .A1(n6368), .A2(EAX_REG_11__SCAN_IN), .ZN(n4529) );
  OAI211_X1 U5543 ( .C1(n6313), .C2(n7001), .A(n4530), .B(n4529), .ZN(U2950)
         );
  INV_X1 U5544 ( .A(n6654), .ZN(n4531) );
  OR2_X1 U5545 ( .A1(n4639), .A2(n4531), .ZN(n4532) );
  NAND2_X1 U5546 ( .A1(n6373), .A2(n4532), .ZN(n4534) );
  NAND2_X1 U5547 ( .A1(n6685), .A2(n4628), .ZN(n6301) );
  INV_X1 U5548 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n7113) );
  INV_X1 U5549 ( .A(EAX_REG_23__SCAN_IN), .ZN(n7043) );
  INV_X1 U5550 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n7098) );
  OAI222_X1 U5551 ( .A1(n6302), .A2(n7113), .B1(n6287), .B2(n7043), .C1(n6301), 
        .C2(n7098), .ZN(U2900) );
  INV_X1 U5552 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7057) );
  INV_X1 U5553 ( .A(n4535), .ZN(n4539) );
  NAND2_X1 U5554 ( .A1(n3452), .A2(n6702), .ZN(n4536) );
  NAND3_X1 U5555 ( .A1(n4536), .A2(n4640), .A3(n4700), .ZN(n4537) );
  OAI211_X1 U5556 ( .C1(n4540), .C2(n4539), .A(n4538), .B(n4537), .ZN(n4541)
         );
  NAND2_X1 U5557 ( .A1(n4541), .A2(n6673), .ZN(n4548) );
  NAND3_X1 U5558 ( .A1(n4492), .A2(n4542), .A3(n6795), .ZN(n4544) );
  NAND3_X1 U5559 ( .A1(n4544), .A2(n3448), .A3(n4543), .ZN(n4545) );
  NAND2_X1 U5560 ( .A1(n4545), .A2(n3462), .ZN(n4546) );
  INV_X1 U5561 ( .A(n4549), .ZN(n4550) );
  NAND2_X1 U5562 ( .A1(n4561), .A2(n4550), .ZN(n4868) );
  NAND2_X1 U5563 ( .A1(n5792), .A2(n4868), .ZN(n5948) );
  NAND2_X1 U5564 ( .A1(n7057), .A2(n5948), .ZN(n4869) );
  XOR2_X1 U5565 ( .A(n4551), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4568) );
  AOI22_X1 U5566 ( .A1(n4492), .A2(n4861), .B1(n4552), .B2(n3419), .ZN(n4553)
         );
  NAND3_X1 U5567 ( .A1(n4554), .A2(n4553), .A3(n3198), .ZN(n4555) );
  INV_X1 U5568 ( .A(n4556), .ZN(n4557) );
  OAI21_X1 U5569 ( .B1(n4558), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4557), 
        .ZN(n5268) );
  NAND2_X1 U5570 ( .A1(n4552), .A2(n3573), .ZN(n4559) );
  NAND2_X1 U5571 ( .A1(n6677), .A2(n4559), .ZN(n4560) );
  NAND2_X1 U5572 ( .A1(n4561), .A2(n6654), .ZN(n5945) );
  INV_X1 U5573 ( .A(n5945), .ZN(n6495) );
  NOR2_X1 U5574 ( .A1(n4561), .A2(n6471), .ZN(n4870) );
  OAI21_X1 U5575 ( .B1(n6495), .B2(n4870), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4562) );
  NAND2_X1 U5576 ( .A1(n6471), .A2(REIP_REG_0__SCAN_IN), .ZN(n4570) );
  OAI211_X1 U5577 ( .C1(n5268), .C2(n6463), .A(n4562), .B(n4570), .ZN(n4563)
         );
  AOI21_X1 U5578 ( .B1(n4568), .B2(n6477), .A(n4563), .ZN(n4564) );
  NAND2_X1 U5579 ( .A1(n4869), .A2(n4564), .ZN(U3018) );
  OAI21_X1 U5580 ( .B1(n4567), .B2(n4566), .A(n4565), .ZN(n6286) );
  NAND2_X1 U5581 ( .A1(n4568), .A2(n6402), .ZN(n4574) );
  NAND2_X1 U5582 ( .A1(n4569), .A2(n5780), .ZN(n4572) );
  INV_X1 U5583 ( .A(n4570), .ZN(n4571) );
  AOI21_X1 U5584 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4572), .A(n4571), 
        .ZN(n4573) );
  OAI211_X1 U5585 ( .C1(n6286), .C2(n5766), .A(n4574), .B(n4573), .ZN(U2986)
         );
  AOI22_X1 U5586 ( .A1(n6796), .A2(UWORD_REG_14__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5587 ( .B1(n4140), .B2(n6287), .A(n4575), .ZN(U2893) );
  INV_X1 U5588 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6312) );
  AOI22_X1 U5589 ( .A1(n6796), .A2(UWORD_REG_0__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4576) );
  OAI21_X1 U5590 ( .B1(n6312), .B2(n6287), .A(n4576), .ZN(U2907) );
  INV_X1 U5591 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6315) );
  AOI22_X1 U5592 ( .A1(n6796), .A2(UWORD_REG_1__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5593 ( .B1(n6315), .B2(n6287), .A(n4577), .ZN(U2906) );
  INV_X1 U5594 ( .A(EAX_REG_18__SCAN_IN), .ZN(n7122) );
  AOI22_X1 U5595 ( .A1(n6796), .A2(UWORD_REG_2__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5596 ( .B1(n7122), .B2(n6287), .A(n4578), .ZN(U2905) );
  AOI22_X1 U5597 ( .A1(n4587), .A2(UWORD_REG_3__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5598 ( .B1(n3922), .B2(n6287), .A(n4579), .ZN(U2904) );
  INV_X1 U5599 ( .A(EAX_REG_20__SCAN_IN), .ZN(n7146) );
  AOI22_X1 U5600 ( .A1(n4587), .A2(UWORD_REG_4__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4580) );
  OAI21_X1 U5601 ( .B1(n7146), .B2(n6287), .A(n4580), .ZN(U2903) );
  INV_X1 U5602 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U5603 ( .A1(n4587), .A2(UWORD_REG_5__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4581) );
  OAI21_X1 U5604 ( .B1(n6320), .B2(n6287), .A(n4581), .ZN(U2902) );
  AOI22_X1 U5605 ( .A1(n6796), .A2(UWORD_REG_12__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4582) );
  OAI21_X1 U5606 ( .B1(n4094), .B2(n6287), .A(n4582), .ZN(U2895) );
  AOI22_X1 U5607 ( .A1(n4587), .A2(UWORD_REG_8__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4583) );
  OAI21_X1 U5608 ( .B1(n4018), .B2(n6287), .A(n4583), .ZN(U2899) );
  INV_X1 U5609 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U5610 ( .A1(n4587), .A2(UWORD_REG_9__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4584) );
  OAI21_X1 U5611 ( .B1(n6932), .B2(n6287), .A(n4584), .ZN(U2898) );
  INV_X1 U5612 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6330) );
  AOI22_X1 U5613 ( .A1(n4587), .A2(UWORD_REG_10__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4585) );
  OAI21_X1 U5614 ( .B1(n6330), .B2(n6287), .A(n4585), .ZN(U2897) );
  INV_X1 U5615 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6333) );
  AOI22_X1 U5616 ( .A1(n6796), .A2(UWORD_REG_11__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4586) );
  OAI21_X1 U5617 ( .B1(n6333), .B2(n6287), .A(n4586), .ZN(U2896) );
  INV_X1 U5618 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U5619 ( .A1(n4587), .A2(UWORD_REG_6__SCAN_IN), .B1(
        DATAO_REG_22__SCAN_IN), .B2(n6308), .ZN(n4588) );
  OAI21_X1 U5620 ( .B1(n7007), .B2(n6287), .A(n4588), .ZN(U2901) );
  NAND2_X1 U5621 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7090), .ZN(n4620) );
  INV_X1 U5622 ( .A(n4593), .ZN(n4619) );
  NAND2_X1 U5623 ( .A1(n3200), .A2(n6652), .ZN(n4603) );
  INV_X1 U5624 ( .A(n4638), .ZN(n4590) );
  OR2_X1 U5625 ( .A1(n4656), .A2(n4590), .ZN(n4612) );
  MUX2_X1 U5626 ( .A(n4592), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4591), 
        .Z(n4594) );
  NOR2_X1 U5627 ( .A1(n4594), .A2(n4593), .ZN(n4601) );
  AOI21_X1 U5628 ( .B1(n4591), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3632), 
        .ZN(n4595) );
  NOR2_X1 U5629 ( .A1(n4596), .A2(n4595), .ZN(n6772) );
  NAND2_X1 U5630 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4597) );
  XNOR2_X1 U5631 ( .A(n4597), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4598)
         );
  NAND2_X1 U5632 ( .A1(n6654), .A2(n4598), .ZN(n4599) );
  OAI21_X1 U5633 ( .B1(n6772), .B2(n4609), .A(n4599), .ZN(n4600) );
  AOI21_X1 U5634 ( .B1(n4612), .B2(n4601), .A(n4600), .ZN(n4602) );
  NAND2_X1 U5635 ( .A1(n4603), .A2(n4602), .ZN(n6770) );
  MUX2_X1 U5636 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6770), .S(n6655), 
        .Z(n6670) );
  OR2_X1 U5637 ( .A1(n4605), .A2(n4606), .ZN(n4614) );
  XNOR2_X1 U5638 ( .A(n4591), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4611)
         );
  XNOR2_X1 U5639 ( .A(n3604), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4607)
         );
  NAND2_X1 U5640 ( .A1(n6654), .A2(n4607), .ZN(n4608) );
  OAI21_X1 U5641 ( .B1(n4611), .B2(n4609), .A(n4608), .ZN(n4610) );
  AOI21_X1 U5642 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4613) );
  NAND2_X1 U5643 ( .A1(n4614), .A2(n4613), .ZN(n5450) );
  NAND2_X1 U5644 ( .A1(n5450), .A2(n6655), .ZN(n4617) );
  NAND2_X1 U5645 ( .A1(n4615), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5646 ( .A1(n4617), .A2(n4616), .ZN(n6665) );
  NAND3_X1 U5647 ( .A1(n6670), .A2(n6776), .A3(n6665), .ZN(n4618) );
  OAI21_X1 U5648 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n6650) );
  INV_X1 U5649 ( .A(n4621), .ZN(n4622) );
  NAND2_X1 U5650 ( .A1(n6650), .A2(n4622), .ZN(n4626) );
  INV_X1 U5651 ( .A(n5099), .ZN(n6501) );
  NOR2_X1 U5652 ( .A1(n3611), .A2(n6501), .ZN(n4623) );
  XNOR2_X1 U5653 ( .A(n4623), .B(n6115), .ZN(n5551) );
  INV_X1 U5654 ( .A(n4499), .ZN(n4624) );
  AND2_X1 U5655 ( .A1(n5551), .A2(n4624), .ZN(n6114) );
  AOI211_X1 U5656 ( .C1(n6776), .C2(n6655), .A(FLUSH_REG_SCAN_IN), .B(n6115), 
        .ZN(n4625) );
  AOI21_X1 U5657 ( .B1(n6114), .B2(n6776), .A(n4625), .ZN(n6648) );
  NAND2_X1 U5658 ( .A1(n4626), .A2(n6648), .ZN(n4630) );
  NOR2_X1 U5659 ( .A1(n4630), .A2(FLUSH_REG_SCAN_IN), .ZN(n4627) );
  INV_X1 U5660 ( .A(n6694), .ZN(n6799) );
  OAI21_X1 U5661 ( .B1(n4627), .B2(n6767), .A(n5283), .ZN(n6498) );
  INV_X1 U5662 ( .A(n4628), .ZN(n4629) );
  OR2_X1 U5663 ( .A1(n4630), .A2(n4629), .ZN(n6681) );
  INV_X1 U5664 ( .A(n6681), .ZN(n4632) );
  NOR2_X1 U5665 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6776), .ZN(n5971) );
  OAI22_X1 U5666 ( .A1(n5108), .A2(n6559), .B1(n3595), .B2(n5971), .ZN(n4631)
         );
  OAI21_X1 U5667 ( .B1(n4632), .B2(n4631), .A(n6498), .ZN(n4633) );
  OAI21_X1 U5668 ( .B1(n6498), .B2(n6504), .A(n4633), .ZN(U3465) );
  NOR2_X1 U5669 ( .A1(n4635), .A2(n4634), .ZN(n4636) );
  OR2_X1 U5670 ( .A1(n4637), .A2(n4636), .ZN(n4863) );
  OR2_X1 U5671 ( .A1(n4639), .A2(n4638), .ZN(n4649) );
  NAND2_X1 U5672 ( .A1(n6673), .A2(n4640), .ZN(n4646) );
  INV_X1 U5673 ( .A(n4641), .ZN(n4645) );
  NOR2_X1 U5674 ( .A1(n3483), .A2(n6682), .ZN(n4643) );
  NOR2_X1 U5675 ( .A1(n3585), .A2(n4700), .ZN(n4642) );
  NAND4_X1 U5676 ( .A1(n4645), .A2(n4644), .A3(n4643), .A4(n4642), .ZN(n4658)
         );
  OAI22_X1 U5677 ( .A1(n3198), .A2(n4646), .B1(n3491), .B2(n4658), .ZN(n4647)
         );
  INV_X1 U5678 ( .A(n4647), .ZN(n4648) );
  NAND2_X1 U5679 ( .A1(n3450), .A2(n3585), .ZN(n4651) );
  INV_X1 U5680 ( .A(n4651), .ZN(n4652) );
  INV_X1 U5681 ( .A(DATAI_1_), .ZN(n4711) );
  INV_X1 U5682 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6342) );
  OAI222_X1 U5683 ( .A1(n4863), .A2(n6054), .B1(n6284), .B2(n4711), .C1(n6285), 
        .C2(n6342), .ZN(U2890) );
  INV_X1 U5684 ( .A(n4654), .ZN(n4666) );
  OAI21_X1 U5685 ( .B1(n4655), .B2(n4653), .A(n4666), .ZN(n6399) );
  INV_X1 U5686 ( .A(DATAI_2_), .ZN(n4701) );
  INV_X1 U5687 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6345) );
  OAI222_X1 U5688 ( .A1(n6399), .A2(n6054), .B1(n6284), .B2(n4701), .C1(n6285), 
        .C2(n6345), .ZN(U2889) );
  NAND3_X1 U5689 ( .A1(n4657), .A2(n4656), .A3(n6673), .ZN(n4661) );
  INV_X1 U5690 ( .A(n4658), .ZN(n4659) );
  NAND2_X1 U5691 ( .A1(n4659), .A2(n4861), .ZN(n4660) );
  INV_X1 U5692 ( .A(n3585), .ZN(n5628) );
  NAND2_X2 U5693 ( .A1(n6272), .A2(n5628), .ZN(n5627) );
  AND2_X1 U5694 ( .A1(n6272), .A2(n3585), .ZN(n6270) );
  INV_X2 U5695 ( .A(n6270), .ZN(n5626) );
  OAI222_X1 U5696 ( .A1(n5268), .A2(n5627), .B1(n6272), .B2(n5270), .C1(n6286), 
        .C2(n5626), .ZN(U2859) );
  OAI21_X1 U5697 ( .B1(n4664), .B2(n4663), .A(n3272), .ZN(n6470) );
  OAI222_X1 U5698 ( .A1(n6470), .A2(n5627), .B1(n4665), .B2(n6272), .C1(n5626), 
        .C2(n6399), .ZN(U2857) );
  XNOR2_X1 U5699 ( .A(n4666), .B(n4688), .ZN(n6391) );
  INV_X1 U5700 ( .A(n6391), .ZN(n4668) );
  INV_X1 U5701 ( .A(DATAI_3_), .ZN(n4727) );
  INV_X1 U5702 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6348) );
  OAI222_X1 U5703 ( .A1(n4668), .A2(n6054), .B1(n6284), .B2(n4727), .C1(n6285), 
        .C2(n6348), .ZN(U2888) );
  OAI21_X1 U5704 ( .B1(n4662), .B2(n4667), .A(n4879), .ZN(n6462) );
  INV_X1 U5705 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6232) );
  OAI222_X1 U5706 ( .A1(n6462), .A2(n5627), .B1(n6272), .B2(n6232), .C1(n5626), 
        .C2(n4668), .ZN(U2856) );
  INV_X1 U5707 ( .A(n3595), .ZN(n6653) );
  AND2_X1 U5708 ( .A1(n3200), .A2(n6653), .ZN(n4952) );
  NOR2_X1 U5709 ( .A1(n4605), .A2(n4512), .ZN(n6512) );
  INV_X1 U5710 ( .A(n4781), .ZN(n4669) );
  AOI21_X1 U5711 ( .B1(n4952), .B2(n6512), .A(n4669), .ZN(n4680) );
  INV_X1 U5712 ( .A(n4680), .ZN(n4670) );
  NAND2_X1 U5713 ( .A1(n4670), .A2(n6567), .ZN(n4672) );
  NAND2_X1 U5714 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4683), .ZN(n4671) );
  INV_X1 U5715 ( .A(DATAI_0_), .ZN(n6283) );
  NAND2_X1 U5716 ( .A1(n6400), .A2(DATAI_24_), .ZN(n6632) );
  INV_X1 U5717 ( .A(n6632), .ZN(n6517) );
  INV_X1 U5718 ( .A(n3641), .ZN(n4674) );
  INV_X1 U5719 ( .A(n4859), .ZN(n4827) );
  INV_X1 U5720 ( .A(DATAI_16_), .ZN(n7031) );
  NOR2_X1 U5721 ( .A1(n5766), .A2(n7031), .ZN(n6569) );
  INV_X1 U5722 ( .A(n6569), .ZN(n6627) );
  NAND2_X1 U5723 ( .A1(n4754), .A2(n3448), .ZN(n6626) );
  OAI22_X1 U5724 ( .A1(n4769), .A2(n6627), .B1(n6626), .B2(n4781), .ZN(n4678)
         );
  AOI21_X1 U5725 ( .B1(n6517), .B2(n4827), .A(n4678), .ZN(n4685) );
  AND2_X1 U5726 ( .A1(n6567), .A2(n6124), .ZN(n6509) );
  INV_X1 U5727 ( .A(n6509), .ZN(n5974) );
  OAI21_X1 U5728 ( .B1(n4679), .B2(n5766), .A(n5974), .ZN(n4681) );
  NAND2_X1 U5729 ( .A1(n4681), .A2(n4680), .ZN(n4682) );
  OAI211_X1 U5730 ( .C1(n6567), .C2(n4683), .A(n4682), .B(n6565), .ZN(n4779)
         );
  NAND2_X1 U5731 ( .A1(n4779), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4684)
         );
  OAI211_X1 U5732 ( .C1(n4780), .C2(n6572), .A(n4685), .B(n4684), .ZN(U3140)
         );
  AOI21_X1 U5733 ( .B1(n4654), .B2(n4688), .A(n4687), .ZN(n4689) );
  NOR2_X1 U5734 ( .A1(n4686), .A2(n4689), .ZN(n5550) );
  INV_X1 U5735 ( .A(n5550), .ZN(n4882) );
  INV_X1 U5736 ( .A(DATAI_4_), .ZN(n4706) );
  INV_X1 U5737 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6351) );
  OAI222_X1 U5738 ( .A1(n4882), .A2(n6054), .B1(n6284), .B2(n4706), .C1(n6285), 
        .C2(n6351), .ZN(U2887) );
  INV_X1 U5739 ( .A(DATAI_29_), .ZN(n4690) );
  NOR2_X1 U5740 ( .A1(n5766), .A2(n4690), .ZN(n6600) );
  INV_X1 U5741 ( .A(n6600), .ZN(n5290) );
  NAND2_X1 U5742 ( .A1(n4779), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4694)
         );
  NAND2_X1 U5743 ( .A1(n6400), .A2(DATAI_21_), .ZN(n6597) );
  INV_X1 U5744 ( .A(n6597), .ZN(n5288) );
  NAND2_X1 U5745 ( .A1(n4754), .A2(n4691), .ZN(n6598) );
  INV_X1 U5746 ( .A(DATAI_5_), .ZN(n7078) );
  NOR2_X1 U5747 ( .A1(n7078), .A2(n5283), .ZN(n6538) );
  OAI22_X1 U5748 ( .A1(n6598), .A2(n4781), .B1(n4780), .B2(n6603), .ZN(n4692)
         );
  AOI21_X1 U5749 ( .B1(n5288), .B2(n4783), .A(n4692), .ZN(n4693) );
  OAI211_X1 U5750 ( .C1(n4859), .C2(n5290), .A(n4694), .B(n4693), .ZN(U3145)
         );
  INV_X1 U5751 ( .A(DATAI_30_), .ZN(n4695) );
  NOR2_X1 U5752 ( .A1(n5766), .A2(n4695), .ZN(n6609) );
  INV_X1 U5753 ( .A(n6609), .ZN(n5295) );
  NAND2_X1 U5754 ( .A1(n4779), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4698)
         );
  NAND2_X1 U5755 ( .A1(n6400), .A2(DATAI_22_), .ZN(n6604) );
  INV_X1 U5756 ( .A(n6604), .ZN(n5293) );
  NAND2_X1 U5757 ( .A1(n4754), .A2(n3393), .ZN(n6606) );
  INV_X1 U5758 ( .A(DATAI_6_), .ZN(n4790) );
  NOR2_X1 U5759 ( .A1(n4790), .A2(n5283), .ZN(n6542) );
  OAI22_X1 U5760 ( .A1(n6606), .A2(n4781), .B1(n4780), .B2(n6612), .ZN(n4696)
         );
  AOI21_X1 U5761 ( .B1(n5293), .B2(n4783), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5762 ( .C1(n4859), .C2(n5295), .A(n4698), .B(n4697), .ZN(U3146)
         );
  INV_X1 U5763 ( .A(DATAI_26_), .ZN(n4699) );
  NOR2_X1 U5764 ( .A1(n5766), .A2(n4699), .ZN(n6583) );
  INV_X1 U5765 ( .A(n6583), .ZN(n5303) );
  NAND2_X1 U5766 ( .A1(n4779), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4704)
         );
  NAND2_X1 U5767 ( .A1(n6400), .A2(DATAI_18_), .ZN(n6580) );
  INV_X1 U5768 ( .A(n6580), .ZN(n5301) );
  NAND2_X1 U5769 ( .A1(n4754), .A2(n4700), .ZN(n6581) );
  NOR2_X1 U5770 ( .A1(n4701), .A2(n5283), .ZN(n6526) );
  OAI22_X1 U5771 ( .A1(n6581), .A2(n4781), .B1(n4780), .B2(n6586), .ZN(n4702)
         );
  AOI21_X1 U5772 ( .B1(n5301), .B2(n4783), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5773 ( .C1(n4859), .C2(n5303), .A(n4704), .B(n4703), .ZN(U3142)
         );
  INV_X1 U5774 ( .A(DATAI_28_), .ZN(n4705) );
  NOR2_X1 U5775 ( .A1(n5766), .A2(n4705), .ZN(n6594) );
  INV_X1 U5776 ( .A(n6594), .ZN(n7209) );
  NAND2_X1 U5777 ( .A1(n4779), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4709)
         );
  NAND2_X1 U5778 ( .A1(n6400), .A2(DATAI_20_), .ZN(n6592) );
  INV_X1 U5779 ( .A(n6592), .ZN(n7206) );
  NAND2_X1 U5780 ( .A1(n4754), .A2(n3419), .ZN(n7203) );
  NOR2_X1 U5781 ( .A1(n4706), .A2(n5283), .ZN(n6534) );
  OAI22_X1 U5782 ( .A1(n7203), .A2(n4781), .B1(n4780), .B2(n7200), .ZN(n4707)
         );
  AOI21_X1 U5783 ( .B1(n7206), .B2(n4783), .A(n4707), .ZN(n4708) );
  OAI211_X1 U5784 ( .C1(n4859), .C2(n7209), .A(n4709), .B(n4708), .ZN(U3144)
         );
  NAND2_X1 U5785 ( .A1(n6400), .A2(DATAI_25_), .ZN(n6573) );
  NAND2_X1 U5786 ( .A1(n4779), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4714)
         );
  INV_X1 U5787 ( .A(DATAI_17_), .ZN(n4710) );
  NOR2_X1 U5788 ( .A1(n5766), .A2(n4710), .ZN(n6576) );
  NAND2_X1 U5789 ( .A1(n4754), .A2(n3452), .ZN(n6574) );
  NOR2_X1 U5790 ( .A1(n4711), .A2(n5283), .ZN(n6520) );
  OAI22_X1 U5791 ( .A1(n6574), .A2(n4781), .B1(n4780), .B2(n6579), .ZN(n4712)
         );
  AOI21_X1 U5792 ( .B1(n6576), .B2(n4783), .A(n4712), .ZN(n4713) );
  OAI211_X1 U5793 ( .C1(n4859), .C2(n6573), .A(n4714), .B(n4713), .ZN(U3141)
         );
  INV_X1 U5794 ( .A(n4673), .ZN(n5024) );
  OAI21_X1 U5795 ( .B1(n5197), .B2(n6559), .A(n5974), .ZN(n5190) );
  NAND2_X1 U5796 ( .A1(n4605), .A2(n4512), .ZN(n5147) );
  OR2_X1 U5797 ( .A1(n3200), .A2(n5147), .ZN(n5186) );
  OAI211_X1 U5798 ( .C1(n6509), .C2(n4769), .A(n5190), .B(n5186), .ZN(n4718)
         );
  NAND3_X1 U5799 ( .A1(n6669), .A2(n6662), .A3(n6658), .ZN(n5189) );
  NOR2_X1 U5800 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5189), .ZN(n4744)
         );
  INV_X1 U5801 ( .A(n4744), .ZN(n4755) );
  INV_X1 U5802 ( .A(n5283), .ZN(n4753) );
  OAI21_X1 U5803 ( .B1(n3304), .B2(n6680), .A(n4753), .ZN(n4915) );
  AOI21_X1 U5804 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4755), .A(n4915), .ZN(
        n4717) );
  INV_X1 U5805 ( .A(n4720), .ZN(n4716) );
  NAND2_X1 U5806 ( .A1(n4716), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6503) );
  INV_X1 U5807 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4725) );
  NOR2_X2 U5808 ( .A1(n4719), .A2(n5196), .ZN(n5223) );
  INV_X1 U5809 ( .A(n6606), .ZN(n6543) );
  AND2_X1 U5810 ( .A1(n4720), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U5811 ( .A1(n5339), .A2(n3304), .ZN(n4721) );
  OAI21_X1 U5812 ( .B1(n5186), .B2(n6559), .A(n4721), .ZN(n4757) );
  AOI22_X1 U5813 ( .A1(n6543), .A2(n4744), .B1(n6542), .B2(n4757), .ZN(n4722)
         );
  OAI21_X1 U5814 ( .B1(n5295), .B2(n4769), .A(n4722), .ZN(n4723) );
  AOI21_X1 U5815 ( .B1(n5293), .B2(n5223), .A(n4723), .ZN(n4724) );
  OAI21_X1 U5816 ( .B1(n4761), .B2(n4725), .A(n4724), .ZN(U3026) );
  INV_X1 U5817 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4731) );
  INV_X1 U5818 ( .A(DATAI_19_), .ZN(n4726) );
  NOR2_X1 U5819 ( .A1(n5766), .A2(n4726), .ZN(n6588) );
  NAND2_X1 U5820 ( .A1(n6400), .A2(DATAI_27_), .ZN(n6643) );
  NAND2_X1 U5821 ( .A1(n4754), .A2(n3483), .ZN(n6634) );
  INV_X1 U5822 ( .A(n6634), .ZN(n6530) );
  NOR2_X1 U5823 ( .A1(n4727), .A2(n5283), .ZN(n6638) );
  AOI22_X1 U5824 ( .A1(n6530), .A2(n4744), .B1(n6638), .B2(n4757), .ZN(n4728)
         );
  OAI21_X1 U5825 ( .B1(n6643), .B2(n4769), .A(n4728), .ZN(n4729) );
  AOI21_X1 U5826 ( .B1(n6588), .B2(n5223), .A(n4729), .ZN(n4730) );
  OAI21_X1 U5827 ( .B1(n4761), .B2(n4731), .A(n4730), .ZN(U3023) );
  INV_X1 U5828 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4735) );
  INV_X1 U5829 ( .A(n6581), .ZN(n6527) );
  AOI22_X1 U5830 ( .A1(n6527), .A2(n4744), .B1(n6526), .B2(n4757), .ZN(n4732)
         );
  OAI21_X1 U5831 ( .B1(n5303), .B2(n4769), .A(n4732), .ZN(n4733) );
  AOI21_X1 U5832 ( .B1(n5301), .B2(n5223), .A(n4733), .ZN(n4734) );
  OAI21_X1 U5833 ( .B1(n4761), .B2(n4735), .A(n4734), .ZN(U3022) );
  INV_X1 U5834 ( .A(n6574), .ZN(n6521) );
  AOI22_X1 U5835 ( .A1(n6521), .A2(n4744), .B1(n6520), .B2(n4757), .ZN(n4736)
         );
  OAI21_X1 U5836 ( .B1(n6573), .B2(n4769), .A(n4736), .ZN(n4737) );
  AOI21_X1 U5837 ( .B1(n6576), .B2(n5223), .A(n4737), .ZN(n4738) );
  OAI21_X1 U5838 ( .B1(n4761), .B2(n4739), .A(n4738), .ZN(U3021) );
  INV_X1 U5839 ( .A(n7203), .ZN(n6535) );
  AOI22_X1 U5840 ( .A1(n6535), .A2(n4744), .B1(n6534), .B2(n4757), .ZN(n4740)
         );
  OAI21_X1 U5841 ( .B1(n7209), .B2(n4769), .A(n4740), .ZN(n4741) );
  AOI21_X1 U5842 ( .B1(n7206), .B2(n5223), .A(n4741), .ZN(n4742) );
  OAI21_X1 U5843 ( .B1(n4761), .B2(n4743), .A(n4742), .ZN(U3024) );
  INV_X1 U5844 ( .A(n6598), .ZN(n6539) );
  AOI22_X1 U5845 ( .A1(n6539), .A2(n4744), .B1(n6538), .B2(n4757), .ZN(n4745)
         );
  OAI21_X1 U5846 ( .B1(n5290), .B2(n4769), .A(n4745), .ZN(n4746) );
  AOI21_X1 U5847 ( .B1(n5288), .B2(n5223), .A(n4746), .ZN(n4747) );
  OAI21_X1 U5848 ( .B1(n4761), .B2(n4748), .A(n4747), .ZN(U3025) );
  OAI22_X1 U5849 ( .A1(n4769), .A2(n6632), .B1(n6626), .B2(n4755), .ZN(n4749)
         );
  AOI21_X1 U5850 ( .B1(n6629), .B2(n4757), .A(n4749), .ZN(n4751) );
  NAND2_X1 U5851 ( .A1(n5223), .A2(n6569), .ZN(n4750) );
  OAI211_X1 U5852 ( .C1(n4761), .C2(n4752), .A(n4751), .B(n4750), .ZN(U3020)
         );
  INV_X1 U5853 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U5854 ( .A1(DATAI_7_), .A2(n4753), .ZN(n6623) );
  NAND2_X1 U5855 ( .A1(n6400), .A2(DATAI_31_), .ZN(n6613) );
  NAND2_X1 U5856 ( .A1(n4754), .A2(n3585), .ZN(n6616) );
  OAI22_X1 U5857 ( .A1(n4769), .A2(n6613), .B1(n6616), .B2(n4755), .ZN(n4756)
         );
  AOI21_X1 U5858 ( .B1(n6549), .B2(n4757), .A(n4756), .ZN(n4759) );
  INV_X1 U5859 ( .A(DATAI_23_), .ZN(n7012) );
  NOR2_X1 U5860 ( .A1(n5766), .A2(n7012), .ZN(n6619) );
  NAND2_X1 U5861 ( .A1(n5223), .A2(n6619), .ZN(n4758) );
  OAI211_X1 U5862 ( .C1(n4761), .C2(n4760), .A(n4759), .B(n4758), .ZN(U3027)
         );
  XNOR2_X1 U5863 ( .A(n4762), .B(n4763), .ZN(n6490) );
  INV_X1 U5864 ( .A(n4863), .ZN(n6254) );
  INV_X1 U5865 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U5866 ( .A1(n6461), .A2(n6998), .ZN(n6485) );
  AOI21_X1 U5867 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6485), 
        .ZN(n4764) );
  OAI21_X1 U5868 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6406), .A(n4764), 
        .ZN(n4765) );
  AOI21_X1 U5869 ( .B1(n6254), .B2(n6400), .A(n4765), .ZN(n4766) );
  OAI21_X1 U5870 ( .B1(n6490), .B2(n6125), .A(n4766), .ZN(U2985) );
  INV_X1 U5871 ( .A(n4767), .ZN(n4768) );
  XNOR2_X1 U5872 ( .A(n4686), .B(n4768), .ZN(n6382) );
  INV_X1 U5873 ( .A(n6382), .ZN(n4794) );
  INV_X1 U5874 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6355) );
  OAI222_X1 U5875 ( .A1(n6054), .A2(n4794), .B1(n6284), .B2(n7078), .C1(n6285), 
        .C2(n6355), .ZN(U2886) );
  INV_X1 U5876 ( .A(n6619), .ZN(n6555) );
  OAI22_X1 U5877 ( .A1(n4769), .A2(n6555), .B1(n6616), .B2(n4781), .ZN(n4771)
         );
  OAI22_X1 U5878 ( .A1(n6623), .A2(n4780), .B1(n6613), .B2(n4859), .ZN(n4770)
         );
  AOI211_X1 U5879 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4779), .A(n4771), 
        .B(n4770), .ZN(n4772) );
  INV_X1 U5880 ( .A(n4772), .ZN(U3147) );
  OAI21_X1 U5881 ( .B1(n4775), .B2(n4774), .A(n4773), .ZN(n6452) );
  AOI22_X1 U5882 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6471), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4776) );
  OAI21_X1 U5883 ( .B1(n5555), .B2(n6406), .A(n4776), .ZN(n4777) );
  AOI21_X1 U5884 ( .B1(n5550), .B2(n6400), .A(n4777), .ZN(n4778) );
  OAI21_X1 U5885 ( .B1(n6452), .B2(n6125), .A(n4778), .ZN(U2982) );
  NAND2_X1 U5886 ( .A1(n4779), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4785)
         );
  OAI22_X1 U5887 ( .A1(n6634), .A2(n4781), .B1(n4780), .B2(n6591), .ZN(n4782)
         );
  AOI21_X1 U5888 ( .B1(n6588), .B2(n4783), .A(n4782), .ZN(n4784) );
  OAI211_X1 U5889 ( .C1(n4859), .C2(n6643), .A(n4785), .B(n4784), .ZN(U3143)
         );
  AOI21_X1 U5890 ( .B1(n4686), .B2(n4767), .A(n4788), .ZN(n4789) );
  OR2_X1 U5891 ( .A1(n4787), .A2(n4789), .ZN(n5254) );
  OAI222_X1 U5892 ( .A1(n5254), .A2(n6054), .B1(n6284), .B2(n4790), .C1(n6285), 
        .C2(n3702), .ZN(U2885) );
  NAND2_X1 U5893 ( .A1(n4877), .A2(n4791), .ZN(n4792) );
  NAND2_X1 U5894 ( .A1(n4883), .A2(n4792), .ZN(n6225) );
  INV_X1 U5895 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4793) );
  OAI222_X1 U5896 ( .A1(n6225), .A2(n5627), .B1(n5626), .B2(n4794), .C1(n4793), 
        .C2(n6272), .ZN(U2854) );
  NAND2_X1 U5897 ( .A1(n4676), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5968) );
  OAI21_X1 U5898 ( .B1(n5022), .B2(n5968), .A(n6567), .ZN(n4800) );
  INV_X1 U5899 ( .A(n4512), .ZN(n6241) );
  NAND2_X1 U5900 ( .A1(n4605), .A2(n6241), .ZN(n5026) );
  INV_X1 U5901 ( .A(n5026), .ZN(n4795) );
  AND2_X1 U5902 ( .A1(n4795), .A2(n3200), .ZN(n5342) );
  NOR2_X1 U5903 ( .A1(n5027), .A2(n6669), .ZN(n6625) );
  AOI21_X1 U5904 ( .B1(n5342), .B2(n6653), .A(n6625), .ZN(n4796) );
  NAND3_X1 U5905 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6662), .ZN(n5341) );
  OAI22_X1 U5906 ( .A1(n4800), .A2(n4796), .B1(n5341), .B2(n6680), .ZN(n6637)
         );
  INV_X1 U5907 ( .A(n6637), .ZN(n4819) );
  INV_X1 U5908 ( .A(n4796), .ZN(n4799) );
  INV_X1 U5909 ( .A(n6565), .ZN(n4797) );
  AOI21_X1 U5910 ( .B1(n6559), .B2(n5341), .A(n4797), .ZN(n4798) );
  OAI21_X1 U5911 ( .B1(n4800), .B2(n4799), .A(n4798), .ZN(n6639) );
  NAND2_X1 U5912 ( .A1(n4676), .A2(n5108), .ZN(n6499) );
  NAND2_X1 U5913 ( .A1(n4676), .A2(n5196), .ZN(n5138) );
  AOI22_X1 U5914 ( .A1(n5019), .A2(n6619), .B1(n6547), .B2(n6625), .ZN(n4801)
         );
  OAI21_X1 U5915 ( .B1(n6613), .B2(n6642), .A(n4801), .ZN(n4802) );
  AOI21_X1 U5916 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6639), .A(n4802), 
        .ZN(n4803) );
  OAI21_X1 U5917 ( .B1(n4819), .B2(n6623), .A(n4803), .ZN(U3115) );
  AOI22_X1 U5918 ( .A1(n5019), .A2(n6576), .B1(n6521), .B2(n6625), .ZN(n4804)
         );
  OAI21_X1 U5919 ( .B1(n6573), .B2(n6642), .A(n4804), .ZN(n4805) );
  AOI21_X1 U5920 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(n6639), .A(n4805), 
        .ZN(n4806) );
  OAI21_X1 U5921 ( .B1(n4819), .B2(n6579), .A(n4806), .ZN(U3109) );
  AOI22_X1 U5922 ( .A1(n5019), .A2(n5293), .B1(n6543), .B2(n6625), .ZN(n4807)
         );
  OAI21_X1 U5923 ( .B1(n5295), .B2(n6642), .A(n4807), .ZN(n4808) );
  AOI21_X1 U5924 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6639), .A(n4808), 
        .ZN(n4809) );
  OAI21_X1 U5925 ( .B1(n4819), .B2(n6612), .A(n4809), .ZN(U3114) );
  AOI22_X1 U5926 ( .A1(n5019), .A2(n7206), .B1(n6535), .B2(n6625), .ZN(n4810)
         );
  OAI21_X1 U5927 ( .B1(n7209), .B2(n6642), .A(n4810), .ZN(n4811) );
  AOI21_X1 U5928 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6639), .A(n4811), 
        .ZN(n4812) );
  OAI21_X1 U5929 ( .B1(n4819), .B2(n7200), .A(n4812), .ZN(U3112) );
  AOI22_X1 U5930 ( .A1(n5019), .A2(n5288), .B1(n6539), .B2(n6625), .ZN(n4813)
         );
  OAI21_X1 U5931 ( .B1(n5290), .B2(n6642), .A(n4813), .ZN(n4814) );
  AOI21_X1 U5932 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n6639), .A(n4814), 
        .ZN(n4815) );
  OAI21_X1 U5933 ( .B1(n4819), .B2(n6603), .A(n4815), .ZN(U3113) );
  AOI22_X1 U5934 ( .A1(n5019), .A2(n5301), .B1(n6527), .B2(n6625), .ZN(n4816)
         );
  OAI21_X1 U5935 ( .B1(n5303), .B2(n6642), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5936 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n6639), .A(n4817), 
        .ZN(n4818) );
  OAI21_X1 U5937 ( .B1(n4819), .B2(n6586), .A(n4818), .ZN(U3110) );
  NAND3_X1 U5938 ( .A1(n4978), .A2(n4859), .A3(n6567), .ZN(n4821) );
  AOI22_X1 U5939 ( .A1(n4821), .A2(n5974), .B1(n6512), .B2(n3200), .ZN(n4824)
         );
  NOR2_X1 U5940 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4822), .ZN(n4832)
         );
  INV_X1 U5941 ( .A(n5339), .ZN(n6507) );
  NAND2_X1 U5942 ( .A1(n5277), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5337) );
  AOI21_X1 U5943 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5337), .A(n5283), .ZN(
        n5347) );
  OAI211_X1 U5944 ( .C1(n4832), .C2(n6769), .A(n6507), .B(n5347), .ZN(n4823)
         );
  INV_X1 U5945 ( .A(n4852), .ZN(n4831) );
  INV_X1 U5946 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4830) );
  INV_X1 U5947 ( .A(n6613), .ZN(n6551) );
  AOI22_X1 U5948 ( .A1(n4856), .A2(n6551), .B1(n6547), .B2(n4832), .ZN(n4829)
         );
  AND2_X1 U5949 ( .A1(n3200), .A2(n6567), .ZN(n5145) );
  NOR2_X1 U5950 ( .A1(n6503), .A2(n5337), .ZN(n4825) );
  AOI21_X1 U5951 ( .B1(n5145), .B2(n6512), .A(n4825), .ZN(n4853) );
  INV_X1 U5952 ( .A(n4853), .ZN(n4826) );
  AOI22_X1 U5953 ( .A1(n6619), .A2(n4827), .B1(n6549), .B2(n4826), .ZN(n4828)
         );
  OAI211_X1 U5954 ( .C1(n4831), .C2(n4830), .A(n4829), .B(n4828), .ZN(U3139)
         );
  NAND2_X1 U5955 ( .A1(n4852), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4835)
         );
  INV_X1 U5956 ( .A(n4832), .ZN(n4854) );
  OAI22_X1 U5957 ( .A1(n6581), .A2(n4854), .B1(n4853), .B2(n6586), .ZN(n4833)
         );
  AOI21_X1 U5958 ( .B1(n6583), .B2(n4856), .A(n4833), .ZN(n4834) );
  OAI211_X1 U5959 ( .C1(n4859), .C2(n6580), .A(n4835), .B(n4834), .ZN(U3134)
         );
  NAND2_X1 U5960 ( .A1(n4852), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4838)
         );
  OAI22_X1 U5961 ( .A1(n6598), .A2(n4854), .B1(n4853), .B2(n6603), .ZN(n4836)
         );
  AOI21_X1 U5962 ( .B1(n6600), .B2(n4856), .A(n4836), .ZN(n4837) );
  OAI211_X1 U5963 ( .C1(n4859), .C2(n6597), .A(n4838), .B(n4837), .ZN(U3137)
         );
  NAND2_X1 U5964 ( .A1(n4852), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4841)
         );
  OAI22_X1 U5965 ( .A1(n6606), .A2(n4854), .B1(n4853), .B2(n6612), .ZN(n4839)
         );
  AOI21_X1 U5966 ( .B1(n6609), .B2(n4856), .A(n4839), .ZN(n4840) );
  OAI211_X1 U5967 ( .C1(n4859), .C2(n6604), .A(n4841), .B(n4840), .ZN(U3138)
         );
  INV_X1 U5968 ( .A(n6576), .ZN(n6525) );
  NAND2_X1 U5969 ( .A1(n4852), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4844)
         );
  INV_X1 U5970 ( .A(n6573), .ZN(n6522) );
  OAI22_X1 U5971 ( .A1(n6574), .A2(n4854), .B1(n4853), .B2(n6579), .ZN(n4842)
         );
  AOI21_X1 U5972 ( .B1(n6522), .B2(n4856), .A(n4842), .ZN(n4843) );
  OAI211_X1 U5973 ( .C1(n4859), .C2(n6525), .A(n4844), .B(n4843), .ZN(U3133)
         );
  NAND2_X1 U5974 ( .A1(n4852), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4848)
         );
  OAI22_X1 U5975 ( .A1(n4978), .A2(n6632), .B1(n6626), .B2(n4854), .ZN(n4846)
         );
  NOR2_X1 U5976 ( .A1(n4859), .A2(n6627), .ZN(n4845) );
  NOR2_X1 U5977 ( .A1(n4846), .A2(n4845), .ZN(n4847) );
  OAI211_X1 U5978 ( .C1(n4853), .C2(n6572), .A(n4848), .B(n4847), .ZN(U3132)
         );
  INV_X1 U5979 ( .A(n6588), .ZN(n6635) );
  NAND2_X1 U5980 ( .A1(n4852), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4851)
         );
  INV_X1 U5981 ( .A(n6643), .ZN(n6531) );
  OAI22_X1 U5982 ( .A1(n6634), .A2(n4854), .B1(n4853), .B2(n6591), .ZN(n4849)
         );
  AOI21_X1 U5983 ( .B1(n6531), .B2(n4856), .A(n4849), .ZN(n4850) );
  OAI211_X1 U5984 ( .C1(n4859), .C2(n6635), .A(n4851), .B(n4850), .ZN(U3135)
         );
  NAND2_X1 U5985 ( .A1(n4852), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4858)
         );
  OAI22_X1 U5986 ( .A1(n7203), .A2(n4854), .B1(n4853), .B2(n7200), .ZN(n4855)
         );
  AOI21_X1 U5987 ( .B1(n6594), .B2(n4856), .A(n4855), .ZN(n4857) );
  OAI211_X1 U5988 ( .C1(n4859), .C2(n6592), .A(n4858), .B(n4857), .ZN(U3136)
         );
  XNOR2_X1 U5989 ( .A(n4860), .B(n4861), .ZN(n6486) );
  INV_X1 U5990 ( .A(n6272), .ZN(n5263) );
  AOI22_X1 U5991 ( .A1(n6259), .A2(n6486), .B1(n5263), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4862) );
  OAI21_X1 U5992 ( .B1(n4863), .B2(n5626), .A(n4862), .ZN(U2858) );
  OR2_X1 U5993 ( .A1(n4865), .A2(n4864), .ZN(n4866) );
  AND2_X1 U5994 ( .A1(n4867), .A2(n4866), .ZN(n6383) );
  INV_X1 U5995 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6717) );
  OAI22_X1 U5996 ( .A1(n6463), .A2(n6225), .B1(n6717), .B2(n6461), .ZN(n4875)
         );
  NOR2_X1 U5997 ( .A1(n7097), .A2(n6494), .ZN(n4872) );
  NOR2_X1 U5998 ( .A1(n7057), .A2(n4868), .ZN(n5893) );
  AOI21_X1 U5999 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6475) );
  NOR2_X1 U6000 ( .A1(n6475), .A2(n5792), .ZN(n5384) );
  AOI21_X1 U6001 ( .B1(n4872), .B2(n6479), .A(n5384), .ZN(n6469) );
  NAND2_X1 U6002 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U6003 ( .A1(n5935), .A2(n5792), .ZN(n6493) );
  NAND3_X1 U6004 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6445) );
  INV_X1 U6005 ( .A(n4869), .ZN(n4871) );
  NOR2_X1 U6006 ( .A1(n4871), .A2(n4870), .ZN(n6484) );
  INV_X1 U6007 ( .A(n5792), .ZN(n6473) );
  OAI22_X1 U6008 ( .A1(n6484), .A2(n6473), .B1(n5935), .B2(n4872), .ZN(n6478)
         );
  AOI221_X1 U6009 ( .B1(n6475), .B2(n6493), .C1(n6445), .C2(n6493), .A(n6478), 
        .ZN(n6451) );
  AOI221_X1 U6010 ( .B1(n6469), .B2(n4873), .C1(n6456), .C2(n4873), .A(n6451), 
        .ZN(n4874) );
  AOI211_X1 U6011 ( .C1(n6477), .C2(n6383), .A(n4875), .B(n4874), .ZN(n4876)
         );
  INV_X1 U6012 ( .A(n4876), .ZN(U3013) );
  INV_X1 U6013 ( .A(n4877), .ZN(n4878) );
  AOI21_X1 U6014 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n6453) );
  AOI22_X1 U6015 ( .A1(n6453), .A2(n6259), .B1(n5263), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4881) );
  OAI21_X1 U6016 ( .B1(n4882), .B2(n5626), .A(n4881), .ZN(U2855) );
  AOI21_X1 U6017 ( .B1(n4884), .B2(n4883), .A(n6206), .ZN(n6443) );
  AOI22_X1 U6018 ( .A1(n6443), .A2(n6259), .B1(n5263), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4885) );
  OAI21_X1 U6019 ( .B1(n5254), .B2(n5626), .A(n4885), .ZN(U2853) );
  OAI21_X1 U6020 ( .B1(n4888), .B2(n4887), .A(n3197), .ZN(n6444) );
  INV_X1 U6021 ( .A(n5254), .ZN(n4891) );
  NAND2_X1 U6022 ( .A1(n6471), .A2(REIP_REG_6__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U6023 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4889)
         );
  OAI211_X1 U6024 ( .C1(n6406), .C2(n5255), .A(n6441), .B(n4889), .ZN(n4890)
         );
  AOI21_X1 U6025 ( .B1(n4891), .B2(n6400), .A(n4890), .ZN(n4892) );
  OAI21_X1 U6026 ( .B1(n6444), .B2(n6125), .A(n4892), .ZN(U2980) );
  INV_X1 U6027 ( .A(n5147), .ZN(n4893) );
  NAND3_X1 U6028 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6662), .A3(n6658), .ZN(n5141) );
  NOR2_X1 U6029 ( .A1(n6504), .A2(n5141), .ZN(n4900) );
  AOI21_X1 U6030 ( .B1(n4952), .B2(n4893), .A(n4900), .ZN(n4897) );
  OR3_X1 U6031 ( .A1(n5022), .A2(n4676), .A3(n6124), .ZN(n4894) );
  AOI22_X1 U6032 ( .A1(n4897), .A2(n4896), .B1(n6559), .B2(n5141), .ZN(n4895)
         );
  NAND2_X1 U6033 ( .A1(n6565), .A2(n4895), .ZN(n4997) );
  INV_X1 U6034 ( .A(n4896), .ZN(n4898) );
  OAI22_X1 U6035 ( .A1(n4898), .A2(n4897), .B1(n6680), .B2(n5141), .ZN(n4996)
         );
  AOI22_X1 U6036 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4997), .B1(n6538), 
        .B2(n4996), .ZN(n4903) );
  INV_X1 U6037 ( .A(n4900), .ZN(n4998) );
  OAI22_X1 U6038 ( .A1(n5340), .A2(n6597), .B1(n4998), .B2(n6598), .ZN(n4901)
         );
  AOI21_X1 U6039 ( .B1(n5139), .B2(n6600), .A(n4901), .ZN(n4902) );
  NAND2_X1 U6040 ( .A1(n4903), .A2(n4902), .ZN(U3097) );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4997), .B1(n6526), 
        .B2(n4996), .ZN(n4906) );
  OAI22_X1 U6042 ( .A1(n5340), .A2(n6580), .B1(n4998), .B2(n6581), .ZN(n4904)
         );
  AOI21_X1 U6043 ( .B1(n5139), .B2(n6583), .A(n4904), .ZN(n4905) );
  NAND2_X1 U6044 ( .A1(n4906), .A2(n4905), .ZN(U3094) );
  AOI22_X1 U6045 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4997), .B1(n6534), 
        .B2(n4996), .ZN(n4909) );
  OAI22_X1 U6046 ( .A1(n5340), .A2(n6592), .B1(n4998), .B2(n7203), .ZN(n4907)
         );
  AOI21_X1 U6047 ( .B1(n5139), .B2(n6594), .A(n4907), .ZN(n4908) );
  NAND2_X1 U6048 ( .A1(n4909), .A2(n4908), .ZN(U3096) );
  AOI22_X1 U6049 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4997), .B1(n6542), 
        .B2(n4996), .ZN(n4912) );
  OAI22_X1 U6050 ( .A1(n5340), .A2(n6604), .B1(n4998), .B2(n6606), .ZN(n4910)
         );
  AOI21_X1 U6051 ( .B1(n5139), .B2(n6609), .A(n4910), .ZN(n4911) );
  NAND2_X1 U6052 ( .A1(n4912), .A2(n4911), .ZN(U3098) );
  INV_X1 U6053 ( .A(n5030), .ZN(n4914) );
  OR2_X1 U6054 ( .A1(n4605), .A2(n6241), .ZN(n5008) );
  OR2_X1 U6055 ( .A1(n4673), .A2(n3641), .ZN(n6500) );
  AOI21_X1 U6056 ( .B1(n4922), .B2(STATEBS16_REG_SCAN_IN), .A(n6559), .ZN(
        n5104) );
  OAI21_X1 U6057 ( .B1(n5099), .B2(n5008), .A(n5104), .ZN(n4918) );
  NOR2_X1 U6058 ( .A1(n5057), .A2(n6509), .ZN(n4917) );
  NAND3_X1 U6059 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6669), .A3(n6658), .ZN(n5105) );
  OR2_X1 U6060 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5105), .ZN(n4947)
         );
  AOI21_X1 U6061 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4947), .A(n4915), .ZN(
        n4916) );
  NAND2_X1 U6062 ( .A1(n4945), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4925) );
  INV_X1 U6063 ( .A(n3200), .ZN(n5970) );
  NAND3_X1 U6064 ( .A1(n5970), .A2(n6567), .A3(n5101), .ZN(n4921) );
  INV_X1 U6065 ( .A(n6503), .ZN(n4919) );
  NAND2_X1 U6066 ( .A1(n4919), .A2(n3304), .ZN(n4920) );
  AND2_X1 U6067 ( .A1(n4921), .A2(n4920), .ZN(n4946) );
  INV_X1 U6068 ( .A(n4946), .ZN(n4936) );
  OAI22_X1 U6069 ( .A1(n5180), .A2(n6555), .B1(n6616), .B2(n4947), .ZN(n4923)
         );
  AOI21_X1 U6070 ( .B1(n6549), .B2(n4936), .A(n4923), .ZN(n4924) );
  OAI211_X1 U6071 ( .C1(n5057), .C2(n6613), .A(n4925), .B(n4924), .ZN(U3059)
         );
  NAND2_X1 U6072 ( .A1(n4945), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4928) );
  OAI22_X1 U6073 ( .A1(n6598), .A2(n4947), .B1(n4946), .B2(n6603), .ZN(n4926)
         );
  AOI21_X1 U6074 ( .B1(n5288), .B2(n4949), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6075 ( .C1(n5057), .C2(n5290), .A(n4928), .B(n4927), .ZN(U3057)
         );
  NAND2_X1 U6076 ( .A1(n4945), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6077 ( .A1(n6606), .A2(n4947), .B1(n4946), .B2(n6612), .ZN(n4929)
         );
  AOI21_X1 U6078 ( .B1(n5293), .B2(n4949), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6079 ( .C1(n5057), .C2(n5295), .A(n4931), .B(n4930), .ZN(U3058)
         );
  NAND2_X1 U6080 ( .A1(n4945), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6081 ( .A1(n6634), .A2(n4947), .B1(n4946), .B2(n6591), .ZN(n4932)
         );
  AOI21_X1 U6082 ( .B1(n6588), .B2(n4949), .A(n4932), .ZN(n4933) );
  OAI211_X1 U6083 ( .C1(n5057), .C2(n6643), .A(n4934), .B(n4933), .ZN(U3055)
         );
  NAND2_X1 U6084 ( .A1(n4945), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4938) );
  OAI22_X1 U6085 ( .A1(n5180), .A2(n6627), .B1(n6626), .B2(n4947), .ZN(n4935)
         );
  AOI21_X1 U6086 ( .B1(n6629), .B2(n4936), .A(n4935), .ZN(n4937) );
  OAI211_X1 U6087 ( .C1(n5057), .C2(n6632), .A(n4938), .B(n4937), .ZN(U3052)
         );
  NAND2_X1 U6088 ( .A1(n4945), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4941) );
  OAI22_X1 U6089 ( .A1(n6574), .A2(n4947), .B1(n4946), .B2(n6579), .ZN(n4939)
         );
  AOI21_X1 U6090 ( .B1(n6576), .B2(n4949), .A(n4939), .ZN(n4940) );
  OAI211_X1 U6091 ( .C1(n5057), .C2(n6573), .A(n4941), .B(n4940), .ZN(U3053)
         );
  NAND2_X1 U6092 ( .A1(n4945), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4944) );
  OAI22_X1 U6093 ( .A1(n7203), .A2(n4947), .B1(n4946), .B2(n7200), .ZN(n4942)
         );
  AOI21_X1 U6094 ( .B1(n7206), .B2(n4949), .A(n4942), .ZN(n4943) );
  OAI211_X1 U6095 ( .C1(n5057), .C2(n7209), .A(n4944), .B(n4943), .ZN(U3056)
         );
  NAND2_X1 U6096 ( .A1(n4945), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4951) );
  OAI22_X1 U6097 ( .A1(n6581), .A2(n4947), .B1(n4946), .B2(n6586), .ZN(n4948)
         );
  AOI21_X1 U6098 ( .B1(n5301), .B2(n4949), .A(n4948), .ZN(n4950) );
  OAI211_X1 U6099 ( .C1(n5057), .C2(n5303), .A(n4951), .B(n4950), .ZN(U3054)
         );
  NAND3_X1 U6100 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6658), .ZN(n5012) );
  INV_X1 U6101 ( .A(n5012), .ZN(n4955) );
  NOR2_X1 U6102 ( .A1(n6504), .A2(n5012), .ZN(n4975) );
  AOI21_X1 U6103 ( .B1(n4952), .B2(n5101), .A(n4975), .ZN(n4957) );
  NAND2_X1 U6104 ( .A1(n4953), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5023) );
  NAND3_X1 U6105 ( .A1(n6567), .A2(n4957), .A3(n5023), .ZN(n4954) );
  OAI211_X1 U6106 ( .C1(n6567), .C2(n4955), .A(n6565), .B(n4954), .ZN(n4974)
         );
  NAND2_X1 U6107 ( .A1(n6567), .A2(n5023), .ZN(n4956) );
  OAI22_X1 U6108 ( .A1(n4957), .A2(n4956), .B1(n6680), .B2(n5012), .ZN(n4973)
         );
  AOI22_X1 U6109 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4974), .B1(n6534), 
        .B2(n4973), .ZN(n4960) );
  AOI22_X1 U6110 ( .A1(n6594), .A2(n7205), .B1(n6535), .B2(n4975), .ZN(n4959)
         );
  OAI211_X1 U6111 ( .C1(n6592), .C2(n4978), .A(n4960), .B(n4959), .ZN(U3128)
         );
  AOI22_X1 U6112 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4974), .B1(n6538), 
        .B2(n4973), .ZN(n4962) );
  AOI22_X1 U6113 ( .A1(n6600), .A2(n7205), .B1(n6539), .B2(n4975), .ZN(n4961)
         );
  OAI211_X1 U6114 ( .C1(n6597), .C2(n4978), .A(n4962), .B(n4961), .ZN(U3129)
         );
  AOI22_X1 U6115 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4974), .B1(n6542), 
        .B2(n4973), .ZN(n4964) );
  AOI22_X1 U6116 ( .A1(n6609), .A2(n7205), .B1(n6543), .B2(n4975), .ZN(n4963)
         );
  OAI211_X1 U6117 ( .C1(n6604), .C2(n4978), .A(n4964), .B(n4963), .ZN(U3130)
         );
  AOI22_X1 U6118 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4974), .B1(n6549), 
        .B2(n4973), .ZN(n4966) );
  AOI22_X1 U6119 ( .A1(n6551), .A2(n7205), .B1(n6547), .B2(n4975), .ZN(n4965)
         );
  OAI211_X1 U6120 ( .C1(n6555), .C2(n4978), .A(n4966), .B(n4965), .ZN(U3131)
         );
  AOI22_X1 U6121 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4974), .B1(n6629), 
        .B2(n4973), .ZN(n4968) );
  INV_X1 U6122 ( .A(n6626), .ZN(n6505) );
  AOI22_X1 U6123 ( .A1(n6517), .A2(n7205), .B1(n6505), .B2(n4975), .ZN(n4967)
         );
  OAI211_X1 U6124 ( .C1(n6627), .C2(n4978), .A(n4968), .B(n4967), .ZN(U3124)
         );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4974), .B1(n6526), 
        .B2(n4973), .ZN(n4970) );
  AOI22_X1 U6126 ( .A1(n6583), .A2(n7205), .B1(n6527), .B2(n4975), .ZN(n4969)
         );
  OAI211_X1 U6127 ( .C1(n6580), .C2(n4978), .A(n4970), .B(n4969), .ZN(U3126)
         );
  AOI22_X1 U6128 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4974), .B1(n6638), 
        .B2(n4973), .ZN(n4972) );
  AOI22_X1 U6129 ( .A1(n6531), .A2(n7205), .B1(n6530), .B2(n4975), .ZN(n4971)
         );
  OAI211_X1 U6130 ( .C1(n6635), .C2(n4978), .A(n4972), .B(n4971), .ZN(U3127)
         );
  AOI22_X1 U6131 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4974), .B1(n6520), 
        .B2(n4973), .ZN(n4977) );
  AOI22_X1 U6132 ( .A1(n6522), .A2(n7205), .B1(n6521), .B2(n4975), .ZN(n4976)
         );
  OAI211_X1 U6133 ( .C1(n6525), .C2(n4978), .A(n4977), .B(n4976), .ZN(U3125)
         );
  NAND2_X1 U6134 ( .A1(n4980), .A2(n4981), .ZN(n4982) );
  NAND2_X1 U6135 ( .A1(n4979), .A2(n4982), .ZN(n5244) );
  INV_X1 U6136 ( .A(n4983), .ZN(n6205) );
  NAND2_X1 U6137 ( .A1(n6206), .A2(n6205), .ZN(n4984) );
  AOI21_X1 U6138 ( .B1(n4985), .B2(n4984), .A(n5391), .ZN(n6425) );
  AOI22_X1 U6139 ( .A1(n6425), .A2(n6259), .B1(n5263), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4986) );
  OAI21_X1 U6140 ( .B1(n5244), .B2(n5626), .A(n4986), .ZN(U2851) );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4997), .B1(n6520), 
        .B2(n4996), .ZN(n4989) );
  OAI22_X1 U6142 ( .A1(n5340), .A2(n6525), .B1(n4998), .B2(n6574), .ZN(n4987)
         );
  INV_X1 U6143 ( .A(n4987), .ZN(n4988) );
  OAI211_X1 U6144 ( .C1(n5177), .C2(n6573), .A(n4989), .B(n4988), .ZN(U3093)
         );
  AOI22_X1 U6145 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4997), .B1(n6638), 
        .B2(n4996), .ZN(n4992) );
  OAI22_X1 U6146 ( .A1(n5340), .A2(n6635), .B1(n4998), .B2(n6634), .ZN(n4990)
         );
  INV_X1 U6147 ( .A(n4990), .ZN(n4991) );
  OAI211_X1 U6148 ( .C1(n5177), .C2(n6643), .A(n4992), .B(n4991), .ZN(U3095)
         );
  AOI22_X1 U6149 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4997), .B1(n6629), 
        .B2(n4996), .ZN(n4995) );
  OAI22_X1 U6150 ( .A1(n5340), .A2(n6627), .B1(n6626), .B2(n4998), .ZN(n4993)
         );
  INV_X1 U6151 ( .A(n4993), .ZN(n4994) );
  OAI211_X1 U6152 ( .C1(n5177), .C2(n6632), .A(n4995), .B(n4994), .ZN(U3092)
         );
  AOI22_X1 U6153 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4997), .B1(n6549), 
        .B2(n4996), .ZN(n5001) );
  OAI22_X1 U6154 ( .A1(n5340), .A2(n6555), .B1(n4998), .B2(n6616), .ZN(n4999)
         );
  INV_X1 U6155 ( .A(n4999), .ZN(n5000) );
  OAI211_X1 U6156 ( .C1(n5177), .C2(n6613), .A(n5001), .B(n5000), .ZN(U3099)
         );
  INV_X1 U6157 ( .A(DATAI_8_), .ZN(n5002) );
  INV_X1 U6158 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7116) );
  OAI222_X1 U6159 ( .A1(n5244), .A2(n6054), .B1(n6284), .B2(n5002), .C1(n6285), 
        .C2(n7116), .ZN(U2883) );
  INV_X1 U6160 ( .A(n5003), .ZN(n5004) );
  XNOR2_X1 U6161 ( .A(n4787), .B(n5004), .ZN(n6378) );
  INV_X1 U6162 ( .A(n6378), .ZN(n5006) );
  OAI222_X1 U6163 ( .A1(n5007), .A2(n6284), .B1(n6054), .B2(n5006), .C1(n5005), 
        .C2(n6285), .ZN(U2884) );
  NOR3_X1 U6164 ( .A1(n5019), .A2(n7205), .A3(n6559), .ZN(n5009) );
  OAI22_X1 U6165 ( .A1(n5009), .A2(n6509), .B1(n5970), .B2(n5008), .ZN(n5014)
         );
  INV_X1 U6166 ( .A(n5277), .ZN(n5011) );
  NAND2_X1 U6167 ( .A1(n5011), .A2(n5010), .ZN(n5146) );
  AOI21_X1 U6168 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5146), .A(n5283), .ZN(
        n5143) );
  NOR2_X1 U6169 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5012), .ZN(n5093)
         );
  INV_X1 U6170 ( .A(n5093), .ZN(n7202) );
  NAND2_X1 U6171 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7202), .ZN(n5013) );
  NAND4_X1 U6172 ( .A1(n5014), .A2(n5143), .A3(n6507), .A4(n5013), .ZN(n7199)
         );
  INV_X1 U6173 ( .A(n7199), .ZN(n5021) );
  INV_X1 U6174 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U6175 ( .A1(n5145), .A2(n5101), .ZN(n5016) );
  OR2_X1 U6176 ( .A1(n6503), .A2(n5146), .ZN(n5015) );
  AOI22_X1 U6177 ( .A1(n6619), .A2(n7205), .B1(n6547), .B2(n5093), .ZN(n5017)
         );
  OAI21_X1 U6178 ( .B1(n6623), .B2(n7201), .A(n5017), .ZN(n5018) );
  AOI21_X1 U6179 ( .B1(n6551), .B2(n5019), .A(n5018), .ZN(n5020) );
  OAI21_X1 U6180 ( .B1(n5021), .B2(n6949), .A(n5020), .ZN(U3123) );
  NAND2_X1 U6181 ( .A1(n5023), .A2(n5022), .ZN(n5969) );
  NOR3_X1 U6182 ( .A1(n5969), .A2(n5024), .A3(n5968), .ZN(n5025) );
  NOR2_X1 U6183 ( .A1(n5025), .A2(n6559), .ZN(n5032) );
  OR2_X1 U6184 ( .A1(n3200), .A2(n5026), .ZN(n5282) );
  INV_X1 U6185 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6186 ( .A1(n5028), .A2(n6669), .ZN(n5056) );
  OAI21_X1 U6187 ( .B1(n5282), .B2(n3595), .A(n5056), .ZN(n5034) );
  NAND3_X1 U6188 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6669), .A3(n6662), .ZN(n5276) );
  INV_X1 U6189 ( .A(n5276), .ZN(n5029) );
  AOI22_X1 U6190 ( .A1(n5032), .A2(n5034), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5029), .ZN(n5062) );
  OAI22_X1 U6191 ( .A1(n5057), .A2(n6627), .B1(n6626), .B2(n5056), .ZN(n5031)
         );
  AOI21_X1 U6192 ( .B1(n6517), .B2(n5986), .A(n5031), .ZN(n5037) );
  INV_X1 U6193 ( .A(n5032), .ZN(n5035) );
  NAND2_X1 U6194 ( .A1(n6559), .A2(n5276), .ZN(n5033) );
  NAND2_X1 U6195 ( .A1(n5059), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5036) );
  OAI211_X1 U6196 ( .C1(n5062), .C2(n6572), .A(n5037), .B(n5036), .ZN(U3044)
         );
  OAI22_X1 U6197 ( .A1(n5057), .A2(n6604), .B1(n6606), .B2(n5056), .ZN(n5038)
         );
  AOI21_X1 U6198 ( .B1(n6609), .B2(n5986), .A(n5038), .ZN(n5040) );
  NAND2_X1 U6199 ( .A1(n5059), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5039) );
  OAI211_X1 U6200 ( .C1(n5062), .C2(n6612), .A(n5040), .B(n5039), .ZN(U3050)
         );
  OAI22_X1 U6201 ( .A1(n5057), .A2(n6555), .B1(n6616), .B2(n5056), .ZN(n5041)
         );
  AOI21_X1 U6202 ( .B1(n6551), .B2(n5986), .A(n5041), .ZN(n5043) );
  NAND2_X1 U6203 ( .A1(n5059), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5042) );
  OAI211_X1 U6204 ( .C1(n5062), .C2(n6623), .A(n5043), .B(n5042), .ZN(U3051)
         );
  OAI22_X1 U6205 ( .A1(n5057), .A2(n6592), .B1(n7203), .B2(n5056), .ZN(n5044)
         );
  AOI21_X1 U6206 ( .B1(n6594), .B2(n5986), .A(n5044), .ZN(n5046) );
  NAND2_X1 U6207 ( .A1(n5059), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5045) );
  OAI211_X1 U6208 ( .C1(n5062), .C2(n7200), .A(n5046), .B(n5045), .ZN(U3048)
         );
  OAI22_X1 U6209 ( .A1(n5057), .A2(n6597), .B1(n6598), .B2(n5056), .ZN(n5047)
         );
  AOI21_X1 U6210 ( .B1(n6600), .B2(n5986), .A(n5047), .ZN(n5049) );
  NAND2_X1 U6211 ( .A1(n5059), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5048) );
  OAI211_X1 U6212 ( .C1(n5062), .C2(n6603), .A(n5049), .B(n5048), .ZN(U3049)
         );
  OAI22_X1 U6213 ( .A1(n5057), .A2(n6580), .B1(n6581), .B2(n5056), .ZN(n5050)
         );
  AOI21_X1 U6214 ( .B1(n6583), .B2(n5986), .A(n5050), .ZN(n5052) );
  NAND2_X1 U6215 ( .A1(n5059), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5051) );
  OAI211_X1 U6216 ( .C1(n5062), .C2(n6586), .A(n5052), .B(n5051), .ZN(U3046)
         );
  OAI22_X1 U6217 ( .A1(n5057), .A2(n6525), .B1(n6574), .B2(n5056), .ZN(n5053)
         );
  AOI21_X1 U6218 ( .B1(n6522), .B2(n5986), .A(n5053), .ZN(n5055) );
  NAND2_X1 U6219 ( .A1(n5059), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5054) );
  OAI211_X1 U6220 ( .C1(n5062), .C2(n6579), .A(n5055), .B(n5054), .ZN(U3045)
         );
  OAI22_X1 U6221 ( .A1(n5057), .A2(n6635), .B1(n6634), .B2(n5056), .ZN(n5058)
         );
  AOI21_X1 U6222 ( .B1(n6531), .B2(n5986), .A(n5058), .ZN(n5061) );
  NAND2_X1 U6223 ( .A1(n5059), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5060) );
  OAI211_X1 U6224 ( .C1(n5062), .C2(n6591), .A(n5061), .B(n5060), .ZN(U3047)
         );
  AOI22_X1 U6225 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6244), .B1(n6249), 
        .B2(n6425), .ZN(n5064) );
  NAND2_X1 U6226 ( .A1(n5548), .A2(n5063), .ZN(n6226) );
  OAI211_X1 U6227 ( .C1(n6251), .C2(n5065), .A(n5064), .B(n6226), .ZN(n5066)
         );
  AOI21_X1 U6228 ( .B1(n6212), .B2(n5247), .A(n5066), .ZN(n5072) );
  INV_X1 U6229 ( .A(n5067), .ZN(n5226) );
  OAI21_X1 U6230 ( .B1(n5226), .B2(n6247), .A(n5548), .ZN(n5070) );
  NOR2_X1 U6231 ( .A1(n5226), .A2(n6247), .ZN(n5068) );
  AOI22_X1 U6232 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5070), .B1(n5069), .B2(n5068), .ZN(n5071) );
  OAI211_X1 U6233 ( .C1(n6198), .C2(n5244), .A(n5072), .B(n5071), .ZN(U2819)
         );
  AOI21_X1 U6234 ( .B1(n5074), .B2(n4979), .A(n5073), .ZN(n5326) );
  INV_X1 U6235 ( .A(n5326), .ZN(n5077) );
  XNOR2_X1 U6236 ( .A(n5391), .B(n5389), .ZN(n6417) );
  AOI22_X1 U6237 ( .A1(n6417), .A2(n6259), .B1(n5263), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5075) );
  OAI21_X1 U6238 ( .B1(n5077), .B2(n5626), .A(n5075), .ZN(U2850) );
  INV_X1 U6239 ( .A(n6284), .ZN(n5645) );
  AOI22_X1 U6240 ( .A1(n5645), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6279), .ZN(n5076) );
  OAI21_X1 U6241 ( .B1(n5077), .B2(n6054), .A(n5076), .ZN(U2882) );
  NAND2_X1 U6242 ( .A1(n7199), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5080)
         );
  OAI22_X1 U6243 ( .A1(n6606), .A2(n7202), .B1(n7201), .B2(n6612), .ZN(n5078)
         );
  AOI21_X1 U6244 ( .B1(n5293), .B2(n7205), .A(n5078), .ZN(n5079) );
  OAI211_X1 U6245 ( .C1(n7210), .C2(n5295), .A(n5080), .B(n5079), .ZN(U3122)
         );
  NAND2_X1 U6246 ( .A1(n7199), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5083)
         );
  OAI22_X1 U6247 ( .A1(n6634), .A2(n7202), .B1(n7201), .B2(n6591), .ZN(n5081)
         );
  AOI21_X1 U6248 ( .B1(n6588), .B2(n7205), .A(n5081), .ZN(n5082) );
  OAI211_X1 U6249 ( .C1(n7210), .C2(n6643), .A(n5083), .B(n5082), .ZN(U3119)
         );
  NAND2_X1 U6250 ( .A1(n7199), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5086)
         );
  OAI22_X1 U6251 ( .A1(n6581), .A2(n7202), .B1(n7201), .B2(n6586), .ZN(n5084)
         );
  AOI21_X1 U6252 ( .B1(n5301), .B2(n7205), .A(n5084), .ZN(n5085) );
  OAI211_X1 U6253 ( .C1(n7210), .C2(n5303), .A(n5086), .B(n5085), .ZN(U3118)
         );
  NAND2_X1 U6254 ( .A1(n7199), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5089)
         );
  OAI22_X1 U6255 ( .A1(n6574), .A2(n7202), .B1(n7201), .B2(n6579), .ZN(n5087)
         );
  AOI21_X1 U6256 ( .B1(n6576), .B2(n7205), .A(n5087), .ZN(n5088) );
  OAI211_X1 U6257 ( .C1(n7210), .C2(n6573), .A(n5089), .B(n5088), .ZN(U3117)
         );
  NAND2_X1 U6258 ( .A1(n7199), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5092)
         );
  OAI22_X1 U6259 ( .A1(n6598), .A2(n7202), .B1(n7201), .B2(n6603), .ZN(n5090)
         );
  AOI21_X1 U6260 ( .B1(n5288), .B2(n7205), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6261 ( .C1(n7210), .C2(n5290), .A(n5092), .B(n5091), .ZN(U3121)
         );
  AOI22_X1 U6262 ( .A1(n6569), .A2(n7205), .B1(n6505), .B2(n5093), .ZN(n5096)
         );
  INV_X1 U6263 ( .A(n7201), .ZN(n5094) );
  NAND2_X1 U6264 ( .A1(n6629), .A2(n5094), .ZN(n5095) );
  OAI211_X1 U6265 ( .C1(n7210), .C2(n6632), .A(n5096), .B(n5095), .ZN(n5097)
         );
  AOI21_X1 U6266 ( .B1(n7199), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n5097), 
        .ZN(n5098) );
  INV_X1 U6267 ( .A(n5098), .ZN(U3116) );
  NOR2_X1 U6268 ( .A1(n3595), .A2(n5099), .ZN(n5100) );
  NOR2_X1 U6269 ( .A1(n6504), .A2(n5105), .ZN(n5178) );
  AOI21_X1 U6270 ( .B1(n5101), .B2(n5100), .A(n5178), .ZN(n5106) );
  INV_X1 U6271 ( .A(n5105), .ZN(n5102) );
  OAI21_X1 U6272 ( .B1(n6567), .B2(n5102), .A(n6565), .ZN(n5103) );
  INV_X1 U6273 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5113) );
  INV_X1 U6274 ( .A(n5104), .ZN(n5107) );
  OAI22_X1 U6275 ( .A1(n5107), .A2(n5106), .B1(n5105), .B2(n6680), .ZN(n5182)
         );
  NOR2_X2 U6276 ( .A1(n5109), .A2(n5108), .ZN(n6550) );
  AOI22_X1 U6277 ( .A1(n6550), .A2(n6619), .B1(n6547), .B2(n5178), .ZN(n5110)
         );
  OAI21_X1 U6278 ( .B1(n6613), .B2(n5180), .A(n5110), .ZN(n5111) );
  AOI21_X1 U6279 ( .B1(n6549), .B2(n5182), .A(n5111), .ZN(n5112) );
  OAI21_X1 U6280 ( .B1(n5185), .B2(n5113), .A(n5112), .ZN(U3067) );
  INV_X1 U6281 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U6282 ( .A1(n6550), .A2(n5288), .B1(n6539), .B2(n5178), .ZN(n5114)
         );
  OAI21_X1 U6283 ( .B1(n5290), .B2(n5180), .A(n5114), .ZN(n5115) );
  AOI21_X1 U6284 ( .B1(n6538), .B2(n5182), .A(n5115), .ZN(n5116) );
  OAI21_X1 U6285 ( .B1(n5185), .B2(n5117), .A(n5116), .ZN(U3065) );
  INV_X1 U6286 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5121) );
  AOI22_X1 U6287 ( .A1(n6550), .A2(n5301), .B1(n6527), .B2(n5178), .ZN(n5118)
         );
  OAI21_X1 U6288 ( .B1(n5303), .B2(n5180), .A(n5118), .ZN(n5119) );
  AOI21_X1 U6289 ( .B1(n6526), .B2(n5182), .A(n5119), .ZN(n5120) );
  OAI21_X1 U6290 ( .B1(n5185), .B2(n5121), .A(n5120), .ZN(U3062) );
  INV_X1 U6291 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5125) );
  AOI22_X1 U6292 ( .A1(n6550), .A2(n5293), .B1(n6543), .B2(n5178), .ZN(n5122)
         );
  OAI21_X1 U6293 ( .B1(n5295), .B2(n5180), .A(n5122), .ZN(n5123) );
  AOI21_X1 U6294 ( .B1(n6542), .B2(n5182), .A(n5123), .ZN(n5124) );
  OAI21_X1 U6295 ( .B1(n5185), .B2(n5125), .A(n5124), .ZN(U3066) );
  INV_X1 U6296 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5129) );
  AOI22_X1 U6297 ( .A1(n6550), .A2(n7206), .B1(n6535), .B2(n5178), .ZN(n5126)
         );
  OAI21_X1 U6298 ( .B1(n7209), .B2(n5180), .A(n5126), .ZN(n5127) );
  AOI21_X1 U6299 ( .B1(n6534), .B2(n5182), .A(n5127), .ZN(n5128) );
  OAI21_X1 U6300 ( .B1(n5185), .B2(n5129), .A(n5128), .ZN(U3064) );
  INV_X1 U6301 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U6302 ( .A1(n6550), .A2(n6576), .B1(n6521), .B2(n5178), .ZN(n5130)
         );
  OAI21_X1 U6303 ( .B1(n6573), .B2(n5180), .A(n5130), .ZN(n5131) );
  AOI21_X1 U6304 ( .B1(n6520), .B2(n5182), .A(n5131), .ZN(n5132) );
  OAI21_X1 U6305 ( .B1(n5185), .B2(n5133), .A(n5132), .ZN(U3061) );
  INV_X1 U6306 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5137) );
  AOI22_X1 U6307 ( .A1(n6550), .A2(n6588), .B1(n6530), .B2(n5178), .ZN(n5134)
         );
  OAI21_X1 U6308 ( .B1(n6643), .B2(n5180), .A(n5134), .ZN(n5135) );
  AOI21_X1 U6309 ( .B1(n6638), .B2(n5182), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6310 ( .B1(n5185), .B2(n5137), .A(n5136), .ZN(U3063) );
  OAI21_X1 U6311 ( .B1(n5139), .B2(n6618), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5140) );
  OAI211_X1 U6312 ( .C1(n5970), .C2(n5147), .A(n5140), .B(n6567), .ZN(n5144)
         );
  NOR2_X1 U6313 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5141), .ZN(n5148)
         );
  OR2_X1 U6314 ( .A1(n6769), .A2(n5148), .ZN(n5142) );
  NAND4_X1 U6315 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n6503), .ZN(n5171)
         );
  NAND2_X1 U6316 ( .A1(n5171), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5151) );
  INV_X1 U6317 ( .A(n5145), .ZN(n6511) );
  OAI22_X1 U6318 ( .A1(n6511), .A2(n5147), .B1(n6507), .B2(n5146), .ZN(n5165)
         );
  INV_X1 U6319 ( .A(n5148), .ZN(n5173) );
  OAI22_X1 U6320 ( .A1(n6616), .A2(n5173), .B1(n6605), .B2(n6613), .ZN(n5149)
         );
  AOI21_X1 U6321 ( .B1(n6549), .B2(n5165), .A(n5149), .ZN(n5150) );
  OAI211_X1 U6322 ( .C1(n6555), .C2(n5177), .A(n5151), .B(n5150), .ZN(U3091)
         );
  NAND2_X1 U6323 ( .A1(n5171), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5154) );
  INV_X1 U6324 ( .A(n5165), .ZN(n5172) );
  OAI22_X1 U6325 ( .A1(n6574), .A2(n5173), .B1(n5172), .B2(n6579), .ZN(n5152)
         );
  AOI21_X1 U6326 ( .B1(n6522), .B2(n6618), .A(n5152), .ZN(n5153) );
  OAI211_X1 U6327 ( .C1(n6525), .C2(n5177), .A(n5154), .B(n5153), .ZN(U3085)
         );
  NAND2_X1 U6328 ( .A1(n5171), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6329 ( .A1(n6606), .A2(n5173), .B1(n5172), .B2(n6612), .ZN(n5155)
         );
  AOI21_X1 U6330 ( .B1(n6609), .B2(n6618), .A(n5155), .ZN(n5156) );
  OAI211_X1 U6331 ( .C1(n6604), .C2(n5177), .A(n5157), .B(n5156), .ZN(U3090)
         );
  NAND2_X1 U6332 ( .A1(n5171), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5160) );
  OAI22_X1 U6333 ( .A1(n6598), .A2(n5173), .B1(n5172), .B2(n6603), .ZN(n5158)
         );
  AOI21_X1 U6334 ( .B1(n6600), .B2(n6618), .A(n5158), .ZN(n5159) );
  OAI211_X1 U6335 ( .C1(n6597), .C2(n5177), .A(n5160), .B(n5159), .ZN(U3089)
         );
  NAND2_X1 U6336 ( .A1(n5171), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5163) );
  OAI22_X1 U6337 ( .A1(n6634), .A2(n5173), .B1(n5172), .B2(n6591), .ZN(n5161)
         );
  AOI21_X1 U6338 ( .B1(n6531), .B2(n6618), .A(n5161), .ZN(n5162) );
  OAI211_X1 U6339 ( .C1(n6635), .C2(n5177), .A(n5163), .B(n5162), .ZN(U3087)
         );
  NAND2_X1 U6340 ( .A1(n5171), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5167) );
  OAI22_X1 U6341 ( .A1(n6626), .A2(n5173), .B1(n6605), .B2(n6632), .ZN(n5164)
         );
  AOI21_X1 U6342 ( .B1(n6629), .B2(n5165), .A(n5164), .ZN(n5166) );
  OAI211_X1 U6343 ( .C1(n6627), .C2(n5177), .A(n5167), .B(n5166), .ZN(U3084)
         );
  NAND2_X1 U6344 ( .A1(n5171), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5170) );
  OAI22_X1 U6345 ( .A1(n6581), .A2(n5173), .B1(n5172), .B2(n6586), .ZN(n5168)
         );
  AOI21_X1 U6346 ( .B1(n6583), .B2(n6618), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6347 ( .C1(n6580), .C2(n5177), .A(n5170), .B(n5169), .ZN(U3086)
         );
  NAND2_X1 U6348 ( .A1(n5171), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5176) );
  OAI22_X1 U6349 ( .A1(n7203), .A2(n5173), .B1(n5172), .B2(n7200), .ZN(n5174)
         );
  AOI21_X1 U6350 ( .B1(n6594), .B2(n6618), .A(n5174), .ZN(n5175) );
  OAI211_X1 U6351 ( .C1(n6592), .C2(n5177), .A(n5176), .B(n5175), .ZN(U3088)
         );
  INV_X1 U6352 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5184) );
  AOI22_X1 U6353 ( .A1(n6550), .A2(n6569), .B1(n6505), .B2(n5178), .ZN(n5179)
         );
  OAI21_X1 U6354 ( .B1(n6632), .B2(n5180), .A(n5179), .ZN(n5181) );
  AOI21_X1 U6355 ( .B1(n6629), .B2(n5182), .A(n5181), .ZN(n5183) );
  OAI21_X1 U6356 ( .B1(n5185), .B2(n5184), .A(n5183), .ZN(U3060) );
  NOR2_X1 U6357 ( .A1(n6504), .A2(n5189), .ZN(n5220) );
  INV_X1 U6358 ( .A(n5220), .ZN(n5195) );
  OAI21_X1 U6359 ( .B1(n5186), .B2(n3595), .A(n5195), .ZN(n5188) );
  INV_X1 U6360 ( .A(n5189), .ZN(n5187) );
  AOI22_X1 U6361 ( .A1(n5190), .A2(n5188), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5187), .ZN(n5225) );
  INV_X1 U6362 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5194) );
  INV_X1 U6363 ( .A(n5188), .ZN(n5191) );
  AOI22_X1 U6364 ( .A1(n5191), .A2(n5190), .B1(n5189), .B2(n6559), .ZN(n5192)
         );
  NAND2_X1 U6365 ( .A1(n6565), .A2(n5192), .ZN(n5219) );
  INV_X1 U6366 ( .A(n5219), .ZN(n5193) );
  OAI22_X1 U6367 ( .A1(n6626), .A2(n5195), .B1(n5194), .B2(n5193), .ZN(n5199)
         );
  NOR2_X1 U6368 ( .A1(n5989), .A2(n6627), .ZN(n5198) );
  AOI211_X1 U6369 ( .C1(n5223), .C2(n6517), .A(n5199), .B(n5198), .ZN(n5200)
         );
  OAI21_X1 U6370 ( .B1(n5225), .B2(n6572), .A(n5200), .ZN(U3028) );
  AOI22_X1 U6371 ( .A1(n6539), .A2(n5220), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5219), .ZN(n5201) );
  OAI21_X1 U6372 ( .B1(n6597), .B2(n5989), .A(n5201), .ZN(n5202) );
  AOI21_X1 U6373 ( .B1(n6600), .B2(n5223), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6374 ( .B1(n5225), .B2(n6603), .A(n5203), .ZN(U3033) );
  AOI22_X1 U6375 ( .A1(n6543), .A2(n5220), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5219), .ZN(n5204) );
  OAI21_X1 U6376 ( .B1(n6604), .B2(n5989), .A(n5204), .ZN(n5205) );
  AOI21_X1 U6377 ( .B1(n6609), .B2(n5223), .A(n5205), .ZN(n5206) );
  OAI21_X1 U6378 ( .B1(n5225), .B2(n6612), .A(n5206), .ZN(U3034) );
  AOI22_X1 U6379 ( .A1(n6527), .A2(n5220), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5219), .ZN(n5207) );
  OAI21_X1 U6380 ( .B1(n6580), .B2(n5989), .A(n5207), .ZN(n5208) );
  AOI21_X1 U6381 ( .B1(n6583), .B2(n5223), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6382 ( .B1(n5225), .B2(n6586), .A(n5209), .ZN(U3030) );
  AOI22_X1 U6383 ( .A1(n6530), .A2(n5220), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5219), .ZN(n5210) );
  OAI21_X1 U6384 ( .B1(n6635), .B2(n5989), .A(n5210), .ZN(n5211) );
  AOI21_X1 U6385 ( .B1(n6531), .B2(n5223), .A(n5211), .ZN(n5212) );
  OAI21_X1 U6386 ( .B1(n5225), .B2(n6591), .A(n5212), .ZN(U3031) );
  AOI22_X1 U6387 ( .A1(n6535), .A2(n5220), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5219), .ZN(n5213) );
  OAI21_X1 U6388 ( .B1(n6592), .B2(n5989), .A(n5213), .ZN(n5214) );
  AOI21_X1 U6389 ( .B1(n6594), .B2(n5223), .A(n5214), .ZN(n5215) );
  OAI21_X1 U6390 ( .B1(n5225), .B2(n7200), .A(n5215), .ZN(U3032) );
  AOI22_X1 U6391 ( .A1(n6521), .A2(n5220), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5219), .ZN(n5216) );
  OAI21_X1 U6392 ( .B1(n6525), .B2(n5989), .A(n5216), .ZN(n5217) );
  AOI21_X1 U6393 ( .B1(n6522), .B2(n5223), .A(n5217), .ZN(n5218) );
  OAI21_X1 U6394 ( .B1(n5225), .B2(n6579), .A(n5218), .ZN(U3029) );
  AOI22_X1 U6395 ( .A1(n6547), .A2(n5220), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5219), .ZN(n5221) );
  OAI21_X1 U6396 ( .B1(n6555), .B2(n5989), .A(n5221), .ZN(n5222) );
  AOI21_X1 U6397 ( .B1(n6551), .B2(n5223), .A(n5222), .ZN(n5224) );
  OAI21_X1 U6398 ( .B1(n5225), .B2(n6623), .A(n5224), .ZN(U3035) );
  NAND2_X1 U6399 ( .A1(n5326), .A2(n6210), .ZN(n5235) );
  INV_X1 U6400 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U6401 ( .A1(n6217), .A2(n5226), .ZN(n6193) );
  NAND2_X1 U6402 ( .A1(n6725), .A2(n6193), .ZN(n5233) );
  NAND2_X1 U6403 ( .A1(n5226), .A2(REIP_REG_9__SCAN_IN), .ZN(n5227) );
  INV_X1 U6404 ( .A(n5548), .ZN(n6243) );
  AOI21_X1 U6405 ( .B1(n6217), .B2(n5227), .A(n6243), .ZN(n6197) );
  INV_X1 U6406 ( .A(n6197), .ZN(n5232) );
  OAI21_X1 U6407 ( .B1(n6227), .B2(n7009), .A(n6226), .ZN(n5228) );
  AOI21_X1 U6408 ( .B1(n6249), .B2(n6417), .A(n5228), .ZN(n5229) );
  OAI21_X1 U6409 ( .B1(n6251), .B2(n5230), .A(n5229), .ZN(n5231) );
  AOI21_X1 U6410 ( .B1(n5233), .B2(n5232), .A(n5231), .ZN(n5234) );
  OAI211_X1 U6411 ( .C1(n6257), .C2(n5324), .A(n5235), .B(n5234), .ZN(U2818)
         );
  CLKBUF_X1 U6412 ( .A(n5236), .Z(n5260) );
  NOR2_X1 U6413 ( .A1(n5073), .A2(n5237), .ZN(n5238) );
  OR2_X1 U6414 ( .A1(n5260), .A2(n5238), .ZN(n6265) );
  AOI22_X1 U6415 ( .A1(n5645), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6279), .ZN(n5239) );
  OAI21_X1 U6416 ( .B1(n6265), .B2(n6054), .A(n5239), .ZN(U2881) );
  OAI21_X1 U6417 ( .B1(n5242), .B2(n5241), .A(n5240), .ZN(n6426) );
  INV_X1 U6418 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6419 ( .A1(n6471), .A2(REIP_REG_8__SCAN_IN), .ZN(n6423) );
  OAI21_X1 U6420 ( .B1(n5780), .B2(n5243), .A(n6423), .ZN(n5246) );
  NOR2_X1 U6421 ( .A1(n5244), .A2(n5766), .ZN(n5245) );
  AOI211_X1 U6422 ( .C1(n5782), .C2(n5247), .A(n5246), .B(n5245), .ZN(n5248)
         );
  OAI21_X1 U6423 ( .B1(n6426), .B2(n6125), .A(n5248), .ZN(U2978) );
  AOI21_X1 U6424 ( .B1(n6217), .B2(n5249), .A(n6243), .ZN(n6221) );
  NAND2_X1 U6425 ( .A1(n6249), .A2(n6443), .ZN(n5250) );
  OAI211_X1 U6426 ( .C1(n6227), .C2(n5251), .A(n5250), .B(n6226), .ZN(n5252)
         );
  AOI21_X1 U6427 ( .B1(EBX_REG_6__SCAN_IN), .B2(n6224), .A(n5252), .ZN(n5253)
         );
  NAND4_X1 U6428 ( .A1(n6217), .A2(REIP_REG_5__SCAN_IN), .A3(n6216), .A4(n6720), .ZN(n6204) );
  OAI211_X1 U6429 ( .C1(n6221), .C2(n6720), .A(n5253), .B(n6204), .ZN(n5257)
         );
  OAI22_X1 U6430 ( .A1(n6257), .A2(n5255), .B1(n6198), .B2(n5254), .ZN(n5256)
         );
  OR2_X1 U6431 ( .A1(n5257), .A2(n5256), .ZN(U2821) );
  OR2_X1 U6432 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U6433 ( .A1(n5258), .A2(n5261), .ZN(n5415) );
  AOI21_X1 U6434 ( .B1(n5262), .B2(n5394), .A(n3266), .ZN(n6408) );
  AOI22_X1 U6435 ( .A1(n6408), .A2(n6259), .B1(n5263), .B2(EBX_REG_11__SCAN_IN), .ZN(n5264) );
  OAI21_X1 U6436 ( .B1(n5415), .B2(n5626), .A(n5264), .ZN(U2848) );
  INV_X1 U6437 ( .A(n5267), .ZN(n5265) );
  AOI21_X1 U6438 ( .B1(n3463), .B2(n5265), .A(n6210), .ZN(n5547) );
  NOR2_X1 U6439 ( .A1(n5267), .A2(n5266), .ZN(n6242) );
  INV_X1 U6440 ( .A(n6242), .ZN(n5269) );
  OAI22_X1 U6441 ( .A1(n3595), .A2(n5269), .B1(n6234), .B2(n5268), .ZN(n5272)
         );
  NOR2_X1 U6442 ( .A1(n6251), .A2(n5270), .ZN(n5271) );
  AOI211_X1 U6443 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5273), .A(n5272), .B(n5271), 
        .ZN(n5275) );
  OAI21_X1 U6444 ( .B1(n6212), .B2(n6244), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5274) );
  OAI211_X1 U6445 ( .C1(n5547), .C2(n6286), .A(n5275), .B(n5274), .ZN(U2827)
         );
  NOR2_X1 U6446 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5276), .ZN(n5285)
         );
  INV_X1 U6447 ( .A(n5285), .ZN(n5983) );
  NAND2_X1 U6448 ( .A1(n5277), .A2(n6669), .ZN(n6502) );
  INV_X1 U6449 ( .A(n6502), .ZN(n5278) );
  NAND2_X1 U6450 ( .A1(n5339), .A2(n5278), .ZN(n5279) );
  OAI21_X1 U6451 ( .B1(n5282), .B2(n6559), .A(n5279), .ZN(n5985) );
  INV_X1 U6452 ( .A(n5989), .ZN(n5280) );
  OAI21_X1 U6453 ( .B1(n5986), .B2(n5280), .A(n5974), .ZN(n5281) );
  NAND2_X1 U6454 ( .A1(n5282), .A2(n5281), .ZN(n5284) );
  AOI21_X1 U6455 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6502), .A(n5283), .ZN(
        n6506) );
  OAI221_X1 U6456 ( .B1(n5285), .B2(n6769), .C1(n5285), .C2(n5284), .A(n6506), 
        .ZN(n5976) );
  AOI22_X1 U6457 ( .A1(n5985), .A2(n6538), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n5976), .ZN(n5286) );
  OAI21_X1 U6458 ( .B1(n6598), .B2(n5983), .A(n5286), .ZN(n5287) );
  AOI21_X1 U6459 ( .B1(n5288), .B2(n5986), .A(n5287), .ZN(n5289) );
  OAI21_X1 U6460 ( .B1(n5290), .B2(n5989), .A(n5289), .ZN(U3041) );
  AOI22_X1 U6461 ( .A1(n5985), .A2(n6542), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n5976), .ZN(n5291) );
  OAI21_X1 U6462 ( .B1(n6606), .B2(n5983), .A(n5291), .ZN(n5292) );
  AOI21_X1 U6463 ( .B1(n5293), .B2(n5986), .A(n5292), .ZN(n5294) );
  OAI21_X1 U6464 ( .B1(n5295), .B2(n5989), .A(n5294), .ZN(U3042) );
  AOI22_X1 U6465 ( .A1(n5985), .A2(n6534), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n5976), .ZN(n5296) );
  OAI21_X1 U6466 ( .B1(n7203), .B2(n5983), .A(n5296), .ZN(n5297) );
  AOI21_X1 U6467 ( .B1(n7206), .B2(n5986), .A(n5297), .ZN(n5298) );
  OAI21_X1 U6468 ( .B1(n7209), .B2(n5989), .A(n5298), .ZN(U3040) );
  AOI22_X1 U6469 ( .A1(n5985), .A2(n6526), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n5976), .ZN(n5299) );
  OAI21_X1 U6470 ( .B1(n6581), .B2(n5983), .A(n5299), .ZN(n5300) );
  AOI21_X1 U6471 ( .B1(n5301), .B2(n5986), .A(n5300), .ZN(n5302) );
  OAI21_X1 U6472 ( .B1(n5303), .B2(n5989), .A(n5302), .ZN(U3038) );
  AOI22_X1 U6473 ( .A1(n5985), .A2(n6520), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n5976), .ZN(n5304) );
  OAI21_X1 U6474 ( .B1(n6574), .B2(n5983), .A(n5304), .ZN(n5305) );
  AOI21_X1 U6475 ( .B1(n6576), .B2(n5986), .A(n5305), .ZN(n5306) );
  OAI21_X1 U6476 ( .B1(n6573), .B2(n5989), .A(n5306), .ZN(U3037) );
  AOI22_X1 U6477 ( .A1(n5985), .A2(n6638), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n5976), .ZN(n5307) );
  OAI21_X1 U6478 ( .B1(n6634), .B2(n5983), .A(n5307), .ZN(n5308) );
  AOI21_X1 U6479 ( .B1(n6588), .B2(n5986), .A(n5308), .ZN(n5309) );
  OAI21_X1 U6480 ( .B1(n6643), .B2(n5989), .A(n5309), .ZN(U3039) );
  INV_X1 U6481 ( .A(DATAI_11_), .ZN(n5310) );
  INV_X1 U6482 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6922) );
  OAI222_X1 U6483 ( .A1(n5415), .A2(n6054), .B1(n6284), .B2(n5310), .C1(n6285), 
        .C2(n6922), .ZN(U2880) );
  OAI21_X1 U6484 ( .B1(n5311), .B2(n6193), .A(n6728), .ZN(n5317) );
  OAI21_X1 U6485 ( .B1(n5425), .B2(n6247), .A(n5548), .ZN(n6185) );
  NAND2_X1 U6486 ( .A1(n6408), .A2(n6249), .ZN(n5312) );
  OAI211_X1 U6487 ( .C1(n5313), .C2(n6227), .A(n5312), .B(n6226), .ZN(n5314)
         );
  AOI21_X1 U6488 ( .B1(EBX_REG_11__SCAN_IN), .B2(n6224), .A(n5314), .ZN(n5315)
         );
  OAI21_X1 U6489 ( .B1(n6257), .B2(n5410), .A(n5315), .ZN(n5316) );
  AOI21_X1 U6490 ( .B1(n5317), .B2(n6185), .A(n5316), .ZN(n5318) );
  OAI21_X1 U6491 ( .B1(n6198), .B2(n5415), .A(n5318), .ZN(U2816) );
  NAND2_X1 U6492 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  XNOR2_X1 U6493 ( .A(n5319), .B(n5322), .ZN(n6419) );
  INV_X1 U6494 ( .A(n6419), .ZN(n5328) );
  NAND2_X1 U6495 ( .A1(n6471), .A2(REIP_REG_9__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U6496 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5323)
         );
  OAI211_X1 U6497 ( .C1(n6406), .C2(n5324), .A(n6415), .B(n5323), .ZN(n5325)
         );
  AOI21_X1 U6498 ( .B1(n5326), .B2(n6400), .A(n5325), .ZN(n5327) );
  OAI21_X1 U6499 ( .B1(n5328), .B2(n6125), .A(n5327), .ZN(U2977) );
  INV_X1 U6500 ( .A(n4605), .ZN(n5329) );
  AOI22_X1 U6501 ( .A1(n6242), .A2(n5329), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6244), .ZN(n5330) );
  OAI21_X1 U6502 ( .B1(n6234), .B2(n6470), .A(n5330), .ZN(n5332) );
  NOR2_X1 U6503 ( .A1(n6257), .A2(n6405), .ZN(n5331) );
  AOI211_X1 U6504 ( .C1(EBX_REG_2__SCAN_IN), .C2(n6224), .A(n5332), .B(n5331), 
        .ZN(n5335) );
  INV_X1 U6505 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6715) );
  AOI211_X1 U6506 ( .C1(n6217), .C2(n6998), .A(n6243), .B(n6715), .ZN(n6238)
         );
  AOI221_X1 U6507 ( .B1(n6998), .B2(n6715), .C1(n6247), .C2(n6715), .A(n6238), 
        .ZN(n5333) );
  INV_X1 U6508 ( .A(n5333), .ZN(n5334) );
  OAI211_X1 U6509 ( .C1(n5547), .C2(n6399), .A(n5335), .B(n5334), .ZN(U2825)
         );
  NAND2_X1 U6510 ( .A1(n5340), .A2(n6642), .ZN(n5336) );
  AOI21_X1 U6511 ( .B1(n5336), .B2(STATEBS16_REG_SCAN_IN), .A(n6559), .ZN(
        n5345) );
  INV_X1 U6512 ( .A(n5337), .ZN(n5338) );
  NOR2_X1 U6513 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5341), .ZN(n5370)
         );
  INV_X1 U6514 ( .A(n5342), .ZN(n5344) );
  INV_X1 U6515 ( .A(n5370), .ZN(n5343) );
  AOI22_X1 U6516 ( .A1(n5345), .A2(n5344), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5343), .ZN(n5346) );
  NAND3_X1 U6517 ( .A1(n5347), .A2(n5346), .A3(n6503), .ZN(n5369) );
  AOI22_X1 U6518 ( .A1(n6530), .A2(n5370), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5369), .ZN(n5348) );
  OAI21_X1 U6519 ( .B1(n6635), .B2(n6642), .A(n5348), .ZN(n5349) );
  AOI21_X1 U6520 ( .B1(n5373), .B2(n6531), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6521 ( .B1(n5375), .B2(n6591), .A(n5350), .ZN(U3103) );
  AOI22_X1 U6522 ( .A1(n6505), .A2(n5370), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5369), .ZN(n5351) );
  OAI21_X1 U6523 ( .B1(n6627), .B2(n6642), .A(n5351), .ZN(n5352) );
  AOI21_X1 U6524 ( .B1(n6517), .B2(n5373), .A(n5352), .ZN(n5353) );
  OAI21_X1 U6525 ( .B1(n5375), .B2(n6572), .A(n5353), .ZN(U3100) );
  AOI22_X1 U6526 ( .A1(n6535), .A2(n5370), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5369), .ZN(n5354) );
  OAI21_X1 U6527 ( .B1(n6592), .B2(n6642), .A(n5354), .ZN(n5355) );
  AOI21_X1 U6528 ( .B1(n5373), .B2(n6594), .A(n5355), .ZN(n5356) );
  OAI21_X1 U6529 ( .B1(n5375), .B2(n7200), .A(n5356), .ZN(U3104) );
  AOI22_X1 U6530 ( .A1(n6539), .A2(n5370), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5369), .ZN(n5357) );
  OAI21_X1 U6531 ( .B1(n6597), .B2(n6642), .A(n5357), .ZN(n5358) );
  AOI21_X1 U6532 ( .B1(n5373), .B2(n6600), .A(n5358), .ZN(n5359) );
  OAI21_X1 U6533 ( .B1(n5375), .B2(n6603), .A(n5359), .ZN(U3105) );
  AOI22_X1 U6534 ( .A1(n6527), .A2(n5370), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5369), .ZN(n5360) );
  OAI21_X1 U6535 ( .B1(n6580), .B2(n6642), .A(n5360), .ZN(n5361) );
  AOI21_X1 U6536 ( .B1(n5373), .B2(n6583), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6537 ( .B1(n5375), .B2(n6586), .A(n5362), .ZN(U3102) );
  AOI22_X1 U6538 ( .A1(n6543), .A2(n5370), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5369), .ZN(n5363) );
  OAI21_X1 U6539 ( .B1(n6604), .B2(n6642), .A(n5363), .ZN(n5364) );
  AOI21_X1 U6540 ( .B1(n5373), .B2(n6609), .A(n5364), .ZN(n5365) );
  OAI21_X1 U6541 ( .B1(n5375), .B2(n6612), .A(n5365), .ZN(U3106) );
  AOI22_X1 U6542 ( .A1(n6521), .A2(n5370), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5369), .ZN(n5366) );
  OAI21_X1 U6543 ( .B1(n6525), .B2(n6642), .A(n5366), .ZN(n5367) );
  AOI21_X1 U6544 ( .B1(n5373), .B2(n6522), .A(n5367), .ZN(n5368) );
  OAI21_X1 U6545 ( .B1(n5375), .B2(n6579), .A(n5368), .ZN(U3101) );
  AOI22_X1 U6546 ( .A1(n6547), .A2(n5370), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5369), .ZN(n5371) );
  OAI21_X1 U6547 ( .B1(n6555), .B2(n6642), .A(n5371), .ZN(n5372) );
  AOI21_X1 U6548 ( .B1(n5373), .B2(n6551), .A(n5372), .ZN(n5374) );
  OAI21_X1 U6549 ( .B1(n5375), .B2(n6623), .A(n5374), .ZN(U3107) );
  AOI21_X1 U6550 ( .B1(n5377), .B2(n5258), .A(n5376), .ZN(n6260) );
  INV_X1 U6551 ( .A(n6260), .ZN(n5380) );
  INV_X1 U6552 ( .A(DATAI_12_), .ZN(n5378) );
  OAI222_X1 U6553 ( .A1(n5380), .A2(n6054), .B1(n6285), .B2(n5379), .C1(n5378), 
        .C2(n6284), .ZN(U2879) );
  NAND2_X1 U6554 ( .A1(n5405), .A2(n5382), .ZN(n5383) );
  XNOR2_X1 U6555 ( .A(n5381), .B(n5383), .ZN(n5399) );
  INV_X1 U6556 ( .A(n5399), .ZN(n5398) );
  NOR2_X1 U6557 ( .A1(n6439), .A2(n6432), .ZN(n6427) );
  INV_X1 U6558 ( .A(n5937), .ZN(n5791) );
  NOR2_X1 U6559 ( .A1(n6450), .A2(n6445), .ZN(n5385) );
  NAND2_X1 U6560 ( .A1(n5384), .A2(n5385), .ZN(n5786) );
  INV_X1 U6561 ( .A(n5935), .ZN(n5790) );
  NAND3_X1 U6562 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5385), .ZN(n5787) );
  AOI22_X1 U6563 ( .A1(n5791), .A2(n5786), .B1(n5790), .B2(n5787), .ZN(n6440)
         );
  OAI21_X1 U6564 ( .B1(n5906), .B2(n6427), .A(n6440), .ZN(n6418) );
  INV_X1 U6565 ( .A(n6469), .ZN(n6455) );
  NAND2_X1 U6566 ( .A1(n6427), .A2(n6435), .ZN(n6422) );
  AOI221_X1 U6567 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5387), .C2(n5386), .A(n6422), 
        .ZN(n5388) );
  AOI21_X1 U6568 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6418), .A(n5388), 
        .ZN(n5397) );
  INV_X1 U6569 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6570 ( .A1(n5391), .A2(n5390), .ZN(n5393) );
  NAND2_X1 U6571 ( .A1(n5393), .A2(n5392), .ZN(n5395) );
  AND2_X1 U6572 ( .A1(n5395), .A2(n5394), .ZN(n6263) );
  AND2_X1 U6573 ( .A1(n6471), .A2(REIP_REG_10__SCAN_IN), .ZN(n5402) );
  AOI21_X1 U6574 ( .B1(n6263), .B2(n6487), .A(n5402), .ZN(n5396) );
  OAI211_X1 U6575 ( .C1(n5398), .C2(n6489), .A(n5397), .B(n5396), .ZN(U3008)
         );
  NAND2_X1 U6576 ( .A1(n5399), .A2(n6402), .ZN(n5404) );
  NOR2_X1 U6577 ( .A1(n6406), .A2(n5400), .ZN(n5401) );
  AOI211_X1 U6578 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5402), 
        .B(n5401), .ZN(n5403) );
  OAI211_X1 U6579 ( .C1(n5766), .C2(n6265), .A(n5404), .B(n5403), .ZN(U2976)
         );
  NAND2_X1 U6580 ( .A1(n5406), .A2(n5405), .ZN(n5409) );
  XNOR2_X1 U6581 ( .A(n3194), .B(n5407), .ZN(n5408) );
  XNOR2_X1 U6582 ( .A(n5409), .B(n5408), .ZN(n6411) );
  NAND2_X1 U6583 ( .A1(n6411), .A2(n6402), .ZN(n5414) );
  INV_X1 U6584 ( .A(n5410), .ZN(n5412) );
  OAI22_X1 U6585 ( .A1(n5780), .A2(n5313), .B1(n6461), .B2(n6728), .ZN(n5411)
         );
  AOI21_X1 U6586 ( .B1(n5782), .B2(n5412), .A(n5411), .ZN(n5413) );
  OAI211_X1 U6587 ( .C1(n5766), .C2(n5415), .A(n5414), .B(n5413), .ZN(U2975)
         );
  OAI21_X1 U6588 ( .B1(n5416), .B2(n5419), .A(n5418), .ZN(n5769) );
  NOR2_X1 U6589 ( .A1(n6257), .A2(n5771), .ZN(n5430) );
  NOR3_X1 U6590 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6247), .A3(n5420), .ZN(n5429) );
  AND2_X1 U6591 ( .A1(n5956), .A2(n5421), .ZN(n5422) );
  NOR2_X1 U6592 ( .A1(n5441), .A2(n5422), .ZN(n5952) );
  AOI22_X1 U6593 ( .A1(n5952), .A2(n6249), .B1(EBX_REG_13__SCAN_IN), .B2(n6224), .ZN(n5423) );
  OAI211_X1 U6594 ( .C1(n6227), .C2(n5424), .A(n5423), .B(n6226), .ZN(n5428)
         );
  INV_X1 U6595 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6729) );
  AND3_X1 U6596 ( .A1(n6217), .A2(n6729), .A3(n5425), .ZN(n6186) );
  OAI21_X1 U6597 ( .B1(n6185), .B2(n6186), .A(REIP_REG_13__SCAN_IN), .ZN(n5426) );
  INV_X1 U6598 ( .A(n5426), .ZN(n5427) );
  NOR4_X1 U6599 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n5431)
         );
  OAI21_X1 U6600 ( .B1(n5769), .B2(n6198), .A(n5431), .ZN(U2814) );
  INV_X1 U6601 ( .A(DATAI_13_), .ZN(n5432) );
  INV_X1 U6602 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7091) );
  OAI222_X1 U6603 ( .A1(n5769), .A2(n6054), .B1(n6284), .B2(n5432), .C1(n7091), 
        .C2(n6285), .ZN(U2878) );
  INV_X1 U6604 ( .A(n5952), .ZN(n5433) );
  INV_X1 U6605 ( .A(EBX_REG_13__SCAN_IN), .ZN(n7049) );
  OAI222_X1 U6606 ( .A1(n5433), .A2(n5627), .B1(n6272), .B2(n7049), .C1(n5626), 
        .C2(n5769), .ZN(U2846) );
  INV_X1 U6607 ( .A(n5434), .ZN(n5438) );
  NAND3_X1 U6608 ( .A1(n5418), .A2(n5436), .A3(n5435), .ZN(n5437) );
  NAND2_X1 U6609 ( .A1(n5438), .A2(n5437), .ZN(n6178) );
  INV_X1 U6610 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5443) );
  NOR2_X1 U6611 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  OR2_X1 U6612 ( .A1(n5439), .A2(n5442), .ZN(n6176) );
  OAI222_X1 U6613 ( .A1(n6178), .A2(n5626), .B1(n6272), .B2(n5443), .C1(n5627), 
        .C2(n6176), .ZN(U2845) );
  INV_X1 U6614 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5445) );
  INV_X1 U6615 ( .A(DATAI_14_), .ZN(n5444) );
  OAI222_X1 U6616 ( .A1(n6178), .A2(n6054), .B1(n6285), .B2(n5445), .C1(n5444), 
        .C2(n6284), .ZN(U2877) );
  NOR2_X1 U6617 ( .A1(n5447), .A2(n5446), .ZN(n5449) );
  INV_X1 U6618 ( .A(n4591), .ZN(n5452) );
  NOR3_X1 U6619 ( .A1(n5452), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6771), 
        .ZN(n5448) );
  AOI211_X1 U6620 ( .C1(n5450), .C2(n6113), .A(n5449), .B(n5448), .ZN(n5454)
         );
  AOI21_X1 U6621 ( .B1(n5452), .B2(n5451), .A(n6774), .ZN(n5453) );
  OAI22_X1 U6622 ( .A1(n6774), .A2(n5454), .B1(n5453), .B2(n3604), .ZN(U3459)
         );
  AOI22_X1 U6623 ( .A1(n6276), .A2(DATAI_30_), .B1(n6279), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5459) );
  AND2_X1 U6624 ( .A1(n3460), .A2(n3585), .ZN(n5457) );
  NAND2_X1 U6625 ( .A1(n6280), .A2(DATAI_14_), .ZN(n5458) );
  OAI211_X1 U6626 ( .C1(n5455), .C2(n6054), .A(n5459), .B(n5458), .ZN(U2861)
         );
  INV_X1 U6627 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5460) );
  OAI222_X1 U6628 ( .A1(n5626), .A2(n5455), .B1(n6272), .B2(n5460), .C1(n5812), 
        .C2(n5627), .ZN(U2829) );
  AOI21_X1 U6629 ( .B1(n5462), .B2(n3217), .A(n5461), .ZN(n5665) );
  INV_X1 U6630 ( .A(n5665), .ZN(n5633) );
  INV_X1 U6631 ( .A(n5463), .ZN(n5474) );
  INV_X1 U6632 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6934) );
  OAI211_X1 U6633 ( .C1(n5599), .C2(n5465), .A(n5569), .B(n5464), .ZN(n5466)
         );
  INV_X1 U6634 ( .A(n5466), .ZN(n5467) );
  AOI22_X1 U6635 ( .A1(n6224), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6244), .ZN(n5471) );
  INV_X1 U6636 ( .A(n5663), .ZN(n5469) );
  NAND2_X1 U6637 ( .A1(n6212), .A2(n5469), .ZN(n5470) );
  OAI211_X1 U6638 ( .C1(n5817), .C2(n6234), .A(n5471), .B(n5470), .ZN(n5473)
         );
  NOR3_X1 U6639 ( .A1(n5990), .A2(n5991), .A3(n6934), .ZN(n5472) );
  AOI211_X1 U6640 ( .C1(n5474), .C2(n6934), .A(n5473), .B(n5472), .ZN(n5475)
         );
  OAI21_X1 U6641 ( .B1(n5633), .B2(n6198), .A(n5475), .ZN(U2798) );
  NAND2_X1 U6642 ( .A1(n5477), .A2(n5478), .ZN(n5479) );
  AND2_X1 U6643 ( .A1(n5573), .A2(n5479), .ZN(n6058) );
  INV_X1 U6644 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6746) );
  NOR3_X1 U6645 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6026), .A3(n6746), .ZN(n5489) );
  INV_X1 U6646 ( .A(n5578), .ZN(n5482) );
  NAND2_X1 U6647 ( .A1(n5587), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U6648 ( .A1(n5482), .A2(n5481), .ZN(n5854) );
  OAI21_X1 U6649 ( .B1(REIP_REG_24__SCAN_IN), .B2(n6026), .A(n6037), .ZN(n5485) );
  OAI22_X1 U6650 ( .A1(n5483), .A2(n6227), .B1(n5694), .B2(n6257), .ZN(n5484)
         );
  AOI21_X1 U6651 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5485), .A(n5484), .ZN(n5487) );
  NAND2_X1 U6652 ( .A1(n6224), .A2(EBX_REG_25__SCAN_IN), .ZN(n5486) );
  OAI211_X1 U6653 ( .C1(n5854), .C2(n6234), .A(n5487), .B(n5486), .ZN(n5488)
         );
  AOI211_X1 U6654 ( .C1(n6058), .C2(n6210), .A(n5489), .B(n5488), .ZN(n5490)
         );
  INV_X1 U6655 ( .A(n5490), .ZN(U2802) );
  INV_X1 U6656 ( .A(n5491), .ZN(n5510) );
  AND2_X1 U6657 ( .A1(n5510), .A2(n5492), .ZN(n5494) );
  OR2_X1 U6658 ( .A1(n5494), .A2(n5493), .ZN(n5721) );
  INV_X1 U6659 ( .A(n5721), .ZN(n6064) );
  NAND2_X1 U6660 ( .A1(n6064), .A2(n6210), .ZN(n5505) );
  INV_X1 U6661 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7075) );
  AND2_X1 U6662 ( .A1(n7075), .A2(n6028), .ZN(n5517) );
  OAI21_X1 U6663 ( .B1(n5517), .B2(n6038), .A(REIP_REG_22__SCAN_IN), .ZN(n5504) );
  INV_X1 U6664 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6743) );
  NAND3_X1 U6665 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6028), .A3(n6743), .ZN(
        n5503) );
  OR2_X1 U6666 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  NAND2_X1 U6667 ( .A1(n5495), .A2(n5498), .ZN(n5879) );
  AOI22_X1 U6668 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6244), .B1(n5724), 
        .B2(n6212), .ZN(n5500) );
  NAND2_X1 U6669 ( .A1(n6224), .A2(EBX_REG_22__SCAN_IN), .ZN(n5499) );
  OAI211_X1 U6670 ( .C1(n5879), .C2(n6234), .A(n5500), .B(n5499), .ZN(n5501)
         );
  INV_X1 U6671 ( .A(n5501), .ZN(n5502) );
  NAND4_X1 U6672 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(U2805)
         );
  NAND2_X1 U6673 ( .A1(n5507), .A2(n5508), .ZN(n5509) );
  NAND2_X1 U6674 ( .A1(n5510), .A2(n5509), .ZN(n6067) );
  INV_X1 U6675 ( .A(n5729), .ZN(n5516) );
  XNOR2_X1 U6676 ( .A(n5512), .B(n5511), .ZN(n5885) );
  AOI22_X1 U6677 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6224), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6244), .ZN(n5513) );
  OAI21_X1 U6678 ( .B1(n5885), .B2(n6234), .A(n5513), .ZN(n5515) );
  AND2_X1 U6679 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6038), .ZN(n5514) );
  AOI211_X1 U6680 ( .C1(n5516), .C2(n6212), .A(n5515), .B(n5514), .ZN(n5519)
         );
  INV_X1 U6681 ( .A(n5517), .ZN(n5518) );
  OAI211_X1 U6682 ( .C1(n6067), .C2(n6198), .A(n5519), .B(n5518), .ZN(U2806)
         );
  AND2_X1 U6683 ( .A1(n5521), .A2(n5522), .ZN(n5523) );
  NOR2_X1 U6684 ( .A1(n5520), .A2(n5523), .ZN(n6073) );
  INV_X1 U6685 ( .A(n6073), .ZN(n5604) );
  OAI21_X1 U6686 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5540), .A(n6150), .ZN(n5535) );
  INV_X1 U6687 ( .A(n5524), .ZN(n5600) );
  MUX2_X1 U6688 ( .A(n5600), .B(n5605), .S(n5599), .Z(n5541) );
  INV_X1 U6689 ( .A(n5541), .ZN(n5527) );
  OR2_X1 U6690 ( .A1(n5598), .A2(n5527), .ZN(n5529) );
  OAI21_X1 U6691 ( .B1(n5525), .B2(n5527), .A(n5526), .ZN(n5528) );
  NAND2_X1 U6692 ( .A1(n5529), .A2(n5528), .ZN(n5916) );
  INV_X1 U6693 ( .A(n6226), .ZN(n6194) );
  AOI21_X1 U6694 ( .B1(n6244), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6194), 
        .ZN(n5530) );
  OAI21_X1 U6695 ( .B1(n5916), .B2(n6234), .A(n5530), .ZN(n5534) );
  AOI22_X1 U6696 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6224), .B1(n5531), .B2(n6736), .ZN(n5532) );
  OAI21_X1 U6697 ( .B1(n6077), .B2(n6257), .A(n5532), .ZN(n5533) );
  AOI211_X1 U6698 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5535), .A(n5534), .B(n5533), .ZN(n5536) );
  OAI21_X1 U6699 ( .B1(n5604), .B2(n6198), .A(n5536), .ZN(U2808) );
  INV_X1 U6700 ( .A(n5537), .ZN(n5538) );
  OAI21_X1 U6701 ( .B1(n5538), .B2(n3230), .A(n5521), .ZN(n5746) );
  AOI22_X1 U6702 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6224), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6244), .ZN(n5539) );
  OAI21_X1 U6703 ( .B1(n6150), .B2(n6738), .A(n5539), .ZN(n5545) );
  NOR2_X1 U6704 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5540), .ZN(n5544) );
  XNOR2_X1 U6705 ( .A(n5525), .B(n5541), .ZN(n6084) );
  INV_X1 U6706 ( .A(n6084), .ZN(n5606) );
  NAND2_X1 U6707 ( .A1(n6212), .A2(n5743), .ZN(n5542) );
  OAI211_X1 U6708 ( .C1(n5606), .C2(n6234), .A(n5542), .B(n6226), .ZN(n5543)
         );
  NOR3_X1 U6709 ( .A1(n5545), .A2(n5544), .A3(n5543), .ZN(n5546) );
  OAI21_X1 U6710 ( .B1(n5746), .B2(n6198), .A(n5546), .ZN(U2809) );
  INV_X1 U6711 ( .A(n5547), .ZN(n6255) );
  INV_X1 U6712 ( .A(n5557), .ZN(n5549) );
  OAI21_X1 U6713 ( .B1(n5549), .B2(n6247), .A(n5548), .ZN(n6237) );
  AOI22_X1 U6714 ( .A1(n6255), .A2(n5550), .B1(REIP_REG_4__SCAN_IN), .B2(n6237), .ZN(n5561) );
  AOI22_X1 U6715 ( .A1(n6249), .A2(n6453), .B1(n6242), .B2(n5551), .ZN(n5552)
         );
  OAI211_X1 U6716 ( .C1(n6227), .C2(n5553), .A(n5552), .B(n6226), .ZN(n5554)
         );
  AOI21_X1 U6717 ( .B1(n6224), .B2(EBX_REG_4__SCAN_IN), .A(n5554), .ZN(n5560)
         );
  INV_X1 U6718 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U6719 ( .A1(n6212), .A2(n5556), .ZN(n5559) );
  OR3_X1 U6720 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6247), .A3(n5557), .ZN(n5558)
         );
  NAND4_X1 U6721 ( .A1(n5561), .A2(n5560), .A3(n5559), .A4(n5558), .ZN(U2823)
         );
  OAI22_X1 U6722 ( .A1(n5785), .A2(n5627), .B1(n5562), .B2(n6272), .ZN(U2828)
         );
  OAI222_X1 U6723 ( .A1(n5563), .A2(n6272), .B1(n5627), .B2(n5817), .C1(n5633), 
        .C2(n5626), .ZN(U2830) );
  OR2_X1 U6724 ( .A1(n5564), .A2(n5565), .ZN(n5566) );
  OR2_X1 U6725 ( .A1(n5835), .A2(n5567), .ZN(n5568) );
  NAND2_X1 U6726 ( .A1(n5569), .A2(n5568), .ZN(n5994) );
  OAI22_X1 U6727 ( .A1(n5994), .A2(n5627), .B1(n5570), .B2(n6272), .ZN(n5571)
         );
  INV_X1 U6728 ( .A(n5571), .ZN(n5572) );
  OAI21_X1 U6729 ( .B1(n5636), .B2(n5626), .A(n5572), .ZN(U2831) );
  INV_X1 U6730 ( .A(n5573), .ZN(n5575) );
  INV_X1 U6731 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5580) );
  NOR2_X1 U6732 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  OR2_X1 U6733 ( .A1(n5576), .A2(n5579), .ZN(n6011) );
  OAI222_X1 U6734 ( .A1(n5626), .A2(n6012), .B1(n6272), .B2(n5580), .C1(n6011), 
        .C2(n5627), .ZN(U2833) );
  INV_X1 U6735 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5582) );
  INV_X1 U6736 ( .A(n6058), .ZN(n5581) );
  OAI222_X1 U6737 ( .A1(n5854), .A2(n5627), .B1(n5582), .B2(n6272), .C1(n5581), 
        .C2(n5626), .ZN(U2834) );
  OAI21_X1 U6738 ( .B1(n5583), .B2(n5584), .A(n5477), .ZN(n6022) );
  INV_X1 U6739 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U6740 ( .A1(n5592), .A2(n5585), .ZN(n5586) );
  NAND2_X1 U6741 ( .A1(n5587), .A2(n5586), .ZN(n6021) );
  OAI222_X1 U6742 ( .A1(n5626), .A2(n6022), .B1(n6272), .B2(n6946), .C1(n6021), 
        .C2(n5627), .ZN(U2835) );
  NOR2_X1 U6743 ( .A1(n5493), .A2(n5588), .ZN(n5589) );
  OR2_X1 U6744 ( .A1(n5583), .A2(n5589), .ZN(n6032) );
  INV_X1 U6745 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U6746 ( .A1(n5495), .A2(n5590), .ZN(n5591) );
  NAND2_X1 U6747 ( .A1(n5592), .A2(n5591), .ZN(n6031) );
  OAI222_X1 U6748 ( .A1(n5626), .A2(n6032), .B1(n6272), .B2(n5593), .C1(n6031), 
        .C2(n5627), .ZN(U2836) );
  OAI22_X1 U6749 ( .A1(n5879), .A2(n5627), .B1(n5594), .B2(n6272), .ZN(n5595)
         );
  INV_X1 U6750 ( .A(n5595), .ZN(n5596) );
  OAI21_X1 U6751 ( .B1(n5721), .B2(n5626), .A(n5596), .ZN(U2837) );
  INV_X1 U6752 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5597) );
  OAI222_X1 U6753 ( .A1(n6067), .A2(n5626), .B1(n6272), .B2(n5597), .C1(n5885), 
        .C2(n5627), .ZN(U2838) );
  MUX2_X1 U6754 ( .A(n5600), .B(n5599), .S(n5598), .Z(n5602) );
  XNOR2_X1 U6755 ( .A(n5602), .B(n5601), .ZN(n5900) );
  INV_X1 U6756 ( .A(n5900), .ZN(n6041) );
  OAI21_X1 U6757 ( .B1(n5520), .B2(n5603), .A(n5507), .ZN(n6042) );
  OAI222_X1 U6758 ( .A1(n5627), .A2(n6041), .B1(n6272), .B2(n6040), .C1(n5626), 
        .C2(n6042), .ZN(U2839) );
  INV_X1 U6759 ( .A(EBX_REG_19__SCAN_IN), .ZN(n7073) );
  OAI222_X1 U6760 ( .A1(n5916), .A2(n5627), .B1(n6272), .B2(n7073), .C1(n5626), 
        .C2(n5604), .ZN(U2840) );
  OAI222_X1 U6761 ( .A1(n5746), .A2(n5626), .B1(n5627), .B2(n5606), .C1(n5605), 
        .C2(n6272), .ZN(U2841) );
  NAND2_X1 U6762 ( .A1(n5608), .A2(n5609), .ZN(n5610) );
  AND2_X1 U6763 ( .A1(n5537), .A2(n5610), .ZN(n6273) );
  INV_X1 U6764 ( .A(n6273), .ZN(n5615) );
  INV_X1 U6765 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5614) );
  OR2_X1 U6766 ( .A1(n5611), .A2(n5612), .ZN(n5613) );
  NAND2_X1 U6767 ( .A1(n5525), .A2(n5613), .ZN(n6145) );
  OAI222_X1 U6768 ( .A1(n5615), .A2(n5626), .B1(n6272), .B2(n5614), .C1(n5627), 
        .C2(n6145), .ZN(U2842) );
  OAI21_X1 U6769 ( .B1(n5616), .B2(n5617), .A(n5608), .ZN(n6155) );
  INV_X1 U6770 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5620) );
  AND2_X1 U6771 ( .A1(n5623), .A2(n5618), .ZN(n5619) );
  OR2_X1 U6772 ( .A1(n5611), .A2(n5619), .ZN(n6152) );
  OAI222_X1 U6773 ( .A1(n6155), .A2(n5626), .B1(n6272), .B2(n5620), .C1(n5627), 
        .C2(n6152), .ZN(U2843) );
  OR2_X1 U6774 ( .A1(n5439), .A2(n5621), .ZN(n5622) );
  NAND2_X1 U6775 ( .A1(n5623), .A2(n5622), .ZN(n6165) );
  INV_X1 U6776 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7033) );
  INV_X1 U6777 ( .A(n5616), .ZN(n5624) );
  OAI21_X1 U6778 ( .B1(n5434), .B2(n5625), .A(n5624), .ZN(n6164) );
  OAI222_X1 U6779 ( .A1(n6165), .A2(n5627), .B1(n6272), .B2(n7033), .C1(n5626), 
        .C2(n6164), .ZN(U2844) );
  NAND3_X1 U6780 ( .A1(n5656), .A2(n5628), .A3(n6285), .ZN(n5630) );
  AOI22_X1 U6781 ( .A1(n6276), .A2(DATAI_31_), .B1(n6279), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U6782 ( .A1(n5630), .A2(n5629), .ZN(U2860) );
  AOI22_X1 U6783 ( .A1(n6276), .A2(DATAI_29_), .B1(n6279), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U6784 ( .A1(n6280), .A2(DATAI_13_), .ZN(n5631) );
  OAI211_X1 U6785 ( .C1(n5633), .C2(n6054), .A(n5632), .B(n5631), .ZN(U2862)
         );
  AOI22_X1 U6786 ( .A1(n6280), .A2(DATAI_12_), .B1(n6279), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6787 ( .A1(n6276), .A2(DATAI_28_), .ZN(n5634) );
  OAI211_X1 U6788 ( .C1(n5636), .C2(n6054), .A(n5635), .B(n5634), .ZN(U2863)
         );
  AOI22_X1 U6789 ( .A1(n6280), .A2(DATAI_10_), .B1(n6279), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6790 ( .A1(n6276), .A2(DATAI_26_), .ZN(n5637) );
  OAI211_X1 U6791 ( .C1(n6012), .C2(n6054), .A(n5638), .B(n5637), .ZN(U2865)
         );
  AOI22_X1 U6792 ( .A1(n6280), .A2(DATAI_8_), .B1(n6279), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U6793 ( .A1(n6276), .A2(DATAI_24_), .ZN(n5639) );
  OAI211_X1 U6794 ( .C1(n6022), .C2(n6054), .A(n5640), .B(n5639), .ZN(U2867)
         );
  AOI22_X1 U6795 ( .A1(n6280), .A2(DATAI_4_), .B1(n6279), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U6796 ( .A1(n6276), .A2(DATAI_20_), .ZN(n5641) );
  OAI211_X1 U6797 ( .C1(n6042), .C2(n6054), .A(n5642), .B(n5641), .ZN(U2871)
         );
  AOI22_X1 U6798 ( .A1(n6276), .A2(DATAI_18_), .B1(n6279), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U6799 ( .A1(n6280), .A2(DATAI_2_), .ZN(n5643) );
  OAI211_X1 U6800 ( .C1(n5746), .C2(n6054), .A(n5644), .B(n5643), .ZN(U2873)
         );
  AOI22_X1 U6801 ( .A1(n5645), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6279), .ZN(n5646) );
  OAI21_X1 U6802 ( .B1(n6164), .B2(n6054), .A(n5646), .ZN(U2876) );
  NAND2_X1 U6803 ( .A1(n5658), .A2(n3302), .ZN(n5651) );
  INV_X1 U6804 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5809) );
  NAND3_X1 U6805 ( .A1(n5648), .A2(n5809), .A3(n4414), .ZN(n5649) );
  NAND2_X1 U6806 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  XNOR2_X1 U6807 ( .A(n5652), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5808)
         );
  NOR2_X1 U6808 ( .A1(n6461), .A2(n6759), .ZN(n5795) );
  AOI21_X1 U6809 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5795), 
        .ZN(n5653) );
  OAI21_X1 U6810 ( .B1(n5808), .B2(n6125), .A(n5657), .ZN(U2955) );
  INV_X1 U6811 ( .A(n5658), .ZN(n5660) );
  NAND2_X1 U6812 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  XNOR2_X1 U6813 ( .A(n5661), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5824)
         );
  NOR2_X1 U6814 ( .A1(n6461), .A2(n6934), .ZN(n5819) );
  AOI21_X1 U6815 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5819), 
        .ZN(n5662) );
  OAI21_X1 U6816 ( .B1(n5663), .B2(n6406), .A(n5662), .ZN(n5664) );
  AOI21_X1 U6817 ( .B1(n5665), .B2(n6400), .A(n5664), .ZN(n5666) );
  OAI21_X1 U6818 ( .B1(n5824), .B2(n6125), .A(n5666), .ZN(U2957) );
  NOR3_X1 U6819 ( .A1(n4413), .A2(n4396), .A3(n7106), .ZN(n5669) );
  OR2_X1 U6820 ( .A1(n5684), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5668)
         );
  NOR2_X1 U6821 ( .A1(n5667), .A2(n5668), .ZN(n5675) );
  OAI22_X1 U6822 ( .A1(n5669), .A2(n5675), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n7106), .ZN(n5670) );
  XNOR2_X1 U6823 ( .A(n5670), .B(n7066), .ZN(n5832) );
  INV_X1 U6824 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6825 ( .A1(n5993), .A2(n5782), .ZN(n5671) );
  NAND2_X1 U6826 ( .A1(n6471), .A2(REIP_REG_28__SCAN_IN), .ZN(n5825) );
  OAI211_X1 U6827 ( .C1(n5780), .C2(n5672), .A(n5671), .B(n5825), .ZN(n5673)
         );
  AOI21_X1 U6828 ( .B1(n5996), .B2(n6400), .A(n5673), .ZN(n5674) );
  OAI21_X1 U6829 ( .B1(n5832), .B2(n6125), .A(n5674), .ZN(U2958) );
  INV_X1 U6830 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U6831 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  XNOR2_X1 U6832 ( .A(n5678), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5842)
         );
  AND2_X1 U6833 ( .A1(n5574), .A2(n5679), .ZN(n5680) );
  INV_X1 U6834 ( .A(n6050), .ZN(n6055) );
  INV_X1 U6835 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U6836 ( .A1(n6461), .A2(n6749), .ZN(n5837) );
  AOI21_X1 U6837 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5837), 
        .ZN(n5681) );
  OAI21_X1 U6838 ( .B1(n6002), .B2(n6406), .A(n5681), .ZN(n5682) );
  AOI21_X1 U6839 ( .B1(n6055), .B2(n6400), .A(n5682), .ZN(n5683) );
  OAI21_X1 U6840 ( .B1(n5842), .B2(n6125), .A(n5683), .ZN(U2959) );
  INV_X1 U6841 ( .A(n5684), .ZN(n5685) );
  NOR2_X1 U6842 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  XNOR2_X1 U6843 ( .A(n4413), .B(n5687), .ZN(n5849) );
  NAND2_X1 U6844 ( .A1(n6471), .A2(REIP_REG_26__SCAN_IN), .ZN(n5846) );
  OAI21_X1 U6845 ( .B1(n5780), .B2(n6018), .A(n5846), .ZN(n5689) );
  NOR2_X1 U6846 ( .A1(n6012), .A2(n5766), .ZN(n5688) );
  AOI211_X1 U6847 ( .C1(n5782), .C2(n6008), .A(n5689), .B(n5688), .ZN(n5690)
         );
  OAI21_X1 U6848 ( .B1(n5849), .B2(n6125), .A(n5690), .ZN(U2960) );
  AOI21_X1 U6849 ( .B1(n5692), .B2(n5667), .A(n5691), .ZN(n5857) );
  NAND2_X1 U6850 ( .A1(n6471), .A2(REIP_REG_25__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U6851 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5693)
         );
  OAI211_X1 U6852 ( .C1(n5694), .C2(n6406), .A(n5853), .B(n5693), .ZN(n5695)
         );
  AOI21_X1 U6853 ( .B1(n6058), .B2(n6400), .A(n5695), .ZN(n5696) );
  OAI21_X1 U6854 ( .B1(n5857), .B2(n6125), .A(n5696), .ZN(U2961) );
  INV_X1 U6855 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5913) );
  NOR2_X1 U6856 ( .A1(n3194), .A2(n5913), .ZN(n5697) );
  NOR2_X1 U6857 ( .A1(n5698), .A2(n3300), .ZN(n5734) );
  INV_X1 U6858 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6859 ( .A1(n3194), .A2(n5699), .ZN(n5701) );
  NOR2_X1 U6860 ( .A1(n3194), .A2(n5699), .ZN(n5700) );
  XNOR2_X1 U6861 ( .A(n3194), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5728)
         );
  NAND2_X1 U6862 ( .A1(n5727), .A2(n5728), .ZN(n5726) );
  NOR2_X1 U6863 ( .A1(n3194), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5717)
         );
  NAND2_X1 U6864 ( .A1(n3187), .A2(n5717), .ZN(n5711) );
  OAI21_X1 U6865 ( .B1(n4396), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5726), 
        .ZN(n5719) );
  NAND3_X1 U6866 ( .A1(n3194), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U6867 ( .A(n5703), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5865)
         );
  NAND2_X1 U6868 ( .A1(n6471), .A2(REIP_REG_24__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U6869 ( .B1(n5780), .B2(n5704), .A(n5860), .ZN(n5706) );
  NOR2_X1 U6870 ( .A1(n6022), .A2(n5766), .ZN(n5705) );
  AOI211_X1 U6871 ( .C1(n5782), .C2(n6019), .A(n5706), .B(n5705), .ZN(n5707)
         );
  OAI21_X1 U6872 ( .B1(n5865), .B2(n6125), .A(n5707), .ZN(U2962) );
  INV_X1 U6873 ( .A(n5912), .ZN(n5709) );
  NAND2_X1 U6874 ( .A1(n5709), .A2(n5896), .ZN(n5797) );
  INV_X1 U6875 ( .A(n5797), .ZN(n5710) );
  NAND3_X1 U6876 ( .A1(n3194), .A2(n5873), .A3(n5710), .ZN(n5712) );
  OAI21_X1 U6877 ( .B1(n5708), .B2(n5712), .A(n5711), .ZN(n5713) );
  XNOR2_X1 U6878 ( .A(n5713), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5872)
         );
  INV_X1 U6879 ( .A(n6032), .ZN(n6061) );
  NAND2_X1 U6880 ( .A1(n6471), .A2(REIP_REG_23__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6881 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5714)
         );
  OAI211_X1 U6882 ( .C1(n6029), .C2(n6406), .A(n5867), .B(n5714), .ZN(n5715)
         );
  AOI21_X1 U6883 ( .B1(n6061), .B2(n6400), .A(n5715), .ZN(n5716) );
  OAI21_X1 U6884 ( .B1(n5872), .B2(n6125), .A(n5716), .ZN(U2963) );
  AOI21_X1 U6885 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3194), .A(n5717), 
        .ZN(n5718) );
  XNOR2_X1 U6886 ( .A(n5719), .B(n5718), .ZN(n5883) );
  NAND2_X1 U6887 ( .A1(n6471), .A2(REIP_REG_22__SCAN_IN), .ZN(n5877) );
  OAI21_X1 U6888 ( .B1(n5780), .B2(n5720), .A(n5877), .ZN(n5723) );
  NOR2_X1 U6889 ( .A1(n5721), .A2(n5766), .ZN(n5722) );
  AOI211_X1 U6890 ( .C1(n5782), .C2(n5724), .A(n5723), .B(n5722), .ZN(n5725)
         );
  OAI21_X1 U6891 ( .B1(n5883), .B2(n6125), .A(n5725), .ZN(U2964) );
  OAI21_X1 U6892 ( .B1(n5728), .B2(n5727), .A(n3199), .ZN(n5884) );
  NAND2_X1 U6893 ( .A1(n5884), .A2(n6402), .ZN(n5732) );
  NOR2_X1 U6894 ( .A1(n6461), .A2(n7075), .ZN(n5886) );
  NOR2_X1 U6895 ( .A1(n5729), .A2(n6406), .ZN(n5730) );
  AOI211_X1 U6896 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5886), 
        .B(n5730), .ZN(n5731) );
  OAI211_X1 U6897 ( .C1(n5766), .C2(n6067), .A(n5732), .B(n5731), .ZN(U2965)
         );
  XNOR2_X1 U6898 ( .A(n3194), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733)
         );
  XNOR2_X1 U6899 ( .A(n5734), .B(n5733), .ZN(n5909) );
  INV_X1 U6900 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5735) );
  NOR2_X1 U6901 ( .A1(n6461), .A2(n5735), .ZN(n5899) );
  NOR2_X1 U6902 ( .A1(n5780), .A2(n6039), .ZN(n5736) );
  AOI211_X1 U6903 ( .C1(n6045), .C2(n5782), .A(n5899), .B(n5736), .ZN(n5739)
         );
  INV_X1 U6904 ( .A(n6042), .ZN(n5737) );
  NAND2_X1 U6905 ( .A1(n5737), .A2(n6400), .ZN(n5738) );
  OAI211_X1 U6906 ( .C1(n5909), .C2(n6125), .A(n5739), .B(n5738), .ZN(U2966)
         );
  NOR3_X1 U6907 ( .A1(n5708), .A2(n4396), .A3(n6082), .ZN(n5927) );
  OR2_X1 U6908 ( .A1(n3194), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5922)
         );
  NOR3_X1 U6909 ( .A1(n5740), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5922), 
        .ZN(n5924) );
  NOR2_X1 U6910 ( .A1(n5927), .A2(n5924), .ZN(n5741) );
  XNOR2_X1 U6911 ( .A(n5741), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6085)
         );
  NAND2_X1 U6912 ( .A1(n6085), .A2(n6402), .ZN(n5745) );
  OAI22_X1 U6913 ( .A1(n5780), .A2(n3906), .B1(n6461), .B2(n6738), .ZN(n5742)
         );
  AOI21_X1 U6914 ( .B1(n5782), .B2(n5743), .A(n5742), .ZN(n5744) );
  OAI211_X1 U6915 ( .C1(n5766), .C2(n5746), .A(n5745), .B(n5744), .ZN(U2968)
         );
  MUX2_X1 U6916 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n6098), .S(n3194), 
        .Z(n5748) );
  AOI21_X1 U6917 ( .B1(n4396), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5708), 
        .ZN(n5747) );
  AOI21_X1 U6918 ( .B1(n5749), .B2(n5748), .A(n5747), .ZN(n6095) );
  NAND2_X1 U6919 ( .A1(n6095), .A2(n6402), .ZN(n5753) );
  INV_X1 U6920 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5750) );
  NOR2_X1 U6921 ( .A1(n6461), .A2(n5750), .ZN(n6089) );
  NOR2_X1 U6922 ( .A1(n6406), .A2(n6151), .ZN(n5751) );
  AOI211_X1 U6923 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6089), 
        .B(n5751), .ZN(n5752) );
  OAI211_X1 U6924 ( .C1(n5766), .C2(n6155), .A(n5753), .B(n5752), .ZN(U2970)
         );
  NAND2_X1 U6925 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  NAND2_X1 U6926 ( .A1(n5740), .A2(n5756), .ZN(n5939) );
  NAND2_X1 U6927 ( .A1(n5939), .A2(n6402), .ZN(n5760) );
  INV_X1 U6928 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5757) );
  NOR2_X1 U6929 ( .A1(n6461), .A2(n5757), .ZN(n5941) );
  NOR2_X1 U6930 ( .A1(n6406), .A2(n6166), .ZN(n5758) );
  AOI211_X1 U6931 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5941), 
        .B(n5758), .ZN(n5759) );
  OAI211_X1 U6932 ( .C1(n5766), .C2(n6164), .A(n5760), .B(n5759), .ZN(U2971)
         );
  XNOR2_X1 U6933 ( .A(n3194), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5762)
         );
  XNOR2_X1 U6934 ( .A(n5761), .B(n5762), .ZN(n6106) );
  NAND2_X1 U6935 ( .A1(n6106), .A2(n6402), .ZN(n5765) );
  NOR2_X1 U6936 ( .A1(n6461), .A2(n6732), .ZN(n6100) );
  NOR2_X1 U6937 ( .A1(n6406), .A2(n6179), .ZN(n5763) );
  AOI211_X1 U6938 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6100), 
        .B(n5763), .ZN(n5764) );
  OAI211_X1 U6939 ( .C1(n5766), .C2(n6178), .A(n5765), .B(n5764), .ZN(U2972)
         );
  XOR2_X1 U6940 ( .A(n5767), .B(n5768), .Z(n5954) );
  INV_X1 U6941 ( .A(n5769), .ZN(n5773) );
  NOR2_X1 U6942 ( .A1(n6461), .A2(n6906), .ZN(n5951) );
  AOI21_X1 U6943 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5951), 
        .ZN(n5770) );
  OAI21_X1 U6944 ( .B1(n5771), .B2(n6406), .A(n5770), .ZN(n5772) );
  AOI21_X1 U6945 ( .B1(n5773), .B2(n6400), .A(n5772), .ZN(n5774) );
  OAI21_X1 U6946 ( .B1(n5954), .B2(n6125), .A(n5774), .ZN(U2973) );
  NOR2_X1 U6947 ( .A1(n5777), .A2(n3244), .ZN(n5778) );
  XNOR2_X1 U6948 ( .A(n5775), .B(n5778), .ZN(n5963) );
  NOR2_X1 U6949 ( .A1(n6461), .A2(n6729), .ZN(n5960) );
  INV_X1 U6950 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U6951 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  AOI211_X1 U6952 ( .C1(n5782), .C2(n6187), .A(n5960), .B(n5781), .ZN(n5784)
         );
  NAND2_X1 U6953 ( .A1(n6260), .A2(n6400), .ZN(n5783) );
  OAI211_X1 U6954 ( .C1(n5963), .C2(n6125), .A(n5784), .B(n5783), .ZN(U2974)
         );
  INV_X1 U6955 ( .A(n5785), .ZN(n5806) );
  NOR2_X1 U6956 ( .A1(n7109), .A2(n5850), .ZN(n5800) );
  NAND3_X1 U6957 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6427), .ZN(n5788) );
  NOR2_X1 U6958 ( .A1(n5786), .A2(n5788), .ZN(n5936) );
  NAND2_X1 U6959 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5947) );
  NOR2_X1 U6960 ( .A1(n5949), .A2(n5947), .ZN(n6109) );
  NAND2_X1 U6961 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6109), .ZN(n6091) );
  NAND2_X1 U6962 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6093) );
  NOR2_X1 U6963 ( .A1(n6091), .A2(n6093), .ZN(n5895) );
  NAND2_X1 U6964 ( .A1(n5936), .A2(n5895), .ZN(n5902) );
  NOR2_X1 U6965 ( .A1(n5788), .A2(n5787), .ZN(n5934) );
  NAND2_X1 U6966 ( .A1(n5895), .A2(n5934), .ZN(n5796) );
  NAND2_X1 U6967 ( .A1(n5937), .A2(n5935), .ZN(n5789) );
  AOI222_X1 U6968 ( .A1(n5902), .A2(n5791), .B1(n5790), .B2(n5796), .C1(n5789), 
        .C2(n5797), .ZN(n5892) );
  OAI21_X1 U6969 ( .B1(n5873), .B2(n5906), .A(n5892), .ZN(n5870) );
  INV_X1 U6970 ( .A(n6479), .ZN(n5793) );
  AOI21_X1 U6971 ( .B1(n5793), .B2(n5792), .A(n5798), .ZN(n5794) );
  NOR2_X1 U6972 ( .A1(n5870), .A2(n5794), .ZN(n5843) );
  OAI21_X1 U6973 ( .B1(n5906), .B2(n5800), .A(n5843), .ZN(n5839) );
  AOI21_X1 U6974 ( .B1(n5801), .B2(n6493), .A(n5839), .ZN(n5821) );
  OAI21_X1 U6975 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5906), .A(n5821), 
        .ZN(n5814) );
  AOI21_X1 U6976 ( .B1(n5809), .B2(n6493), .A(n5814), .ZN(n5804) );
  INV_X1 U6977 ( .A(n5795), .ZN(n5803) );
  INV_X1 U6978 ( .A(n5796), .ZN(n5903) );
  NAND2_X1 U6979 ( .A1(n6479), .A2(n5903), .ZN(n5901) );
  AOI21_X1 U6980 ( .B1(n5902), .B2(n5901), .A(n5797), .ZN(n5888) );
  NAND2_X1 U6981 ( .A1(n5888), .A2(n5873), .ZN(n5866) );
  INV_X1 U6982 ( .A(n5798), .ZN(n5799) );
  NOR2_X1 U6983 ( .A1(n5866), .A2(n5799), .ZN(n5851) );
  NAND2_X1 U6984 ( .A1(n5851), .A2(n5800), .ZN(n5829) );
  NOR2_X1 U6985 ( .A1(n5829), .A2(n5801), .ZN(n5820) );
  NAND4_X1 U6986 ( .A1(n5820), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4511), .ZN(n5802) );
  OAI211_X1 U6987 ( .C1(n5804), .C2(n4511), .A(n5803), .B(n5802), .ZN(n5805)
         );
  AOI21_X1 U6988 ( .B1(n6487), .B2(n5806), .A(n5805), .ZN(n5807) );
  OAI21_X1 U6989 ( .B1(n5808), .B2(n6489), .A(n5807), .ZN(U2987) );
  NAND3_X1 U6990 ( .A1(n5820), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5809), .ZN(n5811) );
  OAI211_X1 U6991 ( .C1(n5812), .C2(n6463), .A(n5811), .B(n5810), .ZN(n5813)
         );
  AOI21_X1 U6992 ( .B1(n5814), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5813), 
        .ZN(n5815) );
  OAI21_X1 U6993 ( .B1(n5816), .B2(n6489), .A(n5815), .ZN(U2988) );
  NOR2_X1 U6994 ( .A1(n5817), .A2(n6463), .ZN(n5818) );
  AOI211_X1 U6995 ( .C1(n5820), .C2(n4414), .A(n5819), .B(n5818), .ZN(n5823)
         );
  OR2_X1 U6996 ( .A1(n5821), .A2(n4414), .ZN(n5822) );
  OAI211_X1 U6997 ( .C1(n5824), .C2(n6489), .A(n5823), .B(n5822), .ZN(U2989)
         );
  INV_X1 U6998 ( .A(n5994), .ZN(n5828) );
  INV_X1 U6999 ( .A(n5825), .ZN(n5827) );
  NOR3_X1 U7000 ( .A1(n5829), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n7106), 
        .ZN(n5826) );
  AOI211_X1 U7001 ( .C1(n6487), .C2(n5828), .A(n5827), .B(n5826), .ZN(n5831)
         );
  NOR2_X1 U7002 ( .A1(n5829), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5836)
         );
  OAI21_X1 U7003 ( .B1(n5839), .B2(n5836), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5830) );
  OAI211_X1 U7004 ( .C1(n5832), .C2(n6489), .A(n5831), .B(n5830), .ZN(U2990)
         );
  NOR2_X1 U7005 ( .A1(n5576), .A2(n5833), .ZN(n5834) );
  INV_X1 U7006 ( .A(n6049), .ZN(n5838) );
  AOI211_X1 U7007 ( .C1(n6487), .C2(n5838), .A(n5837), .B(n5836), .ZN(n5841)
         );
  NAND2_X1 U7008 ( .A1(n5839), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5840) );
  OAI211_X1 U7009 ( .C1(n5842), .C2(n6489), .A(n5841), .B(n5840), .ZN(U2991)
         );
  INV_X1 U7010 ( .A(n5843), .ZN(n5863) );
  XNOR2_X1 U7011 ( .A(n5850), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5844)
         );
  NAND2_X1 U7012 ( .A1(n5851), .A2(n5844), .ZN(n5845) );
  OAI211_X1 U7013 ( .C1(n6011), .C2(n6463), .A(n5846), .B(n5845), .ZN(n5847)
         );
  AOI21_X1 U7014 ( .B1(n5863), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5847), 
        .ZN(n5848) );
  OAI21_X1 U7015 ( .B1(n5849), .B2(n6489), .A(n5848), .ZN(U2992) );
  NAND2_X1 U7016 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  OAI211_X1 U7017 ( .C1(n5854), .C2(n6463), .A(n5853), .B(n5852), .ZN(n5855)
         );
  AOI21_X1 U7018 ( .B1(n5863), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5855), 
        .ZN(n5856) );
  OAI21_X1 U7019 ( .B1(n5857), .B2(n6489), .A(n5856), .ZN(U2993) );
  OAI21_X1 U7020 ( .B1(n5866), .B2(n5859), .A(n5858), .ZN(n5862) );
  OAI21_X1 U7021 ( .B1(n6021), .B2(n6463), .A(n5860), .ZN(n5861) );
  AOI21_X1 U7022 ( .B1(n5863), .B2(n5862), .A(n5861), .ZN(n5864) );
  OAI21_X1 U7023 ( .B1(n5865), .B2(n6489), .A(n5864), .ZN(U2994) );
  NOR2_X1 U7024 ( .A1(n5866), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5869)
         );
  OAI21_X1 U7025 ( .B1(n6031), .B2(n6463), .A(n5867), .ZN(n5868) );
  AOI211_X1 U7026 ( .C1(n5870), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5869), .B(n5868), .ZN(n5871) );
  OAI21_X1 U7027 ( .B1(n5872), .B2(n6489), .A(n5871), .ZN(U2995) );
  INV_X1 U7028 ( .A(n5892), .ZN(n5881) );
  INV_X1 U7029 ( .A(n5873), .ZN(n5876) );
  INV_X1 U7030 ( .A(n5874), .ZN(n5875) );
  NAND3_X1 U7031 ( .A1(n5888), .A2(n5876), .A3(n5875), .ZN(n5878) );
  OAI211_X1 U7032 ( .C1(n6463), .C2(n5879), .A(n5878), .B(n5877), .ZN(n5880)
         );
  AOI21_X1 U7033 ( .B1(n5881), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5880), 
        .ZN(n5882) );
  OAI21_X1 U7034 ( .B1(n5883), .B2(n6489), .A(n5882), .ZN(U2996) );
  INV_X1 U7035 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7036 ( .A1(n5884), .A2(n6477), .ZN(n5890) );
  NOR2_X1 U7037 ( .A1(n5885), .A2(n6463), .ZN(n5887) );
  AOI211_X1 U7038 ( .C1(n5888), .C2(n5891), .A(n5887), .B(n5886), .ZN(n5889)
         );
  OAI211_X1 U7039 ( .C1(n5892), .C2(n5891), .A(n5890), .B(n5889), .ZN(U2997)
         );
  INV_X1 U7040 ( .A(n5934), .ZN(n5894) );
  AOI21_X1 U7041 ( .B1(n5934), .B2(n5893), .A(n5936), .ZN(n6104) );
  OAI21_X1 U7042 ( .B1(n5945), .B2(n5894), .A(n6104), .ZN(n6107) );
  NAND2_X1 U7043 ( .A1(n5895), .A2(n6107), .ZN(n6081) );
  NOR4_X1 U7044 ( .A1(n5897), .A2(n5896), .A3(n5912), .A4(n6081), .ZN(n5898)
         );
  AOI211_X1 U7045 ( .C1(n5900), .C2(n6487), .A(n5899), .B(n5898), .ZN(n5908)
         );
  INV_X1 U7046 ( .A(n5901), .ZN(n5905) );
  NOR2_X1 U7047 ( .A1(n6082), .A2(n5902), .ZN(n5904) );
  OAI22_X1 U7048 ( .A1(n5937), .A2(n5904), .B1(n5935), .B2(n5903), .ZN(n5931)
         );
  AOI21_X1 U7049 ( .B1(n5905), .B2(n6082), .A(n5931), .ZN(n6088) );
  OAI21_X1 U7050 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5906), .A(n6088), 
        .ZN(n5918) );
  NAND2_X1 U7051 ( .A1(n5918), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5907) );
  OAI211_X1 U7052 ( .C1(n5909), .C2(n6489), .A(n5908), .B(n5907), .ZN(U2998)
         );
  XNOR2_X1 U7053 ( .A(n3194), .B(n5913), .ZN(n5911) );
  XNOR2_X1 U7054 ( .A(n5910), .B(n5911), .ZN(n6074) );
  INV_X1 U7055 ( .A(n6074), .ZN(n5920) );
  NOR2_X1 U7056 ( .A1(n5912), .A2(n6081), .ZN(n5914) );
  AOI22_X1 U7057 ( .A1(n6471), .A2(REIP_REG_19__SCAN_IN), .B1(n5914), .B2(
        n5913), .ZN(n5915) );
  OAI21_X1 U7058 ( .B1(n5916), .B2(n6463), .A(n5915), .ZN(n5917) );
  AOI21_X1 U7059 ( .B1(n5918), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5917), 
        .ZN(n5919) );
  OAI21_X1 U7060 ( .B1(n5920), .B2(n6489), .A(n5919), .ZN(U2999) );
  INV_X1 U7061 ( .A(n5708), .ZN(n5923) );
  AOI21_X1 U7062 ( .B1(n4396), .B2(n6098), .A(n6082), .ZN(n5921) );
  AOI21_X1 U7063 ( .B1(n5923), .B2(n5922), .A(n5921), .ZN(n5926) );
  INV_X1 U7064 ( .A(n5924), .ZN(n5925) );
  OAI21_X1 U7065 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n6078) );
  INV_X1 U7066 ( .A(n6078), .ZN(n5933) );
  INV_X1 U7067 ( .A(n6081), .ZN(n5928) );
  AOI22_X1 U7068 ( .A1(n6471), .A2(REIP_REG_17__SCAN_IN), .B1(n5928), .B2(
        n6082), .ZN(n5929) );
  OAI21_X1 U7069 ( .B1(n6145), .B2(n6463), .A(n5929), .ZN(n5930) );
  AOI21_X1 U7070 ( .B1(n5931), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5930), 
        .ZN(n5932) );
  OAI21_X1 U7071 ( .B1(n5933), .B2(n6489), .A(n5932), .ZN(U3001) );
  OAI22_X1 U7072 ( .A1(n5937), .A2(n5936), .B1(n5935), .B2(n5934), .ZN(n6407)
         );
  AND2_X1 U7073 ( .A1(n6493), .A2(n6091), .ZN(n5938) );
  NOR2_X1 U7074 ( .A1(n6407), .A2(n5938), .ZN(n6099) );
  NAND2_X1 U7075 ( .A1(n5939), .A2(n6477), .ZN(n5944) );
  INV_X1 U7076 ( .A(n6107), .ZN(n6414) );
  NOR2_X1 U7077 ( .A1(n6414), .A2(n6091), .ZN(n5942) );
  NOR2_X1 U7078 ( .A1(n6165), .A2(n6463), .ZN(n5940) );
  AOI211_X1 U7079 ( .C1(n5942), .C2(n6092), .A(n5941), .B(n5940), .ZN(n5943)
         );
  OAI211_X1 U7080 ( .C1(n6099), .C2(n6092), .A(n5944), .B(n5943), .ZN(U3003)
         );
  OR2_X1 U7081 ( .A1(n5947), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6103)
         );
  NOR2_X1 U7082 ( .A1(n6109), .A2(n5945), .ZN(n5946) );
  AOI211_X1 U7083 ( .C1(n5948), .C2(n5947), .A(n5946), .B(n6407), .ZN(n6102)
         );
  OAI22_X1 U7084 ( .A1(n6414), .A2(n6103), .B1(n6102), .B2(n5949), .ZN(n5950)
         );
  AOI211_X1 U7085 ( .C1(n6487), .C2(n5952), .A(n5951), .B(n5950), .ZN(n5953)
         );
  OAI21_X1 U7086 ( .B1(n5954), .B2(n6489), .A(n5953), .ZN(U3005) );
  XNOR2_X1 U7087 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n5407), .ZN(n5955)
         );
  AOI22_X1 U7088 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6407), .B1(n6107), .B2(n5955), .ZN(n5962) );
  INV_X1 U7089 ( .A(n5956), .ZN(n5957) );
  AOI21_X1 U7090 ( .B1(n5959), .B2(n5958), .A(n5957), .ZN(n6258) );
  AOI21_X1 U7091 ( .B1(n6258), .B2(n6487), .A(n5960), .ZN(n5961) );
  OAI211_X1 U7092 ( .C1(n5963), .C2(n6489), .A(n5962), .B(n5961), .ZN(U3006)
         );
  OAI211_X1 U7093 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4676), .A(n5968), .B(
        n6567), .ZN(n5964) );
  OAI21_X1 U7094 ( .B1(n5971), .B2(n4512), .A(n5964), .ZN(n5965) );
  MUX2_X1 U7095 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5965), .S(n6498), 
        .Z(U3464) );
  XNOR2_X1 U7096 ( .A(n4673), .B(n5968), .ZN(n5966) );
  OAI22_X1 U7097 ( .A1(n5966), .A2(n6559), .B1(n4605), .B2(n5971), .ZN(n5967)
         );
  MUX2_X1 U7098 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5967), .S(n6498), 
        .Z(U3463) );
  INV_X1 U7099 ( .A(n4715), .ZN(n5973) );
  NOR2_X1 U7100 ( .A1(n6500), .A2(n5968), .ZN(n6562) );
  NOR2_X1 U7101 ( .A1(n5969), .A2(n6562), .ZN(n5972) );
  OAI222_X1 U7102 ( .A1(n5974), .A2(n5973), .B1(n6559), .B2(n5972), .C1(n5971), 
        .C2(n5970), .ZN(n5975) );
  MUX2_X1 U7103 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5975), .S(n6498), 
        .Z(U3462) );
  INV_X1 U7104 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5977) );
  INV_X1 U7105 ( .A(n5976), .ZN(n5981) );
  OAI22_X1 U7106 ( .A1(n6626), .A2(n5983), .B1(n5977), .B2(n5981), .ZN(n5978)
         );
  AOI21_X1 U7107 ( .B1(n6629), .B2(n5985), .A(n5978), .ZN(n5980) );
  NAND2_X1 U7108 ( .A1(n5986), .A2(n6569), .ZN(n5979) );
  OAI211_X1 U7109 ( .C1(n5989), .C2(n6632), .A(n5980), .B(n5979), .ZN(U3036)
         );
  INV_X1 U7110 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5982) );
  OAI22_X1 U7111 ( .A1(n6616), .A2(n5983), .B1(n5982), .B2(n5981), .ZN(n5984)
         );
  AOI21_X1 U7112 ( .B1(n6549), .B2(n5985), .A(n5984), .ZN(n5988) );
  NAND2_X1 U7113 ( .A1(n5986), .A2(n6619), .ZN(n5987) );
  OAI211_X1 U7114 ( .C1(n5989), .C2(n6613), .A(n5988), .B(n5987), .ZN(U3043)
         );
  AND2_X1 U7115 ( .A1(n6308), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7116 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6224), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6244), .ZN(n6000) );
  NOR2_X1 U7117 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  AOI22_X1 U7118 ( .A1(n5993), .A2(n6212), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5992), .ZN(n5999) );
  NOR2_X1 U7119 ( .A1(n5994), .A2(n6234), .ZN(n5995) );
  AOI21_X1 U7120 ( .B1(n5996), .B2(n6210), .A(n5995), .ZN(n5998) );
  INV_X1 U7121 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6752) );
  NAND3_X1 U7122 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6004), .A3(n6752), .ZN(
        n5997) );
  NAND4_X1 U7123 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(U2799)
         );
  AOI22_X1 U7124 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6224), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6244), .ZN(n6001) );
  OAI21_X1 U7125 ( .B1(n6002), .B2(n6257), .A(n6001), .ZN(n6003) );
  AOI221_X1 U7126 ( .B1(n6004), .B2(n6749), .C1(n6015), .C2(
        REIP_REG_27__SCAN_IN), .A(n6003), .ZN(n6007) );
  OAI22_X1 U7127 ( .A1(n6050), .A2(n6198), .B1(n6049), .B2(n6234), .ZN(n6005)
         );
  INV_X1 U7128 ( .A(n6005), .ZN(n6006) );
  NAND2_X1 U7129 ( .A1(n6007), .A2(n6006), .ZN(U2800) );
  AOI22_X1 U7130 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6224), .B1(n6008), .B2(n6212), .ZN(n6017) );
  NAND2_X1 U7131 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6010) );
  INV_X1 U7132 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6009) );
  OAI21_X1 U7133 ( .B1(n6026), .B2(n6010), .A(n6009), .ZN(n6014) );
  OAI22_X1 U7134 ( .A1(n6012), .A2(n6198), .B1(n6011), .B2(n6234), .ZN(n6013)
         );
  AOI21_X1 U7135 ( .B1(n6015), .B2(n6014), .A(n6013), .ZN(n6016) );
  OAI211_X1 U7136 ( .C1(n6018), .C2(n6227), .A(n6017), .B(n6016), .ZN(U2801)
         );
  AOI22_X1 U7137 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6244), .B1(n6019), 
        .B2(n6212), .ZN(n6020) );
  OAI21_X1 U7138 ( .B1(n6037), .B2(n6746), .A(n6020), .ZN(n6024) );
  OAI22_X1 U7139 ( .A1(n6022), .A2(n6198), .B1(n6021), .B2(n6234), .ZN(n6023)
         );
  AOI211_X1 U7140 ( .C1(EBX_REG_24__SCAN_IN), .C2(n6224), .A(n6024), .B(n6023), 
        .ZN(n6025) );
  OAI21_X1 U7141 ( .B1(REIP_REG_24__SCAN_IN), .B2(n6026), .A(n6025), .ZN(U2803) );
  NOR2_X1 U7142 ( .A1(n6743), .A2(n7075), .ZN(n6027) );
  AOI21_X1 U7143 ( .B1(n6028), .B2(n6027), .A(REIP_REG_23__SCAN_IN), .ZN(n6036) );
  OAI22_X1 U7144 ( .A1(n3998), .A2(n6227), .B1(n6029), .B2(n6257), .ZN(n6030)
         );
  AOI21_X1 U7145 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6224), .A(n6030), .ZN(n6035)
         );
  OAI22_X1 U7146 ( .A1(n6032), .A2(n6198), .B1(n6031), .B2(n6234), .ZN(n6033)
         );
  INV_X1 U7147 ( .A(n6033), .ZN(n6034) );
  OAI211_X1 U7148 ( .C1(n6037), .C2(n6036), .A(n6035), .B(n6034), .ZN(U2804)
         );
  INV_X1 U7149 ( .A(n6038), .ZN(n6048) );
  OAI22_X1 U7150 ( .A1(n6251), .A2(n6040), .B1(n6039), .B2(n6227), .ZN(n6044)
         );
  OAI22_X1 U7151 ( .A1(n6042), .A2(n6198), .B1(n6234), .B2(n6041), .ZN(n6043)
         );
  AOI211_X1 U7152 ( .C1(n6045), .C2(n6212), .A(n6044), .B(n6043), .ZN(n6046)
         );
  OAI221_X1 U7153 ( .B1(n6048), .B2(n5735), .C1(n6048), .C2(n6047), .A(n6046), 
        .ZN(U2807) );
  OAI22_X1 U7154 ( .A1(n6050), .A2(n5626), .B1(n6049), .B2(n5627), .ZN(n6051)
         );
  INV_X1 U7155 ( .A(n6051), .ZN(n6052) );
  OAI21_X1 U7156 ( .B1(n6053), .B2(n6272), .A(n6052), .ZN(U2832) );
  AOI22_X1 U7157 ( .A1(n6055), .A2(n6277), .B1(n6276), .B2(DATAI_27_), .ZN(
        n6057) );
  AOI22_X1 U7158 ( .A1(n6280), .A2(DATAI_11_), .B1(n6279), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7159 ( .A1(n6057), .A2(n6056), .ZN(U2864) );
  AOI22_X1 U7160 ( .A1(n6058), .A2(n6277), .B1(n6276), .B2(DATAI_25_), .ZN(
        n6060) );
  AOI22_X1 U7161 ( .A1(n6280), .A2(DATAI_9_), .B1(n6279), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7162 ( .A1(n6060), .A2(n6059), .ZN(U2866) );
  AOI22_X1 U7163 ( .A1(n6061), .A2(n6277), .B1(n6276), .B2(DATAI_23_), .ZN(
        n6063) );
  AOI22_X1 U7164 ( .A1(n6280), .A2(DATAI_7_), .B1(n6279), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7165 ( .A1(n6063), .A2(n6062), .ZN(U2868) );
  AOI22_X1 U7166 ( .A1(n6064), .A2(n6277), .B1(n6276), .B2(DATAI_22_), .ZN(
        n6066) );
  AOI22_X1 U7167 ( .A1(n6280), .A2(DATAI_6_), .B1(n6279), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7168 ( .A1(n6066), .A2(n6065), .ZN(U2869) );
  INV_X1 U7169 ( .A(n6067), .ZN(n6068) );
  AOI22_X1 U7170 ( .A1(n6068), .A2(n6277), .B1(n6276), .B2(DATAI_21_), .ZN(
        n6070) );
  AOI22_X1 U7171 ( .A1(n6280), .A2(DATAI_5_), .B1(n6279), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7172 ( .A1(n6070), .A2(n6069), .ZN(U2870) );
  AOI22_X1 U7173 ( .A1(n6073), .A2(n6277), .B1(n6276), .B2(DATAI_19_), .ZN(
        n6072) );
  AOI22_X1 U7174 ( .A1(n6280), .A2(DATAI_3_), .B1(n6279), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7175 ( .A1(n6072), .A2(n6071), .ZN(U2872) );
  AOI22_X1 U7176 ( .A1(n6471), .A2(REIP_REG_19__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6076) );
  AOI22_X1 U7177 ( .A1(n6074), .A2(n6402), .B1(n6400), .B2(n6073), .ZN(n6075)
         );
  OAI211_X1 U7178 ( .C1(n6406), .C2(n6077), .A(n6076), .B(n6075), .ZN(U2967)
         );
  AOI22_X1 U7179 ( .A1(n6471), .A2(REIP_REG_17__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6080) );
  AOI22_X1 U7180 ( .A1(n6078), .A2(n6402), .B1(n6400), .B2(n6273), .ZN(n6079)
         );
  OAI211_X1 U7181 ( .C1(n6406), .C2(n6142), .A(n6080), .B(n6079), .ZN(U2969)
         );
  NOR3_X1 U7182 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6082), .A3(n6081), 
        .ZN(n6083) );
  AOI21_X1 U7183 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6471), .A(n6083), .ZN(n6087) );
  AOI22_X1 U7184 ( .A1(n6085), .A2(n6477), .B1(n6487), .B2(n6084), .ZN(n6086)
         );
  OAI211_X1 U7185 ( .C1(n6088), .C2(n4402), .A(n6087), .B(n6086), .ZN(U3000)
         );
  INV_X1 U7186 ( .A(n6152), .ZN(n6090) );
  AOI21_X1 U7187 ( .B1(n6090), .B2(n6487), .A(n6089), .ZN(n6097) );
  AOI211_X1 U7188 ( .C1(n6092), .C2(n6098), .A(n6414), .B(n6091), .ZN(n6094)
         );
  AOI22_X1 U7189 ( .A1(n6095), .A2(n6477), .B1(n6094), .B2(n6093), .ZN(n6096)
         );
  OAI211_X1 U7190 ( .C1(n6099), .C2(n6098), .A(n6097), .B(n6096), .ZN(U3002)
         );
  INV_X1 U7191 ( .A(n6176), .ZN(n6101) );
  AOI21_X1 U7192 ( .B1(n6101), .B2(n6487), .A(n6100), .ZN(n6112) );
  OAI21_X1 U7193 ( .B1(n6104), .B2(n6103), .A(n6102), .ZN(n6105) );
  AOI22_X1 U7194 ( .A1(n6106), .A2(n6477), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6105), .ZN(n6111) );
  NAND3_X1 U7195 ( .A1(n6109), .A2(n6108), .A3(n6107), .ZN(n6110) );
  NAND3_X1 U7196 ( .A1(n6112), .A2(n6111), .A3(n6110), .ZN(U3004) );
  NAND2_X1 U7197 ( .A1(n6114), .A2(n6113), .ZN(n6116) );
  OAI22_X1 U7198 ( .A1(n6117), .A2(n6116), .B1(n6115), .B2(n6780), .ZN(U3455)
         );
  INV_X1 U7199 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6713) );
  AOI21_X1 U7200 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6713), .A(n6707), .ZN(n6122) );
  INV_X1 U7201 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6118) );
  INV_X1 U7202 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6703) );
  NOR2_X2 U7203 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6703), .ZN(n6804) );
  AOI21_X1 U7204 ( .B1(n6122), .B2(n6118), .A(n6804), .ZN(U2789) );
  OAI21_X1 U7205 ( .B1(n6119), .B2(n6690), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6120) );
  OAI21_X1 U7206 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6689), .A(n6120), .ZN(
        U2790) );
  INV_X1 U7207 ( .A(n6804), .ZN(n6792) );
  CLKBUF_X1 U7208 ( .A(n6792), .Z(n6760) );
  NOR2_X1 U7209 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6123) );
  OAI21_X1 U7210 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6123), .A(n6760), .ZN(n6121)
         );
  OAI21_X1 U7211 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6760), .A(n6121), .ZN(
        U2791) );
  NOR2_X1 U7212 ( .A1(n6804), .A2(n6122), .ZN(n6765) );
  OAI21_X1 U7213 ( .B1(n6123), .B2(BS16_N), .A(n6765), .ZN(n6763) );
  OAI21_X1 U7214 ( .B1(n6765), .B2(n6124), .A(n6763), .ZN(U2792) );
  OAI21_X1 U7215 ( .B1(n6126), .B2(n7090), .A(n6125), .ZN(U2793) );
  NOR4_X1 U7216 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6130) );
  NOR4_X1 U7217 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6129)
         );
  NOR4_X1 U7218 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6128) );
  NOR4_X1 U7219 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6127) );
  NAND4_X1 U7220 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n6136)
         );
  NOR4_X1 U7221 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6134) );
  AOI211_X1 U7222 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_6__SCAN_IN), .B(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6133) );
  NOR4_X1 U7223 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6132) );
  NOR4_X1 U7224 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6131) );
  NAND4_X1 U7225 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n6135)
         );
  NOR2_X1 U7226 ( .A1(n6136), .A2(n6135), .ZN(n6790) );
  INV_X1 U7227 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6138) );
  NOR3_X1 U7228 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6139) );
  OAI21_X1 U7229 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6139), .A(n6790), .ZN(n6137)
         );
  OAI21_X1 U7230 ( .B1(n6790), .B2(n6138), .A(n6137), .ZN(U2794) );
  INV_X1 U7231 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6764) );
  AOI21_X1 U7232 ( .B1(n6998), .B2(n6764), .A(n6139), .ZN(n6141) );
  INV_X1 U7233 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6140) );
  INV_X1 U7234 ( .A(n6790), .ZN(n6785) );
  AOI22_X1 U7235 ( .A1(n6790), .A2(n6141), .B1(n6140), .B2(n6785), .ZN(U2795)
         );
  NOR2_X1 U7236 ( .A1(n5750), .A2(n5757), .ZN(n6157) );
  AOI21_X1 U7237 ( .B1(n6163), .B2(n6157), .A(REIP_REG_17__SCAN_IN), .ZN(n6149) );
  INV_X1 U7238 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6143) );
  OAI22_X1 U7239 ( .A1(n6143), .A2(n6227), .B1(n6142), .B2(n6257), .ZN(n6144)
         );
  AOI211_X1 U7240 ( .C1(EBX_REG_17__SCAN_IN), .C2(n6224), .A(n6194), .B(n6144), 
        .ZN(n6148) );
  NOR2_X1 U7241 ( .A1(n6145), .A2(n6234), .ZN(n6146) );
  AOI21_X1 U7242 ( .B1(n6273), .B2(n6210), .A(n6146), .ZN(n6147) );
  OAI211_X1 U7243 ( .C1(n6150), .C2(n6149), .A(n6148), .B(n6147), .ZN(U2810)
         );
  AOI22_X1 U7244 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6224), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6174), .ZN(n6162) );
  INV_X1 U7245 ( .A(n6151), .ZN(n6154) );
  NOR2_X1 U7246 ( .A1(n6152), .A2(n6234), .ZN(n6153) );
  AOI21_X1 U7247 ( .B1(n6212), .B2(n6154), .A(n6153), .ZN(n6161) );
  INV_X1 U7248 ( .A(n6155), .ZN(n6278) );
  OAI21_X1 U7249 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n6163), .ZN(n6158) );
  AOI21_X1 U7250 ( .B1(n6244), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6194), 
        .ZN(n6156) );
  OAI21_X1 U7251 ( .B1(n6158), .B2(n6157), .A(n6156), .ZN(n6159) );
  AOI21_X1 U7252 ( .B1(n6278), .B2(n6210), .A(n6159), .ZN(n6160) );
  NAND3_X1 U7253 ( .A1(n6162), .A2(n6161), .A3(n6160), .ZN(U2811) );
  AOI22_X1 U7254 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6224), .B1(n6163), .B2(n5757), .ZN(n6171) );
  AOI22_X1 U7255 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6244), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6174), .ZN(n6170) );
  INV_X1 U7256 ( .A(n6164), .ZN(n6168) );
  OAI22_X1 U7257 ( .A1(n6257), .A2(n6166), .B1(n6165), .B2(n6234), .ZN(n6167)
         );
  AOI21_X1 U7258 ( .B1(n6168), .B2(n6210), .A(n6167), .ZN(n6169) );
  NAND4_X1 U7259 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6226), .ZN(U2812)
         );
  NAND2_X1 U7260 ( .A1(n6732), .A2(n6172), .ZN(n6173) );
  AOI22_X1 U7261 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6224), .B1(n6174), .B2(n6173), .ZN(n6184) );
  INV_X1 U7262 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6175) );
  OAI22_X1 U7263 ( .A1(n6176), .A2(n6234), .B1(n6175), .B2(n6227), .ZN(n6177)
         );
  INV_X1 U7264 ( .A(n6177), .ZN(n6183) );
  INV_X1 U7265 ( .A(n6178), .ZN(n6181) );
  INV_X1 U7266 ( .A(n6179), .ZN(n6180) );
  AOI22_X1 U7267 ( .A1(n6181), .A2(n6210), .B1(n6180), .B2(n6212), .ZN(n6182)
         );
  NAND4_X1 U7268 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6226), .ZN(U2813)
         );
  AOI22_X1 U7269 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6224), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6185), .ZN(n6191) );
  AOI211_X1 U7270 ( .C1(n6258), .C2(n6249), .A(n6194), .B(n6186), .ZN(n6190)
         );
  AOI22_X1 U7271 ( .A1(n6260), .A2(n6210), .B1(n6187), .B2(n6212), .ZN(n6189)
         );
  NAND2_X1 U7272 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6244), .ZN(n6188)
         );
  NAND4_X1 U7273 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(U2815)
         );
  AOI22_X1 U7274 ( .A1(n6249), .A2(n6263), .B1(n6224), .B2(EBX_REG_10__SCAN_IN), .ZN(n6203) );
  AOI22_X1 U7275 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n6244), .B1(n6192), 
        .B2(n6212), .ZN(n6202) );
  NOR2_X1 U7276 ( .A1(n6193), .A2(REIP_REG_10__SCAN_IN), .ZN(n6195) );
  AOI21_X1 U7277 ( .B1(n6195), .B2(REIP_REG_9__SCAN_IN), .A(n6194), .ZN(n6201)
         );
  INV_X1 U7278 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6196) );
  OAI22_X1 U7279 ( .A1(n6265), .A2(n6198), .B1(n6197), .B2(n6196), .ZN(n6199)
         );
  INV_X1 U7280 ( .A(n6199), .ZN(n6200) );
  NAND4_X1 U7281 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(U2817)
         );
  AOI21_X1 U7282 ( .B1(n6221), .B2(n6204), .A(n6722), .ZN(n6209) );
  XNOR2_X1 U7283 ( .A(n6206), .B(n6205), .ZN(n6433) );
  NAND2_X1 U7284 ( .A1(n6244), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6207)
         );
  OAI211_X1 U7285 ( .C1(n6234), .C2(n6433), .A(n6226), .B(n6207), .ZN(n6208)
         );
  NOR2_X1 U7286 ( .A1(n6209), .A2(n6208), .ZN(n6215) );
  NAND2_X1 U7287 ( .A1(n6210), .A2(n6378), .ZN(n6214) );
  INV_X1 U7288 ( .A(n6381), .ZN(n6211) );
  NAND2_X1 U7289 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  AND3_X1 U7290 ( .A1(n6215), .A2(n6214), .A3(n6213), .ZN(n6220) );
  NAND2_X1 U7291 ( .A1(n6217), .A2(n6216), .ZN(n6222) );
  NOR2_X1 U7292 ( .A1(n6717), .A2(n6222), .ZN(n6218) );
  NAND3_X1 U7293 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6218), .A3(n6722), .ZN(n6219) );
  OAI211_X1 U7294 ( .C1(n6251), .C2(n7076), .A(n6220), .B(n6219), .ZN(U2820)
         );
  AOI21_X1 U7295 ( .B1(n6717), .B2(n6222), .A(n6221), .ZN(n6223) );
  AOI21_X1 U7296 ( .B1(EBX_REG_5__SCAN_IN), .B2(n6224), .A(n6223), .ZN(n6231)
         );
  NOR2_X1 U7297 ( .A1(n6234), .A2(n6225), .ZN(n6229) );
  OAI21_X1 U7298 ( .B1(n6227), .B2(n3683), .A(n6226), .ZN(n6228) );
  AOI211_X1 U7299 ( .C1(n6255), .C2(n6382), .A(n6229), .B(n6228), .ZN(n6230)
         );
  OAI211_X1 U7300 ( .C1(n6386), .C2(n6257), .A(n6231), .B(n6230), .ZN(U2822)
         );
  NOR2_X1 U7301 ( .A1(n6251), .A2(n6232), .ZN(n6236) );
  AOI22_X1 U7302 ( .A1(n6242), .A2(n3200), .B1(n6244), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6233) );
  OAI21_X1 U7303 ( .B1(n6234), .B2(n6462), .A(n6233), .ZN(n6235) );
  AOI211_X1 U7304 ( .C1(n6255), .C2(n6391), .A(n6236), .B(n6235), .ZN(n6240)
         );
  OAI21_X1 U7305 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6238), .A(n6237), .ZN(n6239)
         );
  OAI211_X1 U7306 ( .C1(n6257), .C2(n6394), .A(n6240), .B(n6239), .ZN(U2824)
         );
  NAND2_X1 U7307 ( .A1(n6242), .A2(n6241), .ZN(n6246) );
  AOI22_X1 U7308 ( .A1(n6244), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6243), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6245) );
  OAI211_X1 U7309 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6247), .A(n6246), .B(n6245), 
        .ZN(n6248) );
  AOI21_X1 U7310 ( .B1(n6249), .B2(n6486), .A(n6248), .ZN(n6250) );
  OAI21_X1 U7311 ( .B1(n6252), .B2(n6251), .A(n6250), .ZN(n6253) );
  AOI21_X1 U7312 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(n6256) );
  OAI21_X1 U7313 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6257), .A(n6256), 
        .ZN(U2826) );
  AOI22_X1 U7314 ( .A1(n6260), .A2(n6270), .B1(n6259), .B2(n6258), .ZN(n6261)
         );
  OAI21_X1 U7315 ( .B1(n6262), .B2(n6272), .A(n6261), .ZN(U2847) );
  INV_X1 U7316 ( .A(n6263), .ZN(n6264) );
  OAI22_X1 U7317 ( .A1(n6265), .A2(n5626), .B1(n5627), .B2(n6264), .ZN(n6266)
         );
  INV_X1 U7318 ( .A(n6266), .ZN(n6267) );
  OAI21_X1 U7319 ( .B1(n6268), .B2(n6272), .A(n6267), .ZN(U2849) );
  NOR2_X1 U7320 ( .A1(n6433), .A2(n5627), .ZN(n6269) );
  AOI21_X1 U7321 ( .B1(n6378), .B2(n6270), .A(n6269), .ZN(n6271) );
  OAI21_X1 U7322 ( .B1(n7076), .B2(n6272), .A(n6271), .ZN(U2852) );
  AOI22_X1 U7323 ( .A1(n6273), .A2(n6277), .B1(n6276), .B2(DATAI_17_), .ZN(
        n6275) );
  AOI22_X1 U7324 ( .A1(n6280), .A2(DATAI_1_), .B1(n6279), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7325 ( .A1(n6275), .A2(n6274), .ZN(U2874) );
  AOI22_X1 U7326 ( .A1(n6278), .A2(n6277), .B1(n6276), .B2(DATAI_16_), .ZN(
        n6282) );
  AOI22_X1 U7327 ( .A1(n6280), .A2(DATAI_0_), .B1(n6279), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7328 ( .A1(n6282), .A2(n6281), .ZN(U2875) );
  INV_X1 U7329 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6943) );
  OAI222_X1 U7330 ( .A1(n6286), .A2(n6054), .B1(n6285), .B2(n6943), .C1(n6284), 
        .C2(n6283), .ZN(U2891) );
  INV_X1 U7331 ( .A(n6287), .ZN(n6288) );
  AOI22_X1 U7332 ( .A1(n6308), .A2(DATAO_REG_29__SCAN_IN), .B1(n6288), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6289) );
  OAI21_X1 U7333 ( .B1(n6301), .B2(n7138), .A(n6289), .ZN(U2894) );
  INV_X1 U7334 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7128) );
  AOI22_X1 U7335 ( .A1(n6796), .A2(LWORD_REG_15__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7336 ( .B1(n7128), .B2(n6310), .A(n6290), .ZN(U2908) );
  AOI22_X1 U7337 ( .A1(n6796), .A2(LWORD_REG_14__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6291) );
  OAI21_X1 U7338 ( .B1(n5445), .B2(n6310), .A(n6291), .ZN(U2909) );
  INV_X1 U7339 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n7063) );
  INV_X1 U7340 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6292) );
  OAI222_X1 U7341 ( .A1(n6302), .A2(n7063), .B1(n6310), .B2(n7091), .C1(n6301), 
        .C2(n6292), .ZN(U2910) );
  AOI22_X1 U7342 ( .A1(n6796), .A2(LWORD_REG_12__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7343 ( .B1(n5379), .B2(n6310), .A(n6293), .ZN(U2911) );
  INV_X1 U7344 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6294) );
  OAI222_X1 U7345 ( .A1(n6302), .A2(n6294), .B1(n6310), .B2(n6922), .C1(n6301), 
        .C2(n7001), .ZN(U2912) );
  INV_X1 U7346 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n7129) );
  INV_X1 U7347 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6362) );
  INV_X1 U7348 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6295) );
  OAI222_X1 U7349 ( .A1(n6302), .A2(n7129), .B1(n6310), .B2(n6362), .C1(n6301), 
        .C2(n6295), .ZN(U2913) );
  AOI22_X1 U7350 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6298), .B1(n6308), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7351 ( .B1(n6301), .B2(n7029), .A(n6296), .ZN(U2914) );
  INV_X1 U7352 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n7110) );
  INV_X1 U7353 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6297) );
  OAI222_X1 U7354 ( .A1(n6302), .A2(n7110), .B1(n6310), .B2(n7116), .C1(n6301), 
        .C2(n6297), .ZN(U2915) );
  AOI22_X1 U7355 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6298), .B1(n6308), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6299) );
  OAI21_X1 U7356 ( .B1(n6301), .B2(n7145), .A(n6299), .ZN(U2916) );
  INV_X1 U7357 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n7011) );
  INV_X1 U7358 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6300) );
  OAI222_X1 U7359 ( .A1(n6302), .A2(n7011), .B1(n6310), .B2(n3702), .C1(n6301), 
        .C2(n6300), .ZN(U2917) );
  AOI22_X1 U7360 ( .A1(n6796), .A2(LWORD_REG_5__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6303) );
  OAI21_X1 U7361 ( .B1(n6355), .B2(n6310), .A(n6303), .ZN(U2918) );
  AOI22_X1 U7362 ( .A1(n6796), .A2(LWORD_REG_4__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7363 ( .B1(n6351), .B2(n6310), .A(n6304), .ZN(U2919) );
  AOI22_X1 U7364 ( .A1(n6796), .A2(LWORD_REG_3__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6305) );
  OAI21_X1 U7365 ( .B1(n6348), .B2(n6310), .A(n6305), .ZN(U2920) );
  AOI22_X1 U7366 ( .A1(n6796), .A2(LWORD_REG_2__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7367 ( .B1(n6345), .B2(n6310), .A(n6306), .ZN(U2921) );
  AOI22_X1 U7368 ( .A1(n6796), .A2(LWORD_REG_1__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6307) );
  OAI21_X1 U7369 ( .B1(n6342), .B2(n6310), .A(n6307), .ZN(U2922) );
  AOI22_X1 U7370 ( .A1(n6796), .A2(LWORD_REG_0__SCAN_IN), .B1(n6308), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6309) );
  OAI21_X1 U7371 ( .B1(n6943), .B2(n6310), .A(n6309), .ZN(U2923) );
  AND2_X1 U7372 ( .A1(n6371), .A2(DATAI_0_), .ZN(n6338) );
  AOI21_X1 U7373 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6353), .A(n6338), .ZN(n6311) );
  OAI21_X1 U7374 ( .B1(n6312), .B2(n6373), .A(n6311), .ZN(U2924) );
  AND2_X1 U7375 ( .A1(n6371), .A2(DATAI_1_), .ZN(n6340) );
  AOI21_X1 U7376 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6366), .A(n6340), .ZN(n6314) );
  OAI21_X1 U7377 ( .B1(n6315), .B2(n6373), .A(n6314), .ZN(U2925) );
  AND2_X1 U7378 ( .A1(n6371), .A2(DATAI_2_), .ZN(n6343) );
  AOI21_X1 U7379 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6366), .A(n6343), .ZN(n6316) );
  OAI21_X1 U7380 ( .B1(n7122), .B2(n6373), .A(n6316), .ZN(U2926) );
  AND2_X1 U7381 ( .A1(n6371), .A2(DATAI_3_), .ZN(n6346) );
  AOI21_X1 U7382 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6366), .A(n6346), .ZN(n6317) );
  OAI21_X1 U7383 ( .B1(n3922), .B2(n6373), .A(n6317), .ZN(U2927) );
  AND2_X1 U7384 ( .A1(n6371), .A2(DATAI_4_), .ZN(n6349) );
  AOI21_X1 U7385 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6366), .A(n6349), .ZN(n6318) );
  OAI21_X1 U7386 ( .B1(n7146), .B2(n6373), .A(n6318), .ZN(U2928) );
  AND2_X1 U7387 ( .A1(n6371), .A2(DATAI_5_), .ZN(n6352) );
  AOI21_X1 U7388 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6366), .A(n6352), .ZN(n6319) );
  OAI21_X1 U7389 ( .B1(n6320), .B2(n6373), .A(n6319), .ZN(U2929) );
  AND2_X1 U7390 ( .A1(n6371), .A2(DATAI_6_), .ZN(n6356) );
  AOI21_X1 U7391 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6366), .A(n6356), .ZN(n6321) );
  OAI21_X1 U7392 ( .B1(n7007), .B2(n6373), .A(n6321), .ZN(U2930) );
  AOI21_X1 U7393 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6353), .A(n6322), .ZN(n6323) );
  OAI21_X1 U7394 ( .B1(n7043), .B2(n6373), .A(n6323), .ZN(U2931) );
  AND2_X1 U7395 ( .A1(n6371), .A2(DATAI_8_), .ZN(n6358) );
  AOI21_X1 U7396 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6353), .A(n6358), .ZN(n6324) );
  OAI21_X1 U7397 ( .B1(n4018), .B2(n6373), .A(n6324), .ZN(U2932) );
  AOI21_X1 U7398 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6353), .A(n6325), .ZN(n6326) );
  OAI21_X1 U7399 ( .B1(n6932), .B2(n6373), .A(n6326), .ZN(U2933) );
  INV_X1 U7400 ( .A(DATAI_10_), .ZN(n6327) );
  NOR2_X1 U7401 ( .A1(n6328), .A2(n6327), .ZN(n6360) );
  AOI21_X1 U7402 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6353), .A(n6360), .ZN(
        n6329) );
  OAI21_X1 U7403 ( .B1(n6330), .B2(n6373), .A(n6329), .ZN(U2934) );
  AOI21_X1 U7404 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6353), .A(n6331), .ZN(
        n6332) );
  OAI21_X1 U7405 ( .B1(n6333), .B2(n6373), .A(n6332), .ZN(U2935) );
  NAND2_X1 U7406 ( .A1(n6371), .A2(DATAI_12_), .ZN(n6363) );
  INV_X1 U7407 ( .A(n6363), .ZN(n6334) );
  AOI21_X1 U7408 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6353), .A(n6334), .ZN(
        n6335) );
  OAI21_X1 U7409 ( .B1(n4094), .B2(n6373), .A(n6335), .ZN(U2936) );
  NAND2_X1 U7410 ( .A1(n6371), .A2(DATAI_14_), .ZN(n6369) );
  INV_X1 U7411 ( .A(n6369), .ZN(n6336) );
  AOI21_X1 U7412 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6353), .A(n6336), .ZN(
        n6337) );
  OAI21_X1 U7413 ( .B1(n4140), .B2(n6373), .A(n6337), .ZN(U2938) );
  AOI21_X1 U7414 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6353), .A(n6338), .ZN(n6339) );
  OAI21_X1 U7415 ( .B1(n6943), .B2(n6373), .A(n6339), .ZN(U2939) );
  AOI21_X1 U7416 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6353), .A(n6340), .ZN(n6341) );
  OAI21_X1 U7417 ( .B1(n6342), .B2(n6373), .A(n6341), .ZN(U2940) );
  AOI21_X1 U7418 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6366), .A(n6343), .ZN(n6344) );
  OAI21_X1 U7419 ( .B1(n6345), .B2(n6373), .A(n6344), .ZN(U2941) );
  AOI21_X1 U7420 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6353), .A(n6346), .ZN(n6347) );
  OAI21_X1 U7421 ( .B1(n6348), .B2(n6373), .A(n6347), .ZN(U2942) );
  AOI21_X1 U7422 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6353), .A(n6349), .ZN(n6350) );
  OAI21_X1 U7423 ( .B1(n6351), .B2(n6373), .A(n6350), .ZN(U2943) );
  AOI21_X1 U7424 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6353), .A(n6352), .ZN(n6354) );
  OAI21_X1 U7425 ( .B1(n6355), .B2(n6373), .A(n6354), .ZN(U2944) );
  AOI21_X1 U7426 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6353), .A(n6356), .ZN(n6357) );
  OAI21_X1 U7427 ( .B1(n3702), .B2(n6373), .A(n6357), .ZN(U2945) );
  AOI21_X1 U7428 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6366), .A(n6358), .ZN(n6359) );
  OAI21_X1 U7429 ( .B1(n7116), .B2(n6373), .A(n6359), .ZN(U2947) );
  AOI21_X1 U7430 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6366), .A(n6360), .ZN(
        n6361) );
  OAI21_X1 U7431 ( .B1(n6362), .B2(n6373), .A(n6361), .ZN(U2949) );
  AOI22_X1 U7432 ( .A1(n6353), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6368), .ZN(n6364) );
  NAND2_X1 U7433 ( .A1(n6364), .A2(n6363), .ZN(U2951) );
  AOI21_X1 U7434 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6366), .A(n6365), .ZN(
        n6367) );
  OAI21_X1 U7435 ( .B1(n7091), .B2(n6373), .A(n6367), .ZN(U2952) );
  AOI22_X1 U7436 ( .A1(n6353), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6368), .ZN(n6370) );
  NAND2_X1 U7437 ( .A1(n6370), .A2(n6369), .ZN(U2953) );
  AOI22_X1 U7438 ( .A1(n6353), .A2(LWORD_REG_15__SCAN_IN), .B1(n6371), .B2(
        DATAI_15_), .ZN(n6372) );
  OAI21_X1 U7439 ( .B1(n7128), .B2(n6373), .A(n6372), .ZN(U2954) );
  AOI22_X1 U7440 ( .A1(n6471), .A2(REIP_REG_7__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6380) );
  OAI21_X1 U7441 ( .B1(n3196), .B2(n6375), .A(n6374), .ZN(n6377) );
  INV_X1 U7442 ( .A(n6377), .ZN(n6436) );
  AOI22_X1 U7443 ( .A1(n6436), .A2(n6402), .B1(n6400), .B2(n6378), .ZN(n6379)
         );
  OAI211_X1 U7444 ( .C1(n6406), .C2(n6381), .A(n6380), .B(n6379), .ZN(U2979)
         );
  AOI22_X1 U7445 ( .A1(n6471), .A2(REIP_REG_5__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6385) );
  AOI22_X1 U7446 ( .A1(n6383), .A2(n6402), .B1(n6400), .B2(n6382), .ZN(n6384)
         );
  OAI211_X1 U7447 ( .C1(n6406), .C2(n6386), .A(n6385), .B(n6384), .ZN(U2981)
         );
  AOI22_X1 U7448 ( .A1(n6471), .A2(REIP_REG_3__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6393) );
  OAI21_X1 U7449 ( .B1(n6389), .B2(n6387), .A(n6388), .ZN(n6390) );
  INV_X1 U7450 ( .A(n6390), .ZN(n6465) );
  AOI22_X1 U7451 ( .A1(n6465), .A2(n6402), .B1(n6391), .B2(n6400), .ZN(n6392)
         );
  OAI211_X1 U7452 ( .C1(n6406), .C2(n6394), .A(n6393), .B(n6392), .ZN(U2983)
         );
  AOI22_X1 U7453 ( .A1(n6471), .A2(REIP_REG_2__SCAN_IN), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6404) );
  XOR2_X1 U7454 ( .A(n6396), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6397) );
  XNOR2_X1 U7455 ( .A(n6398), .B(n6397), .ZN(n6476) );
  INV_X1 U7456 ( .A(n6399), .ZN(n6401) );
  AOI22_X1 U7457 ( .A1(n6402), .A2(n6476), .B1(n6401), .B2(n6400), .ZN(n6403)
         );
  OAI211_X1 U7458 ( .C1(n6406), .C2(n6405), .A(n6404), .B(n6403), .ZN(U2984)
         );
  INV_X1 U7459 ( .A(n6407), .ZN(n6413) );
  INV_X1 U7460 ( .A(n6408), .ZN(n6409) );
  OAI22_X1 U7461 ( .A1(n6409), .A2(n6463), .B1(n6728), .B2(n6461), .ZN(n6410)
         );
  AOI21_X1 U7462 ( .B1(n6477), .B2(n6411), .A(n6410), .ZN(n6412) );
  OAI221_X1 U7463 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6414), .C1(
        n5407), .C2(n6413), .A(n6412), .ZN(U3007) );
  INV_X1 U7464 ( .A(n6415), .ZN(n6416) );
  AOI21_X1 U7465 ( .B1(n6417), .B2(n6487), .A(n6416), .ZN(n6421) );
  AOI22_X1 U7466 ( .A1(n6419), .A2(n6477), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6418), .ZN(n6420) );
  OAI211_X1 U7467 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6422), .A(n6421), 
        .B(n6420), .ZN(U3009) );
  INV_X1 U7468 ( .A(n6423), .ZN(n6424) );
  AOI21_X1 U7469 ( .B1(n6425), .B2(n6487), .A(n6424), .ZN(n6431) );
  INV_X1 U7470 ( .A(n6426), .ZN(n6429) );
  AOI21_X1 U7471 ( .B1(n6439), .B2(n6432), .A(n6427), .ZN(n6428) );
  AOI22_X1 U7472 ( .A1(n6429), .A2(n6477), .B1(n6435), .B2(n6428), .ZN(n6430)
         );
  OAI211_X1 U7473 ( .C1(n6440), .C2(n6432), .A(n6431), .B(n6430), .ZN(U3010)
         );
  INV_X1 U7474 ( .A(n6433), .ZN(n6434) );
  AOI22_X1 U7475 ( .A1(n6434), .A2(n6487), .B1(n6471), .B2(REIP_REG_7__SCAN_IN), .ZN(n6438) );
  AOI22_X1 U7476 ( .A1(n6436), .A2(n6477), .B1(n6435), .B2(n6439), .ZN(n6437)
         );
  OAI211_X1 U7477 ( .C1(n6440), .C2(n6439), .A(n6438), .B(n6437), .ZN(U3011)
         );
  INV_X1 U7478 ( .A(n6441), .ZN(n6442) );
  AOI21_X1 U7479 ( .B1(n6443), .B2(n6487), .A(n6442), .ZN(n6449) );
  INV_X1 U7480 ( .A(n6444), .ZN(n6447) );
  NOR3_X1 U7481 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6469), .A3(n6445), 
        .ZN(n6446) );
  AOI21_X1 U7482 ( .B1(n6447), .B2(n6477), .A(n6446), .ZN(n6448) );
  OAI211_X1 U7483 ( .C1(n6451), .C2(n6450), .A(n6449), .B(n6448), .ZN(U3012)
         );
  INV_X1 U7484 ( .A(n6452), .ZN(n6454) );
  AOI22_X1 U7485 ( .A1(n6454), .A2(n6477), .B1(n6487), .B2(n6453), .ZN(n6460)
         );
  AOI21_X1 U7486 ( .B1(n6473), .B2(n6475), .A(n6478), .ZN(n6467) );
  NAND2_X1 U7487 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  OAI21_X1 U7488 ( .B1(n6467), .B2(n7065), .A(n6457), .ZN(n6458) );
  OAI21_X1 U7489 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6458), .ZN(n6459) );
  OAI211_X1 U7490 ( .C1(n6718), .C2(n6461), .A(n6460), .B(n6459), .ZN(U3014)
         );
  INV_X1 U7491 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6714) );
  OAI22_X1 U7492 ( .A1(n6463), .A2(n6462), .B1(n6714), .B2(n6461), .ZN(n6464)
         );
  AOI21_X1 U7493 ( .B1(n6465), .B2(n6477), .A(n6464), .ZN(n6466) );
  OAI221_X1 U7494 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6469), .C1(n6468), .C2(n6467), .A(n6466), .ZN(U3015) );
  INV_X1 U7495 ( .A(n6470), .ZN(n6472) );
  AOI22_X1 U7496 ( .A1(n6487), .A2(n6472), .B1(n6471), .B2(REIP_REG_2__SCAN_IN), .ZN(n6483) );
  OAI221_X1 U7497 ( .B1(n6475), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n6475), .C2(n6474), .A(n6473), .ZN(n6482) );
  AOI22_X1 U7498 ( .A1(n6478), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6477), 
        .B2(n6476), .ZN(n6481) );
  NAND3_X1 U7499 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7097), .A3(n6479), 
        .ZN(n6480) );
  NAND4_X1 U7500 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(U3016)
         );
  INV_X1 U7501 ( .A(n6484), .ZN(n6492) );
  AOI21_X1 U7502 ( .B1(n6487), .B2(n6486), .A(n6485), .ZN(n6488) );
  OAI21_X1 U7503 ( .B1(n6490), .B2(n6489), .A(n6488), .ZN(n6491) );
  AOI21_X1 U7504 ( .B1(n6492), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n6491), 
        .ZN(n6497) );
  OAI211_X1 U7505 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6495), .A(n6494), 
        .B(n6493), .ZN(n6496) );
  NAND2_X1 U7506 ( .A1(n6497), .A2(n6496), .ZN(U3017) );
  NOR2_X1 U7507 ( .A1(n7080), .A2(n6498), .ZN(U3019) );
  NAND2_X1 U7508 ( .A1(n6512), .A2(n6501), .ZN(n6556) );
  OAI22_X1 U7509 ( .A1(n6556), .A2(n6559), .B1(n6503), .B2(n6502), .ZN(n6548)
         );
  AND2_X1 U7510 ( .A1(n6504), .A2(n6568), .ZN(n6546) );
  AOI22_X1 U7511 ( .A1(n6629), .A2(n6548), .B1(n6505), .B2(n6546), .ZN(n6519)
         );
  INV_X1 U7512 ( .A(n6512), .ZN(n6510) );
  OAI211_X1 U7513 ( .C1(n6546), .C2(n6769), .A(n6507), .B(n6506), .ZN(n6508)
         );
  AOI21_X1 U7514 ( .B1(n6510), .B2(n6509), .A(n6508), .ZN(n6516) );
  INV_X1 U7515 ( .A(n6550), .ZN(n6514) );
  OAI21_X1 U7516 ( .B1(n6512), .B2(n6559), .A(n6511), .ZN(n6513) );
  NAND3_X1 U7517 ( .A1(n6514), .A2(n6513), .A3(n6614), .ZN(n6515) );
  NAND2_X1 U7518 ( .A1(n6516), .A2(n6515), .ZN(n6552) );
  AOI22_X1 U7519 ( .A1(n6552), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6517), 
        .B2(n6550), .ZN(n6518) );
  OAI211_X1 U7520 ( .C1(n6627), .C2(n6614), .A(n6519), .B(n6518), .ZN(U3068)
         );
  AOI22_X1 U7521 ( .A1(n6521), .A2(n6546), .B1(n6520), .B2(n6548), .ZN(n6524)
         );
  AOI22_X1 U7522 ( .A1(n6552), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6522), 
        .B2(n6550), .ZN(n6523) );
  OAI211_X1 U7523 ( .C1(n6525), .C2(n6614), .A(n6524), .B(n6523), .ZN(U3069)
         );
  AOI22_X1 U7524 ( .A1(n6527), .A2(n6546), .B1(n6526), .B2(n6548), .ZN(n6529)
         );
  AOI22_X1 U7525 ( .A1(n6552), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6583), 
        .B2(n6550), .ZN(n6528) );
  OAI211_X1 U7526 ( .C1(n6580), .C2(n6614), .A(n6529), .B(n6528), .ZN(U3070)
         );
  AOI22_X1 U7527 ( .A1(n6530), .A2(n6546), .B1(n6638), .B2(n6548), .ZN(n6533)
         );
  AOI22_X1 U7528 ( .A1(n6552), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6531), 
        .B2(n6550), .ZN(n6532) );
  OAI211_X1 U7529 ( .C1(n6635), .C2(n6614), .A(n6533), .B(n6532), .ZN(U3071)
         );
  AOI22_X1 U7530 ( .A1(n6535), .A2(n6546), .B1(n6534), .B2(n6548), .ZN(n6537)
         );
  AOI22_X1 U7531 ( .A1(n6552), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6594), 
        .B2(n6550), .ZN(n6536) );
  OAI211_X1 U7532 ( .C1(n6592), .C2(n6614), .A(n6537), .B(n6536), .ZN(U3072)
         );
  AOI22_X1 U7533 ( .A1(n6539), .A2(n6546), .B1(n6538), .B2(n6548), .ZN(n6541)
         );
  AOI22_X1 U7534 ( .A1(n6552), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6600), 
        .B2(n6550), .ZN(n6540) );
  OAI211_X1 U7535 ( .C1(n6597), .C2(n6614), .A(n6541), .B(n6540), .ZN(U3073)
         );
  AOI22_X1 U7536 ( .A1(n6543), .A2(n6546), .B1(n6542), .B2(n6548), .ZN(n6545)
         );
  AOI22_X1 U7537 ( .A1(n6552), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6609), 
        .B2(n6550), .ZN(n6544) );
  OAI211_X1 U7538 ( .C1(n6604), .C2(n6614), .A(n6545), .B(n6544), .ZN(U3074)
         );
  AOI22_X1 U7539 ( .A1(n6549), .A2(n6548), .B1(n6547), .B2(n6546), .ZN(n6554)
         );
  AOI22_X1 U7540 ( .A1(n6552), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6551), 
        .B2(n6550), .ZN(n6553) );
  OAI211_X1 U7541 ( .C1(n6555), .C2(n6614), .A(n6554), .B(n6553), .ZN(U3075)
         );
  INV_X1 U7542 ( .A(n6556), .ZN(n6558) );
  INV_X1 U7543 ( .A(n6615), .ZN(n6557) );
  AOI21_X1 U7544 ( .B1(n6558), .B2(n6653), .A(n6557), .ZN(n6563) );
  NOR2_X1 U7545 ( .A1(n6563), .A2(n6559), .ZN(n6560) );
  AOI21_X1 U7546 ( .B1(n6568), .B2(STATE2_REG_2__SCAN_IN), .A(n6560), .ZN(
        n6624) );
  OAI22_X1 U7547 ( .A1(n6626), .A2(n6615), .B1(n6614), .B2(n6632), .ZN(n6561)
         );
  INV_X1 U7548 ( .A(n6561), .ZN(n6571) );
  INV_X1 U7549 ( .A(n6562), .ZN(n6564) );
  NAND3_X1 U7550 ( .A1(n6564), .A2(n6567), .A3(n6563), .ZN(n6566) );
  OAI211_X1 U7551 ( .C1(n6568), .C2(n6567), .A(n6566), .B(n6565), .ZN(n6620)
         );
  AOI22_X1 U7552 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6620), .B1(n6569), 
        .B2(n6618), .ZN(n6570) );
  OAI211_X1 U7553 ( .C1(n6624), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3076)
         );
  OAI22_X1 U7554 ( .A1(n6574), .A2(n6615), .B1(n6614), .B2(n6573), .ZN(n6575)
         );
  INV_X1 U7555 ( .A(n6575), .ZN(n6578) );
  AOI22_X1 U7556 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6620), .B1(n6576), 
        .B2(n6618), .ZN(n6577) );
  OAI211_X1 U7557 ( .C1(n6624), .C2(n6579), .A(n6578), .B(n6577), .ZN(U3077)
         );
  OAI22_X1 U7558 ( .A1(n6581), .A2(n6615), .B1(n6605), .B2(n6580), .ZN(n6582)
         );
  INV_X1 U7559 ( .A(n6582), .ZN(n6585) );
  INV_X1 U7560 ( .A(n6614), .ZN(n6608) );
  AOI22_X1 U7561 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6620), .B1(n6583), 
        .B2(n6608), .ZN(n6584) );
  OAI211_X1 U7562 ( .C1(n6624), .C2(n6586), .A(n6585), .B(n6584), .ZN(U3078)
         );
  OAI22_X1 U7563 ( .A1(n6634), .A2(n6615), .B1(n6614), .B2(n6643), .ZN(n6587)
         );
  INV_X1 U7564 ( .A(n6587), .ZN(n6590) );
  AOI22_X1 U7565 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6620), .B1(n6588), 
        .B2(n6618), .ZN(n6589) );
  OAI211_X1 U7566 ( .C1(n6624), .C2(n6591), .A(n6590), .B(n6589), .ZN(U3079)
         );
  OAI22_X1 U7567 ( .A1(n7203), .A2(n6615), .B1(n6605), .B2(n6592), .ZN(n6593)
         );
  INV_X1 U7568 ( .A(n6593), .ZN(n6596) );
  AOI22_X1 U7569 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6620), .B1(n6594), 
        .B2(n6608), .ZN(n6595) );
  OAI211_X1 U7570 ( .C1(n6624), .C2(n7200), .A(n6596), .B(n6595), .ZN(U3080)
         );
  OAI22_X1 U7571 ( .A1(n6598), .A2(n6615), .B1(n6605), .B2(n6597), .ZN(n6599)
         );
  INV_X1 U7572 ( .A(n6599), .ZN(n6602) );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6620), .B1(n6600), 
        .B2(n6608), .ZN(n6601) );
  OAI211_X1 U7574 ( .C1(n6624), .C2(n6603), .A(n6602), .B(n6601), .ZN(U3081)
         );
  OAI22_X1 U7575 ( .A1(n6606), .A2(n6615), .B1(n6605), .B2(n6604), .ZN(n6607)
         );
  INV_X1 U7576 ( .A(n6607), .ZN(n6611) );
  AOI22_X1 U7577 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6620), .B1(n6609), 
        .B2(n6608), .ZN(n6610) );
  OAI211_X1 U7578 ( .C1(n6624), .C2(n6612), .A(n6611), .B(n6610), .ZN(U3082)
         );
  OAI22_X1 U7579 ( .A1(n6616), .A2(n6615), .B1(n6614), .B2(n6613), .ZN(n6617)
         );
  INV_X1 U7580 ( .A(n6617), .ZN(n6622) );
  AOI22_X1 U7581 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6620), .B1(n6619), 
        .B2(n6618), .ZN(n6621) );
  OAI211_X1 U7582 ( .C1(n6624), .C2(n6623), .A(n6622), .B(n6621), .ZN(U3083)
         );
  INV_X1 U7583 ( .A(n6625), .ZN(n6633) );
  OAI22_X1 U7584 ( .A1(n7210), .A2(n6627), .B1(n6626), .B2(n6633), .ZN(n6628)
         );
  INV_X1 U7585 ( .A(n6628), .ZN(n6631) );
  AOI22_X1 U7586 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6639), .B1(n6629), 
        .B2(n6637), .ZN(n6630) );
  OAI211_X1 U7587 ( .C1(n6632), .C2(n6642), .A(n6631), .B(n6630), .ZN(U3108)
         );
  OAI22_X1 U7588 ( .A1(n7210), .A2(n6635), .B1(n6634), .B2(n6633), .ZN(n6636)
         );
  INV_X1 U7589 ( .A(n6636), .ZN(n6641) );
  AOI22_X1 U7590 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6639), .B1(n6638), 
        .B2(n6637), .ZN(n6640) );
  OAI211_X1 U7591 ( .C1(n6643), .C2(n6642), .A(n6641), .B(n6640), .ZN(U3111)
         );
  OAI21_X1 U7592 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6644), 
        .ZN(n6645) );
  NAND4_X1 U7593 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6649)
         );
  NOR2_X1 U7594 ( .A1(n6650), .A2(n6649), .ZN(n6672) );
  NAND2_X1 U7595 ( .A1(n6670), .A2(n6669), .ZN(n6667) );
  AOI22_X1 U7596 ( .A1(n6653), .A2(n6652), .B1(n6651), .B2(n3308), .ZN(n6777)
         );
  NAND2_X1 U7597 ( .A1(n6654), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6783) );
  NAND3_X1 U7598 ( .A1(n6777), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6783), .ZN(n6657) );
  OAI211_X1 U7599 ( .C1(n6658), .C2(n6657), .A(n6656), .B(n6655), .ZN(n6660)
         );
  NAND2_X1 U7600 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  NAND2_X1 U7601 ( .A1(n6660), .A2(n6659), .ZN(n6663) );
  INV_X1 U7602 ( .A(n6663), .ZN(n6661) );
  NOR2_X1 U7603 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6661), .ZN(n6664)
         );
  OAI22_X1 U7604 ( .A1(n6665), .A2(n6664), .B1(n6663), .B2(n6662), .ZN(n6666)
         );
  NAND2_X1 U7605 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  OAI211_X1 U7606 ( .C1(n6670), .C2(n6669), .A(n6668), .B(n7080), .ZN(n6671)
         );
  AND2_X1 U7607 ( .A1(n6672), .A2(n6671), .ZN(n6683) );
  NAND2_X1 U7608 ( .A1(n6683), .A2(n6673), .ZN(n6675) );
  NAND2_X1 U7609 ( .A1(READY_N), .A2(n6796), .ZN(n6674) );
  NAND2_X1 U7610 ( .A1(n6675), .A2(n6674), .ZN(n6679) );
  OR2_X1 U7611 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  OAI21_X1 U7612 ( .B1(n6694), .B2(n6771), .A(n6685), .ZN(n6687) );
  AOI21_X1 U7613 ( .B1(READY_N), .B2(n6680), .A(n6766), .ZN(n6688) );
  OAI211_X1 U7614 ( .C1(n6683), .C2(n6682), .A(n6688), .B(n6681), .ZN(n6684)
         );
  AOI21_X1 U7615 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6799), .A(n6684), .ZN(
        n6686) );
  OAI22_X1 U7616 ( .A1(n6766), .A2(n6687), .B1(n6686), .B2(n6685), .ZN(U3148)
         );
  NOR3_X1 U7617 ( .A1(n6697), .A2(n6688), .A3(n6776), .ZN(n6692) );
  AOI221_X1 U7618 ( .B1(READY_N), .B2(n6690), .C1(n6689), .C2(n6690), .A(n6766), .ZN(n6691) );
  OR3_X1 U7619 ( .A1(n6693), .A2(n6692), .A3(n6691), .ZN(U3149) );
  OAI211_X1 U7620 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6795), .A(n6767), .B(
        n6694), .ZN(n6696) );
  OAI21_X1 U7621 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(U3150) );
  AND2_X1 U7622 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6762), .ZN(U3151) );
  AND2_X1 U7623 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6762), .ZN(U3152) );
  AND2_X1 U7624 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6762), .ZN(U3153) );
  AND2_X1 U7625 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6762), .ZN(U3154) );
  AND2_X1 U7626 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6762), .ZN(U3155) );
  AND2_X1 U7627 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6762), .ZN(U3156) );
  AND2_X1 U7628 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6762), .ZN(U3157) );
  AND2_X1 U7629 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6762), .ZN(U3158) );
  AND2_X1 U7630 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6762), .ZN(U3159) );
  INV_X1 U7631 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7050) );
  NOR2_X1 U7632 ( .A1(n6765), .A2(n7050), .ZN(U3160) );
  AND2_X1 U7633 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6762), .ZN(U3161) );
  INV_X1 U7634 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U7635 ( .A1(n6765), .A2(n6918), .ZN(U3162) );
  INV_X1 U7636 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U7637 ( .A1(n6765), .A2(n6983), .ZN(U3163) );
  AND2_X1 U7638 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6762), .ZN(U3164) );
  AND2_X1 U7639 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6762), .ZN(U3165) );
  AND2_X1 U7640 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6762), .ZN(U3166) );
  INV_X1 U7641 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7141) );
  NOR2_X1 U7642 ( .A1(n6765), .A2(n7141), .ZN(U3167) );
  AND2_X1 U7643 ( .A1(n6762), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7644 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6762), .ZN(U3169) );
  AND2_X1 U7645 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6762), .ZN(U3170) );
  INV_X1 U7646 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7093) );
  NOR2_X1 U7647 ( .A1(n6765), .A2(n7093), .ZN(U3171) );
  INV_X1 U7648 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7125) );
  NOR2_X1 U7649 ( .A1(n6765), .A2(n7125), .ZN(U3172) );
  AND2_X1 U7650 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6762), .ZN(U3173) );
  AND2_X1 U7651 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6762), .ZN(U3174) );
  AND2_X1 U7652 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6762), .ZN(U3175) );
  INV_X1 U7653 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6955) );
  NOR2_X1 U7654 ( .A1(n6765), .A2(n6955), .ZN(U3176) );
  INV_X1 U7655 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7139) );
  NOR2_X1 U7656 ( .A1(n6765), .A2(n7139), .ZN(U3177) );
  AND2_X1 U7657 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6762), .ZN(U3178) );
  AND2_X1 U7658 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6762), .ZN(U3179) );
  AND2_X1 U7659 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6762), .ZN(U3180) );
  NOR2_X1 U7660 ( .A1(n6703), .A2(n6713), .ZN(n6704) );
  AOI22_X1 U7661 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6712) );
  AND2_X1 U7662 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6700) );
  INV_X1 U7663 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7144) );
  INV_X1 U7664 ( .A(NA_N), .ZN(n6705) );
  AOI221_X1 U7665 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6705), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6709) );
  AOI221_X1 U7666 ( .B1(n6700), .B2(n6760), .C1(n7144), .C2(n6760), .A(n6709), 
        .ZN(n6698) );
  OAI21_X1 U7667 ( .B1(n6704), .B2(n6712), .A(n6698), .ZN(U3181) );
  NOR2_X1 U7668 ( .A1(n6707), .A2(n7144), .ZN(n6706) );
  NAND2_X1 U7669 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6699) );
  OAI21_X1 U7670 ( .B1(n6706), .B2(n6700), .A(n6699), .ZN(n6701) );
  OAI211_X1 U7671 ( .C1(n6703), .C2(n6795), .A(n6702), .B(n6701), .ZN(U3182)
         );
  AOI21_X1 U7672 ( .B1(n6706), .B2(n6705), .A(n6704), .ZN(n6711) );
  AOI221_X1 U7673 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6795), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6708) );
  AOI221_X1 U7674 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6708), .C2(HOLD), .A(n6707), .ZN(n6710) );
  OAI22_X1 U7675 ( .A1(n6712), .A2(n6711), .B1(n6710), .B2(n6709), .ZN(U3183)
         );
  NAND2_X1 U7676 ( .A1(n6804), .A2(n6713), .ZN(n6758) );
  INV_X1 U7677 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U7678 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6804), .ZN(n6755) );
  OAI222_X1 U7679 ( .A1(n6758), .A2(n6715), .B1(n7094), .B2(n6804), .C1(n6998), 
        .C2(n6755), .ZN(U3184) );
  INV_X1 U7680 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6995) );
  OAI222_X1 U7681 ( .A1(n6755), .A2(n6715), .B1(n6995), .B2(n6804), .C1(n6714), 
        .C2(n6758), .ZN(U3185) );
  INV_X1 U7682 ( .A(n6755), .ZN(n6756) );
  AOI22_X1 U7683 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6792), .ZN(n6716) );
  OAI21_X1 U7684 ( .B1(n6718), .B2(n6758), .A(n6716), .ZN(U3186) );
  INV_X1 U7685 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6971) );
  OAI222_X1 U7686 ( .A1(n6755), .A2(n6718), .B1(n6971), .B2(n6804), .C1(n6717), 
        .C2(n6758), .ZN(U3187) );
  AOI22_X1 U7687 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6792), .ZN(n6719) );
  OAI21_X1 U7688 ( .B1(n6720), .B2(n6758), .A(n6719), .ZN(U3188) );
  AOI22_X1 U7689 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6792), .ZN(n6721) );
  OAI21_X1 U7690 ( .B1(n6722), .B2(n6758), .A(n6721), .ZN(U3189) );
  INV_X1 U7691 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6947) );
  INV_X1 U7692 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6723) );
  OAI222_X1 U7693 ( .A1(n6755), .A2(n6722), .B1(n6947), .B2(n6804), .C1(n6723), 
        .C2(n6758), .ZN(U3190) );
  INV_X1 U7694 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6724) );
  OAI222_X1 U7695 ( .A1(n6758), .A2(n6725), .B1(n6724), .B2(n6804), .C1(n6723), 
        .C2(n6755), .ZN(U3191) );
  INV_X1 U7696 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6989) );
  OAI222_X1 U7697 ( .A1(n6755), .A2(n6725), .B1(n6989), .B2(n6804), .C1(n6196), 
        .C2(n6758), .ZN(U3192) );
  AOI22_X1 U7698 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6792), .ZN(n6726) );
  OAI21_X1 U7699 ( .B1(n6728), .B2(n6758), .A(n6726), .ZN(U3193) );
  INV_X1 U7700 ( .A(n6758), .ZN(n6753) );
  AOI22_X1 U7701 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6760), .ZN(n6727) );
  OAI21_X1 U7702 ( .B1(n6728), .B2(n6755), .A(n6727), .ZN(U3194) );
  INV_X1 U7703 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7056) );
  OAI222_X1 U7704 ( .A1(n6755), .A2(n6729), .B1(n7056), .B2(n6804), .C1(n6906), 
        .C2(n6758), .ZN(U3195) );
  AOI22_X1 U7705 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6792), .ZN(n6730) );
  OAI21_X1 U7706 ( .B1(n6732), .B2(n6758), .A(n6730), .ZN(U3196) );
  AOI22_X1 U7707 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6760), .ZN(n6731) );
  OAI21_X1 U7708 ( .B1(n6732), .B2(n6755), .A(n6731), .ZN(U3197) );
  AOI22_X1 U7709 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6760), .ZN(n6733) );
  OAI21_X1 U7710 ( .B1(n5750), .B2(n6758), .A(n6733), .ZN(U3198) );
  AOI22_X1 U7711 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6792), .ZN(n6734) );
  OAI21_X1 U7712 ( .B1(n5750), .B2(n6755), .A(n6734), .ZN(U3199) );
  AOI22_X1 U7713 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6760), .ZN(n6735) );
  OAI21_X1 U7714 ( .B1(n6738), .B2(n6758), .A(n6735), .ZN(U3200) );
  INV_X1 U7715 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6737) );
  OAI222_X1 U7716 ( .A1(n6755), .A2(n6738), .B1(n6737), .B2(n6804), .C1(n6736), 
        .C2(n6758), .ZN(U3201) );
  AOI22_X1 U7717 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6760), .ZN(n6739) );
  OAI21_X1 U7718 ( .B1(n5735), .B2(n6758), .A(n6739), .ZN(U3202) );
  AOI22_X1 U7719 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6760), .ZN(n6740) );
  OAI21_X1 U7720 ( .B1(n7075), .B2(n6758), .A(n6740), .ZN(U3203) );
  INV_X1 U7721 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6741) );
  OAI222_X1 U7722 ( .A1(n6755), .A2(n7075), .B1(n6741), .B2(n6804), .C1(n6743), 
        .C2(n6758), .ZN(U3204) );
  AOI22_X1 U7723 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6760), .ZN(n6742) );
  OAI21_X1 U7724 ( .B1(n6743), .B2(n6755), .A(n6742), .ZN(U3205) );
  INV_X1 U7725 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6744) );
  INV_X1 U7726 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6986) );
  OAI222_X1 U7727 ( .A1(n6755), .A2(n6744), .B1(n6986), .B2(n6804), .C1(n6746), 
        .C2(n6758), .ZN(U3206) );
  AOI22_X1 U7728 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6760), .ZN(n6745) );
  OAI21_X1 U7729 ( .B1(n6746), .B2(n6755), .A(n6745), .ZN(U3207) );
  AOI222_X1 U7730 ( .A1(n6756), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6760), .C1(REIP_REG_26__SCAN_IN), .C2(
        n6753), .ZN(n6747) );
  INV_X1 U7731 ( .A(n6747), .ZN(U3208) );
  AOI22_X1 U7732 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6760), .ZN(n6748) );
  OAI21_X1 U7733 ( .B1(n6749), .B2(n6758), .A(n6748), .ZN(U3209) );
  AOI22_X1 U7734 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6792), .ZN(n6750) );
  OAI21_X1 U7735 ( .B1(n6752), .B2(n6758), .A(n6750), .ZN(U3210) );
  AOI22_X1 U7736 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6760), .ZN(n6751) );
  OAI21_X1 U7737 ( .B1(n6752), .B2(n6755), .A(n6751), .ZN(U3211) );
  AOI22_X1 U7738 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6753), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6760), .ZN(n6754) );
  OAI21_X1 U7739 ( .B1(n6934), .B2(n6755), .A(n6754), .ZN(U3212) );
  AOI22_X1 U7740 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6756), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6760), .ZN(n6757) );
  OAI21_X1 U7741 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(U3213) );
  MUX2_X1 U7742 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6804), .Z(U3445) );
  MUX2_X1 U7743 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6804), .Z(U3446) );
  MUX2_X1 U7744 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6804), .Z(U3447) );
  INV_X1 U7745 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6789) );
  INV_X1 U7746 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6999) );
  AOI22_X1 U7747 ( .A1(n6804), .A2(n6789), .B1(n6999), .B2(n6760), .ZN(U3448)
         );
  INV_X1 U7748 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7060) );
  INV_X1 U7749 ( .A(n6763), .ZN(n6761) );
  AOI21_X1 U7750 ( .B1(n7060), .B2(n6762), .A(n6761), .ZN(U3451) );
  OAI21_X1 U7751 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(U3452) );
  INV_X1 U7752 ( .A(n6766), .ZN(n6768) );
  OAI221_X1 U7753 ( .B1(n6769), .B2(STATE2_REG_0__SCAN_IN), .C1(n6769), .C2(
        n6768), .A(n6767), .ZN(U3453) );
  INV_X1 U7754 ( .A(n6770), .ZN(n6773) );
  OAI22_X1 U7755 ( .A1(n6773), .A2(n6782), .B1(n6772), .B2(n6771), .ZN(n6775)
         );
  MUX2_X1 U7756 ( .A(n6775), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6774), 
        .Z(U3456) );
  OAI22_X1 U7757 ( .A1(n6777), .A2(n6782), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6776), .ZN(n6779) );
  OAI22_X1 U7758 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6780), .B1(n6779), .B2(n6778), .ZN(n6781) );
  OAI21_X1 U7759 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(U3461) );
  AOI21_X1 U7760 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7761 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6784), .B2(n6998), .ZN(n6787) );
  INV_X1 U7762 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6786) );
  AOI22_X1 U7763 ( .A1(n6790), .A2(n6787), .B1(n6786), .B2(n6785), .ZN(U3468)
         );
  OAI21_X1 U7764 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6790), .ZN(n6788) );
  OAI21_X1 U7765 ( .B1(n6790), .B2(n6789), .A(n6788), .ZN(U3469) );
  NAND2_X1 U7766 ( .A1(n6792), .A2(W_R_N_REG_SCAN_IN), .ZN(n6791) );
  OAI21_X1 U7767 ( .B1(n6792), .B2(READREQUEST_REG_SCAN_IN), .A(n6791), .ZN(
        U3470) );
  AOI211_X1 U7768 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n6793), .ZN(n6803)
         );
  OAI211_X1 U7769 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6798), .A(n6797), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6800) );
  AOI21_X1 U7770 ( .B1(n6800), .B2(STATE2_REG_0__SCAN_IN), .A(n6799), .ZN(
        n6802) );
  NAND2_X1 U7771 ( .A1(n6803), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6801) );
  OAI21_X1 U7772 ( .B1(n6803), .B2(n6802), .A(n6801), .ZN(U3472) );
  MUX2_X1 U7773 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6804), .Z(U3473) );
  OAI22_X1 U7774 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput122), .B1(
        keyinput105), .B2(DATAO_REG_22__SCAN_IN), .ZN(n6805) );
  AOI221_X1 U7775 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput122), .C1(
        DATAO_REG_22__SCAN_IN), .C2(keyinput105), .A(n6805), .ZN(n6812) );
  OAI22_X1 U7776 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(keyinput1), .B1(
        keyinput111), .B2(UWORD_REG_2__SCAN_IN), .ZN(n6806) );
  AOI221_X1 U7777 ( .B1(INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput1), .C1(
        UWORD_REG_2__SCAN_IN), .C2(keyinput111), .A(n6806), .ZN(n6811) );
  OAI22_X1 U7778 ( .A1(UWORD_REG_1__SCAN_IN), .A2(keyinput66), .B1(keyinput88), 
        .B2(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6807) );
  AOI221_X1 U7779 ( .B1(UWORD_REG_1__SCAN_IN), .B2(keyinput66), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput88), .A(n6807), .ZN(n6810) );
  OAI22_X1 U7780 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(keyinput94), .B1(
        EAX_REG_0__SCAN_IN), .B2(keyinput113), .ZN(n6808) );
  AOI221_X1 U7781 ( .B1(INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput94), .C1(
        keyinput113), .C2(EAX_REG_0__SCAN_IN), .A(n6808), .ZN(n6809) );
  NAND4_X1 U7782 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6840)
         );
  OAI22_X1 U7783 ( .A1(ADDRESS_REG_20__SCAN_IN), .A2(keyinput95), .B1(
        keyinput43), .B2(ADDRESS_REG_8__SCAN_IN), .ZN(n6813) );
  AOI221_X1 U7784 ( .B1(ADDRESS_REG_20__SCAN_IN), .B2(keyinput95), .C1(
        ADDRESS_REG_8__SCAN_IN), .C2(keyinput43), .A(n6813), .ZN(n6820) );
  OAI22_X1 U7785 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput123), 
        .B1(EAX_REG_22__SCAN_IN), .B2(keyinput6), .ZN(n6814) );
  AOI221_X1 U7786 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput123), 
        .C1(keyinput6), .C2(EAX_REG_22__SCAN_IN), .A(n6814), .ZN(n6819) );
  OAI22_X1 U7787 ( .A1(EAX_REG_25__SCAN_IN), .A2(keyinput106), .B1(keyinput108), .B2(DATAI_23_), .ZN(n6815) );
  AOI221_X1 U7788 ( .B1(EAX_REG_25__SCAN_IN), .B2(keyinput106), .C1(DATAI_23_), 
        .C2(keyinput108), .A(n6815), .ZN(n6818) );
  OAI22_X1 U7789 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput56), .B1(
        keyinput78), .B2(LWORD_REG_11__SCAN_IN), .ZN(n6816) );
  AOI221_X1 U7790 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput56), .C1(
        LWORD_REG_11__SCAN_IN), .C2(keyinput78), .A(n6816), .ZN(n6817) );
  NAND4_X1 U7791 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6839)
         );
  OAI22_X1 U7792 ( .A1(EBX_REG_18__SCAN_IN), .A2(keyinput101), .B1(
        REIP_REG_4__SCAN_IN), .B2(keyinput87), .ZN(n6821) );
  AOI221_X1 U7793 ( .B1(EBX_REG_18__SCAN_IN), .B2(keyinput101), .C1(keyinput87), .C2(REIP_REG_4__SCAN_IN), .A(n6821), .ZN(n6828) );
  OAI22_X1 U7794 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput76), .B1(
        keyinput102), .B2(DATAO_REG_11__SCAN_IN), .ZN(n6822) );
  AOI221_X1 U7795 ( .B1(INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput76), .C1(
        DATAO_REG_11__SCAN_IN), .C2(keyinput102), .A(n6822), .ZN(n6827) );
  OAI22_X1 U7796 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(keyinput80), .B1(
        keyinput4), .B2(DATAO_REG_6__SCAN_IN), .ZN(n6823) );
  AOI221_X1 U7797 ( .B1(INSTQUEUE_REG_15__4__SCAN_IN), .B2(keyinput80), .C1(
        DATAO_REG_6__SCAN_IN), .C2(keyinput4), .A(n6823), .ZN(n6826) );
  OAI22_X1 U7798 ( .A1(REIP_REG_14__SCAN_IN), .A2(keyinput82), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(keyinput0), .ZN(n6824) );
  AOI221_X1 U7799 ( .B1(REIP_REG_14__SCAN_IN), .B2(keyinput82), .C1(keyinput0), 
        .C2(ADDRESS_REG_3__SCAN_IN), .A(n6824), .ZN(n6825) );
  NAND4_X1 U7800 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n6825), .ZN(n6838)
         );
  OAI22_X1 U7801 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(keyinput54), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput31), .ZN(n6829) );
  AOI221_X1 U7802 ( .B1(INSTQUEUE_REG_12__2__SCAN_IN), .B2(keyinput54), .C1(
        keyinput31), .C2(BE_N_REG_0__SCAN_IN), .A(n6829), .ZN(n6836) );
  OAI22_X1 U7803 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(keyinput107), .B1(
        UWORD_REG_8__SCAN_IN), .B2(keyinput71), .ZN(n6830) );
  AOI221_X1 U7804 ( .B1(INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput107), .C1(
        keyinput71), .C2(UWORD_REG_8__SCAN_IN), .A(n6830), .ZN(n6835) );
  OAI22_X1 U7805 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(keyinput68), .B1(
        keyinput50), .B2(UWORD_REG_9__SCAN_IN), .ZN(n6831) );
  AOI221_X1 U7806 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput68), .C1(
        UWORD_REG_9__SCAN_IN), .C2(keyinput50), .A(n6831), .ZN(n6834) );
  OAI22_X1 U7807 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput64), .B1(keyinput100), .B2(DATAO_REG_29__SCAN_IN), .ZN(n6832) );
  AOI221_X1 U7808 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput64), .C1(
        DATAO_REG_29__SCAN_IN), .C2(keyinput100), .A(n6832), .ZN(n6833) );
  NAND4_X1 U7809 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6837)
         );
  NOR4_X1 U7810 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n7198)
         );
  AOI22_X1 U7811 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(keyinput207), .B1(
        INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput164), .ZN(n6841) );
  OAI221_X1 U7812 ( .B1(INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput207), .C1(
        INSTQUEUE_REG_15__6__SCAN_IN), .C2(keyinput164), .A(n6841), .ZN(n6848)
         );
  AOI22_X1 U7813 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(keyinput131), .B1(
        INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput158), .ZN(n6842) );
  OAI221_X1 U7814 ( .B1(INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput131), .C1(
        INSTQUEUE_REG_10__4__SCAN_IN), .C2(keyinput158), .A(n6842), .ZN(n6847)
         );
  AOI22_X1 U7815 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(keyinput235), .B1(
        INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput224), .ZN(n6843) );
  OAI221_X1 U7816 ( .B1(INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput235), .C1(
        INSTQUEUE_REG_3__0__SCAN_IN), .C2(keyinput224), .A(n6843), .ZN(n6846)
         );
  AOI22_X1 U7817 ( .A1(EBX_REG_19__SCAN_IN), .A2(keyinput212), .B1(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput174), .ZN(n6844) );
  OAI221_X1 U7818 ( .B1(EBX_REG_19__SCAN_IN), .B2(keyinput212), .C1(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(keyinput174), .A(n6844), .ZN(
        n6845) );
  NOR4_X1 U7819 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6876)
         );
  AOI22_X1 U7820 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(keyinput196), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput145), .ZN(n6849) );
  OAI221_X1 U7821 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput196), 
        .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput145), .A(n6849), 
        .ZN(n6856) );
  AOI22_X1 U7822 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput181), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(keyinput223), .ZN(n6850) );
  OAI221_X1 U7823 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput181), .C1(
        ADDRESS_REG_20__SCAN_IN), .C2(keyinput223), .A(n6850), .ZN(n6855) );
  AOI22_X1 U7824 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput250), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput180), .ZN(n6851) );
  OAI221_X1 U7825 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput250), .C1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput180), .A(n6851), .ZN(
        n6854) );
  AOI22_X1 U7826 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput136), .B1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput246), .ZN(n6852) );
  OAI221_X1 U7827 ( .B1(INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput136), .C1(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(keyinput246), .A(n6852), .ZN(
        n6853) );
  NOR4_X1 U7828 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6875)
         );
  AOI22_X1 U7829 ( .A1(EAX_REG_18__SCAN_IN), .A2(keyinput165), .B1(
        INSTQUEUE_REG_14__5__SCAN_IN), .B2(keyinput153), .ZN(n6857) );
  OAI221_X1 U7830 ( .B1(EAX_REG_18__SCAN_IN), .B2(keyinput165), .C1(
        INSTQUEUE_REG_14__5__SCAN_IN), .C2(keyinput153), .A(n6857), .ZN(n6864)
         );
  AOI22_X1 U7831 ( .A1(LWORD_REG_2__SCAN_IN), .A2(keyinput162), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput169), .ZN(n6858) );
  OAI221_X1 U7832 ( .B1(LWORD_REG_2__SCAN_IN), .B2(keyinput162), .C1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput169), .A(n6858), .ZN(
        n6863) );
  AOI22_X1 U7833 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput146), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput225), .ZN(n6859) );
  OAI221_X1 U7834 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput146), .C1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput225), .A(n6859), .ZN(
        n6862) );
  AOI22_X1 U7835 ( .A1(DATAO_REG_22__SCAN_IN), .A2(keyinput233), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput133), .ZN(n6860) );
  OAI221_X1 U7836 ( .B1(DATAO_REG_22__SCAN_IN), .B2(keyinput233), .C1(
        INSTQUEUE_REG_8__6__SCAN_IN), .C2(keyinput133), .A(n6860), .ZN(n6861)
         );
  NOR4_X1 U7837 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n6874)
         );
  AOI22_X1 U7838 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput219), .B1(
        DATAI_31_), .B2(keyinput209), .ZN(n6865) );
  OAI221_X1 U7839 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput219), .C1(
        DATAI_31_), .C2(keyinput209), .A(n6865), .ZN(n6872) );
  AOI22_X1 U7840 ( .A1(REIP_REG_14__SCAN_IN), .A2(keyinput210), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput148), .ZN(n6866) );
  OAI221_X1 U7841 ( .B1(REIP_REG_14__SCAN_IN), .B2(keyinput210), .C1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput148), .A(n6866), .ZN(
        n6871) );
  AOI22_X1 U7842 ( .A1(DATAO_REG_29__SCAN_IN), .A2(keyinput228), .B1(
        INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput141), .ZN(n6867) );
  OAI221_X1 U7843 ( .B1(DATAO_REG_29__SCAN_IN), .B2(keyinput228), .C1(
        INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput141), .A(n6867), .ZN(n6870)
         );
  AOI22_X1 U7844 ( .A1(EAX_REG_3__SCAN_IN), .A2(keyinput214), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput154), .ZN(n6868) );
  OAI221_X1 U7845 ( .B1(EAX_REG_3__SCAN_IN), .B2(keyinput214), .C1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput154), .A(n6868), .ZN(n6869) );
  NOR4_X1 U7846 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6873)
         );
  NAND4_X1 U7847 ( .A1(n6876), .A2(n6875), .A3(n6874), .A4(n6873), .ZN(n7026)
         );
  AOI22_X1 U7848 ( .A1(DATAI_5_), .A2(keyinput144), .B1(
        INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput254), .ZN(n6877) );
  OAI221_X1 U7849 ( .B1(DATAI_5_), .B2(keyinput144), .C1(
        INSTQUEUE_REG_0__3__SCAN_IN), .C2(keyinput254), .A(n6877), .ZN(n6884)
         );
  AOI22_X1 U7850 ( .A1(LWORD_REG_9__SCAN_IN), .A2(keyinput193), .B1(DATAI_28_), 
        .B2(keyinput253), .ZN(n6878) );
  OAI221_X1 U7851 ( .B1(LWORD_REG_9__SCAN_IN), .B2(keyinput193), .C1(DATAI_28_), .C2(keyinput253), .A(n6878), .ZN(n6883) );
  AOI22_X1 U7852 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput163), .B1(
        INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput177), .ZN(n6879) );
  OAI221_X1 U7853 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput163), .C1(
        INSTQUEUE_REG_0__2__SCAN_IN), .C2(keyinput177), .A(n6879), .ZN(n6882)
         );
  AOI22_X1 U7854 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput230), .B1(
        INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput237), .ZN(n6880) );
  OAI221_X1 U7855 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput230), .C1(
        INSTQUEUE_REG_3__2__SCAN_IN), .C2(keyinput237), .A(n6880), .ZN(n6881)
         );
  NOR4_X1 U7856 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6914)
         );
  AOI22_X1 U7857 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput192), .B1(
        EAX_REG_2__SCAN_IN), .B2(keyinput143), .ZN(n6885) );
  OAI221_X1 U7858 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput192), .C1(
        EAX_REG_2__SCAN_IN), .C2(keyinput143), .A(n6885), .ZN(n6892) );
  AOI22_X1 U7859 ( .A1(DATAO_REG_23__SCAN_IN), .A2(keyinput247), .B1(DATAI_10_), .B2(keyinput138), .ZN(n6886) );
  OAI221_X1 U7860 ( .B1(DATAO_REG_23__SCAN_IN), .B2(keyinput247), .C1(
        DATAI_10_), .C2(keyinput138), .A(n6886), .ZN(n6891) );
  AOI22_X1 U7861 ( .A1(UWORD_REG_7__SCAN_IN), .A2(keyinput149), .B1(
        REIP_REG_8__SCAN_IN), .B2(keyinput195), .ZN(n6887) );
  OAI221_X1 U7862 ( .B1(UWORD_REG_7__SCAN_IN), .B2(keyinput149), .C1(
        REIP_REG_8__SCAN_IN), .C2(keyinput195), .A(n6887), .ZN(n6890) );
  AOI22_X1 U7863 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(keyinput172), .B1(
        EAX_REG_15__SCAN_IN), .B2(keyinput166), .ZN(n6888) );
  OAI221_X1 U7864 ( .B1(DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput172), .C1(
        EAX_REG_15__SCAN_IN), .C2(keyinput166), .A(n6888), .ZN(n6889) );
  NOR4_X1 U7865 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6913)
         );
  AOI22_X1 U7866 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput242), .B1(
        INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput204), .ZN(n6893) );
  OAI221_X1 U7867 ( .B1(DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput242), .C1(
        INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput204), .A(n6893), .ZN(n6900)
         );
  AOI22_X1 U7868 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput140), .B1(
        INSTQUEUE_REG_6__2__SCAN_IN), .B2(keyinput168), .ZN(n6894) );
  OAI221_X1 U7869 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput140), .C1(
        INSTQUEUE_REG_6__2__SCAN_IN), .C2(keyinput168), .A(n6894), .ZN(n6899)
         );
  AOI22_X1 U7870 ( .A1(REIP_REG_4__SCAN_IN), .A2(keyinput215), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput200), .ZN(n6895) );
  OAI221_X1 U7871 ( .B1(REIP_REG_4__SCAN_IN), .B2(keyinput215), .C1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput200), .A(n6895), .ZN(n6898) );
  AOI22_X1 U7872 ( .A1(EBX_REG_18__SCAN_IN), .A2(keyinput229), .B1(
        INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput135), .ZN(n6896) );
  OAI221_X1 U7873 ( .B1(EBX_REG_18__SCAN_IN), .B2(keyinput229), .C1(
        INSTQUEUE_REG_6__4__SCAN_IN), .C2(keyinput135), .A(n6896), .ZN(n6897)
         );
  NOR4_X1 U7874 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6912)
         );
  AOI22_X1 U7875 ( .A1(EAX_REG_20__SCAN_IN), .A2(keyinput186), .B1(
        EBX_REG_15__SCAN_IN), .B2(keyinput226), .ZN(n6901) );
  OAI221_X1 U7876 ( .B1(EAX_REG_20__SCAN_IN), .B2(keyinput186), .C1(
        EBX_REG_15__SCAN_IN), .C2(keyinput226), .A(n6901), .ZN(n6910) );
  AOI22_X1 U7877 ( .A1(keyinput176), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .B1(n7129), .B2(keyinput221), .ZN(n6902) );
  OAI221_X1 U7878 ( .B1(keyinput176), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .C1(n7129), .C2(keyinput221), .A(n6902), .ZN(n6909) );
  INV_X1 U7879 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7880 ( .A1(n7115), .A2(keyinput142), .B1(keyinput178), .B2(n6904), 
        .ZN(n6903) );
  OAI221_X1 U7881 ( .B1(n7115), .B2(keyinput142), .C1(n6904), .C2(keyinput178), 
        .A(n6903), .ZN(n6908) );
  AOI22_X1 U7882 ( .A1(n7031), .A2(keyinput213), .B1(n6906), .B2(keyinput183), 
        .ZN(n6905) );
  OAI221_X1 U7883 ( .B1(n7031), .B2(keyinput213), .C1(n6906), .C2(keyinput183), 
        .A(n6905), .ZN(n6907) );
  NOR4_X1 U7884 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6911)
         );
  NAND4_X1 U7885 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n7025)
         );
  INV_X1 U7886 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6916) );
  AOI22_X1 U7887 ( .A1(n6916), .A2(keyinput239), .B1(n7028), .B2(keyinput201), 
        .ZN(n6915) );
  OAI221_X1 U7888 ( .B1(n6916), .B2(keyinput239), .C1(n7028), .C2(keyinput201), 
        .A(n6915), .ZN(n6927) );
  INV_X1 U7889 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U7890 ( .A1(n6919), .A2(keyinput227), .B1(keyinput184), .B2(n6918), 
        .ZN(n6917) );
  OAI221_X1 U7891 ( .B1(n6919), .B2(keyinput227), .C1(n6918), .C2(keyinput184), 
        .A(n6917), .ZN(n6926) );
  INV_X1 U7892 ( .A(DATAI_24_), .ZN(n7062) );
  AOI22_X1 U7893 ( .A1(n7116), .A2(keyinput173), .B1(keyinput160), .B2(n7062), 
        .ZN(n6920) );
  OAI221_X1 U7894 ( .B1(n7116), .B2(keyinput173), .C1(n7062), .C2(keyinput160), 
        .A(n6920), .ZN(n6925) );
  INV_X1 U7895 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6923) );
  AOI22_X1 U7896 ( .A1(n6923), .A2(keyinput222), .B1(keyinput167), .B2(n6922), 
        .ZN(n6921) );
  OAI221_X1 U7897 ( .B1(n6923), .B2(keyinput222), .C1(n6922), .C2(keyinput167), 
        .A(n6921), .ZN(n6924) );
  NOR4_X1 U7898 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n6968)
         );
  INV_X1 U7899 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6929) );
  AOI22_X1 U7900 ( .A1(n7090), .A2(keyinput150), .B1(keyinput199), .B2(n6929), 
        .ZN(n6928) );
  OAI221_X1 U7901 ( .B1(n7090), .B2(keyinput150), .C1(n6929), .C2(keyinput199), 
        .A(n6928), .ZN(n6941) );
  INV_X1 U7902 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7903 ( .A1(n6932), .A2(keyinput234), .B1(n6931), .B2(keyinput208), 
        .ZN(n6930) );
  OAI221_X1 U7904 ( .B1(n6932), .B2(keyinput234), .C1(n6931), .C2(keyinput208), 
        .A(n6930), .ZN(n6940) );
  INV_X1 U7905 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U7906 ( .A1(n6935), .A2(keyinput255), .B1(keyinput220), .B2(n6934), 
        .ZN(n6933) );
  OAI221_X1 U7907 ( .B1(n6935), .B2(keyinput255), .C1(n6934), .C2(keyinput220), 
        .A(n6933), .ZN(n6939) );
  XNOR2_X1 U7908 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .B(keyinput245), .ZN(
        n6937) );
  XNOR2_X1 U7909 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput190), .ZN(n6936) );
  NAND2_X1 U7910 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  NOR4_X1 U7911 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n6967)
         );
  AOI22_X1 U7912 ( .A1(n3702), .A2(keyinput211), .B1(n6943), .B2(keyinput241), 
        .ZN(n6942) );
  OAI221_X1 U7913 ( .B1(n3702), .B2(keyinput211), .C1(n6943), .C2(keyinput241), 
        .A(n6942), .ZN(n6953) );
  AOI22_X1 U7914 ( .A1(n7056), .A2(keyinput187), .B1(n7076), .B2(keyinput191), 
        .ZN(n6944) );
  OAI221_X1 U7915 ( .B1(n7056), .B2(keyinput187), .C1(n7076), .C2(keyinput191), 
        .A(n6944), .ZN(n6952) );
  AOI22_X1 U7916 ( .A1(n6947), .A2(keyinput249), .B1(n6946), .B2(keyinput179), 
        .ZN(n6945) );
  OAI221_X1 U7917 ( .B1(n6947), .B2(keyinput249), .C1(n6946), .C2(keyinput179), 
        .A(n6945), .ZN(n6951) );
  INV_X1 U7918 ( .A(DATAI_18_), .ZN(n7047) );
  AOI22_X1 U7919 ( .A1(n6949), .A2(keyinput129), .B1(keyinput189), .B2(n7047), 
        .ZN(n6948) );
  OAI221_X1 U7920 ( .B1(n6949), .B2(keyinput129), .C1(n7047), .C2(keyinput189), 
        .A(n6948), .ZN(n6950) );
  NOR4_X1 U7921 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n6966)
         );
  INV_X1 U7922 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U7923 ( .A1(n7123), .A2(keyinput238), .B1(keyinput248), .B2(n6955), 
        .ZN(n6954) );
  OAI221_X1 U7924 ( .B1(n7123), .B2(keyinput238), .C1(n6955), .C2(keyinput248), 
        .A(n6954), .ZN(n6964) );
  AOI22_X1 U7925 ( .A1(n7049), .A2(keyinput197), .B1(keyinput152), .B2(n4094), 
        .ZN(n6956) );
  OAI221_X1 U7926 ( .B1(n7049), .B2(keyinput197), .C1(n4094), .C2(keyinput152), 
        .A(n6956), .ZN(n6963) );
  INV_X1 U7927 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U7928 ( .A1(n7093), .A2(keyinput202), .B1(n6958), .B2(keyinput198), 
        .ZN(n6957) );
  OAI221_X1 U7929 ( .B1(n7093), .B2(keyinput202), .C1(n6958), .C2(keyinput198), 
        .A(n6957), .ZN(n6962) );
  INV_X1 U7930 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7931 ( .A1(n6960), .A2(keyinput194), .B1(n7057), .B2(keyinput147), 
        .ZN(n6959) );
  OAI221_X1 U7932 ( .B1(n6960), .B2(keyinput194), .C1(n7057), .C2(keyinput147), 
        .A(n6959), .ZN(n6961) );
  NOR4_X1 U7933 ( .A1(n6964), .A2(n6963), .A3(n6962), .A4(n6961), .ZN(n6965)
         );
  NAND4_X1 U7934 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n7024)
         );
  INV_X1 U7935 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6970) );
  AOI22_X1 U7936 ( .A1(n6971), .A2(keyinput128), .B1(n6970), .B2(keyinput252), 
        .ZN(n6969) );
  OAI221_X1 U7937 ( .B1(n6971), .B2(keyinput128), .C1(n6970), .C2(keyinput252), 
        .A(n6969), .ZN(n6980) );
  AOI22_X1 U7938 ( .A1(n7145), .A2(keyinput157), .B1(keyinput156), .B2(n7139), 
        .ZN(n6972) );
  OAI221_X1 U7939 ( .B1(n7145), .B2(keyinput157), .C1(n7139), .C2(keyinput156), 
        .A(n6972), .ZN(n6979) );
  AOI22_X1 U7940 ( .A1(n7094), .A2(keyinput161), .B1(n6974), .B2(keyinput251), 
        .ZN(n6973) );
  OAI221_X1 U7941 ( .B1(n7094), .B2(keyinput161), .C1(n6974), .C2(keyinput251), 
        .A(n6973), .ZN(n6978) );
  XOR2_X1 U7942 ( .A(n3998), .B(keyinput139), .Z(n6976) );
  XNOR2_X1 U7943 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .B(keyinput170), .ZN(
        n6975) );
  NAND2_X1 U7944 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  NOR4_X1 U7945 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n7022)
         );
  AOI22_X1 U7946 ( .A1(n7109), .A2(keyinput203), .B1(keyinput232), .B2(n7138), 
        .ZN(n6981) );
  OAI221_X1 U7947 ( .B1(n7109), .B2(keyinput203), .C1(n7138), .C2(keyinput232), 
        .A(n6981), .ZN(n6993) );
  INV_X1 U7948 ( .A(DATAI_25_), .ZN(n6984) );
  AOI22_X1 U7949 ( .A1(n6984), .A2(keyinput151), .B1(keyinput216), .B2(n6983), 
        .ZN(n6982) );
  OAI221_X1 U7950 ( .B1(n6984), .B2(keyinput151), .C1(n6983), .C2(keyinput216), 
        .A(n6982), .ZN(n6992) );
  AOI22_X1 U7951 ( .A1(n6986), .A2(keyinput188), .B1(keyinput218), .B2(n7125), 
        .ZN(n6985) );
  OAI221_X1 U7952 ( .B1(n6986), .B2(keyinput188), .C1(n7125), .C2(keyinput218), 
        .A(n6985), .ZN(n6991) );
  INV_X1 U7953 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7954 ( .A1(n6989), .A2(keyinput171), .B1(n6988), .B2(keyinput182), 
        .ZN(n6987) );
  OAI221_X1 U7955 ( .B1(n6989), .B2(keyinput171), .C1(n6988), .C2(keyinput182), 
        .A(n6987), .ZN(n6990) );
  NOR4_X1 U7956 ( .A1(n6993), .A2(n6992), .A3(n6991), .A4(n6990), .ZN(n7021)
         );
  AOI22_X1 U7957 ( .A1(n7110), .A2(keyinput185), .B1(keyinput231), .B2(n6995), 
        .ZN(n6994) );
  OAI221_X1 U7958 ( .B1(n7110), .B2(keyinput185), .C1(n6995), .C2(keyinput231), 
        .A(n6994), .ZN(n7005) );
  AOI22_X1 U7959 ( .A1(n7075), .A2(keyinput130), .B1(n4018), .B2(keyinput175), 
        .ZN(n6996) );
  OAI221_X1 U7960 ( .B1(n7075), .B2(keyinput130), .C1(n4018), .C2(keyinput175), 
        .A(n6996), .ZN(n7004) );
  AOI22_X1 U7961 ( .A1(n6999), .A2(keyinput159), .B1(n6998), .B2(keyinput243), 
        .ZN(n6997) );
  OAI221_X1 U7962 ( .B1(n6999), .B2(keyinput159), .C1(n6998), .C2(keyinput243), 
        .A(n6997), .ZN(n7003) );
  AOI22_X1 U7963 ( .A1(n7001), .A2(keyinput206), .B1(n7091), .B2(keyinput244), 
        .ZN(n7000) );
  OAI221_X1 U7964 ( .B1(n7001), .B2(keyinput206), .C1(n7091), .C2(keyinput244), 
        .A(n7000), .ZN(n7002) );
  NOR4_X1 U7965 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n7020)
         );
  AOI22_X1 U7966 ( .A1(n7007), .A2(keyinput134), .B1(keyinput137), .B2(n7043), 
        .ZN(n7006) );
  OAI221_X1 U7967 ( .B1(n7007), .B2(keyinput134), .C1(n7043), .C2(keyinput137), 
        .A(n7006), .ZN(n7018) );
  INV_X1 U7968 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n7107) );
  AOI22_X1 U7969 ( .A1(n7009), .A2(keyinput240), .B1(n7107), .B2(keyinput217), 
        .ZN(n7008) );
  AOI22_X1 U7970 ( .A1(n7141), .A2(keyinput205), .B1(keyinput132), .B2(n7011), 
        .ZN(n7010) );
  OAI221_X1 U7971 ( .B1(n7141), .B2(keyinput205), .C1(n7011), .C2(keyinput132), 
        .A(n7010), .ZN(n7016) );
  XOR2_X1 U7972 ( .A(n7012), .B(keyinput236), .Z(n7014) );
  XNOR2_X1 U7973 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput155), .ZN(
        n7013) );
  NAND2_X1 U7974 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  NOR4_X1 U7975 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7019)
         );
  NAND4_X1 U7976 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n7023)
         );
  NOR4_X1 U7977 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n7023), .ZN(n7159)
         );
  AOI22_X1 U7978 ( .A1(n7029), .A2(keyinput65), .B1(n7028), .B2(keyinput73), 
        .ZN(n7027) );
  OAI221_X1 U7979 ( .B1(n7029), .B2(keyinput65), .C1(n7028), .C2(keyinput73), 
        .A(n7027), .ZN(n7039) );
  AOI22_X1 U7980 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput12), .B1(n7031), 
        .B2(keyinput85), .ZN(n7030) );
  OAI221_X1 U7981 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput12), .C1(n7031), 
        .C2(keyinput85), .A(n7030), .ZN(n7038) );
  AOI22_X1 U7982 ( .A1(ADDRESS_REG_22__SCAN_IN), .A2(keyinput60), .B1(
        INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput99), .ZN(n7032) );
  OAI221_X1 U7983 ( .B1(ADDRESS_REG_22__SCAN_IN), .B2(keyinput60), .C1(
        INSTQUEUE_REG_1__1__SCAN_IN), .C2(keyinput99), .A(n7032), .ZN(n7037)
         );
  XOR2_X1 U7984 ( .A(n7033), .B(keyinput98), .Z(n7035) );
  XNOR2_X1 U7985 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput46), .ZN(
        n7034) );
  NAND2_X1 U7986 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  NOR4_X1 U7987 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7088)
         );
  INV_X1 U7988 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n7041) );
  AOI22_X1 U7989 ( .A1(n7041), .A2(keyinput13), .B1(keyinput47), .B2(n4018), 
        .ZN(n7040) );
  OAI221_X1 U7990 ( .B1(n7041), .B2(keyinput13), .C1(n4018), .C2(keyinput47), 
        .A(n7040), .ZN(n7054) );
  INV_X1 U7991 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n7044) );
  AOI22_X1 U7992 ( .A1(n7044), .A2(keyinput40), .B1(keyinput9), .B2(n7043), 
        .ZN(n7042) );
  OAI221_X1 U7993 ( .B1(n7044), .B2(keyinput40), .C1(n7043), .C2(keyinput9), 
        .A(n7042), .ZN(n7053) );
  INV_X1 U7994 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U7995 ( .A1(n7047), .A2(keyinput61), .B1(n7046), .B2(keyinput109), 
        .ZN(n7045) );
  OAI221_X1 U7996 ( .B1(n7047), .B2(keyinput61), .C1(n7046), .C2(keyinput109), 
        .A(n7045), .ZN(n7052) );
  AOI22_X1 U7997 ( .A1(n7050), .A2(keyinput114), .B1(n7049), .B2(keyinput69), 
        .ZN(n7048) );
  OAI221_X1 U7998 ( .B1(n7050), .B2(keyinput114), .C1(n7049), .C2(keyinput69), 
        .A(n7048), .ZN(n7051) );
  NOR4_X1 U7999 ( .A1(n7054), .A2(n7053), .A3(n7052), .A4(n7051), .ZN(n7087)
         );
  AOI22_X1 U8000 ( .A1(n7057), .A2(keyinput19), .B1(keyinput59), .B2(n7056), 
        .ZN(n7055) );
  OAI221_X1 U8001 ( .B1(n7057), .B2(keyinput19), .C1(n7056), .C2(keyinput59), 
        .A(n7055), .ZN(n7070) );
  INV_X1 U8002 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U8003 ( .A1(n7060), .A2(keyinput53), .B1(n7059), .B2(keyinput7), 
        .ZN(n7058) );
  OAI221_X1 U8004 ( .B1(n7060), .B2(keyinput53), .C1(n7059), .C2(keyinput7), 
        .A(n7058), .ZN(n7069) );
  AOI22_X1 U8005 ( .A1(n7063), .A2(keyinput18), .B1(n7062), .B2(keyinput32), 
        .ZN(n7061) );
  OAI221_X1 U8006 ( .B1(n7063), .B2(keyinput18), .C1(n7062), .C2(keyinput32), 
        .A(n7061), .ZN(n7068) );
  AOI22_X1 U8007 ( .A1(n7066), .A2(keyinput17), .B1(keyinput117), .B2(n7065), 
        .ZN(n7064) );
  OAI221_X1 U8008 ( .B1(n7066), .B2(keyinput17), .C1(n7065), .C2(keyinput117), 
        .A(n7064), .ZN(n7067) );
  NOR4_X1 U8009 ( .A1(n7070), .A2(n7069), .A3(n7068), .A4(n7067), .ZN(n7086)
         );
  INV_X1 U8010 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n7072) );
  AOI22_X1 U8011 ( .A1(n7073), .A2(keyinput84), .B1(n7072), .B2(keyinput25), 
        .ZN(n7071) );
  OAI221_X1 U8012 ( .B1(n7073), .B2(keyinput84), .C1(n7072), .C2(keyinput25), 
        .A(n7071), .ZN(n7084) );
  AOI22_X1 U8013 ( .A1(n7076), .A2(keyinput63), .B1(keyinput2), .B2(n7075), 
        .ZN(n7074) );
  OAI221_X1 U8014 ( .B1(n7076), .B2(keyinput63), .C1(n7075), .C2(keyinput2), 
        .A(n7074), .ZN(n7083) );
  AOI22_X1 U8015 ( .A1(n7078), .A2(keyinput16), .B1(n3719), .B2(keyinput26), 
        .ZN(n7077) );
  OAI221_X1 U8016 ( .B1(n7078), .B2(keyinput16), .C1(n3719), .C2(keyinput26), 
        .A(n7077), .ZN(n7082) );
  AOI22_X1 U8017 ( .A1(n4705), .A2(keyinput125), .B1(n7080), .B2(keyinput118), 
        .ZN(n7079) );
  OAI221_X1 U8018 ( .B1(n4705), .B2(keyinput125), .C1(n7080), .C2(keyinput118), 
        .A(n7079), .ZN(n7081) );
  NOR4_X1 U8019 ( .A1(n7084), .A2(n7083), .A3(n7082), .A4(n7081), .ZN(n7085)
         );
  NAND4_X1 U8020 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n7158)
         );
  AOI22_X1 U8021 ( .A1(n7091), .A2(keyinput116), .B1(keyinput22), .B2(n7090), 
        .ZN(n7089) );
  OAI221_X1 U8022 ( .B1(n7091), .B2(keyinput116), .C1(n7090), .C2(keyinput22), 
        .A(n7089), .ZN(n7104) );
  AOI22_X1 U8023 ( .A1(n7094), .A2(keyinput33), .B1(n7093), .B2(keyinput74), 
        .ZN(n7092) );
  OAI221_X1 U8024 ( .B1(n7094), .B2(keyinput33), .C1(n7093), .C2(keyinput74), 
        .A(n7092), .ZN(n7103) );
  INV_X1 U8025 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n7096) );
  AOI22_X1 U8026 ( .A1(n7097), .A2(keyinput20), .B1(n7096), .B2(keyinput79), 
        .ZN(n7095) );
  OAI221_X1 U8027 ( .B1(n7097), .B2(keyinput20), .C1(n7096), .C2(keyinput79), 
        .A(n7095), .ZN(n7102) );
  XOR2_X1 U8028 ( .A(n7098), .B(keyinput21), .Z(n7100) );
  XNOR2_X1 U8029 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput126), .ZN(n7099) );
  NAND2_X1 U8030 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  NOR4_X1 U8031 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), .ZN(n7156)
         );
  AOI22_X1 U8032 ( .A1(n7107), .A2(keyinput89), .B1(keyinput97), .B2(n7106), 
        .ZN(n7105) );
  OAI221_X1 U8033 ( .B1(n7107), .B2(keyinput89), .C1(n7106), .C2(keyinput97), 
        .A(n7105), .ZN(n7120) );
  AOI22_X1 U8034 ( .A1(n7110), .A2(keyinput57), .B1(n7109), .B2(keyinput75), 
        .ZN(n7108) );
  OAI221_X1 U8035 ( .B1(n7110), .B2(keyinput57), .C1(n7109), .C2(keyinput75), 
        .A(n7108), .ZN(n7119) );
  INV_X1 U8036 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n7112) );
  AOI22_X1 U8037 ( .A1(n7113), .A2(keyinput119), .B1(n7112), .B2(keyinput96), 
        .ZN(n7111) );
  OAI221_X1 U8038 ( .B1(n7113), .B2(keyinput119), .C1(n7112), .C2(keyinput96), 
        .A(n7111), .ZN(n7118) );
  AOI22_X1 U8039 ( .A1(n7116), .A2(keyinput45), .B1(n7115), .B2(keyinput14), 
        .ZN(n7114) );
  OAI221_X1 U8040 ( .B1(n7116), .B2(keyinput45), .C1(n7115), .C2(keyinput14), 
        .A(n7114), .ZN(n7117) );
  NOR4_X1 U8041 ( .A1(n7120), .A2(n7119), .A3(n7118), .A4(n7117), .ZN(n7155)
         );
  AOI22_X1 U8042 ( .A1(n7123), .A2(keyinput110), .B1(keyinput37), .B2(n7122), 
        .ZN(n7121) );
  OAI221_X1 U8043 ( .B1(n7123), .B2(keyinput110), .C1(n7122), .C2(keyinput37), 
        .A(n7121), .ZN(n7136) );
  AOI22_X1 U8044 ( .A1(n7126), .A2(keyinput52), .B1(keyinput90), .B2(n7125), 
        .ZN(n7124) );
  OAI221_X1 U8045 ( .B1(n7126), .B2(keyinput52), .C1(n7125), .C2(keyinput90), 
        .A(n7124), .ZN(n7135) );
  AOI22_X1 U8046 ( .A1(n7129), .A2(keyinput93), .B1(n7128), .B2(keyinput38), 
        .ZN(n7127) );
  OAI221_X1 U8047 ( .B1(n7129), .B2(keyinput93), .C1(n7128), .C2(keyinput38), 
        .A(n7127), .ZN(n7134) );
  INV_X1 U8048 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n7130) );
  XOR2_X1 U8049 ( .A(n7130), .B(keyinput36), .Z(n7132) );
  XNOR2_X1 U8050 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput27), .ZN(
        n7131) );
  NAND2_X1 U8051 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  NOR4_X1 U8052 ( .A1(n7136), .A2(n7135), .A3(n7134), .A4(n7133), .ZN(n7154)
         );
  AOI22_X1 U8053 ( .A1(n7139), .A2(keyinput28), .B1(keyinput104), .B2(n7138), 
        .ZN(n7137) );
  OAI221_X1 U8054 ( .B1(n7139), .B2(keyinput28), .C1(n7138), .C2(keyinput104), 
        .A(n7137), .ZN(n7152) );
  INV_X1 U8055 ( .A(DATAI_31_), .ZN(n7142) );
  AOI22_X1 U8056 ( .A1(n7142), .A2(keyinput81), .B1(keyinput77), .B2(n7141), 
        .ZN(n7140) );
  OAI221_X1 U8057 ( .B1(n7142), .B2(keyinput81), .C1(n7141), .C2(keyinput77), 
        .A(n7140), .ZN(n7151) );
  AOI22_X1 U8058 ( .A1(n7145), .A2(keyinput29), .B1(n7144), .B2(keyinput91), 
        .ZN(n7143) );
  OAI221_X1 U8059 ( .B1(n7145), .B2(keyinput29), .C1(n7144), .C2(keyinput91), 
        .A(n7143), .ZN(n7150) );
  XOR2_X1 U8060 ( .A(n7146), .B(keyinput58), .Z(n7148) );
  XNOR2_X1 U8061 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .B(keyinput30), .ZN(n7147) );
  NAND2_X1 U8062 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  NOR4_X1 U8063 ( .A1(n7152), .A2(n7151), .A3(n7150), .A4(n7149), .ZN(n7153)
         );
  NAND4_X1 U8064 ( .A1(n7156), .A2(n7155), .A3(n7154), .A4(n7153), .ZN(n7157)
         );
  NOR3_X1 U8065 ( .A1(n7159), .A2(n7158), .A3(n7157), .ZN(n7197) );
  OAI22_X1 U8066 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput8), .B1(
        keyinput5), .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n7160) );
  AOI221_X1 U8067 ( .B1(INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput8), .C1(
        INSTQUEUE_REG_8__6__SCAN_IN), .C2(keyinput5), .A(n7160), .ZN(n7167) );
  OAI22_X1 U8068 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput72), .B1(
        keyinput34), .B2(LWORD_REG_2__SCAN_IN), .ZN(n7161) );
  AOI221_X1 U8069 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput72), .C1(
        LWORD_REG_2__SCAN_IN), .C2(keyinput34), .A(n7161), .ZN(n7166) );
  OAI22_X1 U8070 ( .A1(REIP_REG_13__SCAN_IN), .A2(keyinput55), .B1(keyinput10), 
        .B2(DATAI_10_), .ZN(n7162) );
  AOI221_X1 U8071 ( .B1(REIP_REG_13__SCAN_IN), .B2(keyinput55), .C1(DATAI_10_), 
        .C2(keyinput10), .A(n7162), .ZN(n7165) );
  OAI22_X1 U8072 ( .A1(EBX_REG_24__SCAN_IN), .A2(keyinput51), .B1(keyinput35), 
        .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n7163) );
  AOI221_X1 U8073 ( .B1(EBX_REG_24__SCAN_IN), .B2(keyinput51), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput35), .A(n7163), .ZN(n7164) );
  NAND4_X1 U8074 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n7195)
         );
  OAI22_X1 U8075 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(keyinput49), .B1(
        DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput120), .ZN(n7168) );
  AOI221_X1 U8076 ( .B1(INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput49), .C1(
        keyinput120), .C2(DATAWIDTH_REG_6__SCAN_IN), .A(n7168), .ZN(n7175) );
  OAI22_X1 U8077 ( .A1(REIP_REG_1__SCAN_IN), .A2(keyinput115), .B1(keyinput103), .B2(ADDRESS_REG_1__SCAN_IN), .ZN(n7169) );
  AOI221_X1 U8078 ( .B1(REIP_REG_1__SCAN_IN), .B2(keyinput115), .C1(
        ADDRESS_REG_1__SCAN_IN), .C2(keyinput103), .A(n7169), .ZN(n7174) );
  OAI22_X1 U8079 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(keyinput3), .B1(
        EAX_REG_11__SCAN_IN), .B2(keyinput39), .ZN(n7170) );
  AOI221_X1 U8080 ( .B1(INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput3), .C1(
        keyinput39), .C2(EAX_REG_11__SCAN_IN), .A(n7170), .ZN(n7173) );
  OAI22_X1 U8081 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput92), .B1(
        DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput44), .ZN(n7171) );
  AOI221_X1 U8082 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput92), .C1(keyinput44), .C2(DATAWIDTH_REG_14__SCAN_IN), .A(n7171), .ZN(n7172) );
  NAND4_X1 U8083 ( .A1(n7175), .A2(n7174), .A3(n7173), .A4(n7172), .ZN(n7194)
         );
  OAI22_X1 U8084 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput48), .B1(
        keyinput112), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7176) );
  AOI221_X1 U8085 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput48), 
        .C1(PHYADDRPOINTER_REG_9__SCAN_IN), .C2(keyinput112), .A(n7176), .ZN(
        n7183) );
  OAI22_X1 U8086 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(keyinput70), .B1(
        keyinput121), .B2(ADDRESS_REG_6__SCAN_IN), .ZN(n7177) );
  AOI221_X1 U8087 ( .B1(INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput70), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(keyinput121), .A(n7177), .ZN(n7182) );
  OAI22_X1 U8088 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput41), .B1(
        keyinput23), .B2(DATAI_25_), .ZN(n7178) );
  AOI221_X1 U8089 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput41), 
        .C1(DATAI_25_), .C2(keyinput23), .A(n7178), .ZN(n7181) );
  OAI22_X1 U8090 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(keyinput42), .B1(
        keyinput127), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n7179) );
  AOI221_X1 U8091 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput42), .C1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput127), .A(n7179), .ZN(n7180) );
  NAND4_X1 U8092 ( .A1(n7183), .A2(n7182), .A3(n7181), .A4(n7180), .ZN(n7193)
         );
  OAI22_X1 U8093 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(keyinput124), .B1(
        EAX_REG_28__SCAN_IN), .B2(keyinput24), .ZN(n7184) );
  AOI221_X1 U8094 ( .B1(INSTQUEUE_REG_10__0__SCAN_IN), .B2(keyinput124), .C1(
        keyinput24), .C2(EAX_REG_28__SCAN_IN), .A(n7184), .ZN(n7191) );
  OAI22_X1 U8095 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(keyinput62), .B1(
        EAX_REG_3__SCAN_IN), .B2(keyinput86), .ZN(n7185) );
  AOI221_X1 U8096 ( .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput62), .C1(
        keyinput86), .C2(EAX_REG_3__SCAN_IN), .A(n7185), .ZN(n7190) );
  OAI22_X1 U8097 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput11), .B1(
        EAX_REG_2__SCAN_IN), .B2(keyinput15), .ZN(n7186) );
  AOI221_X1 U8098 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput11), .C1(
        keyinput15), .C2(EAX_REG_2__SCAN_IN), .A(n7186), .ZN(n7189) );
  OAI22_X1 U8099 ( .A1(EAX_REG_6__SCAN_IN), .A2(keyinput83), .B1(keyinput67), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n7187) );
  AOI221_X1 U8100 ( .B1(EAX_REG_6__SCAN_IN), .B2(keyinput83), .C1(
        REIP_REG_8__SCAN_IN), .C2(keyinput67), .A(n7187), .ZN(n7188) );
  NAND4_X1 U8101 ( .A1(n7191), .A2(n7190), .A3(n7189), .A4(n7188), .ZN(n7192)
         );
  NOR4_X1 U8102 ( .A1(n7195), .A2(n7194), .A3(n7193), .A4(n7192), .ZN(n7196)
         );
  NAND3_X1 U8103 ( .A1(n7198), .A2(n7197), .A3(n7196), .ZN(n7212) );
  NAND2_X1 U8104 ( .A1(n7199), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n7208)
         );
  OAI22_X1 U8105 ( .A1(n7203), .A2(n7202), .B1(n7201), .B2(n7200), .ZN(n7204)
         );
  AOI21_X1 U8106 ( .B1(n7206), .B2(n7205), .A(n7204), .ZN(n7207) );
  OAI211_X1 U8107 ( .C1(n7210), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7211)
         );
  XNOR2_X1 U8108 ( .A(n7212), .B(n7211), .ZN(U3120) );
  AND2_X1 U3661 ( .A1(n3321), .A2(n4519), .ZN(n3540) );
  AND2_X2 U4088 ( .A1(n4523), .A2(n3321), .ZN(n3382) );
  CLKBUF_X1 U3669 ( .A(n3439), .Z(n3727) );
  NAND2_X1 U3672 ( .A1(n3464), .A2(n3463), .ZN(n4471) );
  CLKBUF_X1 U3683 ( .A(n4589), .Z(n3200) );
endmodule

