

module b14_C_SARLock_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005;

  INV_X1 U2402 ( .A(n3062), .ZN(n3077) );
  INV_X1 U2405 ( .A(n2866), .ZN(n2849) );
  AND2_X1 U2406 ( .A1(n3130), .A2(n3131), .ZN(n3133) );
  OAI21_X1 U2407 ( .B1(n3570), .B2(n3572), .A(n3571), .ZN(n3878) );
  INV_X2 U2408 ( .A(n3377), .ZN(n3372) );
  NAND2_X2 U2409 ( .A1(n2943), .A2(n2942), .ZN(n3570) );
  INV_X2 U2410 ( .A(n2991), .ZN(n3009) );
  AND4_X1 U2411 ( .A1(n2533), .A2(n2532), .A3(n2531), .A4(n2530), .ZN(n3330)
         );
  INV_X1 U2412 ( .A(n2542), .ZN(n3501) );
  INV_X2 U2413 ( .A(n3311), .ZN(n2850) );
  INV_X1 U2414 ( .A(n4167), .ZN(n3331) );
  NAND4_X1 U2415 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n4165)
         );
  INV_X4 U2416 ( .A(n2713), .ZN(n2159) );
  OR2_X1 U2417 ( .A1(n2476), .A2(IR_REG_28__SCAN_IN), .ZN(n2462) );
  AOI21_X1 U2418 ( .B1(n2476), .B2(IR_REG_27__SCAN_IN), .A(n2353), .ZN(n2461)
         );
  XNOR2_X1 U2419 ( .A(n2395), .B(IR_REG_1__SCAN_IN), .ZN(n2482) );
  MUX2_X1 U2420 ( .A(REG0_REG_28__SCAN_IN), .B(n3137), .S(n4683), .Z(n3138) );
  MUX2_X1 U2421 ( .A(REG1_REG_28__SCAN_IN), .B(n3137), .S(n4688), .Z(n3129) );
  AOI211_X1 U2422 ( .C1(n3904), .C2(n4544), .A(n3903), .B(n3902), .ZN(n3905)
         );
  OR2_X1 U2423 ( .A1(n3937), .A2(n3021), .ZN(n2219) );
  NAND2_X1 U2424 ( .A1(n2333), .A2(n2331), .ZN(n3119) );
  INV_X1 U2425 ( .A(n3895), .ZN(n3134) );
  OR2_X1 U2426 ( .A1(n3133), .A2(n3132), .ZN(n3895) );
  OAI21_X1 U2427 ( .B1(n3842), .B2(n4131), .A(n2674), .ZN(n4372) );
  NAND2_X1 U2428 ( .A1(n2355), .A2(n3114), .ZN(n3115) );
  OAI21_X1 U2429 ( .B1(n3516), .B2(n2785), .A(n4048), .ZN(n3558) );
  NAND2_X1 U2430 ( .A1(n2357), .A2(n2927), .ZN(n3603) );
  OAI21_X1 U2431 ( .B1(n3391), .B2(n2780), .A(n4043), .ZN(n3411) );
  NAND2_X1 U2432 ( .A1(n3397), .A2(n2559), .ZN(n3477) );
  AND2_X1 U2433 ( .A1(n2919), .A2(n2918), .ZN(n3613) );
  INV_X2 U2434 ( .A(n4544), .ZN(n2160) );
  INV_X1 U2435 ( .A(n3591), .ZN(n4164) );
  INV_X1 U2436 ( .A(n3330), .ZN(n3445) );
  INV_X1 U2437 ( .A(n3536), .ZN(n3489) );
  AND4_X1 U2438 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .ZN(n3536)
         );
  AND4_X1 U2439 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n3620)
         );
  AND4_X1 U2440 ( .A1(n2581), .A2(n2580), .A3(n2579), .A4(n2578), .ZN(n3591)
         );
  NAND2_X1 U2441 ( .A1(n3403), .A2(n2857), .ZN(n2991) );
  AND4_X1 U2442 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n2542)
         );
  NAND4_X1 U2443 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n4167)
         );
  AND3_X1 U2444 ( .A1(n2546), .A2(n2545), .A3(n2269), .ZN(n3311) );
  NAND3_X1 U2445 ( .A1(n4531), .A2(n4530), .A3(n2815), .ZN(n2851) );
  OAI21_X1 U2446 ( .B1(n2773), .B2(n2397), .A(n2529), .ZN(n3160) );
  NAND2_X2 U2447 ( .A1(n3102), .A2(n3158), .ZN(n3062) );
  OAI21_X1 U2448 ( .B1(n2773), .B2(n3224), .A(n2535), .ZN(n3421) );
  NAND2_X1 U2449 ( .A1(n2840), .A2(n4532), .ZN(n3158) );
  NOR2_X4 U2450 ( .A1(n2522), .A2(n2524), .ZN(n2608) );
  NAND2_X2 U2451 ( .A1(n2462), .A2(n2461), .ZN(n2773) );
  INV_X1 U2452 ( .A(n2820), .ZN(n4532) );
  NAND2_X1 U2453 ( .A1(n2520), .A2(n2519), .ZN(n2524) );
  AND2_X1 U2454 ( .A1(n2451), .A2(n2460), .ZN(n4530) );
  OAI21_X1 U2455 ( .B1(n2356), .B2(n4918), .A(n2446), .ZN(n2819) );
  AOI21_X1 U2456 ( .B1(n2169), .B2(n2165), .A(n2242), .ZN(n2241) );
  NOR2_X1 U2457 ( .A1(n2440), .A2(n2439), .ZN(n2464) );
  AND2_X1 U2458 ( .A1(n2182), .A2(n2351), .ZN(n2350) );
  XNOR2_X1 U2459 ( .A(n2207), .B(IR_REG_2__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U2460 ( .A1(n2277), .A2(n2276), .ZN(n2693) );
  AND2_X1 U2461 ( .A1(n2313), .A2(n2358), .ZN(n2312) );
  INV_X1 U2462 ( .A(IR_REG_4__SCAN_IN), .ZN(n4966) );
  INV_X1 U2463 ( .A(IR_REG_23__SCAN_IN), .ZN(n2457) );
  INV_X1 U2464 ( .A(IR_REG_2__SCAN_IN), .ZN(n2358) );
  INV_X1 U2465 ( .A(IR_REG_3__SCAN_IN), .ZN(n2389) );
  INV_X1 U2466 ( .A(IR_REG_17__SCAN_IN), .ZN(n2277) );
  INV_X1 U2467 ( .A(IR_REG_18__SCAN_IN), .ZN(n2276) );
  NOR2_X1 U2468 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2363)
         );
  NOR2_X1 U2469 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2362)
         );
  NOR2_X1 U2470 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2361)
         );
  NOR2_X2 U2471 ( .A1(n3729), .A2(n3744), .ZN(n3778) );
  NAND2_X2 U2472 ( .A1(n2851), .A2(n2848), .ZN(n2866) );
  AND2_X1 U2473 ( .A1(n2851), .A2(n3158), .ZN(n2857) );
  NAND2_X2 U2474 ( .A1(n2462), .A2(n2461), .ZN(n2164) );
  NAND2_X1 U2475 ( .A1(n2462), .A2(n2461), .ZN(n2163) );
  MUX2_X1 U2476 ( .A(IR_REG_31__SCAN_IN), .B(n2518), .S(IR_REG_29__SCAN_IN), 
        .Z(n2520) );
  INV_X1 U2477 ( .A(n2228), .ZN(n2227) );
  OAI21_X1 U2478 ( .B1(n2232), .B2(n2229), .A(n3668), .ZN(n2228) );
  AND2_X1 U2479 ( .A1(n2336), .A2(n2185), .ZN(n2332) );
  NOR2_X1 U2480 ( .A1(n2718), .A2(n2348), .ZN(n2347) );
  INV_X1 U2481 ( .A(n2709), .ZN(n2348) );
  NAND2_X1 U2482 ( .A1(n3203), .A2(n2484), .ZN(n2485) );
  NOR2_X1 U2483 ( .A1(n2262), .A2(n4590), .ZN(n2261) );
  INV_X1 U2484 ( .A(n2426), .ZN(n2262) );
  XNOR2_X1 U2485 ( .A(n2500), .B(n3725), .ZN(n3721) );
  OR2_X1 U2486 ( .A1(n4197), .A2(n2762), .ZN(n3896) );
  OR2_X1 U2487 ( .A1(n2746), .A2(n3982), .ZN(n2755) );
  NOR2_X1 U2488 ( .A1(n4305), .A2(n2344), .ZN(n2343) );
  INV_X1 U2489 ( .A(n2346), .ZN(n2344) );
  NAND2_X1 U2490 ( .A1(n2318), .A2(n2316), .ZN(n2322) );
  NOR2_X1 U2491 ( .A1(n2622), .A2(n2317), .ZN(n2316) );
  INV_X1 U2492 ( .A(n2323), .ZN(n2317) );
  NAND2_X1 U2493 ( .A1(n3335), .A2(n3336), .ZN(n3334) );
  INV_X1 U2494 ( .A(IR_REG_6__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U2495 ( .A1(n2180), .A2(n2275), .ZN(n2440) );
  INV_X1 U2496 ( .A(n2693), .ZN(n2275) );
  OAI21_X1 U2497 ( .B1(n4211), .B2(n2713), .A(n2760), .ZN(n4159) );
  INV_X1 U2498 ( .A(n2230), .ZN(n2229) );
  AND2_X1 U2499 ( .A1(n4083), .A2(n2298), .ZN(n2297) );
  NAND2_X1 U2500 ( .A1(n2301), .A2(n2299), .ZN(n2298) );
  AOI21_X1 U2501 ( .B1(n2781), .B2(n4050), .A(n2309), .ZN(n2308) );
  INV_X1 U2502 ( .A(n4051), .ZN(n2309) );
  NOR2_X1 U2503 ( .A1(n2200), .A2(n2201), .ZN(n2198) );
  INV_X1 U2504 ( .A(n4005), .ZN(n2291) );
  NAND2_X1 U2505 ( .A1(n3508), .A2(n4164), .ZN(n4053) );
  AOI21_X1 U2506 ( .B1(n2558), .B2(n3142), .A(n2557), .ZN(n3397) );
  NOR2_X1 U2507 ( .A1(n3390), .A2(n3393), .ZN(n2557) );
  NAND2_X1 U2508 ( .A1(n3732), .A2(n4117), .ZN(n2295) );
  NAND2_X1 U2509 ( .A1(n2247), .A2(n2775), .ZN(n2246) );
  NAND2_X1 U2510 ( .A1(IR_REG_31__SCAN_IN), .A2(n2693), .ZN(n2247) );
  NAND2_X1 U2511 ( .A1(n2246), .A2(n2165), .ZN(n2244) );
  NAND2_X1 U2512 ( .A1(n2443), .A2(n2777), .ZN(n2243) );
  INV_X1 U2513 ( .A(IR_REG_11__SCAN_IN), .ZN(n4745) );
  INV_X1 U2514 ( .A(n2393), .ZN(n2392) );
  NOR2_X1 U2515 ( .A1(n2236), .A2(n2240), .ZN(n2235) );
  NOR2_X1 U2516 ( .A1(n3468), .A2(n3467), .ZN(n2240) );
  INV_X1 U2517 ( .A(n3381), .ZN(n2236) );
  NOR2_X1 U2518 ( .A1(n2893), .A2(n2239), .ZN(n2238) );
  NAND2_X1 U2519 ( .A1(n2233), .A2(n3876), .ZN(n2232) );
  NAND2_X1 U2520 ( .A1(n3875), .A2(n2231), .ZN(n2230) );
  INV_X1 U2521 ( .A(n3876), .ZN(n2231) );
  INV_X1 U2522 ( .A(n3889), .ZN(n3029) );
  NAND2_X1 U2523 ( .A1(n3601), .A2(n2916), .ZN(n3606) );
  AND2_X1 U2524 ( .A1(n3602), .A2(n2928), .ZN(n2916) );
  AND2_X1 U2525 ( .A1(n2986), .A2(n2985), .ZN(n3802) );
  NAND2_X1 U2526 ( .A1(n2218), .A2(n2178), .ZN(n3425) );
  AND2_X1 U2527 ( .A1(n2949), .A2(n2950), .ZN(n3572) );
  INV_X1 U2528 ( .A(n4307), .ZN(n3956) );
  NOR2_X1 U2529 ( .A1(n2651), .A2(n4694), .ZN(n2658) );
  NAND2_X1 U2530 ( .A1(n2394), .A2(n2266), .ZN(n3202) );
  OR2_X1 U2531 ( .A1(n4540), .A2(n2398), .ZN(n2266) );
  NAND2_X1 U2532 ( .A1(n3201), .A2(n3202), .ZN(n3200) );
  NAND2_X1 U2533 ( .A1(n3213), .A2(n2486), .ZN(n2487) );
  XNOR2_X1 U2534 ( .A(n2202), .B(n4536), .ZN(n3233) );
  NOR2_X1 U2535 ( .A1(n3247), .A2(n2175), .ZN(n2405) );
  AOI21_X1 U2536 ( .B1(n3278), .B2(n3274), .A(n3273), .ZN(n2490) );
  NAND2_X1 U2537 ( .A1(n3287), .A2(REG1_REG_8__SCAN_IN), .ZN(n2199) );
  INV_X1 U2538 ( .A(n2491), .ZN(n2196) );
  NAND2_X1 U2539 ( .A1(n4569), .A2(n2496), .ZN(n2497) );
  INV_X1 U2540 ( .A(n4580), .ZN(n2258) );
  NAND2_X1 U2541 ( .A1(n4598), .A2(n2499), .ZN(n2500) );
  NAND2_X1 U2542 ( .A1(n3721), .A2(REG1_REG_14__SCAN_IN), .ZN(n3720) );
  AOI21_X1 U2543 ( .B1(n4580), .B2(n2261), .A(n2192), .ZN(n2433) );
  NAND2_X1 U2544 ( .A1(n4609), .A2(n2502), .ZN(n2503) );
  NOR2_X1 U2545 ( .A1(n4604), .A2(n2264), .ZN(n2437) );
  AND2_X1 U2546 ( .A1(n4661), .A2(REG2_REG_15__SCAN_IN), .ZN(n2264) );
  NOR2_X1 U2547 ( .A1(n2505), .A2(n4633), .ZN(n4180) );
  NAND2_X1 U2548 ( .A1(n3133), .A2(n2212), .ZN(n2213) );
  NOR2_X1 U2549 ( .A1(n4399), .A2(n2811), .ZN(n2212) );
  AND2_X1 U2550 ( .A1(n2761), .A2(REG3_REG_28__SCAN_IN), .ZN(n4197) );
  AND2_X1 U2551 ( .A1(n2288), .A2(n2283), .ZN(n2282) );
  OR2_X1 U2552 ( .A1(n2293), .A2(n4015), .ZN(n2288) );
  NAND2_X1 U2553 ( .A1(n2289), .A2(n2284), .ZN(n2283) );
  AND2_X1 U2554 ( .A1(n4208), .A2(n2294), .ZN(n2293) );
  AOI21_X1 U2555 ( .B1(n2290), .B2(n2284), .A(n4011), .ZN(n2286) );
  NOR2_X1 U2556 ( .A1(n2755), .A2(n3910), .ZN(n2761) );
  NAND2_X1 U2557 ( .A1(n2337), .A2(n2754), .ZN(n2336) );
  NAND2_X1 U2558 ( .A1(n2738), .A2(n2338), .ZN(n2337) );
  NOR2_X1 U2559 ( .A1(n4221), .A2(n4246), .ZN(n2753) );
  AND2_X1 U2560 ( .A1(n2335), .A2(n4100), .ZN(n2334) );
  OR2_X1 U2561 ( .A1(n2336), .A2(n2338), .ZN(n2335) );
  NAND2_X1 U2562 ( .A1(n2340), .A2(n2176), .ZN(n4275) );
  NOR2_X1 U2563 ( .A1(n2172), .A2(n2342), .ZN(n2341) );
  NAND2_X1 U2564 ( .A1(n4337), .A2(n2347), .ZN(n2345) );
  AOI21_X1 U2565 ( .B1(n2347), .B2(n2710), .A(n2186), .ZN(n2346) );
  OR2_X1 U2566 ( .A1(n2719), .A2(n4728), .ZN(n2732) );
  INV_X1 U2567 ( .A(n2327), .ZN(n2326) );
  OAI21_X1 U2568 ( .B1(n2328), .B2(n2657), .A(n2665), .ZN(n2327) );
  NAND2_X1 U2569 ( .A1(n2329), .A2(n2664), .ZN(n2328) );
  NAND2_X1 U2570 ( .A1(n2322), .A2(n2315), .ZN(n3639) );
  AND2_X1 U2571 ( .A1(n2321), .A2(n2621), .ZN(n2315) );
  INV_X1 U2572 ( .A(n4120), .ZN(n2321) );
  NAND2_X1 U2573 ( .A1(n2325), .A2(n2324), .ZN(n2323) );
  NAND2_X1 U2574 ( .A1(n2601), .A2(n2319), .ZN(n2318) );
  NOR2_X1 U2575 ( .A1(n2613), .A2(n2320), .ZN(n2319) );
  INV_X1 U2576 ( .A(n2600), .ZN(n2320) );
  NAND2_X1 U2577 ( .A1(n2773), .A2(DATAI_4_), .ZN(n2535) );
  NAND2_X1 U2578 ( .A1(n3133), .A2(n2839), .ZN(n4398) );
  NAND2_X1 U2579 ( .A1(n3375), .A2(n3372), .ZN(n3404) );
  AND2_X1 U2580 ( .A1(n3239), .A2(n2840), .ZN(n4479) );
  INV_X1 U2581 ( .A(n3151), .ZN(n3302) );
  OR2_X1 U2582 ( .A1(n2444), .A2(n2443), .ZN(n2356) );
  INV_X1 U2583 ( .A(n2371), .ZN(n2465) );
  OR2_X1 U2584 ( .A1(n2431), .A2(IR_REG_14__SCAN_IN), .ZN(n2375) );
  INV_X1 U2585 ( .A(IR_REG_15__SCAN_IN), .ZN(n4748) );
  AND2_X1 U2586 ( .A1(n2420), .A2(n2419), .ZN(n2602) );
  NAND2_X1 U2587 ( .A1(n2267), .A2(n2268), .ZN(n2393) );
  INV_X1 U2588 ( .A(IR_REG_1__SCAN_IN), .ZN(n2268) );
  NAND2_X1 U2589 ( .A1(n3382), .A2(n3381), .ZN(n3380) );
  AND2_X1 U2590 ( .A1(n2755), .A2(n2747), .ZN(n4236) );
  INV_X1 U2591 ( .A(n3821), .ZN(n3986) );
  INV_X1 U2592 ( .A(n3620), .ZN(n3626) );
  NAND2_X1 U2593 ( .A1(n2206), .A2(n2205), .ZN(n3205) );
  OR2_X1 U2594 ( .A1(n4540), .A2(n3434), .ZN(n2206) );
  NAND2_X1 U2595 ( .A1(n4540), .A2(n3434), .ZN(n2205) );
  NAND2_X1 U2596 ( .A1(n3214), .A2(REG1_REG_3__SCAN_IN), .ZN(n3213) );
  NOR2_X1 U2597 ( .A1(n3246), .A2(n3245), .ZN(n3244) );
  XNOR2_X1 U2598 ( .A(n2405), .B(n4536), .ZN(n3229) );
  NOR2_X1 U2599 ( .A1(n3281), .A2(n3280), .ZN(n3279) );
  XNOR2_X1 U2600 ( .A(n2490), .B(n3291), .ZN(n3287) );
  NAND2_X1 U2601 ( .A1(n4617), .A2(n4615), .ZN(n4616) );
  XNOR2_X1 U2602 ( .A(n2437), .B(n2673), .ZN(n4617) );
  NOR2_X1 U2603 ( .A1(n2478), .A2(n2479), .ZN(n4184) );
  NAND2_X1 U2604 ( .A1(n4626), .A2(n2254), .ZN(n2478) );
  NAND2_X1 U2605 ( .A1(n4636), .A2(n4724), .ZN(n2254) );
  AOI21_X1 U2606 ( .B1(n3119), .B2(n4098), .A(n2767), .ZN(n2774) );
  AND2_X1 U2607 ( .A1(n2270), .A2(n2274), .ZN(n2269) );
  NAND2_X1 U2608 ( .A1(n2549), .A2(REG2_REG_1__SCAN_IN), .ZN(n2545) );
  INV_X1 U2609 ( .A(n2482), .ZN(n2544) );
  NAND2_X1 U2610 ( .A1(n2163), .A2(DATAI_1_), .ZN(n2543) );
  INV_X2 U2611 ( .A(n4686), .ZN(n4688) );
  NOR2_X1 U2612 ( .A1(n3904), .A2(n3126), .ZN(n3127) );
  NOR2_X1 U2613 ( .A1(n2473), .A2(n2311), .ZN(n2310) );
  NAND2_X1 U2614 ( .A1(n2351), .A2(n2516), .ZN(n2311) );
  NAND2_X1 U2615 ( .A1(n3605), .A2(n2934), .ZN(n2937) );
  AOI21_X1 U2616 ( .B1(n2227), .B2(n2229), .A(n2225), .ZN(n2224) );
  INV_X1 U2617 ( .A(n3667), .ZN(n2225) );
  AND2_X1 U2618 ( .A1(n2737), .A2(n2339), .ZN(n2338) );
  INV_X1 U2619 ( .A(n4222), .ZN(n2339) );
  AND2_X1 U2620 ( .A1(n4256), .A2(n4108), .ZN(n4084) );
  NAND2_X1 U2621 ( .A1(n4288), .A2(n4267), .ZN(n2737) );
  INV_X1 U2622 ( .A(n2301), .ZN(n2300) );
  INV_X1 U2623 ( .A(n2347), .ZN(n2342) );
  AOI21_X1 U2624 ( .B1(n3996), .B2(n4076), .A(n2302), .ZN(n2301) );
  INV_X1 U2625 ( .A(n4079), .ZN(n2302) );
  NAND2_X1 U2626 ( .A1(n2303), .A2(n2167), .ZN(n2783) );
  AOI21_X1 U2627 ( .B1(n2308), .B2(n2306), .A(n2305), .ZN(n2304) );
  INV_X1 U2628 ( .A(n4044), .ZN(n2305) );
  OR2_X1 U2629 ( .A1(n3411), .A2(n2307), .ZN(n2303) );
  INV_X1 U2630 ( .A(n2308), .ZN(n2307) );
  OAI21_X1 U2631 ( .B1(n2164), .B2(n2583), .A(n2582), .ZN(n2901) );
  NAND2_X1 U2632 ( .A1(n2773), .A2(DATAI_7_), .ZN(n2582) );
  NAND2_X1 U2633 ( .A1(n2837), .A2(n3501), .ZN(n4043) );
  NAND2_X1 U2634 ( .A1(n4043), .A2(n4039), .ZN(n2556) );
  AND2_X1 U2635 ( .A1(n2534), .A2(n3365), .ZN(n3392) );
  NAND2_X1 U2636 ( .A1(n3335), .A2(n2850), .ZN(n4029) );
  INV_X1 U2637 ( .A(n3178), .ZN(n2831) );
  OR2_X1 U2638 ( .A1(n3777), .A2(n3847), .ZN(n3846) );
  OR2_X1 U2639 ( .A1(n3580), .A2(n3627), .ZN(n2215) );
  AND2_X1 U2640 ( .A1(n4149), .A2(n2820), .ZN(n3239) );
  INV_X1 U2641 ( .A(IR_REG_27__SCAN_IN), .ZN(n2470) );
  NOR2_X1 U2642 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2360)
         );
  INV_X1 U2643 ( .A(IR_REG_28__SCAN_IN), .ZN(n2471) );
  AND2_X1 U2644 ( .A1(n2443), .A2(n4918), .ZN(n2445) );
  INV_X1 U2645 ( .A(IR_REG_21__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U2646 ( .A1(n2929), .A2(n2928), .ZN(n3605) );
  INV_X1 U2647 ( .A(n3603), .ZN(n2929) );
  NAND2_X1 U2648 ( .A1(n3059), .A2(n2249), .ZN(n2248) );
  NOR2_X1 U2649 ( .A1(n2250), .A2(n3976), .ZN(n2249) );
  AND2_X1 U2650 ( .A1(n3020), .A2(n3019), .ZN(n3934) );
  NAND2_X1 U2651 ( .A1(n3005), .A2(n3004), .ZN(n3963) );
  NAND2_X1 U2652 ( .A1(n2981), .A2(n2221), .ZN(n2220) );
  NOR2_X1 U2653 ( .A1(n2987), .A2(n2222), .ZN(n2221) );
  INV_X1 U2654 ( .A(n2980), .ZN(n2222) );
  AND3_X1 U2655 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2568) );
  AND3_X1 U2656 ( .A1(n3155), .A2(n3083), .A3(n3152), .ZN(n3105) );
  AND2_X1 U2657 ( .A1(n2658), .A2(REG3_REG_15__SCAN_IN), .ZN(n2666) );
  INV_X1 U2658 ( .A(n3105), .ZN(n3110) );
  OR2_X1 U2659 ( .A1(n4149), .A2(n4533), .ZN(n3102) );
  NAND2_X1 U2660 ( .A1(n3200), .A2(n2179), .ZN(n2399) );
  INV_X1 U2661 ( .A(n2388), .ZN(n2314) );
  NOR2_X1 U2662 ( .A1(n3251), .A2(n2204), .ZN(n2203) );
  NOR2_X1 U2663 ( .A1(n3233), .A2(n3545), .ZN(n3232) );
  NAND2_X1 U2664 ( .A1(n2196), .A2(n4550), .ZN(n2195) );
  NAND2_X1 U2665 ( .A1(n3287), .A2(n2198), .ZN(n2197) );
  NAND2_X1 U2666 ( .A1(n4570), .A2(n4571), .ZN(n4569) );
  NOR2_X1 U2667 ( .A1(n2253), .A2(n4717), .ZN(n2252) );
  INV_X1 U2668 ( .A(n4185), .ZN(n2253) );
  NAND2_X1 U2669 ( .A1(n2281), .A2(n2278), .ZN(n2804) );
  AOI21_X1 U2670 ( .B1(n2282), .B2(n2280), .A(n2279), .ZN(n2278) );
  NAND2_X1 U2671 ( .A1(n2803), .A2(n2177), .ZN(n2281) );
  NOR2_X1 U2672 ( .A1(n2289), .A2(n4012), .ZN(n2280) );
  OR2_X1 U2673 ( .A1(n4004), .A2(n4013), .ZN(n4096) );
  AOI21_X1 U2674 ( .B1(n2334), .B2(n2332), .A(n2187), .ZN(n2331) );
  INV_X1 U2675 ( .A(n4234), .ZN(n4228) );
  AOI21_X1 U2676 ( .B1(n2803), .B2(n4122), .A(n2802), .ZN(n4226) );
  OAI21_X1 U2677 ( .B1(n4255), .B2(n2738), .A(n2737), .ZN(n4244) );
  NAND2_X1 U2678 ( .A1(n2296), .A2(n2301), .ZN(n4276) );
  NAND2_X1 U2679 ( .A1(n3857), .A2(n3996), .ZN(n2296) );
  NAND2_X1 U2680 ( .A1(n2703), .A2(REG3_REG_20__SCAN_IN), .ZN(n2711) );
  AND2_X1 U2681 ( .A1(n2694), .A2(REG3_REG_19__SCAN_IN), .ZN(n2703) );
  OR2_X1 U2682 ( .A1(n3857), .A2(n4076), .ZN(n4332) );
  NAND2_X1 U2683 ( .A1(n3863), .A2(n2692), .ZN(n4350) );
  NOR2_X1 U2684 ( .A1(n2685), .A2(n2684), .ZN(n2694) );
  AND2_X1 U2685 ( .A1(n4077), .A2(n4074), .ZN(n4131) );
  NAND2_X1 U2686 ( .A1(n2641), .A2(n2640), .ZN(n3685) );
  OR2_X1 U2687 ( .A1(n2615), .A2(n4963), .ZN(n2624) );
  OR2_X1 U2688 ( .A1(n2605), .A2(n2604), .ZN(n2615) );
  NAND2_X1 U2689 ( .A1(n2568), .A2(REG3_REG_6__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U2690 ( .A1(n2303), .A2(n2304), .ZN(n3449) );
  INV_X1 U2691 ( .A(n2901), .ZN(n3508) );
  AND2_X1 U2692 ( .A1(n4038), .A2(n4035), .ZN(n4116) );
  NAND2_X1 U2693 ( .A1(n3358), .A2(n3330), .ZN(n3365) );
  NAND2_X1 U2694 ( .A1(n2273), .A2(n2271), .ZN(n2274) );
  NOR2_X1 U2695 ( .A1(n2524), .A2(n2481), .ZN(n2271) );
  NAND2_X1 U2696 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
  AND2_X1 U2697 ( .A1(n2524), .A2(REG0_REG_1__SCAN_IN), .ZN(n2272) );
  INV_X1 U2698 ( .A(n4479), .ZN(n3403) );
  AND2_X1 U2699 ( .A1(n4232), .A2(n4212), .ZN(n3130) );
  NOR2_X1 U2700 ( .A1(n4245), .A2(n4228), .ZN(n4232) );
  OR2_X1 U2701 ( .A1(n4266), .A2(n4417), .ZN(n4245) );
  INV_X1 U2702 ( .A(n4246), .ZN(n4417) );
  NAND2_X1 U2703 ( .A1(n4289), .A2(n2216), .ZN(n4266) );
  NOR2_X1 U2704 ( .A1(n3042), .A2(n4285), .ZN(n2216) );
  AND2_X1 U2705 ( .A1(n4320), .A2(n4298), .ZN(n4289) );
  NOR2_X1 U2706 ( .A1(n4319), .A2(n4437), .ZN(n4320) );
  INV_X1 U2707 ( .A(n4322), .ZN(n4437) );
  NAND2_X1 U2708 ( .A1(n4373), .A2(n2217), .ZN(n4365) );
  NOR2_X1 U2709 ( .A1(n3836), .A2(n4358), .ZN(n2217) );
  AND2_X1 U2710 ( .A1(n4373), .A2(n3867), .ZN(n4363) );
  NOR2_X2 U2711 ( .A1(n3846), .A2(n4464), .ZN(n4373) );
  NAND2_X1 U2712 ( .A1(n2295), .A2(n3990), .ZN(n3782) );
  NAND2_X1 U2713 ( .A1(n2209), .A2(n2208), .ZN(n3729) );
  INV_X1 U2714 ( .A(n3707), .ZN(n2209) );
  NAND2_X1 U2715 ( .A1(n2211), .A2(n2210), .ZN(n3707) );
  INV_X1 U2716 ( .A(n3705), .ZN(n2211) );
  NOR2_X2 U2717 ( .A1(n2215), .A2(n3657), .ZN(n3649) );
  NAND2_X1 U2718 ( .A1(n3485), .A2(n2214), .ZN(n3580) );
  AND2_X1 U2719 ( .A1(n3581), .A2(n3508), .ZN(n2214) );
  NAND2_X1 U2720 ( .A1(n3485), .A2(n3508), .ZN(n3579) );
  AND2_X1 U2721 ( .A1(n3483), .A2(n3482), .ZN(n3485) );
  NAND2_X1 U2722 ( .A1(n3375), .A2(n2174), .ZN(n3416) );
  NOR2_X1 U2723 ( .A1(n3416), .A2(n3415), .ZN(n3483) );
  INV_X1 U2724 ( .A(n4458), .ZN(n4474) );
  INV_X1 U2725 ( .A(n2852), .ZN(n3335) );
  INV_X1 U2726 ( .A(n3313), .ZN(n3336) );
  AND2_X1 U2727 ( .A1(n3239), .A2(n4143), .ZN(n4463) );
  NAND2_X1 U2728 ( .A1(n2182), .A2(n2472), .ZN(n2473) );
  AND4_X1 U2729 ( .A1(n2449), .A2(n4918), .A3(n2471), .A4(n2470), .ZN(n2472)
         );
  AND2_X1 U2730 ( .A1(n2360), .A2(n2466), .ZN(n2351) );
  OR2_X1 U2731 ( .A1(n2246), .A2(IR_REG_20__SCAN_IN), .ZN(n2245) );
  NAND2_X1 U2732 ( .A1(n2244), .A2(n2243), .ZN(n2242) );
  INV_X1 U2733 ( .A(IR_REG_13__SCAN_IN), .ZN(n2428) );
  AND2_X1 U2734 ( .A1(n2381), .A2(n2380), .ZN(n2631) );
  INV_X1 U2735 ( .A(IR_REG_5__SCAN_IN), .ZN(n2313) );
  AOI21_X1 U2736 ( .B1(n2181), .B2(n3468), .A(n2238), .ZN(n2237) );
  NAND2_X1 U2737 ( .A1(n3878), .A2(n2232), .ZN(n2226) );
  NAND2_X1 U2738 ( .A1(n3886), .A2(n3036), .ZN(n3916) );
  AND4_X1 U2739 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .ZN(n3655)
         );
  NAND2_X1 U2740 ( .A1(n2218), .A2(n2880), .ZN(n3427) );
  OAI21_X1 U2741 ( .B1(n2773), .B2(n2267), .A(n2547), .ZN(n3313) );
  NAND2_X1 U2742 ( .A1(n2163), .A2(DATAI_0_), .ZN(n2547) );
  NAND2_X1 U2743 ( .A1(n2219), .A2(n3024), .ZN(n3888) );
  INV_X1 U2744 ( .A(n3642), .ZN(n3648) );
  NAND2_X1 U2745 ( .A1(n2220), .A2(n2184), .ZN(n3835) );
  INV_X1 U2746 ( .A(n3540), .ZN(n3482) );
  NAND2_X1 U2747 ( .A1(n3380), .A2(n2893), .ZN(n3470) );
  INV_X1 U2748 ( .A(n4261), .ZN(n4221) );
  AOI21_X1 U2749 ( .B1(STATE_REG_SCAN_IN), .B2(n3106), .A(n3301), .ZN(n3821)
         );
  INV_X1 U2750 ( .A(n3792), .ZN(n3814) );
  INV_X1 U2751 ( .A(n3929), .ZN(n3981) );
  OAI21_X1 U2752 ( .B1(n3896), .B2(n2713), .A(n2766), .ZN(n4158) );
  NAND2_X1 U2753 ( .A1(n2752), .A2(n2751), .ZN(n4405) );
  NAND2_X1 U2754 ( .A1(n2728), .A2(n2727), .ZN(n4307) );
  AND2_X1 U2755 ( .A1(n2508), .A2(n2507), .ZN(n3183) );
  XNOR2_X1 U2756 ( .A(n2485), .B(n2265), .ZN(n3214) );
  XNOR2_X1 U2757 ( .A(n2399), .B(n2265), .ZN(n3211) );
  AND2_X1 U2758 ( .A1(n3219), .A2(n2488), .ZN(n3246) );
  AND2_X1 U2759 ( .A1(n2256), .A2(n2255), .ZN(n3281) );
  NAND2_X1 U2760 ( .A1(n2406), .A2(n4536), .ZN(n2255) );
  NAND2_X1 U2761 ( .A1(n3229), .A2(REG2_REG_6__SCAN_IN), .ZN(n2256) );
  OAI21_X1 U2762 ( .B1(n3287), .B2(n2196), .A(n2194), .ZN(n4548) );
  NAND2_X1 U2763 ( .A1(n2199), .A2(n2491), .ZN(n4549) );
  AOI21_X1 U2764 ( .B1(n2491), .B2(n2201), .A(n2200), .ZN(n2194) );
  XNOR2_X1 U2765 ( .A(n2497), .B(n4589), .ZN(n4586) );
  NAND2_X1 U2766 ( .A1(n4586), .A2(REG1_REG_12__SCAN_IN), .ZN(n4585) );
  OAI22_X1 U2767 ( .A1(n2258), .A2(n2257), .B1(n2259), .B2(n4534), .ZN(n2263)
         );
  INV_X1 U2768 ( .A(n2260), .ZN(n2259) );
  NAND2_X1 U2769 ( .A1(n2261), .A2(n3725), .ZN(n2257) );
  NAND2_X1 U2770 ( .A1(n3720), .A2(n2501), .ZN(n4610) );
  XNOR2_X1 U2771 ( .A(n2503), .B(n2673), .ZN(n4620) );
  NOR2_X1 U2772 ( .A1(n4620), .A2(REG1_REG_16__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U2773 ( .A1(n4616), .A2(n2438), .ZN(n4625) );
  AND2_X1 U2774 ( .A1(n2509), .A2(n2508), .ZN(n4630) );
  AND2_X1 U2775 ( .A1(n3183), .A2(n3181), .ZN(n4631) );
  XNOR2_X1 U2776 ( .A(n2251), .B(n4187), .ZN(n4192) );
  NOR2_X1 U2777 ( .A1(n4184), .A2(n2252), .ZN(n2251) );
  XNOR2_X1 U2778 ( .A(n2213), .B(n4394), .ZN(n4542) );
  INV_X1 U2779 ( .A(n2213), .ZN(n4397) );
  AND2_X1 U2780 ( .A1(n3122), .A2(n3121), .ZN(n3904) );
  OAI21_X1 U2781 ( .B1(n2803), .B2(n2285), .A(n2282), .ZN(n3120) );
  INV_X1 U2782 ( .A(n2292), .ZN(n4205) );
  OR2_X1 U2783 ( .A1(n2756), .A2(n2761), .ZN(n4211) );
  OAI21_X1 U2784 ( .B1(n4255), .B2(n2336), .A(n2334), .ZN(n4207) );
  NAND2_X1 U2785 ( .A1(n2345), .A2(n2346), .ZN(n4296) );
  OR2_X1 U2786 ( .A1(n4337), .A2(n2710), .ZN(n2349) );
  AND4_X1 U2787 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n3815)
         );
  INV_X1 U2788 ( .A(n4161), .ZN(n3748) );
  NAND2_X1 U2789 ( .A1(n2322), .A2(n2621), .ZN(n3641) );
  NAND2_X1 U2790 ( .A1(n2318), .A2(n2323), .ZN(n3559) );
  NAND2_X1 U2791 ( .A1(n2601), .A2(n2600), .ZN(n3522) );
  INV_X1 U2792 ( .A(n4368), .ZN(n4647) );
  AND2_X1 U2793 ( .A1(n4544), .A2(n4463), .ZN(n4379) );
  NAND2_X1 U2794 ( .A1(n3302), .A2(n3108), .ZN(n4300) );
  OR2_X1 U2795 ( .A1(n2843), .A2(n3153), .ZN(n4686) );
  INV_X1 U2796 ( .A(n3404), .ZN(n2838) );
  INV_X2 U2797 ( .A(n4682), .ZN(n4683) );
  NAND2_X1 U2798 ( .A1(n2519), .A2(IR_REG_31__SCAN_IN), .ZN(n2517) );
  MUX2_X1 U2799 ( .A(IR_REG_31__SCAN_IN), .B(n2447), .S(IR_REG_26__SCAN_IN), 
        .Z(n2451) );
  NAND2_X1 U2800 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2456) );
  XNOR2_X1 U2801 ( .A(n2776), .B(IR_REG_19__SCAN_IN), .ZN(n4533) );
  OAI21_X1 U2802 ( .B1(n2169), .B2(n2693), .A(IR_REG_31__SCAN_IN), .ZN(n2776)
         );
  AND2_X1 U2803 ( .A1(n2435), .A2(n2377), .ZN(n4661) );
  NAND2_X1 U2804 ( .A1(n2393), .A2(IR_REG_31__SCAN_IN), .ZN(n2207) );
  NAND2_X1 U2805 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2395)
         );
  AOI21_X1 U2806 ( .B1(n4185), .B2(n4168), .A(n2511), .ZN(n2512) );
  OR2_X1 U2807 ( .A1(n4199), .A2(n4470), .ZN(n2846) );
  OR2_X1 U2808 ( .A1(n4199), .A2(n4526), .ZN(n2841) );
  NAND2_X1 U2809 ( .A1(n3134), .A2(n3139), .ZN(n3140) );
  AND2_X1 U2810 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2165)
         );
  INV_X1 U2811 ( .A(n3588), .ZN(n2324) );
  AND2_X1 U2812 ( .A1(n4966), .A2(n2389), .ZN(n2166) );
  AND2_X1 U2813 ( .A1(n2304), .A2(n2782), .ZN(n2167) );
  NAND2_X1 U2814 ( .A1(n2314), .A2(n2166), .ZN(n2383) );
  OR2_X1 U2815 ( .A1(n2851), .A2(n2267), .ZN(n2168) );
  INV_X1 U2816 ( .A(n4123), .ZN(n2802) );
  INV_X1 U2817 ( .A(n2550), .ZN(n2713) );
  INV_X1 U2818 ( .A(n4122), .ZN(n2284) );
  INV_X1 U2819 ( .A(n4358), .ZN(n4362) );
  OR2_X1 U2820 ( .A1(n2371), .A2(n2439), .ZN(n2169) );
  AND2_X2 U2821 ( .A1(n2522), .A2(n2524), .ZN(n2549) );
  OR2_X1 U2822 ( .A1(n2263), .A2(n2433), .ZN(n2170) );
  INV_X1 U2823 ( .A(n2161), .ZN(n2905) );
  OR2_X1 U2824 ( .A1(n2474), .A2(n2473), .ZN(n2171) );
  AND2_X1 U2825 ( .A1(n2522), .A2(n3170), .ZN(n2550) );
  NOR2_X1 U2826 ( .A1(n2723), .A2(n4298), .ZN(n2172) );
  AND3_X1 U2827 ( .A1(n2392), .A2(n2166), .A3(n2312), .ZN(n2385) );
  XNOR2_X1 U2828 ( .A(n2517), .B(IR_REG_30__SCAN_IN), .ZN(n2522) );
  INV_X1 U2829 ( .A(n2522), .ZN(n2273) );
  NAND2_X1 U2830 ( .A1(n2349), .A2(n2709), .ZN(n4316) );
  OAI21_X1 U2831 ( .B1(n2773), .B2(n2544), .A(n2543), .ZN(n2852) );
  INV_X1 U2832 ( .A(n3467), .ZN(n2239) );
  AND2_X1 U2833 ( .A1(n2400), .A2(n2391), .ZN(n4539) );
  INV_X1 U2834 ( .A(n4539), .ZN(n2265) );
  AND3_X1 U2835 ( .A1(n2407), .A2(n2464), .A3(n2350), .ZN(n2444) );
  AND2_X1 U2836 ( .A1(n2385), .A2(n2359), .ZN(n2407) );
  NOR2_X1 U2837 ( .A1(n2802), .A2(n2291), .ZN(n2290) );
  INV_X1 U2838 ( .A(n2290), .ZN(n2287) );
  INV_X1 U2839 ( .A(n4014), .ZN(n2279) );
  NOR2_X1 U2840 ( .A1(n4621), .A2(n2504), .ZN(n2173) );
  AND2_X1 U2841 ( .A1(n3372), .A2(n2837), .ZN(n2174) );
  INV_X1 U2842 ( .A(n2289), .ZN(n2285) );
  NOR2_X1 U2843 ( .A1(n4015), .A2(n2287), .ZN(n2289) );
  AND2_X1 U2844 ( .A1(n4537), .A2(REG2_REG_5__SCAN_IN), .ZN(n2175) );
  OR2_X1 U2845 ( .A1(n2343), .A2(n2172), .ZN(n2176) );
  OR2_X1 U2846 ( .A1(n3244), .A2(n2203), .ZN(n2202) );
  AND2_X1 U2847 ( .A1(n2282), .A2(n4016), .ZN(n2177) );
  AND2_X1 U2848 ( .A1(n2883), .A2(n2880), .ZN(n2178) );
  OR2_X1 U2849 ( .A1(n2397), .A2(n2398), .ZN(n2179) );
  NOR2_X1 U2850 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2180)
         );
  NAND2_X1 U2851 ( .A1(n2893), .A2(n2239), .ZN(n2181) );
  NAND2_X1 U2852 ( .A1(n2392), .A2(n2358), .ZN(n2388) );
  NOR2_X1 U2853 ( .A1(n2442), .A2(IR_REG_22__SCAN_IN), .ZN(n2182) );
  AND2_X1 U2854 ( .A1(n2345), .A2(n2343), .ZN(n2183) );
  INV_X1 U2855 ( .A(n3581), .ZN(n3587) );
  INV_X1 U2856 ( .A(IR_REG_0__SCAN_IN), .ZN(n2267) );
  INV_X1 U2857 ( .A(IR_REG_25__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U2858 ( .A1(n4289), .A2(n4290), .ZN(n4265) );
  OR2_X1 U2859 ( .A1(n3803), .A2(n3802), .ZN(n2184) );
  INV_X1 U2860 ( .A(n3713), .ZN(n2210) );
  NAND2_X1 U2861 ( .A1(n2407), .A2(n2360), .ZN(n2371) );
  INV_X1 U2862 ( .A(n3686), .ZN(n2208) );
  INV_X1 U2863 ( .A(IR_REG_20__SCAN_IN), .ZN(n2777) );
  NAND2_X1 U2864 ( .A1(n3735), .A2(n2657), .ZN(n3779) );
  INV_X1 U2865 ( .A(n4050), .ZN(n2306) );
  OR2_X1 U2866 ( .A1(n4159), .A2(n4404), .ZN(n2185) );
  INV_X1 U2867 ( .A(n3996), .ZN(n2299) );
  OR2_X1 U2868 ( .A1(n4365), .A2(n4344), .ZN(n4319) );
  INV_X1 U2869 ( .A(n4550), .ZN(n2200) );
  INV_X1 U2870 ( .A(n2330), .ZN(n3735) );
  AND2_X1 U2871 ( .A1(n3969), .A2(n4322), .ZN(n2186) );
  NOR2_X1 U2872 ( .A1(n4231), .A2(n4212), .ZN(n2187) );
  INV_X1 U2873 ( .A(n4011), .ZN(n2294) );
  AND2_X1 U2874 ( .A1(n2789), .A2(n3990), .ZN(n2188) );
  AND2_X1 U2875 ( .A1(n3029), .A2(n3024), .ZN(n2189) );
  AND2_X1 U2876 ( .A1(n2184), .A2(n2992), .ZN(n2190) );
  XNOR2_X1 U2877 ( .A(n2456), .B(IR_REG_24__SCAN_IN), .ZN(n2815) );
  OAI21_X1 U2878 ( .B1(n2169), .B2(n2245), .A(n2241), .ZN(n2840) );
  NAND2_X1 U2879 ( .A1(n3778), .A2(n3814), .ZN(n3777) );
  NAND2_X1 U2880 ( .A1(n2226), .A2(n2230), .ZN(n3666) );
  NAND2_X1 U2881 ( .A1(n2234), .A2(n2237), .ZN(n3601) );
  INV_X1 U2882 ( .A(n3836), .ZN(n3867) );
  NAND2_X1 U2883 ( .A1(n3606), .A2(n3605), .ZN(n2191) );
  OR2_X1 U2884 ( .A1(n2260), .A2(n3725), .ZN(n2192) );
  NAND2_X1 U2885 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  INV_X1 U2886 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2201) );
  INV_X1 U2887 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2204) );
  INV_X1 U2888 ( .A(n4636), .ZN(n4657) );
  NOR2_X2 U2889 ( .A1(n3194), .A2(n3084), .ZN(n4471) );
  CLKBUF_X1 U2890 ( .A(n3881), .Z(n2193) );
  NOR3_X1 U2891 ( .A1(n3110), .A2(n4529), .A3(n4153), .ZN(n3881) );
  INV_X1 U2892 ( .A(n2193), .ZN(n3983) );
  NAND3_X1 U2893 ( .A1(n2197), .A2(n2493), .A3(n2195), .ZN(n2494) );
  INV_X1 U2894 ( .A(n2215), .ZN(n3562) );
  NAND2_X1 U2895 ( .A1(n3343), .A2(n3342), .ZN(n2218) );
  NAND2_X1 U2896 ( .A1(n2219), .A2(n2189), .ZN(n3886) );
  NAND2_X1 U2897 ( .A1(n2220), .A2(n2190), .ZN(n2997) );
  NAND2_X1 U2898 ( .A1(n2981), .A2(n2980), .ZN(n3805) );
  NAND2_X1 U2899 ( .A1(n3878), .A2(n2227), .ZN(n2223) );
  NAND2_X1 U2900 ( .A1(n2223), .A2(n2224), .ZN(n2970) );
  INV_X1 U2901 ( .A(n3875), .ZN(n2233) );
  NAND2_X1 U2902 ( .A1(n3382), .A2(n2235), .ZN(n2234) );
  NAND2_X1 U2903 ( .A1(n2248), .A2(n3975), .ZN(n3909) );
  NAND2_X1 U2904 ( .A1(n3059), .A2(n3944), .ZN(n3979) );
  INV_X1 U2905 ( .A(n2248), .ZN(n3907) );
  INV_X1 U2906 ( .A(n3944), .ZN(n2250) );
  NAND2_X1 U2907 ( .A1(n4580), .A2(n2426), .ZN(n4594) );
  NOR2_X1 U2908 ( .A1(n4689), .A2(REG2_REG_13__SCAN_IN), .ZN(n2260) );
  NAND2_X2 U2909 ( .A1(n2273), .A2(n2524), .ZN(n3257) );
  INV_X1 U2910 ( .A(n2524), .ZN(n3170) );
  OAI21_X1 U2911 ( .B1(n2803), .B2(n2287), .A(n2286), .ZN(n2292) );
  NAND2_X1 U2912 ( .A1(n2295), .A2(n2188), .ZN(n3783) );
  OAI21_X1 U2913 ( .B1(n3857), .B2(n2300), .A(n2297), .ZN(n2800) );
  INV_X1 U2914 ( .A(n2779), .ZN(n4118) );
  OAI21_X1 U2915 ( .B1(n3411), .B2(n2781), .A(n4050), .ZN(n3481) );
  NAND3_X1 U2916 ( .A1(n2310), .A2(n2407), .A3(n2464), .ZN(n2519) );
  NAND3_X1 U2917 ( .A1(n2464), .A2(n2407), .A3(n2351), .ZN(n2474) );
  INV_X1 U2918 ( .A(n3627), .ZN(n2325) );
  OAI21_X1 U2919 ( .B1(n3736), .B2(n2328), .A(n2326), .ZN(n3842) );
  NAND2_X1 U2920 ( .A1(n4117), .A2(n2657), .ZN(n2329) );
  NOR2_X1 U2921 ( .A1(n3736), .A2(n4117), .ZN(n2330) );
  NAND3_X1 U2922 ( .A1(n4255), .A2(n2334), .A3(n2185), .ZN(n2333) );
  NAND2_X1 U2923 ( .A1(n4337), .A2(n2341), .ZN(n2340) );
  NAND4_X1 U2924 ( .A1(n2407), .A2(n2464), .A3(n2350), .A4(n4918), .ZN(n2448)
         );
  NAND2_X1 U2925 ( .A1(n3649), .A2(n3648), .ZN(n3705) );
  CLKBUF_X1 U2926 ( .A(n3886), .Z(n3919) );
  AOI22_X1 U2927 ( .A1(n2850), .A2(n3009), .B1(n2852), .B2(n2849), .ZN(n2862)
         );
  NAND2_X1 U2928 ( .A1(n3311), .A2(n2852), .ZN(n4032) );
  NAND2_X1 U2929 ( .A1(n2465), .A2(n2464), .ZN(n2352) );
  NAND2_X1 U2930 ( .A1(n3105), .A2(n3087), .ZN(n3988) );
  AND2_X1 U2931 ( .A1(n2470), .A2(IR_REG_28__SCAN_IN), .ZN(n2353) );
  INV_X1 U2932 ( .A(n3421), .ZN(n2837) );
  NAND2_X1 U2933 ( .A1(n3074), .A2(n3975), .ZN(n2354) );
  OR3_X1 U2934 ( .A1(n3097), .A2(n3988), .A3(n3096), .ZN(n2355) );
  OAI211_X1 U2935 ( .C1(n4269), .C2(n2713), .A(n2736), .B(n2735), .ZN(n4418)
         );
  INV_X1 U2936 ( .A(n3781), .ZN(n2789) );
  AND2_X1 U2937 ( .A1(n2805), .A2(n4026), .ZN(n4360) );
  INV_X1 U2938 ( .A(n4360), .ZN(n3121) );
  INV_X1 U2939 ( .A(n4526), .ZN(n3139) );
  INV_X1 U2940 ( .A(n4535), .ZN(n2583) );
  INV_X1 U2941 ( .A(IR_REG_31__SCAN_IN), .ZN(n2443) );
  NOR2_X1 U2942 ( .A1(n2926), .A2(n2925), .ZN(n2357) );
  NAND2_X2 U2943 ( .A1(n3156), .A2(n4300), .ZN(n4544) );
  OR2_X1 U2944 ( .A1(n3125), .A2(n3124), .ZN(n3126) );
  OAI211_X1 U2945 ( .C1(n4301), .C2(n2713), .A(n2722), .B(n2721), .ZN(n4438)
         );
  INV_X1 U2946 ( .A(n4438), .ZN(n2723) );
  INV_X1 U2947 ( .A(IR_REG_24__SCAN_IN), .ZN(n2441) );
  AND2_X1 U2948 ( .A1(n4159), .A2(n4471), .ZN(n3124) );
  AND2_X1 U2949 ( .A1(n3701), .A2(n3676), .ZN(n4068) );
  INV_X1 U2950 ( .A(n3608), .ZN(n2928) );
  NOR2_X1 U2951 ( .A1(n2937), .A2(n3550), .ZN(n2938) );
  AND2_X1 U2952 ( .A1(n4535), .A2(REG2_REG_7__SCAN_IN), .ZN(n2412) );
  INV_X1 U2953 ( .A(n2971), .ZN(n2972) );
  NAND2_X1 U2954 ( .A1(n3606), .A2(n2938), .ZN(n2941) );
  NOR2_X1 U2955 ( .A1(n4099), .A2(n2753), .ZN(n2754) );
  INV_X1 U2956 ( .A(n2556), .ZN(n3390) );
  AND2_X1 U2957 ( .A1(n4158), .A2(n3898), .ZN(n2767) );
  NAND2_X1 U2958 ( .A1(n2997), .A2(n3831), .ZN(n3926) );
  INV_X1 U2959 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U2960 ( .A1(n4540), .A2(n2398), .ZN(n2394) );
  NOR2_X1 U2961 ( .A1(n2732), .A2(n2731), .ZN(n2739) );
  AND2_X1 U2962 ( .A1(n3463), .A2(n2590), .ZN(n2591) );
  INV_X1 U2963 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2574) );
  AND2_X1 U2964 ( .A1(n2164), .A2(DATAI_20_), .ZN(n4344) );
  INV_X1 U2965 ( .A(n2585), .ZN(n3415) );
  INV_X1 U2966 ( .A(IR_REG_29__SCAN_IN), .ZN(n2516) );
  NOR2_X1 U2967 ( .A1(n2419), .A2(n2374), .ZN(n2427) );
  NAND2_X1 U2968 ( .A1(n3297), .A2(n2873), .ZN(n3343) );
  NAND2_X1 U2969 ( .A1(n3097), .A2(n3091), .ZN(n3092) );
  OR2_X1 U2970 ( .A1(n2711), .A2(n3938), .ZN(n2719) );
  NAND2_X1 U2971 ( .A1(n2666), .A2(REG3_REG_16__SCAN_IN), .ZN(n2676) );
  OR2_X1 U2972 ( .A1(n2676), .A2(n2675), .ZN(n2685) );
  INV_X1 U2973 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2604) );
  OR2_X1 U2974 ( .A1(n2644), .A2(n2643), .ZN(n2651) );
  INV_X1 U2975 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2623) );
  INV_X1 U2976 ( .A(n3928), .ZN(n3980) );
  INV_X1 U2977 ( .A(n3257), .ZN(n2734) );
  AND4_X1 U2978 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n4459)
         );
  NAND2_X1 U2979 ( .A1(n2487), .A2(n4538), .ZN(n2488) );
  INV_X1 U2980 ( .A(n4405), .ZN(n4421) );
  AND2_X1 U2981 ( .A1(n4280), .A2(n2796), .ZN(n4305) );
  AOI21_X1 U2982 ( .B1(n4372), .B2(n2683), .A(n2682), .ZN(n3865) );
  AND4_X1 U2983 ( .A1(n2672), .A2(n2671), .A3(n2670), .A4(n2669), .ZN(n4461)
         );
  NOR2_X1 U2984 ( .A1(n2575), .A2(n2574), .ZN(n2592) );
  NAND2_X1 U2985 ( .A1(n2773), .A2(DATAI_2_), .ZN(n2529) );
  MUX2_X1 U2986 ( .A(n2602), .B(DATAI_9_), .S(n2164), .Z(n3627) );
  INV_X1 U2987 ( .A(n4463), .ZN(n4476) );
  OR2_X1 U2988 ( .A1(n2371), .A2(IR_REG_9__SCAN_IN), .ZN(n2419) );
  XNOR2_X1 U2989 ( .A(n3090), .B(n3089), .ZN(n3908) );
  NAND2_X1 U2990 ( .A1(n3320), .A2(n3319), .ZN(n3318) );
  NOR2_X1 U2991 ( .A1(n2624), .A2(n2623), .ZN(n2633) );
  NAND2_X1 U2992 ( .A1(n2745), .A2(n2744), .ZN(n4261) );
  INV_X1 U2993 ( .A(n4461), .ZN(n3817) );
  NOR2_X1 U2994 ( .A1(n4764), .A2(n2170), .ZN(n3726) );
  AND2_X1 U2995 ( .A1(n3183), .A2(n2477), .ZN(n4592) );
  AND2_X1 U2996 ( .A1(n3990), .A2(n3991), .ZN(n4117) );
  AND2_X1 U2997 ( .A1(n4064), .A2(n4063), .ZN(n4120) );
  INV_X1 U2998 ( .A(n4391), .ZN(n4318) );
  INV_X1 U2999 ( .A(n3160), .ZN(n3358) );
  INV_X1 U3000 ( .A(n3657), .ZN(n3561) );
  NAND2_X1 U3001 ( .A1(n4339), .A2(n4449), .ZN(n4676) );
  AND2_X1 U3002 ( .A1(n3351), .A2(n4149), .ZN(n4674) );
  NAND2_X1 U3003 ( .A1(n2817), .A2(n4530), .ZN(n3178) );
  AND2_X1 U3004 ( .A1(n2430), .A2(n2431), .ZN(n4689) );
  INV_X1 U3005 ( .A(U4043), .ZN(n3263) );
  INV_X1 U3006 ( .A(n3655), .ZN(n4163) );
  OR2_X1 U3007 ( .A1(n3870), .A2(n3403), .ZN(n4368) );
  NAND2_X1 U3008 ( .A1(n3134), .A2(n3633), .ZN(n3135) );
  NAND2_X1 U3009 ( .A1(n4479), .A2(n4688), .ZN(n4470) );
  NAND2_X1 U3010 ( .A1(n4683), .A2(n4479), .ZN(n4526) );
  OR2_X1 U3011 ( .A1(n2843), .A2(n3083), .ZN(n4682) );
  INV_X1 U3012 ( .A(n4654), .ZN(n4653) );
  AND2_X1 U3013 ( .A1(n2411), .A2(n2413), .ZN(n4535) );
  INV_X2 U3014 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U3015 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2364)
         );
  NAND4_X1 U3016 ( .A1(n2364), .A2(n2363), .A3(n2362), .A4(n2361), .ZN(n2439)
         );
  OR2_X1 U3017 ( .A1(n2169), .A2(IR_REG_17__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3018 ( .A1(n2368), .A2(IR_REG_31__SCAN_IN), .ZN(n2365) );
  XNOR2_X1 U3019 ( .A(n2365), .B(IR_REG_18__SCAN_IN), .ZN(n4185) );
  INV_X1 U3020 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4717) );
  NOR2_X1 U3021 ( .A1(n4185), .A2(n4717), .ZN(n2366) );
  AOI21_X1 U3022 ( .B1(n4185), .B2(n4717), .A(n2366), .ZN(n2479) );
  NAND2_X1 U3023 ( .A1(n2169), .A2(IR_REG_31__SCAN_IN), .ZN(n2367) );
  MUX2_X1 U3024 ( .A(IR_REG_31__SCAN_IN), .B(n2367), .S(IR_REG_17__SCAN_IN), 
        .Z(n2369) );
  NAND2_X1 U3025 ( .A1(n2369), .A2(n2368), .ZN(n4636) );
  NOR2_X1 U3026 ( .A1(n4657), .A2(REG2_REG_17__SCAN_IN), .ZN(n2370) );
  AOI21_X1 U3027 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4657), .A(n2370), .ZN(n4627) );
  INV_X1 U3028 ( .A(IR_REG_10__SCAN_IN), .ZN(n2373) );
  INV_X1 U3029 ( .A(IR_REG_12__SCAN_IN), .ZN(n2372) );
  NAND3_X1 U3030 ( .A1(n4745), .A2(n2373), .A3(n2372), .ZN(n2374) );
  NAND2_X1 U3031 ( .A1(n2427), .A2(n2428), .ZN(n2431) );
  NAND2_X1 U3032 ( .A1(n2375), .A2(IR_REG_31__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U3033 ( .A1(n2376), .A2(n4748), .ZN(n2435) );
  OR2_X1 U3034 ( .A1(n2376), .A2(n4748), .ZN(n2377) );
  OAI21_X1 U3035 ( .B1(n2419), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2379) );
  NAND2_X1 U3036 ( .A1(n2379), .A2(n4745), .ZN(n2380) );
  NAND2_X1 U3037 ( .A1(n2380), .A2(IR_REG_31__SCAN_IN), .ZN(n2378) );
  XNOR2_X1 U3038 ( .A(n2378), .B(IR_REG_12__SCAN_IN), .ZN(n4663) );
  OR2_X1 U3039 ( .A1(n2379), .A2(n4745), .ZN(n2381) );
  NAND2_X1 U3040 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2631), .ZN(n2424) );
  INV_X1 U3041 ( .A(n2631), .ZN(n4665) );
  INV_X1 U3042 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U3043 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2631), .B1(n4665), .B2(
        n4759), .ZN(n4574) );
  NAND2_X1 U3044 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  XNOR2_X1 U3045 ( .A(n2382), .B(IR_REG_10__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U3046 ( .A1(n2383), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  MUX2_X1 U3047 ( .A(IR_REG_31__SCAN_IN), .B(n2384), .S(IR_REG_5__SCAN_IN), 
        .Z(n2387) );
  INV_X1 U3048 ( .A(n2385), .ZN(n2386) );
  NAND2_X1 U3049 ( .A1(n2387), .A2(n2386), .ZN(n3251) );
  INV_X1 U3050 ( .A(n3251), .ZN(n4537) );
  NAND2_X1 U3051 ( .A1(n2388), .A2(IR_REG_31__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3052 ( .A1(n2390), .A2(n2389), .ZN(n2400) );
  OR2_X1 U3053 ( .A1(n2390), .A2(n2389), .ZN(n2391) );
  INV_X1 U3054 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2398) );
  INV_X1 U3055 ( .A(n4540), .ZN(n2397) );
  INV_X1 U3056 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3438) );
  XNOR2_X1 U3057 ( .A(n2482), .B(n3438), .ZN(n4174) );
  AND2_X1 U3058 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4173)
         );
  NAND2_X1 U3059 ( .A1(n4174), .A2(n4173), .ZN(n4172) );
  NAND2_X1 U3060 ( .A1(n2482), .A2(REG2_REG_1__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3061 ( .A1(n4172), .A2(n2396), .ZN(n3201) );
  AOI22_X1 U3062 ( .A1(n3211), .A2(REG2_REG_3__SCAN_IN), .B1(n4539), .B2(n2399), .ZN(n2402) );
  NAND2_X1 U3063 ( .A1(n2400), .A2(IR_REG_31__SCAN_IN), .ZN(n2401) );
  XNOR2_X1 U3064 ( .A(n2401), .B(IR_REG_4__SCAN_IN), .ZN(n4538) );
  XNOR2_X1 U3065 ( .A(n2402), .B(n4538), .ZN(n3218) );
  INV_X1 U3066 ( .A(n2402), .ZN(n2403) );
  AOI22_X1 U3067 ( .A1(n3218), .A2(REG2_REG_4__SCAN_IN), .B1(n4538), .B2(n2403), .ZN(n3249) );
  INV_X1 U3068 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3497) );
  MUX2_X1 U3069 ( .A(REG2_REG_5__SCAN_IN), .B(n3497), .S(n3251), .Z(n3248) );
  NOR2_X1 U3070 ( .A1(n3249), .A2(n3248), .ZN(n3247) );
  OR2_X1 U3071 ( .A1(n2385), .A2(n2443), .ZN(n2404) );
  XNOR2_X1 U3072 ( .A(n2404), .B(IR_REG_6__SCAN_IN), .ZN(n4536) );
  INV_X1 U3073 ( .A(n2405), .ZN(n2406) );
  INV_X1 U3074 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3453) );
  NOR2_X1 U3075 ( .A1(n2407), .A2(n2443), .ZN(n2408) );
  NAND2_X1 U3076 ( .A1(n2408), .A2(IR_REG_7__SCAN_IN), .ZN(n2411) );
  INV_X1 U3077 ( .A(n2408), .ZN(n2410) );
  INV_X1 U3078 ( .A(IR_REG_7__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3079 ( .A1(n2410), .A2(n2409), .ZN(n2413) );
  MUX2_X1 U3080 ( .A(n3453), .B(REG2_REG_7__SCAN_IN), .S(n4535), .Z(n3280) );
  NOR2_X1 U3081 ( .A1(n3279), .A2(n2412), .ZN(n2416) );
  NAND2_X1 U3082 ( .A1(n2413), .A2(IR_REG_31__SCAN_IN), .ZN(n2415) );
  INV_X1 U3083 ( .A(IR_REG_8__SCAN_IN), .ZN(n2414) );
  XNOR2_X1 U3084 ( .A(n2415), .B(n2414), .ZN(n3291) );
  XNOR2_X1 U3085 ( .A(n2416), .B(n3291), .ZN(n3288) );
  INV_X1 U3086 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2417) );
  OAI22_X1 U3087 ( .A1(n3288), .A2(n2417), .B1(n2416), .B2(n3291), .ZN(n4552)
         );
  NAND2_X1 U3088 ( .A1(n2371), .A2(IR_REG_31__SCAN_IN), .ZN(n2418) );
  MUX2_X1 U3089 ( .A(IR_REG_31__SCAN_IN), .B(n2418), .S(IR_REG_9__SCAN_IN), 
        .Z(n2420) );
  INV_X1 U3090 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3518) );
  INV_X1 U3091 ( .A(n2602), .ZN(n4669) );
  AOI22_X1 U3092 ( .A1(n2602), .A2(REG2_REG_9__SCAN_IN), .B1(n3518), .B2(n4669), .ZN(n4553) );
  NAND2_X1 U3093 ( .A1(n4552), .A2(n4553), .ZN(n4551) );
  NAND2_X1 U3094 ( .A1(n2602), .A2(REG2_REG_9__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3095 ( .A1(n4551), .A2(n2421), .ZN(n2422) );
  NAND2_X1 U3096 ( .A1(n4666), .A2(n2422), .ZN(n2423) );
  INV_X1 U3097 ( .A(n4666), .ZN(n4568) );
  XNOR2_X1 U3098 ( .A(n2422), .B(n4568), .ZN(n4560) );
  NAND2_X1 U3099 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U3100 ( .A1(n2423), .A2(n4559), .ZN(n4573) );
  NAND2_X1 U3101 ( .A1(n4574), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U3102 ( .A1(n2424), .A2(n4572), .ZN(n2425) );
  NAND2_X1 U3103 ( .A1(n4663), .A2(n2425), .ZN(n2426) );
  INV_X1 U3104 ( .A(n4663), .ZN(n4589) );
  XNOR2_X1 U3105 ( .A(n2425), .B(n4589), .ZN(n4581) );
  NAND2_X1 U3106 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4581), .ZN(n4580) );
  INV_X1 U3107 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4591) );
  OR2_X1 U3108 ( .A1(n2427), .A2(n2443), .ZN(n2429) );
  MUX2_X1 U3109 ( .A(n2429), .B(IR_REG_31__SCAN_IN), .S(n2428), .Z(n2430) );
  INV_X1 U3110 ( .A(n4689), .ZN(n4603) );
  NOR2_X1 U3111 ( .A1(n4591), .A2(n4603), .ZN(n4590) );
  NAND2_X1 U3112 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  XNOR2_X1 U3113 ( .A(n2432), .B(IR_REG_14__SCAN_IN), .ZN(n4534) );
  INV_X1 U3114 ( .A(n4534), .ZN(n3725) );
  INV_X1 U3115 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4764) );
  NOR2_X1 U3116 ( .A1(n2433), .A2(n3726), .ZN(n4606) );
  NAND2_X1 U3117 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4661), .ZN(n2434) );
  OAI21_X1 U3118 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4661), .A(n2434), .ZN(n4605) );
  NOR2_X1 U3119 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U3120 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2436) );
  XNOR2_X1 U3121 ( .A(n2436), .B(IR_REG_16__SCAN_IN), .ZN(n2673) );
  INV_X1 U3122 ( .A(n2673), .ZN(n4660) );
  NAND2_X1 U3123 ( .A1(n2437), .A2(n4660), .ZN(n2438) );
  INV_X1 U3124 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U3125 ( .A1(n4627), .A2(n4625), .ZN(n4626) );
  NAND2_X1 U3126 ( .A1(n2441), .A2(n2457), .ZN(n2442) );
  NOR2_X1 U3127 ( .A1(n2450), .A2(n2445), .ZN(n2446) );
  INV_X1 U3128 ( .A(n2819), .ZN(n4531) );
  NAND2_X1 U3129 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  INV_X1 U3130 ( .A(n2448), .ZN(n2450) );
  INV_X1 U3131 ( .A(IR_REG_26__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3132 ( .A1(n2450), .A2(n2449), .ZN(n2460) );
  INV_X1 U3133 ( .A(n2474), .ZN(n2453) );
  INV_X1 U3134 ( .A(IR_REG_22__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3135 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  NAND2_X1 U3136 ( .A1(n2454), .A2(IR_REG_31__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3137 ( .A1(n2458), .A2(n2457), .ZN(n2455) );
  XNOR2_X1 U3138 ( .A(n2458), .B(n2457), .ZN(n3101) );
  NAND2_X1 U3139 ( .A1(n3101), .A2(STATE_REG_SCAN_IN), .ZN(n4655) );
  INV_X1 U3140 ( .A(n4655), .ZN(n2459) );
  NAND2_X1 U3141 ( .A1(n2851), .A2(n2459), .ZN(n3151) );
  NOR2_X1 U3142 ( .A1(n3101), .A2(U3149), .ZN(n4150) );
  INV_X1 U3143 ( .A(n4150), .ZN(n4155) );
  NAND2_X1 U3144 ( .A1(n3151), .A2(n4155), .ZN(n2508) );
  NAND2_X1 U3145 ( .A1(n2474), .A2(IR_REG_31__SCAN_IN), .ZN(n2463) );
  XNOR2_X1 U3146 ( .A(n2463), .B(n2452), .ZN(n4149) );
  INV_X1 U3147 ( .A(n4149), .ZN(n3168) );
  NAND2_X1 U31480 ( .A1(n2352), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U31490 ( .A(n2467), .B(n2466), .ZN(n2820) );
  NAND2_X1 U3150 ( .A1(n3168), .A2(n4532), .ZN(n3084) );
  INV_X1 U3151 ( .A(n3084), .ZN(n2806) );
  NAND2_X1 U3152 ( .A1(n2806), .A2(n3101), .ZN(n2468) );
  AND2_X1 U3153 ( .A1(n2164), .A2(n2468), .ZN(n2507) );
  OAI21_X1 U3154 ( .B1(n2460), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2469) );
  MUX2_X1 U3155 ( .A(n2469), .B(IR_REG_31__SCAN_IN), .S(n2471), .Z(n2475) );
  NAND2_X1 U3156 ( .A1(n2475), .A2(n2171), .ZN(n3194) );
  INV_X1 U3157 ( .A(n3194), .ZN(n4529) );
  XNOR2_X1 U3158 ( .A(n2476), .B(IR_REG_27__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U3159 ( .A1(n4529), .A2(n3193), .ZN(n4152) );
  INV_X1 U3160 ( .A(n4152), .ZN(n2477) );
  INV_X1 U3161 ( .A(n4592), .ZN(n4624) );
  AOI211_X1 U3162 ( .C1(n2479), .C2(n2478), .A(n4184), .B(n4624), .ZN(n2515)
         );
  NOR2_X1 U3163 ( .A1(n4657), .A2(REG1_REG_17__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3164 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4661), .ZN(n2502) );
  INV_X1 U3165 ( .A(n4661), .ZN(n4614) );
  INV_X1 U3166 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U3167 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4661), .B1(n4614), .B2(
        n4699), .ZN(n4611) );
  NAND2_X1 U3168 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4689), .ZN(n2499) );
  INV_X1 U3169 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2480) );
  AOI22_X1 U3170 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4689), .B1(n4603), .B2(
        n2480), .ZN(n4600) );
  NAND2_X1 U3171 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2631), .ZN(n2496) );
  INV_X1 U3172 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U3173 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2631), .B1(n4665), .B2(
        n4697), .ZN(n4571) );
  NAND2_X1 U3174 ( .A1(n2602), .A2(REG1_REG_9__SCAN_IN), .ZN(n2493) );
  INV_X1 U3175 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2481) );
  XNOR2_X1 U3176 ( .A(n2482), .B(n2481), .ZN(n4171) );
  AND2_X1 U3177 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4170)
         );
  NAND2_X1 U3178 ( .A1(n4171), .A2(n4170), .ZN(n4169) );
  NAND2_X1 U3179 ( .A1(n2482), .A2(REG1_REG_1__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3180 ( .A1(n4169), .A2(n2483), .ZN(n3204) );
  NAND2_X1 U3181 ( .A1(n3205), .A2(n3204), .ZN(n3203) );
  NAND2_X1 U3182 ( .A1(n4540), .A2(REG1_REG_2__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3183 ( .A1(n2485), .A2(n4539), .ZN(n2486) );
  INV_X1 U3184 ( .A(n4538), .ZN(n3224) );
  XNOR2_X1 U3185 ( .A(n2487), .B(n3224), .ZN(n3220) );
  NAND2_X1 U3186 ( .A1(n3220), .A2(REG1_REG_4__SCAN_IN), .ZN(n3219) );
  XNOR2_X1 U3187 ( .A(n4537), .B(REG1_REG_5__SCAN_IN), .ZN(n3245) );
  INV_X1 U3188 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3545) );
  AOI21_X1 U3189 ( .B1(n4536), .B2(n2202), .A(n3232), .ZN(n3278) );
  NAND2_X1 U3190 ( .A1(n4535), .A2(REG1_REG_7__SCAN_IN), .ZN(n3274) );
  NOR2_X1 U3191 ( .A1(n4535), .A2(REG1_REG_7__SCAN_IN), .ZN(n3273) );
  INV_X1 U3192 ( .A(n3291), .ZN(n2489) );
  NAND2_X1 U3193 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  INV_X1 U3194 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2492) );
  AOI22_X1 U3195 ( .A1(n2602), .A2(REG1_REG_9__SCAN_IN), .B1(n2492), .B2(n4669), .ZN(n4550) );
  NAND2_X1 U3196 ( .A1(n4666), .A2(n2494), .ZN(n2495) );
  XNOR2_X1 U3197 ( .A(n2494), .B(n4568), .ZN(n4565) );
  NAND2_X1 U3198 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4565), .ZN(n4564) );
  NAND2_X1 U3199 ( .A1(n2495), .A2(n4564), .ZN(n4570) );
  NAND2_X1 U3200 ( .A1(n4663), .A2(n2497), .ZN(n2498) );
  NAND2_X1 U3201 ( .A1(n2498), .A2(n4585), .ZN(n4599) );
  NAND2_X1 U3202 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U3203 ( .A1(n2500), .A2(n4534), .ZN(n2501) );
  NAND2_X1 U3204 ( .A1(n4611), .A2(n4610), .ZN(n4609) );
  NOR2_X1 U3205 ( .A1(n2673), .A2(n2503), .ZN(n2504) );
  INV_X1 U3206 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U3207 ( .A1(n4657), .A2(n4700), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4636), .ZN(n4632) );
  NOR2_X1 U3208 ( .A1(n2173), .A2(n4632), .ZN(n4633) );
  INV_X1 U3209 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U32100 ( .A(n4185), .B(n2506), .ZN(n4179) );
  XNOR2_X1 U32110 ( .A(n4180), .B(n4179), .ZN(n2513) );
  INV_X1 U32120 ( .A(n3193), .ZN(n3181) );
  INV_X1 U32130 ( .A(n4631), .ZN(n4194) );
  NAND2_X1 U32140 ( .A1(n3183), .A2(n3194), .ZN(n4637) );
  INV_X1 U32150 ( .A(n4637), .ZN(n4168) );
  INV_X1 U32160 ( .A(n2507), .ZN(n2509) );
  INV_X1 U32170 ( .A(n4630), .ZN(n3189) );
  INV_X1 U32180 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32190 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3837) );
  OAI21_X1 U32200 ( .B1(n3189), .B2(n2510), .A(n3837), .ZN(n2511) );
  OAI21_X1 U32210 ( .B1(n2513), .B2(n4194), .A(n2512), .ZN(n2514) );
  OR2_X1 U32220 ( .A1(n2515), .A2(n2514), .ZN(U3258) );
  INV_X1 U32230 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2836) );
  MUX2_X1 U32240 ( .A(n4539), .B(DATAI_3_), .S(n2773), .Z(n3377) );
  NAND2_X1 U32250 ( .A1(n2171), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  INV_X1 U32260 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2521) );
  OR2_X1 U32270 ( .A1(n3257), .A2(n2521), .ZN(n2528) );
  INV_X1 U32280 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32290 ( .A1(n2550), .A2(n2523), .ZN(n2527) );
  NAND2_X1 U32300 ( .A1(n2608), .A2(REG1_REG_3__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32310 ( .A1(n2549), .A2(REG2_REG_3__SCAN_IN), .ZN(n2525) );
  INV_X1 U32320 ( .A(n4165), .ZN(n3424) );
  NAND2_X1 U32330 ( .A1(n3372), .A2(n3424), .ZN(n2534) );
  NAND2_X1 U32340 ( .A1(n2159), .A2(REG3_REG_2__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32350 ( .A1(n2608), .A2(REG1_REG_2__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32360 ( .A1(n2549), .A2(REG2_REG_2__SCAN_IN), .ZN(n2531) );
  INV_X1 U32370 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3362) );
  OR2_X1 U32380 ( .A1(n3257), .A2(n3362), .ZN(n2530) );
  NAND2_X1 U32390 ( .A1(n2608), .A2(REG1_REG_4__SCAN_IN), .ZN(n2541) );
  INV_X1 U32400 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U32410 ( .A(n2536), .B(REG3_REG_3__SCAN_IN), .ZN(n3431) );
  NAND2_X1 U32420 ( .A1(n2550), .A2(n3431), .ZN(n2540) );
  NAND2_X1 U32430 ( .A1(n2549), .A2(REG2_REG_4__SCAN_IN), .ZN(n2539) );
  INV_X1 U32440 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2537) );
  OR2_X1 U32450 ( .A1(n3257), .A2(n2537), .ZN(n2538) );
  NAND2_X1 U32460 ( .A1(n2542), .A2(n3421), .ZN(n4039) );
  AND2_X1 U32470 ( .A1(n3392), .A2(n2556), .ZN(n2558) );
  NAND2_X1 U32480 ( .A1(n3330), .A2(n3160), .ZN(n4033) );
  NAND2_X1 U32490 ( .A1(n3358), .A2(n3445), .ZN(n4036) );
  NAND2_X1 U32500 ( .A1(n4033), .A2(n4036), .ZN(n3143) );
  NAND2_X1 U32510 ( .A1(n2550), .A2(REG3_REG_1__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32520 ( .A1(n4029), .A2(n4032), .ZN(n2779) );
  INV_X1 U32530 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2548) );
  OR2_X1 U32540 ( .A1(n3257), .A2(n2548), .ZN(n2554) );
  NAND2_X1 U32550 ( .A1(n2608), .A2(REG1_REG_0__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32560 ( .A1(n2549), .A2(REG2_REG_0__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32570 ( .A1(n2550), .A2(REG3_REG_0__SCAN_IN), .ZN(n2551) );
  AND2_X1 U32580 ( .A1(n3313), .A2(n4167), .ZN(n3325) );
  NAND2_X1 U32590 ( .A1(n2779), .A2(n3325), .ZN(n3324) );
  NAND2_X1 U32600 ( .A1(n2852), .A2(n2850), .ZN(n2555) );
  AND2_X1 U32610 ( .A1(n3324), .A2(n2555), .ZN(n3144) );
  NAND2_X1 U32620 ( .A1(n3143), .A2(n3144), .ZN(n3142) );
  NAND2_X1 U32630 ( .A1(n3377), .A2(n4165), .ZN(n3393) );
  NAND2_X1 U32640 ( .A1(n3421), .A2(n3501), .ZN(n2559) );
  NAND2_X1 U32650 ( .A1(n2608), .A2(REG1_REG_5__SCAN_IN), .ZN(n2565) );
  AOI21_X1 U32660 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2560) );
  NOR2_X1 U32670 ( .A1(n2560), .A2(n2568), .ZN(n3379) );
  NAND2_X1 U32680 ( .A1(n2159), .A2(n3379), .ZN(n2564) );
  NAND2_X1 U32690 ( .A1(n2549), .A2(REG2_REG_5__SCAN_IN), .ZN(n2563) );
  INV_X1 U32700 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2561) );
  OR2_X1 U32710 ( .A1(n3257), .A2(n2561), .ZN(n2562) );
  INV_X1 U32720 ( .A(DATAI_5_), .ZN(n2566) );
  MUX2_X1 U32730 ( .A(n3251), .B(n2566), .S(n2773), .Z(n2585) );
  NAND2_X1 U32740 ( .A1(n3536), .A2(n2585), .ZN(n3476) );
  INV_X1 U32750 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2567) );
  OR2_X1 U32760 ( .A1(n3257), .A2(n2567), .ZN(n2573) );
  NAND2_X1 U32770 ( .A1(n2608), .A2(REG1_REG_6__SCAN_IN), .ZN(n2572) );
  OAI21_X1 U32780 ( .B1(n2568), .B2(REG3_REG_6__SCAN_IN), .A(n2575), .ZN(n3486) );
  INV_X1 U32790 ( .A(n3486), .ZN(n2569) );
  NAND2_X1 U32800 ( .A1(n2159), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U32810 ( .A1(n2549), .A2(REG2_REG_6__SCAN_IN), .ZN(n2570) );
  NAND4_X1 U32820 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n3511)
         );
  INV_X1 U32830 ( .A(n3511), .ZN(n3498) );
  MUX2_X1 U32840 ( .A(n4536), .B(DATAI_6_), .S(n2773), .Z(n3540) );
  NAND2_X1 U32850 ( .A1(n3498), .A2(n3482), .ZN(n2586) );
  AND2_X1 U32860 ( .A1(n3476), .A2(n2586), .ZN(n3456) );
  NAND2_X1 U32870 ( .A1(n2608), .A2(REG1_REG_7__SCAN_IN), .ZN(n2581) );
  AND2_X1 U32880 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  NOR2_X1 U32890 ( .A1(n2592), .A2(n2576), .ZN(n3512) );
  NAND2_X1 U32900 ( .A1(n2159), .A2(n3512), .ZN(n2580) );
  NAND2_X1 U32910 ( .A1(n2549), .A2(REG2_REG_7__SCAN_IN), .ZN(n2579) );
  INV_X1 U32920 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2577) );
  OR2_X1 U32930 ( .A1(n3257), .A2(n2577), .ZN(n2578) );
  NAND2_X1 U32940 ( .A1(n3591), .A2(n2901), .ZN(n2782) );
  NAND2_X1 U32950 ( .A1(n2782), .A2(n4053), .ZN(n3459) );
  AND2_X1 U32960 ( .A1(n3456), .A2(n3459), .ZN(n2584) );
  NAND2_X1 U32970 ( .A1(n3477), .A2(n2584), .ZN(n3464) );
  AND2_X1 U32980 ( .A1(n3540), .A2(n3511), .ZN(n2588) );
  NAND2_X1 U32990 ( .A1(n3415), .A2(n3489), .ZN(n3478) );
  INV_X1 U33000 ( .A(n3478), .ZN(n2587) );
  OAI21_X1 U33010 ( .B1(n2588), .B2(n2587), .A(n2586), .ZN(n3457) );
  INV_X1 U33020 ( .A(n3457), .ZN(n2589) );
  NAND2_X1 U33030 ( .A1(n3459), .A2(n2589), .ZN(n3463) );
  NAND2_X1 U33040 ( .A1(n2901), .A2(n4164), .ZN(n2590) );
  NAND2_X1 U33050 ( .A1(n3464), .A2(n2591), .ZN(n3584) );
  NAND2_X1 U33060 ( .A1(n2608), .A2(REG1_REG_8__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33070 ( .A1(n2592), .A2(REG3_REG_8__SCAN_IN), .ZN(n2605) );
  OR2_X1 U33080 ( .A1(n2592), .A2(REG3_REG_8__SCAN_IN), .ZN(n2593) );
  AND2_X1 U33090 ( .A1(n2605), .A2(n2593), .ZN(n4638) );
  NAND2_X1 U33100 ( .A1(n2159), .A2(n4638), .ZN(n2597) );
  NAND2_X1 U33110 ( .A1(n2549), .A2(REG2_REG_8__SCAN_IN), .ZN(n2596) );
  INV_X1 U33120 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2594) );
  OR2_X1 U33130 ( .A1(n3257), .A2(n2594), .ZN(n2595) );
  INV_X1 U33140 ( .A(DATAI_8_), .ZN(n3166) );
  MUX2_X1 U33150 ( .A(n3291), .B(n3166), .S(n2773), .Z(n3581) );
  NAND2_X1 U33160 ( .A1(n3620), .A2(n3581), .ZN(n2599) );
  NAND2_X1 U33170 ( .A1(n3584), .A2(n2599), .ZN(n2601) );
  NAND2_X1 U33180 ( .A1(n3587), .A2(n3626), .ZN(n2600) );
  INV_X1 U33190 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2603) );
  OR2_X1 U33200 ( .A1(n3257), .A2(n2603), .ZN(n2612) );
  NAND2_X1 U33210 ( .A1(n2605), .A2(n2604), .ZN(n2606) );
  NAND2_X1 U33220 ( .A1(n2615), .A2(n2606), .ZN(n3624) );
  INV_X1 U33230 ( .A(n3624), .ZN(n2607) );
  NAND2_X1 U33240 ( .A1(n2159), .A2(n2607), .ZN(n2611) );
  NAND2_X1 U33250 ( .A1(n2608), .A2(REG1_REG_9__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33260 ( .A1(n2549), .A2(REG2_REG_9__SCAN_IN), .ZN(n2609) );
  NAND4_X1 U33270 ( .A1(n2612), .A2(n2611), .A3(n2610), .A4(n2609), .ZN(n3588)
         );
  AND2_X1 U33280 ( .A1(n3627), .A2(n3588), .ZN(n2613) );
  MUX2_X1 U33290 ( .A(n4666), .B(DATAI_10_), .S(n2164), .Z(n3657) );
  INV_X1 U33300 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2614) );
  OR2_X1 U33310 ( .A1(n3257), .A2(n2614), .ZN(n2620) );
  NAND2_X1 U33320 ( .A1(n2608), .A2(REG1_REG_10__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U33330 ( .A1(n2615), .A2(n4963), .ZN(n2616) );
  AND2_X1 U33340 ( .A1(n2624), .A2(n2616), .ZN(n3611) );
  NAND2_X1 U33350 ( .A1(n2159), .A2(n3611), .ZN(n2618) );
  NAND2_X1 U33360 ( .A1(n2549), .A2(REG2_REG_10__SCAN_IN), .ZN(n2617) );
  NAND4_X1 U33370 ( .A1(n2620), .A2(n2619), .A3(n2618), .A4(n2617), .ZN(n3652)
         );
  NOR2_X1 U33380 ( .A1(n3657), .A2(n3652), .ZN(n2622) );
  NAND2_X1 U33390 ( .A1(n3657), .A2(n3652), .ZN(n2621) );
  AND2_X1 U33400 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  OR2_X1 U33410 ( .A1(n2625), .A2(n2633), .ZN(n3647) );
  INV_X1 U33420 ( .A(n3647), .ZN(n2626) );
  NAND2_X1 U33430 ( .A1(n2159), .A2(n2626), .ZN(n2630) );
  NAND2_X1 U33440 ( .A1(n2608), .A2(REG1_REG_11__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U33450 ( .A1(n2549), .A2(REG2_REG_11__SCAN_IN), .ZN(n2628) );
  INV_X1 U33460 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3695) );
  OR2_X1 U33470 ( .A1(n3257), .A2(n3695), .ZN(n2627) );
  MUX2_X1 U33480 ( .A(n2631), .B(DATAI_11_), .S(n2164), .Z(n3642) );
  NAND2_X1 U33490 ( .A1(n3655), .A2(n3642), .ZN(n4064) );
  NAND2_X1 U33500 ( .A1(n3648), .A2(n4163), .ZN(n4063) );
  NAND2_X1 U33510 ( .A1(n3655), .A2(n3648), .ZN(n2632) );
  NAND2_X1 U33520 ( .A1(n3639), .A2(n2632), .ZN(n3700) );
  MUX2_X1 U3353 ( .A(n4663), .B(DATAI_12_), .S(n2164), .Z(n3713) );
  INV_X1 U33540 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3762) );
  OR2_X1 U3355 ( .A1(n3257), .A2(n3762), .ZN(n2638) );
  NAND2_X1 U3356 ( .A1(n2608), .A2(REG1_REG_12__SCAN_IN), .ZN(n2637) );
  OR2_X1 U3357 ( .A1(n2633), .A2(REG3_REG_12__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3358 ( .A1(n2633), .A2(REG3_REG_12__SCAN_IN), .ZN(n2644) );
  AND2_X1 U3359 ( .A1(n2634), .A2(n2644), .ZN(n3708) );
  NAND2_X1 U3360 ( .A1(n2159), .A2(n3708), .ZN(n2636) );
  NAND2_X1 U3361 ( .A1(n2549), .A2(REG2_REG_12__SCAN_IN), .ZN(n2635) );
  NAND4_X1 U3362 ( .A1(n2638), .A2(n2637), .A3(n2636), .A4(n2635), .ZN(n4162)
         );
  NAND2_X1 U3363 ( .A1(n3713), .A2(n4162), .ZN(n2639) );
  NAND2_X1 U3364 ( .A1(n3700), .A2(n2639), .ZN(n2641) );
  INV_X1 U3365 ( .A(n4162), .ZN(n3879) );
  NAND2_X1 U3366 ( .A1(n3879), .A2(n2210), .ZN(n2640) );
  MUX2_X1 U3367 ( .A(n4689), .B(DATAI_13_), .S(n2164), .Z(n3686) );
  INV_X1 U3368 ( .A(REG0_REG_13__SCAN_IN), .ZN(n2642) );
  OR2_X1 U3369 ( .A1(n3257), .A2(n2642), .ZN(n2649) );
  NAND2_X1 U3370 ( .A1(n2608), .A2(REG1_REG_13__SCAN_IN), .ZN(n2648) );
  INV_X1 U3371 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U3372 ( .A1(n2644), .A2(n2643), .ZN(n2645) );
  AND2_X1 U3373 ( .A1(n2651), .A2(n2645), .ZN(n3882) );
  NAND2_X1 U3374 ( .A1(n2159), .A2(n3882), .ZN(n2647) );
  NAND2_X1 U3375 ( .A1(n2549), .A2(REG2_REG_13__SCAN_IN), .ZN(n2646) );
  NAND4_X1 U3376 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n4161)
         );
  NOR2_X1 U3377 ( .A1(n3686), .A2(n4161), .ZN(n2650) );
  OAI22_X1 U3378 ( .A1(n3685), .A2(n2650), .B1(n3748), .B2(n2208), .ZN(n3736)
         );
  NAND2_X1 U3379 ( .A1(n2608), .A2(REG1_REG_14__SCAN_IN), .ZN(n2656) );
  INV_X1 U3380 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4694) );
  AND2_X1 U3381 ( .A1(n2651), .A2(n4694), .ZN(n2652) );
  NOR2_X1 U3382 ( .A1(n2658), .A2(n2652), .ZN(n3745) );
  NAND2_X1 U3383 ( .A1(n2159), .A2(n3745), .ZN(n2655) );
  NAND2_X1 U3384 ( .A1(n2549), .A2(REG2_REG_14__SCAN_IN), .ZN(n2654) );
  INV_X1 U3385 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4746) );
  OR2_X1 U3386 ( .A1(n3257), .A2(n4746), .ZN(n2653) );
  MUX2_X1 U3387 ( .A(n4534), .B(DATAI_14_), .S(n2164), .Z(n3744) );
  NAND2_X1 U3388 ( .A1(n3815), .A2(n3744), .ZN(n3990) );
  INV_X1 U3389 ( .A(n3744), .ZN(n3734) );
  INV_X1 U3390 ( .A(n3815), .ZN(n4160) );
  NAND2_X1 U3391 ( .A1(n3734), .A2(n4160), .ZN(n3991) );
  NAND2_X1 U3392 ( .A1(n3815), .A2(n3734), .ZN(n2657) );
  MUX2_X1 U3393 ( .A(n4661), .B(DATAI_15_), .S(n2164), .Z(n3792) );
  INV_X1 U3394 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3787) );
  OR2_X1 U3395 ( .A1(n3257), .A2(n3787), .ZN(n2663) );
  NAND2_X1 U3396 ( .A1(n2608), .A2(REG1_REG_15__SCAN_IN), .ZN(n2662) );
  NOR2_X1 U3397 ( .A1(n2658), .A2(REG3_REG_15__SCAN_IN), .ZN(n2659) );
  OR2_X1 U3398 ( .A1(n2666), .A2(n2659), .ZN(n3820) );
  INV_X1 U3399 ( .A(n3820), .ZN(n3793) );
  NAND2_X1 U3400 ( .A1(n2159), .A2(n3793), .ZN(n2661) );
  NAND2_X1 U3401 ( .A1(n2549), .A2(REG2_REG_15__SCAN_IN), .ZN(n2660) );
  NAND4_X1 U3402 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n4472)
         );
  NAND2_X1 U3403 ( .A1(n3792), .A2(n4472), .ZN(n2664) );
  INV_X1 U3404 ( .A(n4472), .ZN(n3851) );
  NAND2_X1 U3405 ( .A1(n3851), .A2(n3814), .ZN(n2665) );
  NAND2_X1 U3406 ( .A1(n2608), .A2(REG1_REG_16__SCAN_IN), .ZN(n2672) );
  OR2_X1 U3407 ( .A1(n2666), .A2(REG3_REG_16__SCAN_IN), .ZN(n2667) );
  AND2_X1 U3408 ( .A1(n2676), .A2(n2667), .ZN(n3848) );
  NAND2_X1 U3409 ( .A1(n2159), .A2(n3848), .ZN(n2671) );
  NAND2_X1 U3410 ( .A1(n2549), .A2(REG2_REG_16__SCAN_IN), .ZN(n2670) );
  INV_X1 U3411 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2668) );
  OR2_X1 U3412 ( .A1(n3257), .A2(n2668), .ZN(n2669) );
  MUX2_X1 U3413 ( .A(n2673), .B(DATAI_16_), .S(n2164), .Z(n3847) );
  NAND2_X1 U3414 ( .A1(n4461), .A2(n3847), .ZN(n4077) );
  INV_X1 U3415 ( .A(n3847), .ZN(n4477) );
  NAND2_X1 U3416 ( .A1(n4477), .A2(n3817), .ZN(n4074) );
  NAND2_X1 U3417 ( .A1(n3847), .A2(n3817), .ZN(n2674) );
  INV_X1 U3418 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4524) );
  OR2_X1 U3419 ( .A1(n3257), .A2(n4524), .ZN(n2681) );
  NAND2_X1 U3420 ( .A1(n2608), .A2(REG1_REG_17__SCAN_IN), .ZN(n2680) );
  INV_X1 U3421 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3422 ( .A1(n2676), .A2(n2675), .ZN(n2677) );
  AND2_X1 U3423 ( .A1(n2685), .A2(n2677), .ZN(n4380) );
  NAND2_X1 U3424 ( .A1(n2159), .A2(n4380), .ZN(n2679) );
  NAND2_X1 U3425 ( .A1(n2549), .A2(REG2_REG_17__SCAN_IN), .ZN(n2678) );
  NAND4_X1 U3426 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n4473)
         );
  INV_X1 U3427 ( .A(n4473), .ZN(n2791) );
  MUX2_X1 U3428 ( .A(n4657), .B(DATAI_17_), .S(n2164), .Z(n4464) );
  INV_X1 U3429 ( .A(n4464), .ZN(n4375) );
  NAND2_X1 U3430 ( .A1(n2791), .A2(n4375), .ZN(n2683) );
  AND2_X1 U3431 ( .A1(n4464), .A2(n4473), .ZN(n2682) );
  NAND2_X1 U3432 ( .A1(n2608), .A2(REG1_REG_18__SCAN_IN), .ZN(n2691) );
  INV_X1 U3433 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2684) );
  AND2_X1 U3434 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  NOR2_X1 U3435 ( .A1(n2694), .A2(n2686), .ZN(n3868) );
  NAND2_X1 U3436 ( .A1(n2159), .A2(n3868), .ZN(n2690) );
  NAND2_X1 U3437 ( .A1(n2549), .A2(REG2_REG_18__SCAN_IN), .ZN(n2689) );
  INV_X1 U3438 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3439 ( .A1(n3257), .A2(n2687), .ZN(n2688) );
  MUX2_X1 U3440 ( .A(n4185), .B(DATAI_18_), .S(n2164), .Z(n3836) );
  NAND2_X1 U3441 ( .A1(n4459), .A2(n3836), .ZN(n4351) );
  INV_X1 U3442 ( .A(n4459), .ZN(n4377) );
  NAND2_X1 U3443 ( .A1(n3867), .A2(n4377), .ZN(n4352) );
  NAND2_X1 U3444 ( .A1(n4351), .A2(n4352), .ZN(n3864) );
  NAND2_X1 U3445 ( .A1(n3865), .A2(n3864), .ZN(n3863) );
  NAND2_X1 U3446 ( .A1(n4459), .A2(n3867), .ZN(n2692) );
  MUX2_X1 U3447 ( .A(n4533), .B(DATAI_19_), .S(n2164), .Z(n4358) );
  INV_X1 U3448 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4519) );
  OR2_X1 U3449 ( .A1(n3257), .A2(n4519), .ZN(n2699) );
  NAND2_X1 U3450 ( .A1(n2608), .A2(REG1_REG_19__SCAN_IN), .ZN(n2698) );
  NOR2_X1 U3451 ( .A1(n2694), .A2(REG3_REG_19__SCAN_IN), .ZN(n2695) );
  NOR2_X1 U3452 ( .A1(n2703), .A2(n2695), .ZN(n4366) );
  NAND2_X1 U3453 ( .A1(n2159), .A2(n4366), .ZN(n2697) );
  NAND2_X1 U3454 ( .A1(n2549), .A2(REG2_REG_19__SCAN_IN), .ZN(n2696) );
  NAND4_X1 U3455 ( .A1(n2699), .A2(n2698), .A3(n2697), .A4(n2696), .ZN(n3859)
         );
  NAND2_X1 U3456 ( .A1(n4358), .A2(n3859), .ZN(n2700) );
  NAND2_X1 U3457 ( .A1(n4350), .A2(n2700), .ZN(n2702) );
  INV_X1 U34580 ( .A(n3859), .ZN(n4336) );
  NAND2_X1 U34590 ( .A1(n4336), .A2(n4362), .ZN(n2701) );
  NAND2_X1 U3460 ( .A1(n2702), .A2(n2701), .ZN(n4337) );
  INV_X1 U3461 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4886) );
  OR2_X1 U3462 ( .A1(n3257), .A2(n4886), .ZN(n2708) );
  NAND2_X1 U3463 ( .A1(n2608), .A2(REG1_REG_20__SCAN_IN), .ZN(n2707) );
  OR2_X1 U3464 ( .A1(n2703), .A2(REG3_REG_20__SCAN_IN), .ZN(n2704) );
  AND2_X1 U3465 ( .A1(n2711), .A2(n2704), .ZN(n4343) );
  NAND2_X1 U3466 ( .A1(n2159), .A2(n4343), .ZN(n2706) );
  NAND2_X1 U34670 ( .A1(n2549), .A2(REG2_REG_20__SCAN_IN), .ZN(n2705) );
  NAND4_X1 U3468 ( .A1(n2708), .A2(n2707), .A3(n2706), .A4(n2705), .ZN(n4103)
         );
  NOR2_X1 U34690 ( .A1(n4103), .A2(n4344), .ZN(n2710) );
  NAND2_X1 U3470 ( .A1(n4103), .A2(n4344), .ZN(n2709) );
  INV_X1 U34710 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4514) );
  OR2_X1 U3472 ( .A1(n3257), .A2(n4514), .ZN(n2717) );
  INV_X1 U34730 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U3474 ( .A1(n2711), .A2(n3938), .ZN(n2712) );
  AND2_X1 U34750 ( .A1(n2719), .A2(n2712), .ZN(n4324) );
  NAND2_X1 U3476 ( .A1(n4324), .A2(n2159), .ZN(n2716) );
  NAND2_X1 U34770 ( .A1(n2608), .A2(REG1_REG_21__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3478 ( .A1(n2549), .A2(REG2_REG_21__SCAN_IN), .ZN(n2714) );
  NAND4_X1 U34790 ( .A1(n2717), .A2(n2716), .A3(n2715), .A4(n2714), .ZN(n4334)
         );
  NAND2_X1 U3480 ( .A1(n2164), .A2(DATAI_21_), .ZN(n4322) );
  AND2_X1 U34810 ( .A1(n4334), .A2(n4437), .ZN(n2718) );
  INV_X1 U3482 ( .A(n4334), .ZN(n3969) );
  INV_X1 U34830 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U3484 ( .A1(n2719), .A2(n4728), .ZN(n2720) );
  NAND2_X1 U34850 ( .A1(n2732), .A2(n2720), .ZN(n4301) );
  AOI22_X1 U3486 ( .A1(n2734), .A2(REG0_REG_22__SCAN_IN), .B1(n2549), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U34870 ( .A1(n2608), .A2(REG1_REG_22__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3488 ( .A1(n2164), .A2(DATAI_22_), .ZN(n4298) );
  OR2_X1 U34890 ( .A1(n4438), .A2(n4298), .ZN(n4280) );
  NAND2_X1 U3490 ( .A1(n4438), .A2(n4298), .ZN(n2796) );
  INV_X1 U34910 ( .A(n4298), .ZN(n4308) );
  XNOR2_X1 U3492 ( .A(n2732), .B(REG3_REG_23__SCAN_IN), .ZN(n4291) );
  NAND2_X1 U34930 ( .A1(n4291), .A2(n2159), .ZN(n2728) );
  INV_X1 U3494 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U34950 ( .A1(n2608), .A2(REG1_REG_23__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3496 ( .A1(n2549), .A2(REG2_REG_23__SCAN_IN), .ZN(n2724) );
  OAI211_X1 U34970 ( .C1(n3257), .C2(n4506), .A(n2725), .B(n2724), .ZN(n2726)
         );
  INV_X1 U3498 ( .A(n2726), .ZN(n2727) );
  NAND2_X1 U34990 ( .A1(n2164), .A2(DATAI_23_), .ZN(n4290) );
  INV_X1 U3500 ( .A(n4290), .ZN(n4285) );
  NOR2_X1 U35010 ( .A1(n4307), .A2(n4285), .ZN(n2729) );
  OAI22_X1 U3502 ( .A1(n4275), .A2(n2729), .B1(n3956), .B2(n4290), .ZN(n4255)
         );
  INV_X1 U35030 ( .A(n2732), .ZN(n2730) );
  AOI21_X1 U3504 ( .B1(n2730), .B2(REG3_REG_23__SCAN_IN), .A(
        REG3_REG_24__SCAN_IN), .ZN(n2733) );
  NAND2_X1 U35050 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .ZN(
        n2731) );
  OR2_X1 U35060 ( .A1(n2733), .A2(n2739), .ZN(n4269) );
  AOI22_X1 U35070 ( .A1(n2734), .A2(REG0_REG_24__SCAN_IN), .B1(n2608), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U35080 ( .A1(n2549), .A2(REG2_REG_24__SCAN_IN), .ZN(n2735) );
  INV_X1 U35090 ( .A(n4418), .ZN(n4288) );
  NAND2_X1 U35100 ( .A1(n2164), .A2(DATAI_24_), .ZN(n4267) );
  NOR2_X1 U35110 ( .A1(n4288), .A2(n4267), .ZN(n2738) );
  INV_X1 U35120 ( .A(n4267), .ZN(n3042) );
  OR2_X1 U35130 ( .A1(n2739), .A2(REG3_REG_25__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U35140 ( .A1(n2739), .A2(REG3_REG_25__SCAN_IN), .ZN(n2746) );
  AND2_X1 U35150 ( .A1(n2740), .A2(n2746), .ZN(n4248) );
  NAND2_X1 U35160 ( .A1(n4248), .A2(n2159), .ZN(n2745) );
  INV_X1 U35170 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4499) );
  NAND2_X1 U35180 ( .A1(n2608), .A2(REG1_REG_25__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U35190 ( .A1(n2549), .A2(REG2_REG_25__SCAN_IN), .ZN(n2741) );
  OAI211_X1 U35200 ( .C1(n4499), .C2(n3257), .A(n2742), .B(n2741), .ZN(n2743)
         );
  INV_X1 U35210 ( .A(n2743), .ZN(n2744) );
  NAND2_X1 U35220 ( .A1(n2164), .A2(DATAI_25_), .ZN(n4246) );
  NOR2_X1 U35230 ( .A1(n4261), .A2(n4417), .ZN(n4222) );
  INV_X1 U35240 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3982) );
  NAND2_X1 U35250 ( .A1(n2746), .A2(n3982), .ZN(n2747) );
  NAND2_X1 U35260 ( .A1(n4236), .A2(n2159), .ZN(n2752) );
  INV_X1 U35270 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U35280 ( .A1(n2608), .A2(REG1_REG_26__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U35290 ( .A1(n2549), .A2(REG2_REG_26__SCAN_IN), .ZN(n2748) );
  OAI211_X1 U35300 ( .C1(n3257), .C2(n4901), .A(n2749), .B(n2748), .ZN(n2750)
         );
  INV_X1 U35310 ( .A(n2750), .ZN(n2751) );
  NAND2_X1 U35320 ( .A1(n2164), .A2(DATAI_26_), .ZN(n4234) );
  AND2_X1 U35330 ( .A1(n4405), .A2(n4228), .ZN(n4099) );
  NAND2_X1 U35340 ( .A1(n4421), .A2(n4234), .ZN(n4100) );
  INV_X1 U35350 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3910) );
  AND2_X1 U35360 ( .A1(n2755), .A2(n3910), .ZN(n2756) );
  INV_X1 U35370 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U35380 ( .A1(n2608), .A2(REG1_REG_27__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U35390 ( .A1(n2549), .A2(REG2_REG_27__SCAN_IN), .ZN(n2757) );
  OAI211_X1 U35400 ( .C1(n3257), .C2(n4492), .A(n2758), .B(n2757), .ZN(n2759)
         );
  INV_X1 U35410 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U35420 ( .A1(n2164), .A2(DATAI_27_), .ZN(n4212) );
  INV_X1 U35430 ( .A(n4212), .ZN(n4404) );
  INV_X1 U35440 ( .A(n4159), .ZN(n4231) );
  NOR2_X1 U35450 ( .A1(n2761), .A2(REG3_REG_28__SCAN_IN), .ZN(n2762) );
  INV_X1 U35460 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U35470 ( .A1(n2549), .A2(REG2_REG_28__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U35480 ( .A1(n2608), .A2(REG1_REG_28__SCAN_IN), .ZN(n2763) );
  OAI211_X1 U35490 ( .C1(n3257), .C2(n4900), .A(n2764), .B(n2763), .ZN(n2765)
         );
  INV_X1 U35500 ( .A(n2765), .ZN(n2766) );
  NAND2_X1 U35510 ( .A1(n2164), .A2(DATAI_28_), .ZN(n3131) );
  OR2_X1 U35520 ( .A1(n4158), .A2(n3131), .ZN(n4014) );
  NAND2_X1 U35530 ( .A1(n4158), .A2(n3131), .ZN(n4016) );
  NAND2_X1 U35540 ( .A1(n4014), .A2(n4016), .ZN(n4098) );
  INV_X1 U35550 ( .A(n3131), .ZN(n3898) );
  NAND2_X1 U35560 ( .A1(n4197), .A2(n2159), .ZN(n2772) );
  NAND2_X1 U35570 ( .A1(n2549), .A2(REG2_REG_29__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U35580 ( .A1(n2608), .A2(REG1_REG_29__SCAN_IN), .ZN(n2768) );
  OAI211_X1 U35590 ( .C1(n3257), .C2(n2836), .A(n2769), .B(n2768), .ZN(n2770)
         );
  INV_X1 U35600 ( .A(n2770), .ZN(n2771) );
  NAND2_X1 U35610 ( .A1(n2772), .A2(n2771), .ZN(n3899) );
  NAND2_X1 U35620 ( .A1(n2164), .A2(DATAI_29_), .ZN(n2839) );
  NOR2_X1 U35630 ( .A1(n3899), .A2(n2839), .ZN(n4004) );
  NAND2_X1 U35640 ( .A1(n3899), .A2(n2839), .ZN(n4017) );
  INV_X1 U35650 ( .A(n4017), .ZN(n4013) );
  XNOR2_X1 U35660 ( .A(n2774), .B(n4096), .ZN(n4196) );
  INV_X1 U35670 ( .A(IR_REG_19__SCAN_IN), .ZN(n2775) );
  XNOR2_X1 U35680 ( .A(n3158), .B(n3168), .ZN(n2778) );
  INV_X1 U35690 ( .A(n4533), .ZN(n4190) );
  NAND2_X1 U35700 ( .A1(n2778), .A2(n4190), .ZN(n4339) );
  AND2_X1 U35710 ( .A1(n2840), .A2(n4533), .ZN(n3351) );
  INV_X1 U35720 ( .A(n4674), .ZN(n4449) );
  AND2_X1 U35730 ( .A1(n3313), .A2(n3331), .ZN(n4031) );
  NAND2_X1 U35740 ( .A1(n4118), .A2(n4031), .ZN(n3326) );
  NAND2_X1 U35750 ( .A1(n3326), .A2(n4032), .ZN(n3146) );
  INV_X1 U35760 ( .A(n3143), .ZN(n4119) );
  NAND2_X1 U35770 ( .A1(n3146), .A2(n4119), .ZN(n3145) );
  NAND2_X1 U35780 ( .A1(n3145), .A2(n4033), .ZN(n3368) );
  NAND2_X1 U35790 ( .A1(n3424), .A2(n3377), .ZN(n4038) );
  NAND2_X1 U35800 ( .A1(n3372), .A2(n4165), .ZN(n4035) );
  NAND2_X1 U35810 ( .A1(n3368), .A2(n4116), .ZN(n3367) );
  NAND2_X1 U3582 ( .A1(n3367), .A2(n4038), .ZN(n3391) );
  INV_X1 U3583 ( .A(n4039), .ZN(n2780) );
  NAND2_X1 U3584 ( .A1(n2585), .A2(n3489), .ZN(n4041) );
  INV_X1 U3585 ( .A(n4041), .ZN(n2781) );
  NAND2_X1 U3586 ( .A1(n3536), .A2(n3415), .ZN(n4050) );
  NAND2_X1 U3587 ( .A1(n3482), .A2(n3511), .ZN(n4051) );
  NAND2_X1 U3588 ( .A1(n3498), .A2(n3540), .ZN(n4044) );
  NAND2_X1 U3589 ( .A1(n2783), .A2(n4053), .ZN(n3586) );
  NAND2_X1 U3590 ( .A1(n3620), .A2(n3587), .ZN(n4047) );
  NAND2_X1 U3591 ( .A1(n3586), .A2(n4047), .ZN(n2784) );
  NAND2_X1 U3592 ( .A1(n3581), .A2(n3626), .ZN(n4052) );
  NAND2_X1 U3593 ( .A1(n2784), .A2(n4052), .ZN(n3516) );
  NAND2_X1 U3594 ( .A1(n2325), .A2(n3588), .ZN(n4060) );
  INV_X1 U3595 ( .A(n4060), .ZN(n2785) );
  NAND2_X1 U3596 ( .A1(n2324), .A2(n3627), .ZN(n4048) );
  NAND2_X1 U3597 ( .A1(n3561), .A2(n3652), .ZN(n4062) );
  NAND2_X1 U3598 ( .A1(n3558), .A2(n4062), .ZN(n2786) );
  INV_X1 U3599 ( .A(n3652), .ZN(n3691) );
  NAND2_X1 U3600 ( .A1(n3691), .A2(n3657), .ZN(n4057) );
  NAND2_X1 U3601 ( .A1(n2786), .A2(n4057), .ZN(n3643) );
  NAND2_X1 U3602 ( .A1(n3643), .A2(n4063), .ZN(n2787) );
  NAND2_X1 U3603 ( .A1(n2787), .A2(n4064), .ZN(n3675) );
  NAND2_X1 U3604 ( .A1(n2210), .A2(n4162), .ZN(n3701) );
  NAND2_X1 U3605 ( .A1(n2208), .A2(n4161), .ZN(n3676) );
  NAND2_X1 U3606 ( .A1(n3675), .A2(n4068), .ZN(n2788) );
  AND2_X1 U3607 ( .A1(n3713), .A2(n3879), .ZN(n3702) );
  AND2_X1 U3608 ( .A1(n3686), .A2(n3748), .ZN(n3677) );
  AOI21_X1 U3609 ( .B1(n4068), .B2(n3702), .A(n3677), .ZN(n4065) );
  NAND2_X1 U3610 ( .A1(n2788), .A2(n4065), .ZN(n3732) );
  NAND2_X1 U3611 ( .A1(n3851), .A2(n3792), .ZN(n3993) );
  NAND2_X1 U3612 ( .A1(n3814), .A2(n4472), .ZN(n3992) );
  NAND2_X1 U3613 ( .A1(n3993), .A2(n3992), .ZN(n3781) );
  NAND2_X1 U3614 ( .A1(n3783), .A2(n3992), .ZN(n3853) );
  NAND2_X1 U3615 ( .A1(n3853), .A2(n4131), .ZN(n3852) );
  NAND2_X1 U3616 ( .A1(n3852), .A2(n4074), .ZN(n3857) );
  NAND2_X1 U3617 ( .A1(n4362), .A2(n3859), .ZN(n2790) );
  AND2_X1 U3618 ( .A1(n4352), .A2(n2790), .ZN(n2794) );
  NAND2_X1 U3619 ( .A1(n4375), .A2(n4473), .ZN(n4104) );
  NAND2_X1 U3620 ( .A1(n2794), .A2(n4104), .ZN(n4076) );
  NAND2_X1 U3621 ( .A1(n2791), .A2(n4464), .ZN(n4105) );
  NAND2_X1 U3622 ( .A1(n4351), .A2(n4105), .ZN(n2793) );
  NOR2_X1 U3623 ( .A1(n4362), .A2(n3859), .ZN(n2792) );
  AOI21_X1 U3624 ( .B1(n2794), .B2(n2793), .A(n2792), .ZN(n4331) );
  INV_X1 U3625 ( .A(n4103), .ZN(n4441) );
  NAND2_X1 U3626 ( .A1(n4441), .A2(n4344), .ZN(n2795) );
  AND2_X1 U3627 ( .A1(n4331), .A2(n2795), .ZN(n3996) );
  INV_X1 U3628 ( .A(n4344), .ZN(n3970) );
  NAND2_X1 U3629 ( .A1(n4103), .A2(n3970), .ZN(n4079) );
  NAND2_X1 U3630 ( .A1(n3969), .A2(n4437), .ZN(n4278) );
  AND2_X1 U3631 ( .A1(n4280), .A2(n4278), .ZN(n4083) );
  NAND2_X1 U3632 ( .A1(n4307), .A2(n4290), .ZN(n4102) );
  NAND2_X1 U3633 ( .A1(n4102), .A2(n2796), .ZN(n4081) );
  INV_X1 U3634 ( .A(n4081), .ZN(n2798) );
  AND2_X1 U3635 ( .A1(n4334), .A2(n4322), .ZN(n4277) );
  NAND2_X1 U3636 ( .A1(n4280), .A2(n4277), .ZN(n2797) );
  NAND2_X1 U3637 ( .A1(n2798), .A2(n2797), .ZN(n3999) );
  INV_X1 U3638 ( .A(n3999), .ZN(n2799) );
  NAND2_X1 U3639 ( .A1(n2800), .A2(n2799), .ZN(n4257) );
  NAND2_X1 U3640 ( .A1(n3956), .A2(n4285), .ZN(n4256) );
  OR2_X1 U3641 ( .A1(n4418), .A2(n4267), .ZN(n4108) );
  NAND2_X1 U3642 ( .A1(n4257), .A2(n4084), .ZN(n2801) );
  NAND2_X1 U3643 ( .A1(n4418), .A2(n4267), .ZN(n4109) );
  NAND2_X1 U3644 ( .A1(n2801), .A2(n4109), .ZN(n4241) );
  INV_X1 U3645 ( .A(n4241), .ZN(n2803) );
  NAND2_X1 U3646 ( .A1(n4261), .A2(n4246), .ZN(n4122) );
  NAND2_X1 U3647 ( .A1(n4221), .A2(n4417), .ZN(n4123) );
  NAND2_X1 U3648 ( .A1(n4421), .A2(n4228), .ZN(n4005) );
  AND2_X1 U3649 ( .A1(n4405), .A2(n4234), .ZN(n4011) );
  XNOR2_X1 U3650 ( .A(n4159), .B(n4404), .ZN(n4208) );
  OR2_X1 U3651 ( .A1(n4159), .A2(n4212), .ZN(n4006) );
  INV_X1 U3652 ( .A(n4006), .ZN(n4015) );
  INV_X1 U3653 ( .A(n4016), .ZN(n4012) );
  XNOR2_X1 U3654 ( .A(n2804), .B(n4096), .ZN(n2814) );
  NAND2_X1 U3655 ( .A1(n3168), .A2(n4533), .ZN(n2805) );
  INV_X1 U3656 ( .A(n2840), .ZN(n4143) );
  NAND2_X1 U3657 ( .A1(n4143), .A2(n4532), .ZN(n4026) );
  NAND2_X1 U3658 ( .A1(n3194), .A2(n2806), .ZN(n4458) );
  AND2_X1 U3659 ( .A1(n3193), .A2(B_REG_SCAN_IN), .ZN(n2807) );
  NOR2_X1 U3660 ( .A1(n4458), .A2(n2807), .ZN(n4393) );
  INV_X1 U3661 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U3662 ( .A1(n2549), .A2(REG2_REG_30__SCAN_IN), .ZN(n2809) );
  NAND2_X1 U3663 ( .A1(n2608), .A2(REG1_REG_30__SCAN_IN), .ZN(n2808) );
  OAI211_X1 U3664 ( .C1(n3257), .C2(n2810), .A(n2809), .B(n2808), .ZN(n4157)
         );
  INV_X1 U3665 ( .A(n2839), .ZN(n2811) );
  AOI22_X1 U3666 ( .A1(n4393), .A2(n4157), .B1(n2811), .B2(n4463), .ZN(n2813)
         );
  NAND2_X1 U3667 ( .A1(n4158), .A2(n4471), .ZN(n2812) );
  OAI211_X1 U3668 ( .C1(n2814), .C2(n4360), .A(n2813), .B(n2812), .ZN(n4201)
         );
  AOI21_X1 U3669 ( .B1(n4196), .B2(n4676), .A(n4201), .ZN(n2844) );
  NAND2_X1 U3670 ( .A1(n2819), .A2(B_REG_SCAN_IN), .ZN(n2816) );
  MUX2_X1 U3671 ( .A(n2816), .B(B_REG_SCAN_IN), .S(n2815), .Z(n2817) );
  INV_X1 U3672 ( .A(D_REG_1__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U3673 ( .A1(n2831), .A2(n3180), .ZN(n3152) );
  INV_X1 U3674 ( .A(n4530), .ZN(n2818) );
  NAND2_X1 U3675 ( .A1(n2819), .A2(n2818), .ZN(n3081) );
  NAND2_X1 U3676 ( .A1(n3152), .A2(n3081), .ZN(n2835) );
  NAND2_X1 U3677 ( .A1(n4674), .A2(n2820), .ZN(n3107) );
  AND2_X1 U3678 ( .A1(n2840), .A2(n4190), .ZN(n2821) );
  OR2_X1 U3679 ( .A1(n3084), .A2(n2821), .ZN(n3099) );
  NAND2_X1 U3680 ( .A1(n3107), .A2(n3099), .ZN(n2822) );
  NOR2_X1 U3681 ( .A1(n3151), .A2(n2822), .ZN(n2834) );
  NOR4_X1 U3682 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2826) );
  NOR4_X1 U3683 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2825) );
  NOR4_X1 U3684 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2824) );
  NOR4_X1 U3685 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2823) );
  NAND4_X1 U3686 ( .A1(n2826), .A2(n2825), .A3(n2824), .A4(n2823), .ZN(n2833)
         );
  NOR2_X1 U3687 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_23__SCAN_IN), .ZN(n2830)
         );
  NOR4_X1 U3688 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2829) );
  NOR4_X1 U3689 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2828) );
  NOR4_X1 U3690 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2827) );
  NAND4_X1 U3691 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .ZN(n2832)
         );
  OAI21_X1 U3692 ( .B1(n2833), .B2(n2832), .A(n2831), .ZN(n3082) );
  NAND3_X1 U3693 ( .A1(n2835), .A2(n2834), .A3(n3082), .ZN(n2843) );
  OAI22_X1 U3694 ( .A1(n3178), .A2(D_REG_0__SCAN_IN), .B1(n4530), .B2(n2815), 
        .ZN(n3153) );
  INV_X1 U3695 ( .A(n3153), .ZN(n3083) );
  MUX2_X1 U3696 ( .A(n2836), .B(n2844), .S(n4683), .Z(n2842) );
  NOR2_X2 U3697 ( .A1(n3334), .A2(n3160), .ZN(n3375) );
  OAI21_X1 U3698 ( .B1(n3133), .B2(n2839), .A(n4398), .ZN(n4199) );
  NAND2_X1 U3699 ( .A1(n2842), .A2(n2841), .ZN(U3515) );
  INV_X1 U3700 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2845) );
  MUX2_X1 U3701 ( .A(n2845), .B(n2844), .S(n4688), .Z(n2847) );
  NAND2_X1 U3702 ( .A1(n2847), .A2(n2846), .ZN(U3547) );
  INV_X1 U3703 ( .A(n3158), .ZN(n2848) );
  NAND2_X1 U3704 ( .A1(n2850), .A2(n2849), .ZN(n2854) );
  NAND2_X1 U3705 ( .A1(n2852), .A2(n2161), .ZN(n2853) );
  NAND2_X1 U3706 ( .A1(n2854), .A2(n2853), .ZN(n2855) );
  XNOR2_X1 U3707 ( .A(n2855), .B(n3062), .ZN(n2864) );
  XNOR2_X1 U3708 ( .A(n2864), .B(n2862), .ZN(n3320) );
  NAND2_X1 U3709 ( .A1(n3313), .A2(n2849), .ZN(n2856) );
  OAI211_X1 U3710 ( .C1(n3331), .C2(n2991), .A(n2856), .B(n2168), .ZN(n3192)
         );
  NAND2_X1 U3711 ( .A1(n3313), .A2(n2162), .ZN(n2860) );
  INV_X1 U3712 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3185) );
  NOR2_X1 U3713 ( .A1(n2851), .A2(n3185), .ZN(n2858) );
  AOI21_X1 U3714 ( .B1(n4167), .B2(n2849), .A(n2858), .ZN(n2859) );
  NAND2_X1 U3715 ( .A1(n2860), .A2(n2859), .ZN(n3191) );
  NAND2_X1 U3716 ( .A1(n3192), .A2(n3191), .ZN(n3190) );
  NAND2_X1 U3717 ( .A1(n2860), .A2(n3077), .ZN(n2861) );
  NAND2_X1 U3718 ( .A1(n3190), .A2(n2861), .ZN(n3319) );
  INV_X1 U3719 ( .A(n2862), .ZN(n2863) );
  NAND2_X1 U3720 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
  NAND2_X1 U3721 ( .A1(n3318), .A2(n2865), .ZN(n3299) );
  INV_X1 U3722 ( .A(n3299), .ZN(n2870) );
  NAND2_X1 U3723 ( .A1(n3160), .A2(n2162), .ZN(n2867) );
  OAI21_X1 U3724 ( .B1(n3330), .B2(n2866), .A(n2867), .ZN(n2868) );
  XNOR2_X1 U3725 ( .A(n2868), .B(n3077), .ZN(n2872) );
  AOI22_X1 U3726 ( .A1(n3445), .A2(n3009), .B1(n3160), .B2(n3104), .ZN(n2871)
         );
  XNOR2_X1 U3727 ( .A(n2872), .B(n2871), .ZN(n3300) );
  INV_X1 U3728 ( .A(n3300), .ZN(n2869) );
  NAND2_X1 U3729 ( .A1(n2870), .A2(n2869), .ZN(n3297) );
  NAND2_X1 U3730 ( .A1(n2872), .A2(n2871), .ZN(n2873) );
  NAND2_X1 U3731 ( .A1(n3377), .A2(n2162), .ZN(n2875) );
  NAND2_X1 U3732 ( .A1(n4165), .A2(n3104), .ZN(n2874) );
  NAND2_X1 U3733 ( .A1(n2875), .A2(n2874), .ZN(n2876) );
  XNOR2_X1 U3734 ( .A(n2876), .B(n3062), .ZN(n2877) );
  BUF_X4 U3735 ( .A(n2849), .Z(n3104) );
  AOI22_X1 U3736 ( .A1(n3377), .A2(n3104), .B1(n3009), .B2(n4165), .ZN(n2878)
         );
  XNOR2_X1 U3737 ( .A(n2877), .B(n2878), .ZN(n3342) );
  INV_X1 U3738 ( .A(n2877), .ZN(n2879) );
  NAND2_X1 U3739 ( .A1(n2879), .A2(n2878), .ZN(n2880) );
  NAND2_X1 U3740 ( .A1(n3421), .A2(n2161), .ZN(n2881) );
  OAI21_X1 U3741 ( .B1(n2542), .B2(n2866), .A(n2881), .ZN(n2882) );
  XNOR2_X1 U3742 ( .A(n2882), .B(n3077), .ZN(n2884) );
  AOI22_X1 U3743 ( .A1(n3501), .A2(n3009), .B1(n3421), .B2(n3104), .ZN(n2885)
         );
  XNOR2_X1 U3744 ( .A(n2884), .B(n2885), .ZN(n3428) );
  INV_X1 U3745 ( .A(n3428), .ZN(n2883) );
  INV_X1 U3746 ( .A(n2884), .ZN(n2887) );
  INV_X1 U3747 ( .A(n2885), .ZN(n2886) );
  NAND2_X1 U3748 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  NAND2_X1 U3749 ( .A1(n3425), .A2(n2888), .ZN(n3382) );
  OAI22_X1 U3750 ( .A1(n3536), .A2(n2866), .B1(n2585), .B2(n2905), .ZN(n2889)
         );
  XNOR2_X1 U3751 ( .A(n2889), .B(n3077), .ZN(n2890) );
  OAI22_X1 U3752 ( .A1(n3536), .A2(n2991), .B1(n2585), .B2(n2866), .ZN(n2891)
         );
  XNOR2_X1 U3753 ( .A(n2890), .B(n2891), .ZN(n3381) );
  INV_X1 U3754 ( .A(n2890), .ZN(n2892) );
  NAND2_X1 U3755 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
  NAND2_X1 U3756 ( .A1(n3540), .A2(n3104), .ZN(n2895) );
  NAND2_X1 U3757 ( .A1(n3009), .A2(n3511), .ZN(n2894) );
  NAND2_X1 U3758 ( .A1(n2895), .A2(n2894), .ZN(n3467) );
  NAND2_X1 U3759 ( .A1(n3540), .A2(n2161), .ZN(n2897) );
  NAND2_X1 U3760 ( .A1(n3511), .A2(n3104), .ZN(n2896) );
  NAND2_X1 U3761 ( .A1(n2897), .A2(n2896), .ZN(n2898) );
  XNOR2_X1 U3762 ( .A(n2898), .B(n3062), .ZN(n3468) );
  NAND2_X1 U3763 ( .A1(n2901), .A2(n2162), .ZN(n2899) );
  OAI21_X1 U3764 ( .B1(n3591), .B2(n2866), .A(n2899), .ZN(n2900) );
  XNOR2_X1 U3765 ( .A(n2900), .B(n3062), .ZN(n2923) );
  AOI22_X1 U3766 ( .A1(n4164), .A2(n3009), .B1(n3104), .B2(n2901), .ZN(n2921)
         );
  XNOR2_X1 U3767 ( .A(n2923), .B(n2921), .ZN(n3526) );
  NAND2_X1 U3768 ( .A1(n3627), .A2(n2162), .ZN(n2903) );
  NAND2_X1 U3769 ( .A1(n3588), .A2(n3104), .ZN(n2902) );
  NAND2_X1 U3770 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  XNOR2_X1 U3771 ( .A(n2904), .B(n3062), .ZN(n2909) );
  AOI22_X1 U3772 ( .A1(n3627), .A2(n3104), .B1(n3009), .B2(n3588), .ZN(n2910)
         );
  XNOR2_X1 U3773 ( .A(n2909), .B(n2910), .ZN(n3618) );
  INV_X1 U3774 ( .A(n3618), .ZN(n2920) );
  OAI22_X1 U3775 ( .A1(n3620), .A2(n2866), .B1(n3581), .B2(n2905), .ZN(n2906)
         );
  XNOR2_X1 U3776 ( .A(n2906), .B(n3062), .ZN(n2919) );
  INV_X1 U3777 ( .A(n2919), .ZN(n2908) );
  OAI22_X1 U3778 ( .A1(n3620), .A2(n2991), .B1(n3581), .B2(n2866), .ZN(n2918)
         );
  INV_X1 U3779 ( .A(n2918), .ZN(n2907) );
  NAND2_X1 U3780 ( .A1(n2908), .A2(n2907), .ZN(n3615) );
  OR2_X1 U3781 ( .A1(n2920), .A2(n3615), .ZN(n2917) );
  AND2_X1 U3782 ( .A1(n3526), .A2(n2917), .ZN(n2912) );
  INV_X1 U3783 ( .A(n2909), .ZN(n2911) );
  NAND2_X1 U3784 ( .A1(n2911), .A2(n2910), .ZN(n2927) );
  AND2_X1 U3785 ( .A1(n2912), .A2(n2927), .ZN(n3602) );
  NAND2_X1 U3786 ( .A1(n3657), .A2(n2161), .ZN(n2914) );
  NAND2_X1 U3787 ( .A1(n3652), .A2(n3104), .ZN(n2913) );
  NAND2_X1 U3788 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  XNOR2_X1 U3789 ( .A(n2915), .B(n3077), .ZN(n2930) );
  AOI22_X1 U3790 ( .A1(n3657), .A2(n3104), .B1(n3009), .B2(n3652), .ZN(n2931)
         );
  XNOR2_X1 U3791 ( .A(n2930), .B(n2931), .ZN(n3608) );
  INV_X1 U3792 ( .A(n2917), .ZN(n2926) );
  NOR2_X1 U3793 ( .A1(n3613), .A2(n2920), .ZN(n2924) );
  INV_X1 U3794 ( .A(n2921), .ZN(n2922) );
  NAND2_X1 U3795 ( .A1(n2923), .A2(n2922), .ZN(n3527) );
  AND2_X1 U3796 ( .A1(n2924), .A2(n3527), .ZN(n2925) );
  INV_X1 U3797 ( .A(n2930), .ZN(n2933) );
  INV_X1 U3798 ( .A(n2931), .ZN(n2932) );
  NAND2_X1 U3799 ( .A1(n2933), .A2(n2932), .ZN(n2934) );
  INV_X1 U3800 ( .A(n2937), .ZN(n2935) );
  NAND2_X1 U3801 ( .A1(n3606), .A2(n2935), .ZN(n3553) );
  NAND2_X1 U3802 ( .A1(n3642), .A2(n3104), .ZN(n2936) );
  OAI21_X1 U3803 ( .B1(n3655), .B2(n2991), .A(n2936), .ZN(n3550) );
  NAND2_X1 U3804 ( .A1(n3553), .A2(n3550), .ZN(n2943) );
  NAND2_X1 U3805 ( .A1(n3642), .A2(n2162), .ZN(n2939) );
  OAI21_X1 U3806 ( .B1(n3655), .B2(n2866), .A(n2939), .ZN(n2940) );
  XNOR2_X1 U3807 ( .A(n2940), .B(n3062), .ZN(n3551) );
  NAND2_X1 U3808 ( .A1(n2941), .A2(n3551), .ZN(n2942) );
  NAND2_X1 U3809 ( .A1(n3713), .A2(n2161), .ZN(n2945) );
  NAND2_X1 U3810 ( .A1(n4162), .A2(n3104), .ZN(n2944) );
  NAND2_X1 U3811 ( .A1(n2945), .A2(n2944), .ZN(n2946) );
  XNOR2_X1 U3812 ( .A(n2946), .B(n3062), .ZN(n2949) );
  NAND2_X1 U3813 ( .A1(n3713), .A2(n3104), .ZN(n2948) );
  NAND2_X1 U3814 ( .A1(n3009), .A2(n4162), .ZN(n2947) );
  NAND2_X1 U3815 ( .A1(n2948), .A2(n2947), .ZN(n2950) );
  INV_X1 U3816 ( .A(n2949), .ZN(n2952) );
  INV_X1 U3817 ( .A(n2950), .ZN(n2951) );
  NAND2_X1 U3818 ( .A1(n2952), .A2(n2951), .ZN(n3571) );
  NAND2_X1 U3819 ( .A1(n3686), .A2(n2162), .ZN(n2954) );
  NAND2_X1 U3820 ( .A1(n4161), .A2(n3104), .ZN(n2953) );
  NAND2_X1 U3821 ( .A1(n2954), .A2(n2953), .ZN(n2955) );
  XNOR2_X1 U3822 ( .A(n2955), .B(n3077), .ZN(n3875) );
  NAND2_X1 U3823 ( .A1(n3686), .A2(n3104), .ZN(n2957) );
  NAND2_X1 U3824 ( .A1(n3009), .A2(n4161), .ZN(n2956) );
  NAND2_X1 U3825 ( .A1(n2957), .A2(n2956), .ZN(n3876) );
  NAND2_X1 U3826 ( .A1(n3744), .A2(n2161), .ZN(n2958) );
  OAI21_X1 U3827 ( .B1(n3815), .B2(n2866), .A(n2958), .ZN(n2959) );
  XNOR2_X1 U3828 ( .A(n2959), .B(n3062), .ZN(n2961) );
  NAND2_X1 U3829 ( .A1(n3744), .A2(n3104), .ZN(n2960) );
  OAI21_X1 U3830 ( .B1(n3815), .B2(n2991), .A(n2960), .ZN(n2962) );
  NAND2_X1 U3831 ( .A1(n2961), .A2(n2962), .ZN(n3668) );
  INV_X1 U3832 ( .A(n2961), .ZN(n2964) );
  INV_X1 U3833 ( .A(n2962), .ZN(n2963) );
  NAND2_X1 U3834 ( .A1(n2964), .A2(n2963), .ZN(n3667) );
  NAND2_X1 U3835 ( .A1(n3792), .A2(n2162), .ZN(n2966) );
  NAND2_X1 U3836 ( .A1(n4472), .A2(n3104), .ZN(n2965) );
  NAND2_X1 U3837 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  XNOR2_X1 U3838 ( .A(n2967), .B(n3077), .ZN(n2971) );
  NAND2_X1 U3839 ( .A1(n2970), .A2(n2971), .ZN(n3811) );
  NAND2_X1 U3840 ( .A1(n3792), .A2(n3104), .ZN(n2969) );
  NAND2_X1 U3841 ( .A1(n3009), .A2(n4472), .ZN(n2968) );
  NAND2_X1 U3842 ( .A1(n2969), .A2(n2968), .ZN(n3822) );
  NAND2_X1 U3843 ( .A1(n3811), .A2(n3822), .ZN(n2976) );
  INV_X1 U3844 ( .A(n2970), .ZN(n2973) );
  NAND2_X1 U3845 ( .A1(n2973), .A2(n2972), .ZN(n3810) );
  NAND2_X1 U3846 ( .A1(n3847), .A2(n2162), .ZN(n2974) );
  OAI21_X1 U3847 ( .B1(n4461), .B2(n2866), .A(n2974), .ZN(n2975) );
  XNOR2_X1 U3848 ( .A(n2975), .B(n3062), .ZN(n2977) );
  AOI22_X1 U3849 ( .A1(n3817), .A2(n3009), .B1(n3847), .B2(n3104), .ZN(n2978)
         );
  XNOR2_X1 U3850 ( .A(n2977), .B(n2978), .ZN(n3825) );
  NAND3_X1 U3851 ( .A1(n2976), .A2(n3810), .A3(n3825), .ZN(n2981) );
  INV_X1 U3852 ( .A(n2977), .ZN(n2979) );
  NAND2_X1 U3853 ( .A1(n2979), .A2(n2978), .ZN(n2980) );
  NAND2_X1 U3854 ( .A1(n4464), .A2(n2161), .ZN(n2983) );
  NAND2_X1 U3855 ( .A1(n4473), .A2(n3104), .ZN(n2982) );
  NAND2_X1 U3856 ( .A1(n2983), .A2(n2982), .ZN(n2984) );
  XNOR2_X1 U3857 ( .A(n2984), .B(n3077), .ZN(n3803) );
  NAND2_X1 U3858 ( .A1(n4464), .A2(n3104), .ZN(n2986) );
  NAND2_X1 U3859 ( .A1(n3009), .A2(n4473), .ZN(n2985) );
  AND2_X1 U3860 ( .A1(n3803), .A2(n3802), .ZN(n2987) );
  NAND2_X1 U3861 ( .A1(n3836), .A2(n2161), .ZN(n2988) );
  OAI21_X1 U3862 ( .B1(n4459), .B2(n2866), .A(n2988), .ZN(n2989) );
  XNOR2_X1 U3863 ( .A(n2989), .B(n3062), .ZN(n2993) );
  NAND2_X1 U3864 ( .A1(n3836), .A2(n3104), .ZN(n2990) );
  OAI21_X1 U3865 ( .B1(n4459), .B2(n2991), .A(n2990), .ZN(n2994) );
  AND2_X1 U3866 ( .A1(n2993), .A2(n2994), .ZN(n3832) );
  INV_X1 U3867 ( .A(n3832), .ZN(n2992) );
  INV_X1 U3868 ( .A(n2993), .ZN(n2996) );
  INV_X1 U3869 ( .A(n2994), .ZN(n2995) );
  NAND2_X1 U3870 ( .A1(n2996), .A2(n2995), .ZN(n3831) );
  NAND2_X1 U3871 ( .A1(n4358), .A2(n2162), .ZN(n2999) );
  NAND2_X1 U3872 ( .A1(n3859), .A2(n3104), .ZN(n2998) );
  NAND2_X1 U3873 ( .A1(n2999), .A2(n2998), .ZN(n3000) );
  XNOR2_X1 U3874 ( .A(n3000), .B(n3062), .ZN(n3001) );
  AOI22_X1 U3875 ( .A1(n4358), .A2(n3104), .B1(n3009), .B2(n3859), .ZN(n3002)
         );
  XNOR2_X1 U3876 ( .A(n3001), .B(n3002), .ZN(n3927) );
  NAND2_X1 U3877 ( .A1(n3926), .A2(n3927), .ZN(n3005) );
  INV_X1 U3878 ( .A(n3001), .ZN(n3003) );
  NAND2_X1 U3879 ( .A1(n3003), .A2(n3002), .ZN(n3004) );
  NAND2_X1 U3880 ( .A1(n4103), .A2(n3104), .ZN(n3007) );
  NAND2_X1 U3881 ( .A1(n4344), .A2(n2161), .ZN(n3006) );
  NAND2_X1 U3882 ( .A1(n3007), .A2(n3006), .ZN(n3008) );
  XNOR2_X1 U3883 ( .A(n3008), .B(n3062), .ZN(n3012) );
  NAND2_X1 U3884 ( .A1(n3009), .A2(n4103), .ZN(n3011) );
  NAND2_X1 U3885 ( .A1(n4344), .A2(n3104), .ZN(n3010) );
  NAND2_X1 U3886 ( .A1(n3011), .A2(n3010), .ZN(n3013) );
  NAND2_X1 U3887 ( .A1(n3012), .A2(n3013), .ZN(n3964) );
  NAND2_X1 U3888 ( .A1(n3963), .A2(n3964), .ZN(n3962) );
  INV_X1 U3889 ( .A(n3012), .ZN(n3015) );
  INV_X1 U3890 ( .A(n3013), .ZN(n3014) );
  NAND2_X1 U3891 ( .A1(n3015), .A2(n3014), .ZN(n3966) );
  NAND2_X1 U3892 ( .A1(n3962), .A2(n3966), .ZN(n3937) );
  NAND2_X1 U3893 ( .A1(n4334), .A2(n3104), .ZN(n3017) );
  NAND2_X1 U3894 ( .A1(n4437), .A2(n2161), .ZN(n3016) );
  NAND2_X1 U3895 ( .A1(n3017), .A2(n3016), .ZN(n3018) );
  XNOR2_X1 U3896 ( .A(n3018), .B(n3077), .ZN(n3935) );
  NAND2_X1 U3897 ( .A1(n4334), .A2(n3009), .ZN(n3020) );
  NAND2_X1 U3898 ( .A1(n4437), .A2(n3104), .ZN(n3019) );
  AND2_X1 U3899 ( .A1(n3935), .A2(n3934), .ZN(n3021) );
  INV_X1 U3900 ( .A(n3935), .ZN(n3023) );
  INV_X1 U3901 ( .A(n3934), .ZN(n3022) );
  NAND2_X1 U3902 ( .A1(n3023), .A2(n3022), .ZN(n3024) );
  NAND2_X1 U3903 ( .A1(n4438), .A2(n3104), .ZN(n3026) );
  NAND2_X1 U3904 ( .A1(n4308), .A2(n2162), .ZN(n3025) );
  NAND2_X1 U3905 ( .A1(n3026), .A2(n3025), .ZN(n3027) );
  XNOR2_X1 U3906 ( .A(n3027), .B(n3077), .ZN(n3035) );
  NOR2_X1 U3907 ( .A1(n4298), .A2(n2866), .ZN(n3028) );
  AOI21_X1 U3908 ( .B1(n4438), .B2(n3009), .A(n3028), .ZN(n3034) );
  XNOR2_X1 U3909 ( .A(n3035), .B(n3034), .ZN(n3889) );
  NAND2_X1 U3910 ( .A1(n4307), .A2(n3104), .ZN(n3031) );
  NAND2_X1 U3911 ( .A1(n4285), .A2(n2162), .ZN(n3030) );
  NAND2_X1 U3912 ( .A1(n3031), .A2(n3030), .ZN(n3032) );
  XNOR2_X1 U3913 ( .A(n3032), .B(n3062), .ZN(n3039) );
  NOR2_X1 U3914 ( .A1(n4290), .A2(n2866), .ZN(n3033) );
  AOI21_X1 U3915 ( .B1(n4307), .B2(n3009), .A(n3033), .ZN(n3037) );
  XNOR2_X1 U3916 ( .A(n3039), .B(n3037), .ZN(n3917) );
  NAND2_X1 U3917 ( .A1(n3035), .A2(n3034), .ZN(n3918) );
  AND2_X1 U3918 ( .A1(n3917), .A2(n3918), .ZN(n3036) );
  INV_X1 U3919 ( .A(n3037), .ZN(n3038) );
  NAND2_X1 U3920 ( .A1(n3039), .A2(n3038), .ZN(n3046) );
  NOR2_X1 U3921 ( .A1(n4267), .A2(n2866), .ZN(n3040) );
  AOI21_X1 U3922 ( .B1(n4418), .B2(n3009), .A(n3040), .ZN(n3047) );
  AND2_X1 U3923 ( .A1(n3046), .A2(n3047), .ZN(n3041) );
  NAND2_X1 U3924 ( .A1(n3916), .A2(n3041), .ZN(n3951) );
  NAND2_X1 U3925 ( .A1(n4418), .A2(n3104), .ZN(n3044) );
  NAND2_X1 U3926 ( .A1(n3042), .A2(n2161), .ZN(n3043) );
  NAND2_X1 U3927 ( .A1(n3044), .A2(n3043), .ZN(n3045) );
  XNOR2_X1 U3928 ( .A(n3045), .B(n3062), .ZN(n3954) );
  NAND2_X1 U3929 ( .A1(n3951), .A2(n3954), .ZN(n3050) );
  NAND2_X1 U3930 ( .A1(n3916), .A2(n3046), .ZN(n3049) );
  INV_X1 U3931 ( .A(n3047), .ZN(n3048) );
  NAND2_X1 U3932 ( .A1(n3049), .A2(n3048), .ZN(n3952) );
  NAND2_X1 U3933 ( .A1(n3050), .A2(n3952), .ZN(n3945) );
  NAND2_X1 U3934 ( .A1(n4261), .A2(n3104), .ZN(n3052) );
  NAND2_X1 U3935 ( .A1(n4417), .A2(n2162), .ZN(n3051) );
  NAND2_X1 U3936 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNOR2_X1 U3937 ( .A(n3053), .B(n3077), .ZN(n3055) );
  NOR2_X1 U3938 ( .A1(n4246), .A2(n2866), .ZN(n3054) );
  AOI21_X1 U3939 ( .B1(n4261), .B2(n3009), .A(n3054), .ZN(n3056) );
  NAND2_X1 U3940 ( .A1(n3055), .A2(n3056), .ZN(n3943) );
  NAND2_X1 U3941 ( .A1(n3945), .A2(n3943), .ZN(n3059) );
  INV_X1 U3942 ( .A(n3055), .ZN(n3058) );
  INV_X1 U3943 ( .A(n3056), .ZN(n3057) );
  NAND2_X1 U3944 ( .A1(n3058), .A2(n3057), .ZN(n3944) );
  NAND2_X1 U3945 ( .A1(n4405), .A2(n3104), .ZN(n3061) );
  NAND2_X1 U3946 ( .A1(n4228), .A2(n2161), .ZN(n3060) );
  NAND2_X1 U3947 ( .A1(n3061), .A2(n3060), .ZN(n3063) );
  XNOR2_X1 U3948 ( .A(n3063), .B(n3062), .ZN(n3070) );
  NAND2_X1 U3949 ( .A1(n4405), .A2(n3009), .ZN(n3065) );
  NAND2_X1 U3950 ( .A1(n4228), .A2(n3104), .ZN(n3064) );
  NAND2_X1 U3951 ( .A1(n3065), .A2(n3064), .ZN(n3071) );
  AND2_X1 U3952 ( .A1(n3070), .A2(n3071), .ZN(n3976) );
  NAND2_X1 U3953 ( .A1(n4159), .A2(n3104), .ZN(n3067) );
  NAND2_X1 U3954 ( .A1(n4404), .A2(n2162), .ZN(n3066) );
  NAND2_X1 U3955 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
  XNOR2_X1 U3956 ( .A(n3068), .B(n3077), .ZN(n3090) );
  NOR2_X1 U3957 ( .A1(n4212), .A2(n2866), .ZN(n3069) );
  AOI21_X1 U3958 ( .B1(n4159), .B2(n3009), .A(n3069), .ZN(n3089) );
  INV_X1 U3959 ( .A(n3908), .ZN(n3074) );
  INV_X1 U3960 ( .A(n3070), .ZN(n3073) );
  INV_X1 U3961 ( .A(n3071), .ZN(n3072) );
  NAND2_X1 U3962 ( .A1(n3073), .A2(n3072), .ZN(n3975) );
  NOR2_X1 U3963 ( .A1(n3907), .A2(n2354), .ZN(n3093) );
  NAND2_X1 U3964 ( .A1(n4158), .A2(n3009), .ZN(n3076) );
  NAND2_X1 U3965 ( .A1(n3898), .A2(n3104), .ZN(n3075) );
  NAND2_X1 U3966 ( .A1(n3076), .A2(n3075), .ZN(n3078) );
  XNOR2_X1 U3967 ( .A(n3078), .B(n3077), .ZN(n3080) );
  AOI22_X1 U3968 ( .A1(n4158), .A2(n3104), .B1(n3898), .B2(n2161), .ZN(n3079)
         );
  XNOR2_X1 U3969 ( .A(n3080), .B(n3079), .ZN(n3094) );
  AND2_X1 U3970 ( .A1(n3082), .A2(n3081), .ZN(n3155) );
  NAND2_X1 U3971 ( .A1(n3239), .A2(n4533), .ZN(n3085) );
  NAND2_X1 U3972 ( .A1(n3085), .A2(n3084), .ZN(n3086) );
  OR2_X1 U3973 ( .A1(n4463), .A2(n3086), .ZN(n3098) );
  NOR2_X1 U3974 ( .A1(n3151), .A2(n3098), .ZN(n3087) );
  INV_X1 U3975 ( .A(n3988), .ZN(n3088) );
  NAND3_X1 U3976 ( .A1(n3093), .A2(n3094), .A3(n3088), .ZN(n3118) );
  NOR2_X1 U3977 ( .A1(n3090), .A2(n3089), .ZN(n3095) );
  NOR2_X1 U3978 ( .A1(n3095), .A2(n3988), .ZN(n3091) );
  NOR2_X1 U3979 ( .A1(n3093), .A2(n3092), .ZN(n3116) );
  INV_X1 U3980 ( .A(n3094), .ZN(n3097) );
  INV_X1 U3981 ( .A(n3095), .ZN(n3096) );
  NAND2_X1 U3982 ( .A1(n3098), .A2(n4476), .ZN(n3100) );
  INV_X1 U3983 ( .A(n3099), .ZN(n3150) );
  AOI21_X1 U3984 ( .B1(n3110), .B2(n3100), .A(n3150), .ZN(n3303) );
  NAND3_X1 U3985 ( .A1(n3303), .A2(n2851), .A3(n3101), .ZN(n3106) );
  NOR2_X1 U3986 ( .A1(n4655), .A2(n3102), .ZN(n3103) );
  NAND2_X1 U3987 ( .A1(n3104), .A2(n3103), .ZN(n4153) );
  NOR2_X1 U3988 ( .A1(n3105), .A2(n4153), .ZN(n3301) );
  AOI22_X1 U3989 ( .A1(n2193), .A2(n3899), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3112) );
  NOR3_X2 U3990 ( .A1(n3110), .A2(n3194), .A3(n4153), .ZN(n3929) );
  NAND2_X1 U3991 ( .A1(n3302), .A2(n4463), .ZN(n3109) );
  INV_X1 U3992 ( .A(n3107), .ZN(n3108) );
  OAI21_X2 U3993 ( .B1(n3110), .B2(n3109), .A(n4300), .ZN(n3928) );
  AOI22_X1 U3994 ( .A1(n3929), .A2(n4159), .B1(n3898), .B2(n3928), .ZN(n3111)
         );
  OAI211_X1 U3995 ( .C1(n3821), .C2(n3896), .A(n3112), .B(n3111), .ZN(n3113)
         );
  INV_X1 U3996 ( .A(n3113), .ZN(n3114) );
  NOR2_X1 U3997 ( .A1(n3116), .A2(n3115), .ZN(n3117) );
  NAND2_X1 U3998 ( .A1(n3118), .A2(n3117), .ZN(U3217) );
  XNOR2_X1 U3999 ( .A(n3119), .B(n4098), .ZN(n3906) );
  INV_X1 U4000 ( .A(n4676), .ZN(n4483) );
  OR2_X1 U4001 ( .A1(n3906), .A2(n4483), .ZN(n3128) );
  XNOR2_X1 U4002 ( .A(n3120), .B(n4098), .ZN(n3122) );
  INV_X1 U4003 ( .A(n3899), .ZN(n3123) );
  OAI22_X1 U4004 ( .A1(n3123), .A2(n4458), .B1(n4476), .B2(n3131), .ZN(n3125)
         );
  NAND2_X1 U4005 ( .A1(n3128), .A2(n3127), .ZN(n3137) );
  INV_X1 U4006 ( .A(n3129), .ZN(n3136) );
  NOR2_X1 U4007 ( .A1(n3130), .A2(n3131), .ZN(n3132) );
  NAND2_X1 U4008 ( .A1(n3136), .A2(n3135), .ZN(U3546) );
  INV_X1 U4009 ( .A(n3138), .ZN(n3141) );
  NAND2_X1 U4010 ( .A1(n3141), .A2(n3140), .ZN(U3514) );
  NOR2_X1 U4011 ( .A1(n2851), .A2(n4655), .ZN(U4043) );
  OAI21_X1 U4012 ( .B1(n3144), .B2(n3143), .A(n3142), .ZN(n3361) );
  INV_X1 U4013 ( .A(n4339), .ZN(n3585) );
  NAND2_X1 U4014 ( .A1(n3361), .A2(n3585), .ZN(n3149) );
  OAI21_X1 U4015 ( .B1(n4119), .B2(n3146), .A(n3145), .ZN(n3147) );
  NAND2_X1 U4016 ( .A1(n3147), .A2(n3121), .ZN(n3148) );
  NAND2_X1 U4017 ( .A1(n3149), .A2(n3148), .ZN(n3359) );
  NOR2_X1 U4018 ( .A1(n3151), .A2(n3150), .ZN(n3154) );
  NAND4_X1 U4019 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3156)
         );
  MUX2_X1 U4020 ( .A(REG2_REG_2__SCAN_IN), .B(n3359), .S(n4544), .Z(n3165) );
  NAND2_X1 U4021 ( .A1(n4544), .A2(n4471), .ZN(n4383) );
  INV_X1 U4022 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3157) );
  OAI22_X1 U4023 ( .A1(n4383), .A2(n3311), .B1(n3157), .B2(n4300), .ZN(n3164)
         );
  AND2_X1 U4024 ( .A1(n4544), .A2(n4474), .ZN(n4378) );
  INV_X1 U4025 ( .A(n4378), .ZN(n4214) );
  INV_X1 U4026 ( .A(n4379), .ZN(n4213) );
  OAI22_X1 U4027 ( .A1(n3424), .A2(n4214), .B1(n4213), .B2(n3358), .ZN(n3163)
         );
  INV_X1 U4028 ( .A(n3361), .ZN(n3161) );
  OR2_X1 U4029 ( .A1(n3158), .A2(n4190), .ZN(n3461) );
  INV_X1 U4030 ( .A(n3461), .ZN(n3159) );
  NAND2_X1 U4031 ( .A1(n4544), .A2(n3159), .ZN(n4347) );
  XNOR2_X1 U4032 ( .A(n3334), .B(n3160), .ZN(n3436) );
  NAND2_X1 U4033 ( .A1(n4544), .A2(n4190), .ZN(n3870) );
  OAI22_X1 U4034 ( .A1(n3161), .A2(n4347), .B1(n3436), .B2(n4368), .ZN(n3162)
         );
  OR4_X1 U4035 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(U3288) );
  MUX2_X1 U4036 ( .A(n3291), .B(n3166), .S(U3149), .Z(n3167) );
  INV_X1 U4037 ( .A(n3167), .ZN(U3344) );
  INV_X1 U4038 ( .A(DATAI_22_), .ZN(n4974) );
  NAND2_X1 U4039 ( .A1(n3168), .A2(STATE_REG_SCAN_IN), .ZN(n3169) );
  OAI21_X1 U4040 ( .B1(STATE_REG_SCAN_IN), .B2(n4974), .A(n3169), .ZN(U3330)
         );
  INV_X1 U4041 ( .A(DATAI_29_), .ZN(n4733) );
  NAND2_X1 U4042 ( .A1(n3170), .A2(STATE_REG_SCAN_IN), .ZN(n3171) );
  OAI21_X1 U40430 ( .B1(STATE_REG_SCAN_IN), .B2(n4733), .A(n3171), .ZN(U3323)
         );
  INV_X1 U4044 ( .A(DATAI_18_), .ZN(n4938) );
  NAND2_X1 U4045 ( .A1(n4185), .A2(STATE_REG_SCAN_IN), .ZN(n3172) );
  OAI21_X1 U4046 ( .B1(STATE_REG_SCAN_IN), .B2(n4938), .A(n3172), .ZN(U3334)
         );
  INV_X1 U4047 ( .A(DATAI_31_), .ZN(n3174) );
  OR4_X1 U4048 ( .A1(n2519), .A2(IR_REG_30__SCAN_IN), .A3(n2443), .A4(U3149), 
        .ZN(n3173) );
  OAI21_X1 U4049 ( .B1(STATE_REG_SCAN_IN), .B2(n3174), .A(n3173), .ZN(U3321)
         );
  INV_X1 U4050 ( .A(DATAI_20_), .ZN(n4732) );
  NAND2_X1 U4051 ( .A1(n4143), .A2(STATE_REG_SCAN_IN), .ZN(n3175) );
  OAI21_X1 U4052 ( .B1(STATE_REG_SCAN_IN), .B2(n4732), .A(n3175), .ZN(U3332)
         );
  INV_X1 U4053 ( .A(DATAI_27_), .ZN(n3177) );
  NAND2_X1 U4054 ( .A1(n3193), .A2(STATE_REG_SCAN_IN), .ZN(n3176) );
  OAI21_X1 U4055 ( .B1(STATE_REG_SCAN_IN), .B2(n3177), .A(n3176), .ZN(U3325)
         );
  NAND2_X1 U4056 ( .A1(n3302), .A2(n3178), .ZN(n4654) );
  NOR3_X1 U4057 ( .A1(n4531), .A2(n4530), .A3(n4655), .ZN(n3179) );
  AOI21_X1 U4058 ( .B1(n4654), .B2(n3180), .A(n3179), .ZN(U3459) );
  INV_X1 U4059 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3188) );
  AOI21_X1 U4060 ( .B1(n3181), .B2(n3185), .A(IR_REG_0__SCAN_IN), .ZN(n3182)
         );
  OAI21_X1 U4061 ( .B1(n3181), .B2(REG2_REG_0__SCAN_IN), .A(n4529), .ZN(n3197)
         );
  MUX2_X1 U4062 ( .A(n3182), .B(IR_REG_0__SCAN_IN), .S(n3197), .Z(n3184) );
  AOI22_X1 U4063 ( .A1(n3184), .A2(n3183), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3187) );
  NAND3_X1 U4064 ( .A1(n4631), .A2(IR_REG_0__SCAN_IN), .A3(n3185), .ZN(n3186)
         );
  OAI211_X1 U4065 ( .C1(n3189), .C2(n3188), .A(n3187), .B(n3186), .ZN(U3240)
         );
  OAI21_X1 U4066 ( .B1(n3192), .B2(n3191), .A(n3190), .ZN(n3310) );
  NOR2_X1 U4067 ( .A1(n3194), .A2(n3193), .ZN(n3199) );
  INV_X1 U4068 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3195) );
  NOR2_X1 U4069 ( .A1(n4152), .A2(n3195), .ZN(n3196) );
  MUX2_X1 U4070 ( .A(n3197), .B(n3196), .S(IR_REG_0__SCAN_IN), .Z(n3198) );
  AOI211_X1 U4071 ( .C1(n3310), .C2(n3199), .A(n3198), .B(n3263), .ZN(n3225)
         );
  NAND2_X1 U4072 ( .A1(n4168), .A2(n4540), .ZN(n3209) );
  OAI211_X1 U4073 ( .C1(n3202), .C2(n3201), .A(n4592), .B(n3200), .ZN(n3208)
         );
  OAI211_X1 U4074 ( .C1(n3205), .C2(n3204), .A(n4631), .B(n3203), .ZN(n3207)
         );
  AOI22_X1 U4075 ( .A1(n4630), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3206) );
  NAND4_X1 U4076 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3210)
         );
  OR2_X1 U4077 ( .A1(n3225), .A2(n3210), .ZN(U3242) );
  XNOR2_X1 U4078 ( .A(n3211), .B(REG2_REG_3__SCAN_IN), .ZN(n3217) );
  NOR2_X1 U4079 ( .A1(STATE_REG_SCAN_IN), .A2(n2523), .ZN(n3341) );
  NOR2_X1 U4080 ( .A1(n4637), .A2(n2265), .ZN(n3212) );
  AOI211_X1 U4081 ( .C1(n4630), .C2(ADDR_REG_3__SCAN_IN), .A(n3341), .B(n3212), 
        .ZN(n3216) );
  OAI211_X1 U4082 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3214), .A(n4631), .B(n3213), 
        .ZN(n3215) );
  OAI211_X1 U4083 ( .C1(n3217), .C2(n4624), .A(n3216), .B(n3215), .ZN(U3243)
         );
  XOR2_X1 U4084 ( .A(REG2_REG_4__SCAN_IN), .B(n3218), .Z(n3227) );
  OAI211_X1 U4085 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3220), .A(n4631), .B(n3219), 
        .ZN(n3223) );
  NAND2_X1 U4086 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3422) );
  INV_X1 U4087 ( .A(n3422), .ZN(n3221) );
  AOI21_X1 U4088 ( .B1(n4630), .B2(ADDR_REG_4__SCAN_IN), .A(n3221), .ZN(n3222)
         );
  OAI211_X1 U4089 ( .C1(n4637), .C2(n3224), .A(n3223), .B(n3222), .ZN(n3226)
         );
  AOI211_X1 U4090 ( .C1(n4592), .C2(n3227), .A(n3226), .B(n3225), .ZN(n3228)
         );
  INV_X1 U4091 ( .A(n3228), .ZN(U3244) );
  XNOR2_X1 U4092 ( .A(n3229), .B(REG2_REG_6__SCAN_IN), .ZN(n3237) );
  INV_X1 U4093 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3230) );
  NOR2_X1 U4094 ( .A1(STATE_REG_SCAN_IN), .A2(n3230), .ZN(n3473) );
  AOI21_X1 U4095 ( .B1(n4630), .B2(ADDR_REG_6__SCAN_IN), .A(n3473), .ZN(n3231)
         );
  INV_X1 U4096 ( .A(n3231), .ZN(n3235) );
  AOI211_X1 U4097 ( .C1(n3545), .C2(n3233), .A(n4194), .B(n3232), .ZN(n3234)
         );
  AOI211_X1 U4098 ( .C1(n4168), .C2(n4536), .A(n3235), .B(n3234), .ZN(n3236)
         );
  OAI21_X1 U4099 ( .B1(n3237), .B2(n4624), .A(n3236), .ZN(U3246) );
  INV_X2 U4100 ( .A(n3263), .ZN(n4166) );
  NOR2_X1 U4101 ( .A1(n4630), .A2(n4166), .ZN(U3148) );
  INV_X1 U4102 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U4103 ( .A1(n3652), .A2(n4166), .ZN(n3238) );
  OAI21_X1 U4104 ( .B1(n4166), .B2(n4933), .A(n3238), .ZN(U3560) );
  NOR2_X1 U4105 ( .A1(n3331), .A2(n3313), .ZN(n4028) );
  NOR2_X1 U4106 ( .A1(n4028), .A2(n4031), .ZN(n4125) );
  INV_X1 U4107 ( .A(n4125), .ZN(n3242) );
  INV_X1 U4108 ( .A(n3239), .ZN(n3240) );
  NOR2_X1 U4109 ( .A1(n3336), .A2(n3240), .ZN(n3347) );
  NOR2_X1 U4110 ( .A1(n3585), .A2(n3121), .ZN(n3241) );
  OAI22_X1 U4111 ( .A1(n4125), .A2(n3241), .B1(n3311), .B2(n4458), .ZN(n3348)
         );
  AOI211_X1 U4112 ( .C1(n4674), .C2(n3242), .A(n3347), .B(n3348), .ZN(n4670)
         );
  NAND2_X1 U4113 ( .A1(n4686), .A2(REG1_REG_0__SCAN_IN), .ZN(n3243) );
  OAI21_X1 U4114 ( .B1(n4670), .B2(n4686), .A(n3243), .ZN(U3518) );
  AOI211_X1 U4115 ( .C1(n3246), .C2(n3245), .A(n3244), .B(n4194), .ZN(n3254)
         );
  AOI211_X1 U4116 ( .C1(n3249), .C2(n3248), .A(n3247), .B(n4624), .ZN(n3253)
         );
  INV_X1 U4117 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U4118 ( .A1(STATE_REG_SCAN_IN), .A2(n4786), .ZN(n3384) );
  AOI21_X1 U4119 ( .B1(n4630), .B2(ADDR_REG_5__SCAN_IN), .A(n3384), .ZN(n3250)
         );
  OAI21_X1 U4120 ( .B1(n3251), .B2(n4637), .A(n3250), .ZN(n3252) );
  OR3_X1 U4121 ( .A1(n3254), .A2(n3253), .A3(n3252), .ZN(U3245) );
  INV_X1 U4122 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4971) );
  INV_X1 U4123 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U4124 ( .A1(n2608), .A2(REG1_REG_31__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U4125 ( .A1(n2549), .A2(REG2_REG_31__SCAN_IN), .ZN(n3255) );
  OAI211_X1 U4126 ( .C1(n3257), .C2(n4485), .A(n3256), .B(n3255), .ZN(n4392)
         );
  NAND2_X1 U4127 ( .A1(n4392), .A2(n4166), .ZN(n3258) );
  OAI21_X1 U4128 ( .B1(U4043), .B2(n4971), .A(n3258), .ZN(U3581) );
  INV_X1 U4129 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U4130 ( .A1(n3445), .A2(n4166), .ZN(n3259) );
  OAI21_X1 U4131 ( .B1(U4043), .B2(n4975), .A(n3259), .ZN(U3552) );
  INV_X1 U4132 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U4133 ( .A1(n3626), .A2(n4166), .ZN(n3260) );
  OAI21_X1 U4134 ( .B1(U4043), .B2(n4923), .A(n3260), .ZN(U3558) );
  INV_X1 U4135 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U4136 ( .A1(n4307), .A2(n4166), .ZN(n3261) );
  OAI21_X1 U4137 ( .B1(n4166), .B2(n4964), .A(n3261), .ZN(U3573) );
  INV_X1 U4138 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U4139 ( .A1(n3501), .A2(n4166), .ZN(n3262) );
  OAI21_X1 U4140 ( .B1(U4043), .B2(n4937), .A(n3262), .ZN(U3554) );
  INV_X1 U4141 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U4142 ( .A1(n4438), .A2(n4166), .ZN(n3264) );
  OAI21_X1 U4143 ( .B1(n4166), .B2(n4942), .A(n3264), .ZN(U3572) );
  INV_X1 U4144 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U4145 ( .A1(n3817), .A2(n4166), .ZN(n3265) );
  OAI21_X1 U4146 ( .B1(U4043), .B2(n4914), .A(n3265), .ZN(U3566) );
  INV_X1 U4147 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U4148 ( .A1(n3588), .A2(n4166), .ZN(n3266) );
  OAI21_X1 U4149 ( .B1(n4166), .B2(n4981), .A(n3266), .ZN(U3559) );
  INV_X1 U4150 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U4151 ( .A1(n3859), .A2(n4166), .ZN(n3267) );
  OAI21_X1 U4152 ( .B1(n4166), .B2(n4965), .A(n3267), .ZN(U3569) );
  INV_X1 U4153 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U4154 ( .A1(n4377), .A2(U4043), .ZN(n3268) );
  OAI21_X1 U4155 ( .B1(U4043), .B2(n4988), .A(n3268), .ZN(U3568) );
  INV_X1 U4156 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U4157 ( .A1(n3511), .A2(n4166), .ZN(n3269) );
  OAI21_X1 U4158 ( .B1(n4166), .B2(n4972), .A(n3269), .ZN(U3556) );
  INV_X1 U4159 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U4160 ( .A1(n4472), .A2(n4166), .ZN(n3270) );
  OAI21_X1 U4161 ( .B1(n4166), .B2(n4951), .A(n3270), .ZN(U3565) );
  INV_X1 U4162 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U4163 ( .A1(n4103), .A2(n4166), .ZN(n3271) );
  OAI21_X1 U4164 ( .B1(n4166), .B2(n4986), .A(n3271), .ZN(U3570) );
  INV_X1 U4165 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U4166 ( .A1(n3489), .A2(U4043), .ZN(n3272) );
  OAI21_X1 U4167 ( .B1(U4043), .B2(n4948), .A(n3272), .ZN(U3555) );
  INV_X1 U4168 ( .A(n3273), .ZN(n3275) );
  NAND2_X1 U4169 ( .A1(n3275), .A2(n3274), .ZN(n3277) );
  OAI21_X1 U4170 ( .B1(n3278), .B2(n3277), .A(n4631), .ZN(n3276) );
  AOI21_X1 U4171 ( .B1(n3278), .B2(n3277), .A(n3276), .ZN(n3285) );
  AOI211_X1 U4172 ( .C1(n3281), .C2(n3280), .A(n4624), .B(n3279), .ZN(n3284)
         );
  NOR2_X1 U4173 ( .A1(STATE_REG_SCAN_IN), .A2(n2574), .ZN(n3510) );
  AOI21_X1 U4174 ( .B1(n4630), .B2(ADDR_REG_7__SCAN_IN), .A(n3510), .ZN(n3282)
         );
  OAI21_X1 U4175 ( .B1(n2583), .B2(n4637), .A(n3282), .ZN(n3283) );
  OR3_X1 U4176 ( .A1(n3285), .A2(n3284), .A3(n3283), .ZN(U3247) );
  INV_X1 U4177 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U4178 ( .A1(n4261), .A2(n4166), .ZN(n3286) );
  OAI21_X1 U4179 ( .B1(n4166), .B2(n4915), .A(n3286), .ZN(U3575) );
  XNOR2_X1 U4180 ( .A(n3287), .B(REG1_REG_8__SCAN_IN), .ZN(n3295) );
  XNOR2_X1 U4181 ( .A(REG2_REG_8__SCAN_IN), .B(n3288), .ZN(n3289) );
  NAND2_X1 U4182 ( .A1(n4592), .A2(n3289), .ZN(n3290) );
  NAND2_X1 U4183 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3531) );
  NAND2_X1 U4184 ( .A1(n3290), .A2(n3531), .ZN(n3293) );
  NOR2_X1 U4185 ( .A1(n4637), .A2(n3291), .ZN(n3292) );
  AOI211_X1 U4186 ( .C1(n4630), .C2(ADDR_REG_8__SCAN_IN), .A(n3293), .B(n3292), 
        .ZN(n3294) );
  OAI21_X1 U4187 ( .B1(n3295), .B2(n4194), .A(n3294), .ZN(U3248) );
  INV_X1 U4188 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U4189 ( .A1(n4418), .A2(n4166), .ZN(n3296) );
  OAI21_X1 U4190 ( .B1(n4166), .B2(n4955), .A(n3296), .ZN(U3574) );
  INV_X1 U4191 ( .A(n3297), .ZN(n3298) );
  AOI21_X1 U4192 ( .B1(n3300), .B2(n3299), .A(n3298), .ZN(n3308) );
  INV_X1 U4193 ( .A(n3301), .ZN(n3304) );
  NAND3_X1 U4194 ( .A1(n3304), .A2(n3303), .A3(n3302), .ZN(n3309) );
  AOI22_X1 U4195 ( .A1(n2193), .A2(n4165), .B1(n3929), .B2(n2850), .ZN(n3305)
         );
  OAI21_X1 U4196 ( .B1(n3980), .B2(n3358), .A(n3305), .ZN(n3306) );
  AOI21_X1 U4197 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3309), .A(n3306), .ZN(n3307)
         );
  OAI21_X1 U4198 ( .B1(n3308), .B2(n3988), .A(n3307), .ZN(U3234) );
  INV_X1 U4199 ( .A(n3309), .ZN(n3323) );
  INV_X1 U4200 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3352) );
  OAI22_X1 U4201 ( .A1(n3983), .A2(n3311), .B1(n3310), .B2(n3988), .ZN(n3312)
         );
  AOI21_X1 U4202 ( .B1(n3313), .B2(n3928), .A(n3312), .ZN(n3314) );
  OAI21_X1 U4203 ( .B1(n3323), .B2(n3352), .A(n3314), .ZN(U3229) );
  INV_X1 U4204 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U4205 ( .A1(n4405), .A2(n4166), .ZN(n3315) );
  OAI21_X1 U4206 ( .B1(U4043), .B2(n4949), .A(n3315), .ZN(U3576) );
  INV_X1 U4207 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3437) );
  OAI22_X1 U4208 ( .A1(n3331), .A2(n3981), .B1(n3983), .B2(n3330), .ZN(n3317)
         );
  AOI21_X1 U4209 ( .B1(n2852), .B2(n3928), .A(n3317), .ZN(n3322) );
  OAI211_X1 U4210 ( .C1(n3320), .C2(n3319), .A(n3318), .B(n3088), .ZN(n3321)
         );
  OAI211_X1 U4211 ( .C1(n3323), .C2(n3437), .A(n3322), .B(n3321), .ZN(U3219)
         );
  OAI21_X1 U4212 ( .B1(n2779), .B2(n3325), .A(n3324), .ZN(n3441) );
  OR2_X1 U4213 ( .A1(n3441), .A2(n4339), .ZN(n3329) );
  OAI21_X1 U4214 ( .B1(n4118), .B2(n4031), .A(n3326), .ZN(n3327) );
  NAND2_X1 U4215 ( .A1(n3327), .A2(n3121), .ZN(n3328) );
  AND2_X1 U4216 ( .A1(n3329), .A2(n3328), .ZN(n3442) );
  INV_X1 U4217 ( .A(n4471), .ZN(n4460) );
  OAI22_X1 U4218 ( .A1(n3331), .A2(n4460), .B1(n3330), .B2(n4458), .ZN(n3332)
         );
  AOI21_X1 U4219 ( .B1(n2852), .B2(n4463), .A(n3332), .ZN(n3333) );
  OAI211_X1 U4220 ( .C1(n4449), .C2(n3441), .A(n3442), .B(n3333), .ZN(n3388)
         );
  OAI21_X1 U4221 ( .B1(n3336), .B2(n3335), .A(n3334), .ZN(n3448) );
  INV_X1 U4222 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3337) );
  OAI22_X1 U4223 ( .A1(n4526), .A2(n3448), .B1(n4683), .B2(n3337), .ZN(n3338)
         );
  AOI21_X1 U4224 ( .B1(n3388), .B2(n4683), .A(n3338), .ZN(n3339) );
  INV_X1 U4225 ( .A(n3339), .ZN(U3469) );
  OAI22_X1 U4226 ( .A1(n3983), .A2(n2542), .B1(n3980), .B2(n3372), .ZN(n3340)
         );
  AOI211_X1 U4227 ( .C1(n3929), .C2(n3445), .A(n3341), .B(n3340), .ZN(n3346)
         );
  XNOR2_X1 U4228 ( .A(n3343), .B(n3342), .ZN(n3344) );
  NAND2_X1 U4229 ( .A1(n3344), .A2(n3088), .ZN(n3345) );
  OAI211_X1 U4230 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3821), .A(n3346), .B(n3345), 
        .ZN(U3215) );
  INV_X1 U4231 ( .A(n3347), .ZN(n3350) );
  INV_X1 U4232 ( .A(n3348), .ZN(n3349) );
  OAI21_X1 U4233 ( .B1(n3351), .B2(n3350), .A(n3349), .ZN(n3354) );
  OAI22_X1 U4234 ( .A1(n4544), .A2(n3195), .B1(n3352), .B2(n4300), .ZN(n3353)
         );
  AOI21_X1 U4235 ( .B1(n3354), .B2(n4544), .A(n3353), .ZN(n3355) );
  OAI21_X1 U4236 ( .B1(n4125), .B2(n4347), .A(n3355), .ZN(U3290) );
  INV_X1 U4237 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U4238 ( .A1(n3899), .A2(n4166), .ZN(n3356) );
  OAI21_X1 U4239 ( .B1(n4166), .B2(n4987), .A(n3356), .ZN(U3579) );
  AOI22_X1 U4240 ( .A1(n2850), .A2(n4471), .B1(n4474), .B2(n4165), .ZN(n3357)
         );
  OAI21_X1 U4241 ( .B1(n3358), .B2(n4476), .A(n3357), .ZN(n3360) );
  AOI211_X1 U4242 ( .C1(n4674), .C2(n3361), .A(n3360), .B(n3359), .ZN(n3433)
         );
  OAI22_X1 U4243 ( .A1(n4526), .A2(n3436), .B1(n4683), .B2(n3362), .ZN(n3363)
         );
  INV_X1 U4244 ( .A(n3363), .ZN(n3364) );
  OAI21_X1 U4245 ( .B1(n3433), .B2(n4682), .A(n3364), .ZN(U3471) );
  NAND2_X1 U4246 ( .A1(n3142), .A2(n3365), .ZN(n3366) );
  XOR2_X1 U4247 ( .A(n4116), .B(n3366), .Z(n4649) );
  OAI21_X1 U4248 ( .B1(n4116), .B2(n3368), .A(n3367), .ZN(n3369) );
  NAND2_X1 U4249 ( .A1(n3369), .A2(n3121), .ZN(n3371) );
  AOI22_X1 U4250 ( .A1(n4471), .A2(n3445), .B1(n3501), .B2(n4474), .ZN(n3370)
         );
  OAI211_X1 U4251 ( .C1(n4476), .C2(n3372), .A(n3371), .B(n3370), .ZN(n3373)
         );
  AOI21_X1 U4252 ( .B1(n4649), .B2(n3585), .A(n3373), .ZN(n4652) );
  INV_X1 U4253 ( .A(n4652), .ZN(n3374) );
  AOI21_X1 U4254 ( .B1(n4674), .B2(n4649), .A(n3374), .ZN(n3410) );
  INV_X1 U4255 ( .A(n3375), .ZN(n3376) );
  AOI21_X1 U4256 ( .B1(n3377), .B2(n3376), .A(n2838), .ZN(n4646) );
  AOI22_X1 U4257 ( .A1(n4646), .A2(n3139), .B1(REG0_REG_3__SCAN_IN), .B2(n4682), .ZN(n3378) );
  OAI21_X1 U4258 ( .B1(n3410), .B2(n4682), .A(n3378), .ZN(U3473) );
  INV_X1 U4259 ( .A(n3379), .ZN(n3496) );
  OAI211_X1 U4260 ( .C1(n3382), .C2(n3381), .A(n3380), .B(n3088), .ZN(n3386)
         );
  OAI22_X1 U4261 ( .A1(n3983), .A2(n3498), .B1(n3980), .B2(n2585), .ZN(n3383)
         );
  AOI211_X1 U4262 ( .C1(n3929), .C2(n3501), .A(n3384), .B(n3383), .ZN(n3385)
         );
  OAI211_X1 U4263 ( .C1(n3821), .C2(n3496), .A(n3386), .B(n3385), .ZN(U3224)
         );
  OAI22_X1 U4264 ( .A1(n4470), .A2(n3448), .B1(n4688), .B2(n2481), .ZN(n3387)
         );
  AOI21_X1 U4265 ( .B1(n3388), .B2(n4688), .A(n3387), .ZN(n3389) );
  INV_X1 U4266 ( .A(n3389), .ZN(U3519) );
  XNOR2_X1 U4267 ( .A(n3390), .B(n3391), .ZN(n3401) );
  NAND2_X1 U4268 ( .A1(n3142), .A2(n3392), .ZN(n3394) );
  AND2_X1 U4269 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  NAND2_X1 U4270 ( .A1(n3395), .A2(n3390), .ZN(n3396) );
  NAND2_X1 U4271 ( .A1(n3397), .A2(n3396), .ZN(n3406) );
  AOI22_X1 U4272 ( .A1(n3489), .A2(n4474), .B1(n4471), .B2(n4165), .ZN(n3399)
         );
  NAND2_X1 U4273 ( .A1(n3421), .A2(n4463), .ZN(n3398) );
  OAI211_X1 U4274 ( .C1(n3406), .C2(n4339), .A(n3399), .B(n3398), .ZN(n3400)
         );
  AOI21_X1 U4275 ( .B1(n3401), .B2(n3121), .A(n3400), .ZN(n4671) );
  INV_X1 U4276 ( .A(n3416), .ZN(n3402) );
  AOI211_X1 U4277 ( .C1(n3421), .C2(n3404), .A(n3403), .B(n3402), .ZN(n4673)
         );
  INV_X1 U4278 ( .A(n4300), .ZN(n4645) );
  AOI22_X1 U4279 ( .A1(n4673), .A2(n4190), .B1(n4645), .B2(n3431), .ZN(n3405)
         );
  AND2_X1 U4280 ( .A1(n4671), .A2(n3405), .ZN(n3408) );
  INV_X1 U4281 ( .A(n3406), .ZN(n4675) );
  INV_X1 U4282 ( .A(n4347), .ZN(n4648) );
  AOI22_X1 U4283 ( .A1(n4675), .A2(n4648), .B1(REG2_REG_4__SCAN_IN), .B2(n2160), .ZN(n3407) );
  OAI21_X1 U4284 ( .B1(n3408), .B2(n2160), .A(n3407), .ZN(U3286) );
  INV_X1 U4285 ( .A(n4470), .ZN(n3633) );
  AOI22_X1 U4286 ( .A1(n4646), .A2(n3633), .B1(REG1_REG_3__SCAN_IN), .B2(n4686), .ZN(n3409) );
  OAI21_X1 U4287 ( .B1(n3410), .B2(n4686), .A(n3409), .ZN(U3521) );
  NAND2_X1 U4288 ( .A1(n4050), .A2(n4041), .ZN(n4110) );
  XOR2_X1 U4289 ( .A(n4110), .B(n3477), .Z(n3505) );
  XNOR2_X1 U4290 ( .A(n3411), .B(n4110), .ZN(n3412) );
  NAND2_X1 U4291 ( .A1(n3412), .A2(n3121), .ZN(n3507) );
  AOI22_X1 U4292 ( .A1(n3501), .A2(n4471), .B1(n4474), .B2(n3511), .ZN(n3413)
         );
  OAI211_X1 U4293 ( .C1(n4476), .C2(n2585), .A(n3507), .B(n3413), .ZN(n3414)
         );
  AOI21_X1 U4294 ( .B1(n3505), .B2(n4676), .A(n3414), .ZN(n3420) );
  AND2_X1 U4295 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  NOR2_X1 U4296 ( .A1(n3483), .A2(n3417), .ZN(n3495) );
  AOI22_X1 U4297 ( .A1(n3495), .A2(n3633), .B1(REG1_REG_5__SCAN_IN), .B2(n4686), .ZN(n3418) );
  OAI21_X1 U4298 ( .B1(n3420), .B2(n4686), .A(n3418), .ZN(U3523) );
  AOI22_X1 U4299 ( .A1(n3495), .A2(n3139), .B1(REG0_REG_5__SCAN_IN), .B2(n4682), .ZN(n3419) );
  OAI21_X1 U4300 ( .B1(n3420), .B2(n4682), .A(n3419), .ZN(U3477) );
  AOI22_X1 U4301 ( .A1(n2193), .A2(n3489), .B1(n3421), .B2(n3928), .ZN(n3423)
         );
  OAI211_X1 U4302 ( .C1(n3981), .C2(n3424), .A(n3423), .B(n3422), .ZN(n3430)
         );
  INV_X1 U4303 ( .A(n3425), .ZN(n3426) );
  AOI211_X1 U4304 ( .C1(n3428), .C2(n3427), .A(n3988), .B(n3426), .ZN(n3429)
         );
  AOI211_X1 U4305 ( .C1(n3431), .C2(n3986), .A(n3430), .B(n3429), .ZN(n3432)
         );
  INV_X1 U4306 ( .A(n3432), .ZN(U3227) );
  INV_X1 U4307 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3434) );
  MUX2_X1 U4308 ( .A(n3434), .B(n3433), .S(n4688), .Z(n3435) );
  OAI21_X1 U4309 ( .B1(n3436), .B2(n4470), .A(n3435), .ZN(U3520) );
  OAI22_X1 U4310 ( .A1(n4544), .A2(n3438), .B1(n3437), .B2(n4300), .ZN(n3439)
         );
  INV_X1 U4311 ( .A(n3439), .ZN(n3440) );
  OAI21_X1 U4312 ( .B1(n4347), .B2(n3441), .A(n3440), .ZN(n3444) );
  NOR2_X1 U4313 ( .A1(n3442), .A2(n2160), .ZN(n3443) );
  AOI211_X1 U4314 ( .C1(n4378), .C2(n3445), .A(n3444), .B(n3443), .ZN(n3447)
         );
  INV_X1 U4315 ( .A(n4383), .ZN(n3712) );
  AOI22_X1 U4316 ( .A1(n3712), .A2(n4167), .B1(n4379), .B2(n2852), .ZN(n3446)
         );
  OAI211_X1 U4317 ( .C1(n4368), .C2(n3448), .A(n3447), .B(n3446), .ZN(U3289)
         );
  INV_X1 U4318 ( .A(n3459), .ZN(n4126) );
  XNOR2_X1 U4319 ( .A(n3449), .B(n4126), .ZN(n3452) );
  AOI22_X1 U4320 ( .A1(n3626), .A2(n4474), .B1(n4471), .B2(n3511), .ZN(n3450)
         );
  OAI21_X1 U4321 ( .B1(n3508), .B2(n4476), .A(n3450), .ZN(n3451) );
  AOI21_X1 U4322 ( .B1(n3452), .B2(n3121), .A(n3451), .ZN(n4681) );
  NOR2_X1 U4323 ( .A1(n4544), .A2(n3453), .ZN(n3455) );
  OAI211_X1 U4324 ( .C1(n3485), .C2(n3508), .A(n4479), .B(n3579), .ZN(n4680)
         );
  NOR2_X1 U4325 ( .A1(n4680), .A2(n3870), .ZN(n3454) );
  AOI211_X1 U4326 ( .C1(n4645), .C2(n3512), .A(n3455), .B(n3454), .ZN(n3466)
         );
  NAND2_X1 U4327 ( .A1(n3477), .A2(n3456), .ZN(n3458) );
  NAND2_X1 U4328 ( .A1(n3458), .A2(n3457), .ZN(n3460) );
  OR2_X1 U4329 ( .A1(n3460), .A2(n3459), .ZN(n4678) );
  NAND2_X1 U4330 ( .A1(n4339), .A2(n3461), .ZN(n3462) );
  NAND2_X1 U4331 ( .A1(n4544), .A2(n3462), .ZN(n4391) );
  AND2_X1 U4332 ( .A1(n3464), .A2(n3463), .ZN(n4677) );
  NAND3_X1 U4333 ( .A1(n4678), .A2(n4318), .A3(n4677), .ZN(n3465) );
  OAI211_X1 U4334 ( .C1(n4681), .C2(n2160), .A(n3466), .B(n3465), .ZN(U3283)
         );
  XNOR2_X1 U4335 ( .A(n3468), .B(n3467), .ZN(n3469) );
  XNOR2_X1 U4336 ( .A(n3470), .B(n3469), .ZN(n3471) );
  NAND2_X1 U4337 ( .A1(n3471), .A2(n3088), .ZN(n3475) );
  OAI22_X1 U4338 ( .A1(n3983), .A2(n3591), .B1(n3980), .B2(n3482), .ZN(n3472)
         );
  AOI211_X1 U4339 ( .C1(n3929), .C2(n3489), .A(n3473), .B(n3472), .ZN(n3474)
         );
  OAI211_X1 U4340 ( .C1(n3821), .C2(n3486), .A(n3475), .B(n3474), .ZN(U3236)
         );
  NAND2_X1 U4341 ( .A1(n3477), .A2(n3476), .ZN(n3479) );
  NAND2_X1 U4342 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  NAND2_X1 U4343 ( .A1(n4044), .A2(n4051), .ZN(n4133) );
  XNOR2_X1 U4344 ( .A(n3480), .B(n4133), .ZN(n3542) );
  XNOR2_X1 U4345 ( .A(n3481), .B(n4133), .ZN(n3537) );
  INV_X1 U4346 ( .A(n3537), .ZN(n3493) );
  NOR2_X1 U4347 ( .A1(n2160), .A2(n4360), .ZN(n3751) );
  NOR2_X1 U4348 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  OR2_X1 U4349 ( .A1(n3485), .A2(n3484), .ZN(n3546) );
  INV_X1 U4350 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3487) );
  OAI22_X1 U4351 ( .A1(n4544), .A2(n3487), .B1(n3486), .B2(n4300), .ZN(n3488)
         );
  AOI21_X1 U4352 ( .B1(n3712), .B2(n3489), .A(n3488), .ZN(n3491) );
  AOI22_X1 U4353 ( .A1(n4379), .A2(n3540), .B1(n4378), .B2(n4164), .ZN(n3490)
         );
  OAI211_X1 U4354 ( .C1(n3546), .C2(n4368), .A(n3491), .B(n3490), .ZN(n3492)
         );
  AOI21_X1 U4355 ( .B1(n3493), .B2(n3751), .A(n3492), .ZN(n3494) );
  OAI21_X1 U4356 ( .B1(n4391), .B2(n3542), .A(n3494), .ZN(U3284) );
  INV_X1 U4357 ( .A(n3495), .ZN(n3503) );
  OAI22_X1 U4358 ( .A1(n4544), .A2(n3497), .B1(n3496), .B2(n4300), .ZN(n3500)
         );
  OAI22_X1 U4359 ( .A1(n3498), .A2(n4214), .B1(n4213), .B2(n2585), .ZN(n3499)
         );
  AOI211_X1 U4360 ( .C1(n3712), .C2(n3501), .A(n3500), .B(n3499), .ZN(n3502)
         );
  OAI21_X1 U4361 ( .B1(n4368), .B2(n3503), .A(n3502), .ZN(n3504) );
  AOI21_X1 U4362 ( .B1(n3505), .B2(n4318), .A(n3504), .ZN(n3506) );
  OAI21_X1 U4363 ( .B1(n2160), .B2(n3507), .A(n3506), .ZN(U3285) );
  XNOR2_X1 U4364 ( .A(n3601), .B(n3526), .ZN(n3515) );
  OAI22_X1 U4365 ( .A1(n3983), .A2(n3620), .B1(n3980), .B2(n3508), .ZN(n3509)
         );
  AOI211_X1 U4366 ( .C1(n3929), .C2(n3511), .A(n3510), .B(n3509), .ZN(n3514)
         );
  NAND2_X1 U4367 ( .A1(n3986), .A2(n3512), .ZN(n3513) );
  OAI211_X1 U4368 ( .C1(n3515), .C2(n3988), .A(n3514), .B(n3513), .ZN(U3210)
         );
  NAND2_X1 U4369 ( .A1(n4048), .A2(n4060), .ZN(n4111) );
  XNOR2_X1 U4370 ( .A(n3516), .B(n4111), .ZN(n3517) );
  NAND2_X1 U4371 ( .A1(n3517), .A2(n3121), .ZN(n3629) );
  AOI21_X1 U4372 ( .B1(n3627), .B2(n3580), .A(n3562), .ZN(n3637) );
  OAI22_X1 U4373 ( .A1(n3624), .A2(n4300), .B1(n3518), .B2(n4544), .ZN(n3521)
         );
  AOI22_X1 U4374 ( .A1(n3712), .A2(n3626), .B1(n4379), .B2(n3627), .ZN(n3519)
         );
  OAI21_X1 U4375 ( .B1(n3691), .B2(n4214), .A(n3519), .ZN(n3520) );
  AOI211_X1 U4376 ( .C1(n3637), .C2(n4647), .A(n3521), .B(n3520), .ZN(n3525)
         );
  INV_X1 U4377 ( .A(n4111), .ZN(n3523) );
  XNOR2_X1 U4378 ( .A(n3522), .B(n3523), .ZN(n3625) );
  NAND2_X1 U4379 ( .A1(n3625), .A2(n4318), .ZN(n3524) );
  OAI211_X1 U4380 ( .C1(n3629), .C2(n2160), .A(n3525), .B(n3524), .ZN(U3281)
         );
  NAND2_X1 U4381 ( .A1(n3601), .A2(n3526), .ZN(n3528) );
  NAND2_X1 U4382 ( .A1(n3528), .A2(n3527), .ZN(n3614) );
  INV_X1 U4383 ( .A(n3615), .ZN(n3529) );
  NOR2_X1 U4384 ( .A1(n3529), .A2(n3613), .ZN(n3530) );
  XNOR2_X1 U4385 ( .A(n3614), .B(n3530), .ZN(n3535) );
  AOI22_X1 U4386 ( .A1(n2193), .A2(n3588), .B1(n3587), .B2(n3928), .ZN(n3532)
         );
  OAI211_X1 U4387 ( .C1(n3981), .C2(n3591), .A(n3532), .B(n3531), .ZN(n3533)
         );
  AOI21_X1 U4388 ( .B1(n4638), .B2(n3986), .A(n3533), .ZN(n3534) );
  OAI21_X1 U4389 ( .B1(n3535), .B2(n3988), .A(n3534), .ZN(U3218) );
  OAI22_X1 U4390 ( .A1(n3536), .A2(n4460), .B1(n3591), .B2(n4458), .ZN(n3539)
         );
  NOR2_X1 U4391 ( .A1(n3537), .A2(n4360), .ZN(n3538) );
  AOI211_X1 U4392 ( .C1(n4463), .C2(n3540), .A(n3539), .B(n3538), .ZN(n3541)
         );
  OAI21_X1 U4393 ( .B1(n4483), .B2(n3542), .A(n3541), .ZN(n3548) );
  OAI22_X1 U4394 ( .A1(n3546), .A2(n4526), .B1(n4683), .B2(n2567), .ZN(n3543)
         );
  AOI21_X1 U4395 ( .B1(n3548), .B2(n4683), .A(n3543), .ZN(n3544) );
  INV_X1 U4396 ( .A(n3544), .ZN(U3479) );
  OAI22_X1 U4397 ( .A1(n3546), .A2(n4470), .B1(n4688), .B2(n3545), .ZN(n3547)
         );
  AOI21_X1 U4398 ( .B1(n3548), .B2(n4688), .A(n3547), .ZN(n3549) );
  INV_X1 U4399 ( .A(n3549), .ZN(U3524) );
  XNOR2_X1 U4400 ( .A(n3551), .B(n3550), .ZN(n3552) );
  XNOR2_X1 U4401 ( .A(n3553), .B(n3552), .ZN(n3554) );
  NAND2_X1 U4402 ( .A1(n3554), .A2(n3088), .ZN(n3557) );
  AND2_X1 U4403 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4578) );
  OAI22_X1 U4404 ( .A1(n3981), .A2(n3691), .B1(n3980), .B2(n3648), .ZN(n3555)
         );
  AOI211_X1 U4405 ( .C1(n2193), .C2(n4162), .A(n4578), .B(n3555), .ZN(n3556)
         );
  OAI211_X1 U4406 ( .C1(n3821), .C2(n3647), .A(n3557), .B(n3556), .ZN(U3233)
         );
  NAND2_X1 U4407 ( .A1(n4057), .A2(n4062), .ZN(n4112) );
  XNOR2_X1 U4408 ( .A(n3558), .B(n4112), .ZN(n3659) );
  INV_X1 U4409 ( .A(n3751), .ZN(n3569) );
  XNOR2_X1 U4410 ( .A(n3559), .B(n4112), .ZN(n3661) );
  NAND2_X1 U4411 ( .A1(n3661), .A2(n4318), .ZN(n3568) );
  INV_X1 U4412 ( .A(n3649), .ZN(n3560) );
  OAI21_X1 U4413 ( .B1(n3562), .B2(n3561), .A(n3560), .ZN(n3665) );
  INV_X1 U4414 ( .A(n3665), .ZN(n3566) );
  AOI22_X1 U4415 ( .A1(n4379), .A2(n3657), .B1(n4378), .B2(n4163), .ZN(n3564)
         );
  AOI22_X1 U4416 ( .A1(n2160), .A2(REG2_REG_10__SCAN_IN), .B1(n3611), .B2(
        n4645), .ZN(n3563) );
  OAI211_X1 U4417 ( .C1(n2324), .C2(n4383), .A(n3564), .B(n3563), .ZN(n3565)
         );
  AOI21_X1 U4418 ( .B1(n3566), .B2(n4647), .A(n3565), .ZN(n3567) );
  OAI211_X1 U4419 ( .C1(n3659), .C2(n3569), .A(n3568), .B(n3567), .ZN(U3280)
         );
  INV_X1 U4420 ( .A(n3571), .ZN(n3573) );
  NOR2_X1 U4421 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  XNOR2_X1 U4422 ( .A(n3570), .B(n3574), .ZN(n3578) );
  AOI22_X1 U4423 ( .A1(n2193), .A2(n4161), .B1(n3713), .B2(n3928), .ZN(n3575)
         );
  NAND2_X1 U4424 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4582) );
  OAI211_X1 U4425 ( .C1(n3981), .C2(n3655), .A(n3575), .B(n4582), .ZN(n3576)
         );
  AOI21_X1 U4426 ( .B1(n3708), .B2(n3986), .A(n3576), .ZN(n3577) );
  OAI21_X1 U4427 ( .B1(n3578), .B2(n3988), .A(n3577), .ZN(U3221) );
  INV_X1 U4428 ( .A(n3579), .ZN(n3582) );
  OAI21_X1 U4429 ( .B1(n3582), .B2(n3581), .A(n3580), .ZN(n4639) );
  NAND2_X1 U4430 ( .A1(n4047), .A2(n4052), .ZN(n4135) );
  INV_X1 U4431 ( .A(n4135), .ZN(n3583) );
  XNOR2_X1 U4432 ( .A(n3584), .B(n3583), .ZN(n4641) );
  NAND2_X1 U4433 ( .A1(n4641), .A2(n3585), .ZN(n3595) );
  XNOR2_X1 U4434 ( .A(n3586), .B(n4135), .ZN(n3593) );
  NAND2_X1 U4435 ( .A1(n3587), .A2(n4463), .ZN(n3590) );
  NAND2_X1 U4436 ( .A1(n3588), .A2(n4474), .ZN(n3589) );
  OAI211_X1 U4437 ( .C1(n3591), .C2(n4460), .A(n3590), .B(n3589), .ZN(n3592)
         );
  AOI21_X1 U4438 ( .B1(n3593), .B2(n3121), .A(n3592), .ZN(n3594) );
  AND2_X1 U4439 ( .A1(n3595), .A2(n3594), .ZN(n4644) );
  NAND2_X1 U4440 ( .A1(n4641), .A2(n4674), .ZN(n3596) );
  AND2_X1 U4441 ( .A1(n4644), .A2(n3596), .ZN(n3598) );
  MUX2_X1 U4442 ( .A(n3598), .B(n2594), .S(n4682), .Z(n3597) );
  OAI21_X1 U4443 ( .B1(n4639), .B2(n4526), .A(n3597), .ZN(U3483) );
  MUX2_X1 U4444 ( .A(n2201), .B(n3598), .S(n4688), .Z(n3599) );
  OAI21_X1 U4445 ( .B1(n4639), .B2(n4470), .A(n3599), .ZN(U3526) );
  AOI22_X1 U4446 ( .A1(n2193), .A2(n4163), .B1(n3657), .B2(n3928), .ZN(n3600)
         );
  NAND2_X1 U4447 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4561) );
  OAI211_X1 U4448 ( .C1(n3981), .C2(n2324), .A(n3600), .B(n4561), .ZN(n3610)
         );
  NAND2_X1 U4449 ( .A1(n3601), .A2(n3602), .ZN(n3604) );
  AND2_X1 U4450 ( .A1(n3604), .A2(n3603), .ZN(n3607) );
  AOI211_X1 U4451 ( .C1(n3608), .C2(n3607), .A(n3988), .B(n2191), .ZN(n3609)
         );
  AOI211_X1 U4452 ( .C1(n3611), .C2(n3986), .A(n3610), .B(n3609), .ZN(n3612)
         );
  INV_X1 U4453 ( .A(n3612), .ZN(U3214) );
  OR2_X1 U4454 ( .A1(n3614), .A2(n3613), .ZN(n3616) );
  NAND2_X1 U4455 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  XNOR2_X1 U4456 ( .A(n3618), .B(n3617), .ZN(n3619) );
  NAND2_X1 U4457 ( .A1(n3619), .A2(n3088), .ZN(n3623) );
  AND2_X1 U4458 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4557) );
  OAI22_X1 U4459 ( .A1(n3981), .A2(n3620), .B1(n3980), .B2(n2325), .ZN(n3621)
         );
  AOI211_X1 U4460 ( .C1(n2193), .C2(n3652), .A(n4557), .B(n3621), .ZN(n3622)
         );
  OAI211_X1 U4461 ( .C1(n3821), .C2(n3624), .A(n3623), .B(n3622), .ZN(U3228)
         );
  NAND2_X1 U4462 ( .A1(n3625), .A2(n4676), .ZN(n3631) );
  AOI22_X1 U4463 ( .A1(n3626), .A2(n4471), .B1(n4474), .B2(n3652), .ZN(n3630)
         );
  NAND2_X1 U4464 ( .A1(n3627), .A2(n4463), .ZN(n3628) );
  NAND4_X1 U4465 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3635)
         );
  MUX2_X1 U4466 ( .A(REG1_REG_9__SCAN_IN), .B(n3635), .S(n4688), .Z(n3632) );
  AOI21_X1 U4467 ( .B1(n3633), .B2(n3637), .A(n3632), .ZN(n3634) );
  INV_X1 U4468 ( .A(n3634), .ZN(U3527) );
  MUX2_X1 U4469 ( .A(REG0_REG_9__SCAN_IN), .B(n3635), .S(n4683), .Z(n3636) );
  AOI21_X1 U4470 ( .B1(n3637), .B2(n3139), .A(n3636), .ZN(n3638) );
  INV_X1 U4471 ( .A(n3638), .ZN(U3485) );
  INV_X1 U4472 ( .A(n3639), .ZN(n3640) );
  AOI21_X1 U4473 ( .B1(n4120), .B2(n3641), .A(n3640), .ZN(n3692) );
  AOI22_X1 U4474 ( .A1(n3642), .A2(n4463), .B1(n4162), .B2(n4474), .ZN(n3646)
         );
  XNOR2_X1 U4475 ( .A(n3643), .B(n4120), .ZN(n3644) );
  NAND2_X1 U4476 ( .A1(n3644), .A2(n3121), .ZN(n3645) );
  OAI211_X1 U4477 ( .C1(n3692), .C2(n4339), .A(n3646), .B(n3645), .ZN(n3694)
         );
  NAND2_X1 U4478 ( .A1(n3694), .A2(n4544), .ZN(n3654) );
  OAI22_X1 U4479 ( .A1(n3647), .A2(n4300), .B1(n4759), .B2(n4544), .ZN(n3651)
         );
  OAI21_X1 U4480 ( .B1(n3649), .B2(n3648), .A(n3705), .ZN(n3699) );
  NOR2_X1 U4481 ( .A1(n3699), .A2(n4368), .ZN(n3650) );
  AOI211_X1 U4482 ( .C1(n3712), .C2(n3652), .A(n3651), .B(n3650), .ZN(n3653)
         );
  OAI211_X1 U4483 ( .C1(n3692), .C2(n4347), .A(n3654), .B(n3653), .ZN(U3279)
         );
  OAI22_X1 U4484 ( .A1(n2324), .A2(n4460), .B1(n3655), .B2(n4458), .ZN(n3656)
         );
  AOI21_X1 U4485 ( .B1(n3657), .B2(n4463), .A(n3656), .ZN(n3658) );
  OAI21_X1 U4486 ( .B1(n3659), .B2(n4360), .A(n3658), .ZN(n3660) );
  AOI21_X1 U4487 ( .B1(n4676), .B2(n3661), .A(n3660), .ZN(n3663) );
  MUX2_X1 U4488 ( .A(n2614), .B(n3663), .S(n4683), .Z(n3662) );
  OAI21_X1 U4489 ( .B1(n3665), .B2(n4526), .A(n3662), .ZN(U3487) );
  INV_X1 U4490 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4750) );
  MUX2_X1 U4491 ( .A(n4750), .B(n3663), .S(n4688), .Z(n3664) );
  OAI21_X1 U4492 ( .B1(n3665), .B2(n4470), .A(n3664), .ZN(U3528) );
  NAND2_X1 U4493 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  XNOR2_X1 U4494 ( .A(n3666), .B(n3669), .ZN(n3674) );
  AOI22_X1 U4495 ( .A1(n2193), .A2(n4472), .B1(n3744), .B2(n3928), .ZN(n3671)
         );
  NOR2_X1 U4496 ( .A1(n4694), .A2(STATE_REG_SCAN_IN), .ZN(n3722) );
  INV_X1 U4497 ( .A(n3722), .ZN(n3670) );
  OAI211_X1 U4498 ( .C1(n3981), .C2(n3748), .A(n3671), .B(n3670), .ZN(n3672)
         );
  AOI21_X1 U4499 ( .B1(n3745), .B2(n3986), .A(n3672), .ZN(n3673) );
  OAI21_X1 U4500 ( .B1(n3674), .B2(n3988), .A(n3673), .ZN(U3212) );
  OAI21_X1 U4501 ( .B1(n3675), .B2(n3702), .A(n3701), .ZN(n3679) );
  INV_X1 U4502 ( .A(n3676), .ZN(n3678) );
  NOR2_X1 U4503 ( .A1(n3678), .A2(n3677), .ZN(n4106) );
  INV_X1 U4504 ( .A(n4106), .ZN(n3684) );
  XNOR2_X1 U4505 ( .A(n3679), .B(n3684), .ZN(n3683) );
  NAND2_X1 U4506 ( .A1(n3686), .A2(n4463), .ZN(n3681) );
  NAND2_X1 U4507 ( .A1(n4162), .A2(n4471), .ZN(n3680) );
  OAI211_X1 U4508 ( .C1(n3815), .C2(n4458), .A(n3681), .B(n3680), .ZN(n3682)
         );
  AOI21_X1 U4509 ( .B1(n3683), .B2(n3121), .A(n3682), .ZN(n3769) );
  XNOR2_X1 U4510 ( .A(n3685), .B(n3684), .ZN(n3768) );
  NAND2_X1 U4511 ( .A1(n3707), .A2(n3686), .ZN(n3687) );
  NAND2_X1 U4512 ( .A1(n3729), .A2(n3687), .ZN(n3776) );
  AOI22_X1 U4513 ( .A1(n2160), .A2(REG2_REG_13__SCAN_IN), .B1(n3882), .B2(
        n4645), .ZN(n3688) );
  OAI21_X1 U4514 ( .B1(n3776), .B2(n4368), .A(n3688), .ZN(n3689) );
  AOI21_X1 U4515 ( .B1(n3768), .B2(n4318), .A(n3689), .ZN(n3690) );
  OAI21_X1 U4516 ( .B1(n2160), .B2(n3769), .A(n3690), .ZN(U3277) );
  OAI22_X1 U4517 ( .A1(n3692), .A2(n4449), .B1(n3691), .B2(n4460), .ZN(n3693)
         );
  NOR2_X1 U4518 ( .A1(n3694), .A2(n3693), .ZN(n3697) );
  MUX2_X1 U4519 ( .A(n3695), .B(n3697), .S(n4683), .Z(n3696) );
  OAI21_X1 U4520 ( .B1(n3699), .B2(n4526), .A(n3696), .ZN(U3489) );
  MUX2_X1 U4521 ( .A(n4697), .B(n3697), .S(n4688), .Z(n3698) );
  OAI21_X1 U4522 ( .B1(n4470), .B2(n3699), .A(n3698), .ZN(U3529) );
  INV_X1 U4523 ( .A(n3701), .ZN(n3703) );
  NOR2_X1 U4524 ( .A1(n3703), .A2(n3702), .ZN(n4107) );
  INV_X1 U4525 ( .A(n4107), .ZN(n3704) );
  XNOR2_X1 U4526 ( .A(n3700), .B(n3704), .ZN(n3758) );
  NAND2_X1 U4527 ( .A1(n3705), .A2(n3713), .ZN(n3706) );
  NAND2_X1 U4528 ( .A1(n3707), .A2(n3706), .ZN(n3767) );
  INV_X1 U4529 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3710) );
  INV_X1 U4530 ( .A(n3708), .ZN(n3709) );
  OAI22_X1 U4531 ( .A1(n4544), .A2(n3710), .B1(n3709), .B2(n4300), .ZN(n3711)
         );
  AOI21_X1 U4532 ( .B1(n3712), .B2(n4163), .A(n3711), .ZN(n3715) );
  AOI22_X1 U4533 ( .A1(n4379), .A2(n3713), .B1(n4378), .B2(n4161), .ZN(n3714)
         );
  OAI211_X1 U4534 ( .C1(n3767), .C2(n4368), .A(n3715), .B(n3714), .ZN(n3718)
         );
  XNOR2_X1 U4535 ( .A(n3675), .B(n4107), .ZN(n3716) );
  NAND2_X1 U4536 ( .A1(n3716), .A2(n3121), .ZN(n3756) );
  NOR2_X1 U4537 ( .A1(n3756), .A2(n2160), .ZN(n3717) );
  AOI211_X1 U4538 ( .C1(n4318), .C2(n3758), .A(n3718), .B(n3717), .ZN(n3719)
         );
  INV_X1 U4539 ( .A(n3719), .ZN(U3278) );
  OAI211_X1 U4540 ( .C1(n3721), .C2(REG1_REG_14__SCAN_IN), .A(n4631), .B(n3720), .ZN(n3724) );
  AOI21_X1 U4541 ( .B1(n4630), .B2(ADDR_REG_14__SCAN_IN), .A(n3722), .ZN(n3723) );
  OAI211_X1 U4542 ( .C1(n4637), .C2(n3725), .A(n3724), .B(n3723), .ZN(n3728)
         );
  AOI211_X1 U4543 ( .C1(n4764), .C2(n2170), .A(n3726), .B(n4624), .ZN(n3727)
         );
  OR2_X1 U4544 ( .A1(n3728), .A2(n3727), .ZN(U3254) );
  INV_X1 U4545 ( .A(n3729), .ZN(n3731) );
  INV_X1 U4546 ( .A(n3778), .ZN(n3730) );
  OAI21_X1 U4547 ( .B1(n3731), .B2(n3734), .A(n3730), .ZN(n3743) );
  INV_X1 U4548 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3739) );
  XNOR2_X1 U4549 ( .A(n3732), .B(n4117), .ZN(n3752) );
  AOI22_X1 U4550 ( .A1(n4474), .A2(n4472), .B1(n4161), .B2(n4471), .ZN(n3733)
         );
  OAI21_X1 U4551 ( .B1(n3734), .B2(n4476), .A(n3733), .ZN(n3738) );
  AOI21_X1 U4552 ( .B1(n4117), .B2(n3736), .A(n2330), .ZN(n3754) );
  NOR2_X1 U4553 ( .A1(n3754), .A2(n4483), .ZN(n3737) );
  AOI211_X1 U4554 ( .C1(n3752), .C2(n3121), .A(n3738), .B(n3737), .ZN(n3741)
         );
  MUX2_X1 U4555 ( .A(n3739), .B(n3741), .S(n4688), .Z(n3740) );
  OAI21_X1 U4556 ( .B1(n4470), .B2(n3743), .A(n3740), .ZN(U3532) );
  MUX2_X1 U4557 ( .A(n4746), .B(n3741), .S(n4683), .Z(n3742) );
  OAI21_X1 U4558 ( .B1(n3743), .B2(n4526), .A(n3742), .ZN(U3495) );
  NOR2_X1 U4559 ( .A1(n3743), .A2(n4368), .ZN(n3750) );
  AOI22_X1 U4560 ( .A1(n3744), .A2(n4379), .B1(n4378), .B2(n4472), .ZN(n3747)
         );
  AOI22_X1 U4561 ( .A1(n2160), .A2(REG2_REG_14__SCAN_IN), .B1(n3745), .B2(
        n4645), .ZN(n3746) );
  OAI211_X1 U4562 ( .C1(n3748), .C2(n4383), .A(n3747), .B(n3746), .ZN(n3749)
         );
  AOI211_X1 U4563 ( .C1(n3752), .C2(n3751), .A(n3750), .B(n3749), .ZN(n3753)
         );
  OAI21_X1 U4564 ( .B1(n3754), .B2(n4391), .A(n3753), .ZN(U3276) );
  AOI22_X1 U4565 ( .A1(n4163), .A2(n4471), .B1(n4474), .B2(n4161), .ZN(n3755)
         );
  OAI211_X1 U4566 ( .C1(n4476), .C2(n2210), .A(n3756), .B(n3755), .ZN(n3757)
         );
  INV_X1 U4567 ( .A(n3757), .ZN(n3760) );
  NAND2_X1 U4568 ( .A1(n3758), .A2(n4676), .ZN(n3759) );
  NAND2_X1 U4569 ( .A1(n3760), .A2(n3759), .ZN(n3764) );
  INV_X1 U4570 ( .A(n3764), .ZN(n3761) );
  MUX2_X1 U4571 ( .A(n3762), .B(n3761), .S(n4683), .Z(n3763) );
  OAI21_X1 U4572 ( .B1(n3767), .B2(n4526), .A(n3763), .ZN(U3491) );
  MUX2_X1 U4573 ( .A(n3764), .B(REG1_REG_12__SCAN_IN), .S(n4686), .Z(n3765) );
  INV_X1 U4574 ( .A(n3765), .ZN(n3766) );
  OAI21_X1 U4575 ( .B1(n4470), .B2(n3767), .A(n3766), .ZN(U3530) );
  NAND2_X1 U4576 ( .A1(n3768), .A2(n4676), .ZN(n3770) );
  NAND2_X1 U4577 ( .A1(n3770), .A2(n3769), .ZN(n3773) );
  MUX2_X1 U4578 ( .A(REG1_REG_13__SCAN_IN), .B(n3773), .S(n4688), .Z(n3771) );
  INV_X1 U4579 ( .A(n3771), .ZN(n3772) );
  OAI21_X1 U4580 ( .B1(n4470), .B2(n3776), .A(n3772), .ZN(U3531) );
  MUX2_X1 U4581 ( .A(REG0_REG_13__SCAN_IN), .B(n3773), .S(n4683), .Z(n3774) );
  INV_X1 U4582 ( .A(n3774), .ZN(n3775) );
  OAI21_X1 U4583 ( .B1(n3776), .B2(n4526), .A(n3775), .ZN(U3493) );
  OAI21_X1 U4584 ( .B1(n3778), .B2(n3814), .A(n3777), .ZN(n3791) );
  XNOR2_X1 U4585 ( .A(n3779), .B(n2789), .ZN(n3801) );
  OAI22_X1 U4586 ( .A1(n3815), .A2(n4460), .B1(n4461), .B2(n4458), .ZN(n3780)
         );
  AOI21_X1 U4587 ( .B1(n3792), .B2(n4463), .A(n3780), .ZN(n3785) );
  AOI21_X1 U4588 ( .B1(n3782), .B2(n3781), .A(n4360), .ZN(n3784) );
  NAND2_X1 U4589 ( .A1(n3784), .A2(n3783), .ZN(n3796) );
  OAI211_X1 U4590 ( .C1(n3801), .C2(n4483), .A(n3785), .B(n3796), .ZN(n3786)
         );
  INV_X1 U4591 ( .A(n3786), .ZN(n3789) );
  MUX2_X1 U4592 ( .A(n3787), .B(n3789), .S(n4683), .Z(n3788) );
  OAI21_X1 U4593 ( .B1(n3791), .B2(n4526), .A(n3788), .ZN(U3497) );
  MUX2_X1 U4594 ( .A(n4699), .B(n3789), .S(n4688), .Z(n3790) );
  OAI21_X1 U4595 ( .B1(n4470), .B2(n3791), .A(n3790), .ZN(U3533) );
  INV_X1 U4596 ( .A(n3791), .ZN(n3799) );
  AOI22_X1 U4597 ( .A1(n4379), .A2(n3792), .B1(n4378), .B2(n3817), .ZN(n3795)
         );
  AOI22_X1 U4598 ( .A1(n2160), .A2(REG2_REG_15__SCAN_IN), .B1(n3793), .B2(
        n4645), .ZN(n3794) );
  OAI211_X1 U4599 ( .C1(n3815), .C2(n4383), .A(n3795), .B(n3794), .ZN(n3798)
         );
  NOR2_X1 U4600 ( .A1(n3796), .A2(n2160), .ZN(n3797) );
  AOI211_X1 U4601 ( .C1(n3799), .C2(n4647), .A(n3798), .B(n3797), .ZN(n3800)
         );
  OAI21_X1 U4602 ( .B1(n3801), .B2(n4391), .A(n3800), .ZN(U3275) );
  XNOR2_X1 U4603 ( .A(n3803), .B(n3802), .ZN(n3804) );
  XNOR2_X1 U4604 ( .A(n3805), .B(n3804), .ZN(n3809) );
  NOR2_X1 U4605 ( .A1(STATE_REG_SCAN_IN), .A2(n2675), .ZN(n4629) );
  OAI22_X1 U4606 ( .A1(n3981), .A2(n4461), .B1(n3980), .B2(n4375), .ZN(n3806)
         );
  AOI211_X1 U4607 ( .C1(n2193), .C2(n4377), .A(n4629), .B(n3806), .ZN(n3808)
         );
  NAND2_X1 U4608 ( .A1(n3986), .A2(n4380), .ZN(n3807) );
  OAI211_X1 U4609 ( .C1(n3809), .C2(n3988), .A(n3808), .B(n3807), .ZN(U3225)
         );
  NAND2_X1 U4610 ( .A1(n3810), .A2(n3811), .ZN(n3812) );
  XNOR2_X1 U4611 ( .A(n3812), .B(n3822), .ZN(n3813) );
  NAND2_X1 U4612 ( .A1(n3813), .A2(n3088), .ZN(n3819) );
  AND2_X1 U4613 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4608) );
  OAI22_X1 U4614 ( .A1(n3981), .A2(n3815), .B1(n3980), .B2(n3814), .ZN(n3816)
         );
  AOI211_X1 U4615 ( .C1(n2193), .C2(n3817), .A(n4608), .B(n3816), .ZN(n3818)
         );
  OAI211_X1 U4616 ( .C1(n3821), .C2(n3820), .A(n3819), .B(n3818), .ZN(U3238)
         );
  INV_X1 U4617 ( .A(n3810), .ZN(n3823) );
  OAI21_X1 U4618 ( .B1(n3823), .B2(n3822), .A(n3811), .ZN(n3824) );
  XOR2_X1 U4619 ( .A(n3825), .B(n3824), .Z(n3830) );
  AOI22_X1 U4620 ( .A1(n2193), .A2(n4473), .B1(n3847), .B2(n3928), .ZN(n3827)
         );
  INV_X1 U4621 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4936) );
  NOR2_X1 U4622 ( .A1(n4936), .A2(STATE_REG_SCAN_IN), .ZN(n4619) );
  INV_X1 U4623 ( .A(n4619), .ZN(n3826) );
  OAI211_X1 U4624 ( .C1(n3981), .C2(n3851), .A(n3827), .B(n3826), .ZN(n3828)
         );
  AOI21_X1 U4625 ( .B1(n3848), .B2(n3986), .A(n3828), .ZN(n3829) );
  OAI21_X1 U4626 ( .B1(n3830), .B2(n3988), .A(n3829), .ZN(U3223) );
  INV_X1 U4627 ( .A(n3831), .ZN(n3833) );
  NOR2_X1 U4628 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  XNOR2_X1 U4629 ( .A(n3835), .B(n3834), .ZN(n3841) );
  AOI22_X1 U4630 ( .A1(n3929), .A2(n4473), .B1(n3836), .B2(n3928), .ZN(n3838)
         );
  OAI211_X1 U4631 ( .C1(n3983), .C2(n4336), .A(n3838), .B(n3837), .ZN(n3839)
         );
  AOI21_X1 U4632 ( .B1(n3868), .B2(n3986), .A(n3839), .ZN(n3840) );
  OAI21_X1 U4633 ( .B1(n3841), .B2(n3988), .A(n3840), .ZN(U3235) );
  INV_X1 U4634 ( .A(n3842), .ZN(n3845) );
  INV_X1 U4635 ( .A(n4131), .ZN(n3844) );
  OR2_X1 U4636 ( .A1(n3842), .A2(n4131), .ZN(n3843) );
  OAI21_X1 U4637 ( .B1(n3845), .B2(n3844), .A(n3843), .ZN(n4484) );
  INV_X1 U4638 ( .A(n3846), .ZN(n4376) );
  AOI21_X1 U4639 ( .B1(n3847), .B2(n3777), .A(n4376), .ZN(n4480) );
  AOI22_X1 U4640 ( .A1(n3847), .A2(n4379), .B1(n4378), .B2(n4473), .ZN(n3850)
         );
  AOI22_X1 U4641 ( .A1(n2160), .A2(REG2_REG_16__SCAN_IN), .B1(n3848), .B2(
        n4645), .ZN(n3849) );
  OAI211_X1 U4642 ( .C1(n3851), .C2(n4383), .A(n3850), .B(n3849), .ZN(n3855)
         );
  OAI211_X1 U4643 ( .C1(n3853), .C2(n4131), .A(n3852), .B(n3121), .ZN(n4481)
         );
  NOR2_X1 U4644 ( .A1(n4481), .A2(n2160), .ZN(n3854) );
  AOI211_X1 U4645 ( .C1(n4480), .C2(n4647), .A(n3855), .B(n3854), .ZN(n3856)
         );
  OAI21_X1 U4646 ( .B1(n4391), .B2(n4484), .A(n3856), .ZN(U3274) );
  INV_X1 U4647 ( .A(n4104), .ZN(n3858) );
  OAI21_X1 U4648 ( .B1(n3857), .B2(n3858), .A(n4105), .ZN(n4354) );
  INV_X1 U4649 ( .A(n3864), .ZN(n4121) );
  XNOR2_X1 U4650 ( .A(n4354), .B(n4121), .ZN(n3862) );
  AOI22_X1 U4651 ( .A1(n4474), .A2(n3859), .B1(n4473), .B2(n4471), .ZN(n3860)
         );
  OAI21_X1 U4652 ( .B1(n3867), .B2(n4476), .A(n3860), .ZN(n3861) );
  AOI21_X1 U4653 ( .B1(n3862), .B2(n3121), .A(n3861), .ZN(n4456) );
  OAI21_X1 U4654 ( .B1(n3865), .B2(n3864), .A(n3863), .ZN(n4454) );
  INV_X1 U4655 ( .A(n4363), .ZN(n3866) );
  OAI211_X1 U4656 ( .C1(n4373), .C2(n3867), .A(n3866), .B(n4479), .ZN(n4455)
         );
  AOI22_X1 U4657 ( .A1(n2160), .A2(REG2_REG_18__SCAN_IN), .B1(n3868), .B2(
        n4645), .ZN(n3869) );
  OAI21_X1 U4658 ( .B1(n4455), .B2(n3870), .A(n3869), .ZN(n3871) );
  AOI21_X1 U4659 ( .B1(n4454), .B2(n4318), .A(n3871), .ZN(n3872) );
  OAI21_X1 U4660 ( .B1(n2160), .B2(n4456), .A(n3872), .ZN(U3272) );
  INV_X1 U4661 ( .A(D_REG_0__SCAN_IN), .ZN(n3874) );
  NOR3_X1 U4662 ( .A1(n4530), .A2(n2815), .A3(n4655), .ZN(n3873) );
  AOI21_X1 U4663 ( .B1(n4654), .B2(n3874), .A(n3873), .ZN(U3458) );
  XOR2_X1 U4664 ( .A(n3876), .B(n3875), .Z(n3877) );
  XNOR2_X1 U4665 ( .A(n3878), .B(n3877), .ZN(n3885) );
  NOR2_X1 U4666 ( .A1(STATE_REG_SCAN_IN), .A2(n2643), .ZN(n4596) );
  OAI22_X1 U4667 ( .A1(n3981), .A2(n3879), .B1(n3980), .B2(n2208), .ZN(n3880)
         );
  AOI211_X1 U4668 ( .C1(n2193), .C2(n4160), .A(n4596), .B(n3880), .ZN(n3884)
         );
  NAND2_X1 U4669 ( .A1(n3986), .A2(n3882), .ZN(n3883) );
  OAI211_X1 U4670 ( .C1(n3885), .C2(n3988), .A(n3884), .B(n3883), .ZN(U3231)
         );
  INV_X1 U4671 ( .A(n3919), .ZN(n3887) );
  AOI21_X1 U4672 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n3894) );
  INV_X1 U4673 ( .A(n4301), .ZN(n3892) );
  OAI22_X1 U4674 ( .A1(n3983), .A2(n3956), .B1(STATE_REG_SCAN_IN), .B2(n4728), 
        .ZN(n3891) );
  OAI22_X1 U4675 ( .A1(n3981), .A2(n3969), .B1(n3980), .B2(n4298), .ZN(n3890)
         );
  AOI211_X1 U4676 ( .C1(n3892), .C2(n3986), .A(n3891), .B(n3890), .ZN(n3893)
         );
  OAI21_X1 U4677 ( .B1(n3894), .B2(n3988), .A(n3893), .ZN(U3232) );
  NOR2_X1 U4678 ( .A1(n3895), .A2(n4368), .ZN(n3903) );
  INV_X1 U4679 ( .A(n3896), .ZN(n3897) );
  AOI22_X1 U4680 ( .A1(n3897), .A2(n4645), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2160), .ZN(n3901) );
  AOI22_X1 U4681 ( .A1(n3899), .A2(n4378), .B1(n4379), .B2(n3898), .ZN(n3900)
         );
  OAI211_X1 U4682 ( .C1(n4231), .C2(n4383), .A(n3901), .B(n3900), .ZN(n3902)
         );
  OAI21_X1 U4683 ( .B1(n3906), .B2(n4391), .A(n3905), .ZN(U3262) );
  XNOR2_X1 U4684 ( .A(n3909), .B(n3908), .ZN(n3915) );
  INV_X1 U4685 ( .A(n4211), .ZN(n3913) );
  OAI22_X1 U4686 ( .A1(n3981), .A2(n4421), .B1(n3980), .B2(n4212), .ZN(n3912)
         );
  INV_X1 U4687 ( .A(n4158), .ZN(n4408) );
  OAI22_X1 U4688 ( .A1(n4408), .A2(n3983), .B1(STATE_REG_SCAN_IN), .B2(n3910), 
        .ZN(n3911) );
  AOI211_X1 U4689 ( .C1(n3913), .C2(n3986), .A(n3912), .B(n3911), .ZN(n3914)
         );
  OAI21_X1 U4690 ( .B1(n3915), .B2(n3988), .A(n3914), .ZN(U3211) );
  NAND2_X1 U4691 ( .A1(n3916), .A2(n3088), .ZN(n3925) );
  AOI21_X1 U4692 ( .B1(n3919), .B2(n3918), .A(n3917), .ZN(n3924) );
  INV_X1 U4693 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3920) );
  OAI22_X1 U4694 ( .A1(n3983), .A2(n4288), .B1(STATE_REG_SCAN_IN), .B2(n3920), 
        .ZN(n3922) );
  OAI22_X1 U4695 ( .A1(n3981), .A2(n2723), .B1(n3980), .B2(n4290), .ZN(n3921)
         );
  AOI211_X1 U4696 ( .C1(n4291), .C2(n3986), .A(n3922), .B(n3921), .ZN(n3923)
         );
  OAI21_X1 U4697 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(U3213) );
  XOR2_X1 U4698 ( .A(n3927), .B(n3926), .Z(n3933) );
  AOI22_X1 U4699 ( .A1(n3929), .A2(n4377), .B1(n4358), .B2(n3928), .ZN(n3930)
         );
  NAND2_X1 U4700 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4189) );
  OAI211_X1 U4701 ( .C1(n3983), .C2(n4441), .A(n3930), .B(n4189), .ZN(n3931)
         );
  AOI21_X1 U4702 ( .B1(n4366), .B2(n3986), .A(n3931), .ZN(n3932) );
  OAI21_X1 U4703 ( .B1(n3933), .B2(n3988), .A(n3932), .ZN(U3216) );
  XNOR2_X1 U4704 ( .A(n3935), .B(n3934), .ZN(n3936) );
  XNOR2_X1 U4705 ( .A(n3937), .B(n3936), .ZN(n3942) );
  OAI22_X1 U4706 ( .A1(n3983), .A2(n2723), .B1(STATE_REG_SCAN_IN), .B2(n3938), 
        .ZN(n3940) );
  OAI22_X1 U4707 ( .A1(n3981), .A2(n4441), .B1(n3980), .B2(n4322), .ZN(n3939)
         );
  AOI211_X1 U4708 ( .C1(n4324), .C2(n3986), .A(n3940), .B(n3939), .ZN(n3941)
         );
  OAI21_X1 U4709 ( .B1(n3942), .B2(n3988), .A(n3941), .ZN(U3220) );
  NAND2_X1 U4710 ( .A1(n3944), .A2(n3943), .ZN(n3946) );
  XOR2_X1 U4711 ( .A(n3946), .B(n3945), .Z(n3950) );
  INV_X1 U4712 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4720) );
  OAI22_X1 U4713 ( .A1(n3983), .A2(n4421), .B1(STATE_REG_SCAN_IN), .B2(n4720), 
        .ZN(n3948) );
  OAI22_X1 U4714 ( .A1(n3981), .A2(n4288), .B1(n3980), .B2(n4246), .ZN(n3947)
         );
  AOI211_X1 U4715 ( .C1(n4248), .C2(n3986), .A(n3948), .B(n3947), .ZN(n3949)
         );
  OAI21_X1 U4716 ( .B1(n3950), .B2(n3988), .A(n3949), .ZN(U3222) );
  NAND2_X1 U4717 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  XOR2_X1 U4718 ( .A(n3954), .B(n3953), .Z(n3961) );
  INV_X1 U4719 ( .A(n4269), .ZN(n3959) );
  INV_X1 U4720 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3955) );
  OAI22_X1 U4721 ( .A1(n3983), .A2(n4221), .B1(STATE_REG_SCAN_IN), .B2(n3955), 
        .ZN(n3958) );
  OAI22_X1 U4722 ( .A1(n3981), .A2(n3956), .B1(n3980), .B2(n4267), .ZN(n3957)
         );
  AOI211_X1 U4723 ( .C1(n3959), .C2(n3986), .A(n3958), .B(n3957), .ZN(n3960)
         );
  OAI21_X1 U4724 ( .B1(n3961), .B2(n3988), .A(n3960), .ZN(U3226) );
  INV_X1 U4725 ( .A(n3962), .ZN(n3967) );
  AOI21_X1 U4726 ( .B1(n3966), .B2(n3964), .A(n3963), .ZN(n3965) );
  AOI21_X1 U4727 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n3974) );
  INV_X1 U4728 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3968) );
  OAI22_X1 U4729 ( .A1(n3983), .A2(n3969), .B1(STATE_REG_SCAN_IN), .B2(n3968), 
        .ZN(n3972) );
  OAI22_X1 U4730 ( .A1(n3981), .A2(n4336), .B1(n3980), .B2(n3970), .ZN(n3971)
         );
  AOI211_X1 U4731 ( .C1(n4343), .C2(n3986), .A(n3972), .B(n3971), .ZN(n3973)
         );
  OAI21_X1 U4732 ( .B1(n3974), .B2(n3988), .A(n3973), .ZN(U3230) );
  INV_X1 U4733 ( .A(n3975), .ZN(n3977) );
  NOR2_X1 U4734 ( .A1(n3977), .A2(n3976), .ZN(n3978) );
  XNOR2_X1 U4735 ( .A(n3979), .B(n3978), .ZN(n3989) );
  OAI22_X1 U4736 ( .A1(n3981), .A2(n4221), .B1(n3980), .B2(n4234), .ZN(n3985)
         );
  OAI22_X1 U4737 ( .A1(n3983), .A2(n4231), .B1(STATE_REG_SCAN_IN), .B2(n3982), 
        .ZN(n3984) );
  AOI211_X1 U4738 ( .C1(n4236), .C2(n3986), .A(n3985), .B(n3984), .ZN(n3987)
         );
  OAI21_X1 U4739 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(U3237) );
  AND2_X1 U4740 ( .A1(n4122), .A2(n4109), .ZN(n4010) );
  NAND2_X1 U4741 ( .A1(n3990), .A2(n3993), .ZN(n4067) );
  NAND2_X1 U4742 ( .A1(n3992), .A2(n3991), .ZN(n4055) );
  NAND2_X1 U4743 ( .A1(n4055), .A2(n3993), .ZN(n4058) );
  OAI21_X1 U4744 ( .B1(n3732), .B2(n4067), .A(n4058), .ZN(n3995) );
  INV_X1 U4745 ( .A(n4074), .ZN(n3994) );
  AOI211_X1 U4746 ( .C1(n3995), .C2(n4077), .A(n3994), .B(n4076), .ZN(n3997)
         );
  OAI21_X1 U4747 ( .B1(n3997), .B2(n2299), .A(n4079), .ZN(n3998) );
  AND2_X1 U4748 ( .A1(n3998), .A2(n4083), .ZN(n4000) );
  OAI21_X1 U4749 ( .B1(n4000), .B2(n3999), .A(n4084), .ZN(n4009) );
  NAND2_X1 U4750 ( .A1(n2164), .A2(DATAI_31_), .ZN(n4394) );
  INV_X1 U4751 ( .A(n4394), .ZN(n4024) );
  INV_X1 U4752 ( .A(n4392), .ZN(n4002) );
  INV_X1 U4753 ( .A(n4157), .ZN(n4001) );
  AND2_X1 U4754 ( .A1(n2164), .A2(DATAI_30_), .ZN(n4399) );
  NAND2_X1 U4755 ( .A1(n4001), .A2(n4399), .ZN(n4129) );
  OAI21_X1 U4756 ( .B1(n4024), .B2(n4002), .A(n4129), .ZN(n4003) );
  NOR2_X1 U4757 ( .A1(n4004), .A2(n4003), .ZN(n4018) );
  INV_X1 U4758 ( .A(n4018), .ZN(n4008) );
  AND2_X1 U4759 ( .A1(n4005), .A2(n4123), .ZN(n4091) );
  NAND3_X1 U4760 ( .A1(n4091), .A2(n4014), .A3(n4006), .ZN(n4007) );
  AOI211_X1 U4761 ( .C1(n4010), .C2(n4009), .A(n4008), .B(n4007), .ZN(n4022)
         );
  NOR3_X1 U4762 ( .A1(n4013), .A2(n4012), .A3(n4011), .ZN(n4087) );
  NOR2_X1 U4763 ( .A1(n2279), .A2(n4015), .ZN(n4020) );
  NAND2_X1 U4764 ( .A1(n4017), .A2(n4016), .ZN(n4019) );
  OAI21_X1 U4765 ( .B1(n4020), .B2(n4019), .A(n4018), .ZN(n4092) );
  AOI21_X1 U4766 ( .B1(n4208), .B2(n4087), .A(n4092), .ZN(n4021) );
  INV_X1 U4767 ( .A(n4399), .ZN(n4023) );
  OAI22_X1 U4768 ( .A1(n4022), .A2(n4021), .B1(n4392), .B2(n4023), .ZN(n4027)
         );
  NAND2_X1 U4769 ( .A1(n4023), .A2(n4157), .ZN(n4130) );
  NAND2_X1 U4770 ( .A1(n4130), .A2(n4392), .ZN(n4025) );
  NAND2_X1 U4771 ( .A1(n4025), .A2(n4024), .ZN(n4094) );
  AOI21_X1 U4772 ( .B1(n4027), .B2(n4094), .A(n4026), .ZN(n4147) );
  INV_X1 U4773 ( .A(n4028), .ZN(n4030) );
  OAI211_X1 U4774 ( .C1(n4532), .C2(n4031), .A(n4030), .B(n4029), .ZN(n4034)
         );
  NAND3_X1 U4775 ( .A1(n4034), .A2(n4033), .A3(n4032), .ZN(n4037) );
  NAND3_X1 U4776 ( .A1(n4037), .A2(n4036), .A3(n4035), .ZN(n4040) );
  NAND3_X1 U4777 ( .A1(n4040), .A2(n4039), .A3(n4038), .ZN(n4042) );
  NAND4_X1 U4778 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4051), .ZN(n4045)
         );
  NAND3_X1 U4779 ( .A1(n4045), .A2(n4126), .A3(n4044), .ZN(n4046) );
  NAND3_X1 U4780 ( .A1(n4046), .A2(n4053), .A3(n4052), .ZN(n4049) );
  AND3_X1 U4781 ( .A1(n4049), .A2(n4048), .A3(n4047), .ZN(n4056) );
  INV_X1 U4782 ( .A(n4058), .ZN(n4071) );
  NAND4_X1 U4783 ( .A1(n2306), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4054)
         );
  OAI22_X1 U4784 ( .A1(n4056), .A2(n4055), .B1(n4071), .B2(n4054), .ZN(n4061)
         );
  INV_X1 U4785 ( .A(n4057), .ZN(n4059) );
  AOI22_X1 U4786 ( .A1(n4061), .A2(n4060), .B1(n4059), .B2(n4058), .ZN(n4073)
         );
  NAND3_X1 U4787 ( .A1(n4068), .A2(n4063), .A3(n4062), .ZN(n4072) );
  INV_X1 U4788 ( .A(n4064), .ZN(n4069) );
  INV_X1 U4789 ( .A(n4065), .ZN(n4066) );
  AOI211_X1 U4790 ( .C1(n4069), .C2(n4068), .A(n4067), .B(n4066), .ZN(n4070)
         );
  OAI22_X1 U4791 ( .A1(n4073), .A2(n4072), .B1(n4071), .B2(n4070), .ZN(n4075)
         );
  NAND2_X1 U4792 ( .A1(n4075), .A2(n4074), .ZN(n4078) );
  AOI21_X1 U4793 ( .B1(n4078), .B2(n4077), .A(n4076), .ZN(n4080) );
  INV_X1 U4794 ( .A(n4277), .ZN(n4128) );
  OAI211_X1 U4795 ( .C1(n4080), .C2(n2299), .A(n4128), .B(n4079), .ZN(n4082)
         );
  AOI21_X1 U4796 ( .B1(n4083), .B2(n4082), .A(n4081), .ZN(n4086) );
  INV_X1 U4797 ( .A(n4084), .ZN(n4085) );
  OAI211_X1 U4798 ( .C1(n4086), .C2(n4085), .A(n4122), .B(n4109), .ZN(n4090)
         );
  NOR2_X1 U4799 ( .A1(n4231), .A2(n4404), .ZN(n4089) );
  INV_X1 U4800 ( .A(n4087), .ZN(n4088) );
  AOI211_X1 U4801 ( .C1(n4091), .C2(n4090), .A(n4089), .B(n4088), .ZN(n4093)
         );
  OR2_X1 U4802 ( .A1(n4093), .A2(n4092), .ZN(n4095) );
  OAI211_X1 U4803 ( .C1(n4130), .C2(n4392), .A(n4095), .B(n4094), .ZN(n4145)
         );
  INV_X1 U4804 ( .A(n4208), .ZN(n4097) );
  XNOR2_X1 U4805 ( .A(n4336), .B(n4358), .ZN(n4356) );
  NOR4_X1 U4806 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4356), .ZN(n4142)
         );
  INV_X1 U4807 ( .A(n4099), .ZN(n4101) );
  NAND2_X1 U4808 ( .A1(n4101), .A2(n4100), .ZN(n4223) );
  INV_X1 U4809 ( .A(n4223), .ZN(n4225) );
  NAND2_X1 U4810 ( .A1(n4256), .A2(n4102), .ZN(n4282) );
  NOR2_X1 U4811 ( .A1(n4225), .A2(n4282), .ZN(n4115) );
  XNOR2_X1 U4812 ( .A(n4103), .B(n4344), .ZN(n4338) );
  AND2_X1 U4813 ( .A1(n4105), .A2(n4104), .ZN(n4384) );
  AND4_X1 U4814 ( .A1(n4107), .A2(n4106), .A3(n4305), .A4(n4384), .ZN(n4114)
         );
  NAND2_X1 U4815 ( .A1(n4109), .A2(n4108), .ZN(n4258) );
  NOR4_X1 U4816 ( .A1(n4258), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4113)
         );
  NAND4_X1 U4817 ( .A1(n4115), .A2(n4338), .A3(n4114), .A4(n4113), .ZN(n4140)
         );
  NAND4_X1 U4818 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4139)
         );
  NAND4_X1 U4819 ( .A1(n4121), .A2(n2789), .A3(n4120), .A4(n3390), .ZN(n4138)
         );
  NAND2_X1 U4820 ( .A1(n4123), .A2(n4122), .ZN(n4243) );
  INV_X1 U4821 ( .A(n4243), .ZN(n4127) );
  XOR2_X1 U4822 ( .A(n4394), .B(n4392), .Z(n4124) );
  NAND4_X1 U4823 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4136)
         );
  NAND2_X1 U4824 ( .A1(n4128), .A2(n4278), .ZN(n4317) );
  INV_X1 U4825 ( .A(n4317), .ZN(n4132) );
  NAND4_X1 U4826 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4134)
         );
  OR4_X1 U4827 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137) );
  NOR4_X1 U4828 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  AOI21_X1 U4829 ( .B1(n4142), .B2(n4141), .A(n4532), .ZN(n4144) );
  MUX2_X1 U4830 ( .A(n4145), .B(n4144), .S(n4143), .Z(n4146) );
  NOR2_X1 U4831 ( .A1(n4147), .A2(n4146), .ZN(n4148) );
  XNOR2_X1 U4832 ( .A(n4148), .B(n4533), .ZN(n4156) );
  INV_X1 U4833 ( .A(B_REG_SCAN_IN), .ZN(n4727) );
  AOI21_X1 U4834 ( .B1(n4150), .B2(n4149), .A(n4727), .ZN(n4151) );
  OAI21_X1 U4835 ( .B1(n4153), .B2(n4152), .A(n4151), .ZN(n4154) );
  OAI21_X1 U4836 ( .B1(n4156), .B2(n4155), .A(n4154), .ZN(U3239) );
  MUX2_X1 U4837 ( .A(DATAO_REG_30__SCAN_IN), .B(n4157), .S(n4166), .Z(U3580)
         );
  MUX2_X1 U4838 ( .A(DATAO_REG_28__SCAN_IN), .B(n4158), .S(n4166), .Z(U3578)
         );
  MUX2_X1 U4839 ( .A(DATAO_REG_27__SCAN_IN), .B(n4159), .S(n4166), .Z(U3577)
         );
  MUX2_X1 U4840 ( .A(DATAO_REG_21__SCAN_IN), .B(n4334), .S(n4166), .Z(U3571)
         );
  MUX2_X1 U4841 ( .A(DATAO_REG_17__SCAN_IN), .B(n4473), .S(n4166), .Z(U3567)
         );
  MUX2_X1 U4842 ( .A(DATAO_REG_14__SCAN_IN), .B(n4160), .S(n4166), .Z(U3564)
         );
  MUX2_X1 U4843 ( .A(DATAO_REG_13__SCAN_IN), .B(n4161), .S(n4166), .Z(U3563)
         );
  MUX2_X1 U4844 ( .A(DATAO_REG_12__SCAN_IN), .B(n4162), .S(n4166), .Z(U3562)
         );
  MUX2_X1 U4845 ( .A(DATAO_REG_11__SCAN_IN), .B(n4163), .S(n4166), .Z(U3561)
         );
  MUX2_X1 U4846 ( .A(DATAO_REG_7__SCAN_IN), .B(n4164), .S(n4166), .Z(U3557) );
  MUX2_X1 U4847 ( .A(DATAO_REG_3__SCAN_IN), .B(n4165), .S(n4166), .Z(U3553) );
  MUX2_X1 U4848 ( .A(DATAO_REG_1__SCAN_IN), .B(n2850), .S(n4166), .Z(U3551) );
  MUX2_X1 U4849 ( .A(DATAO_REG_0__SCAN_IN), .B(n4167), .S(n4166), .Z(U3550) );
  NAND2_X1 U4850 ( .A1(n4168), .A2(n2482), .ZN(n4178) );
  OAI211_X1 U4851 ( .C1(n4171), .C2(n4170), .A(n4631), .B(n4169), .ZN(n4177)
         );
  OAI211_X1 U4852 ( .C1(n4174), .C2(n4173), .A(n4592), .B(n4172), .ZN(n4176)
         );
  AOI22_X1 U4853 ( .A1(n4630), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4175) );
  NAND4_X1 U4854 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(U3241)
         );
  AOI22_X1 U4855 ( .A1(n4180), .A2(n4179), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4185), .ZN(n4183) );
  INV_X1 U4856 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4181) );
  MUX2_X1 U4857 ( .A(n4181), .B(REG1_REG_19__SCAN_IN), .S(n4533), .Z(n4182) );
  XNOR2_X1 U4858 ( .A(n4183), .B(n4182), .ZN(n4195) );
  INV_X1 U4859 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4186) );
  MUX2_X1 U4860 ( .A(REG2_REG_19__SCAN_IN), .B(n4186), .S(n4533), .Z(n4187) );
  NAND2_X1 U4861 ( .A1(n4630), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4188) );
  OAI211_X1 U4862 ( .C1(n4637), .C2(n4190), .A(n4189), .B(n4188), .ZN(n4191)
         );
  AOI21_X1 U4863 ( .B1(n4192), .B2(n4592), .A(n4191), .ZN(n4193) );
  OAI21_X1 U4864 ( .B1(n4195), .B2(n4194), .A(n4193), .ZN(U3259) );
  INV_X1 U4865 ( .A(n4196), .ZN(n4204) );
  INV_X1 U4866 ( .A(n4197), .ZN(n4198) );
  OAI22_X1 U4867 ( .A1(n4199), .A2(n4368), .B1(n4198), .B2(n4300), .ZN(n4200)
         );
  OAI21_X1 U4868 ( .B1(n4201), .B2(n4200), .A(n4544), .ZN(n4203) );
  NAND2_X1 U4869 ( .A1(n2160), .A2(REG2_REG_29__SCAN_IN), .ZN(n4202) );
  OAI211_X1 U4870 ( .C1(n4204), .C2(n4391), .A(n4203), .B(n4202), .ZN(U3354)
         );
  XNOR2_X1 U4871 ( .A(n4205), .B(n4208), .ZN(n4206) );
  NAND2_X1 U4872 ( .A1(n4206), .A2(n3121), .ZN(n4407) );
  XOR2_X1 U4873 ( .A(n4208), .B(n4207), .Z(n4410) );
  NAND2_X1 U4874 ( .A1(n4410), .A2(n4318), .ZN(n4220) );
  INV_X1 U4875 ( .A(n3130), .ZN(n4209) );
  OAI21_X1 U4876 ( .B1(n4232), .B2(n4212), .A(n4209), .ZN(n4494) );
  NOR2_X1 U4877 ( .A1(n4494), .A2(n4368), .ZN(n4218) );
  NOR2_X1 U4878 ( .A1(n4421), .A2(n4383), .ZN(n4217) );
  INV_X1 U4879 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4210) );
  OAI22_X1 U4880 ( .A1(n4211), .A2(n4300), .B1(n4544), .B2(n4210), .ZN(n4216)
         );
  OAI22_X1 U4881 ( .A1(n4408), .A2(n4214), .B1(n4213), .B2(n4212), .ZN(n4215)
         );
  NOR4_X1 U4882 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4219)
         );
  OAI211_X1 U4883 ( .C1(n2160), .C2(n4407), .A(n4220), .B(n4219), .ZN(U3263)
         );
  OAI22_X1 U4884 ( .A1(n4244), .A2(n4222), .B1(n4221), .B2(n4246), .ZN(n4224)
         );
  XNOR2_X1 U4885 ( .A(n4224), .B(n4223), .ZN(n4414) );
  INV_X1 U4886 ( .A(n4414), .ZN(n4240) );
  XNOR2_X1 U4887 ( .A(n4226), .B(n4225), .ZN(n4227) );
  NAND2_X1 U4888 ( .A1(n4227), .A2(n3121), .ZN(n4230) );
  AOI22_X1 U4889 ( .A1(n4261), .A2(n4471), .B1(n4228), .B2(n4463), .ZN(n4229)
         );
  OAI211_X1 U4890 ( .C1(n4231), .C2(n4458), .A(n4230), .B(n4229), .ZN(n4413)
         );
  INV_X1 U4891 ( .A(n4245), .ZN(n4235) );
  INV_X1 U4892 ( .A(n4232), .ZN(n4233) );
  OAI21_X1 U4893 ( .B1(n4235), .B2(n4234), .A(n4233), .ZN(n4497) );
  AOI22_X1 U4894 ( .A1(n2160), .A2(REG2_REG_26__SCAN_IN), .B1(n4236), .B2(
        n4645), .ZN(n4237) );
  OAI21_X1 U4895 ( .B1(n4497), .B2(n4368), .A(n4237), .ZN(n4238) );
  AOI21_X1 U4896 ( .B1(n4413), .B2(n4544), .A(n4238), .ZN(n4239) );
  OAI21_X1 U4897 ( .B1(n4240), .B2(n4391), .A(n4239), .ZN(U3264) );
  XNOR2_X1 U4898 ( .A(n4241), .B(n4243), .ZN(n4242) );
  NAND2_X1 U4899 ( .A1(n4242), .A2(n3121), .ZN(n4420) );
  XNOR2_X1 U4900 ( .A(n4244), .B(n4243), .ZN(n4423) );
  NAND2_X1 U4901 ( .A1(n4423), .A2(n4318), .ZN(n4254) );
  INV_X1 U4902 ( .A(n4266), .ZN(n4247) );
  OAI21_X1 U4903 ( .B1(n4247), .B2(n4246), .A(n4245), .ZN(n4501) );
  INV_X1 U4904 ( .A(n4501), .ZN(n4252) );
  AOI22_X1 U4905 ( .A1(n4379), .A2(n4417), .B1(n4378), .B2(n4405), .ZN(n4250)
         );
  AOI22_X1 U4906 ( .A1(n2160), .A2(REG2_REG_25__SCAN_IN), .B1(n4248), .B2(
        n4645), .ZN(n4249) );
  OAI211_X1 U4907 ( .C1(n4288), .C2(n4383), .A(n4250), .B(n4249), .ZN(n4251)
         );
  AOI21_X1 U4908 ( .B1(n4252), .B2(n4647), .A(n4251), .ZN(n4253) );
  OAI211_X1 U4909 ( .C1(n2160), .C2(n4420), .A(n4254), .B(n4253), .ZN(U3265)
         );
  XOR2_X1 U4910 ( .A(n4258), .B(n4255), .Z(n4427) );
  INV_X1 U4911 ( .A(n4427), .ZN(n4274) );
  NAND2_X1 U4912 ( .A1(n4257), .A2(n4256), .ZN(n4259) );
  XNOR2_X1 U4913 ( .A(n4259), .B(n4258), .ZN(n4264) );
  NOR2_X1 U4914 ( .A1(n4267), .A2(n4476), .ZN(n4260) );
  AOI21_X1 U4915 ( .B1(n4261), .B2(n4474), .A(n4260), .ZN(n4263) );
  NAND2_X1 U4916 ( .A1(n4307), .A2(n4471), .ZN(n4262) );
  OAI211_X1 U4917 ( .C1(n4264), .C2(n4360), .A(n4263), .B(n4262), .ZN(n4426)
         );
  INV_X1 U4918 ( .A(n4265), .ZN(n4268) );
  OAI21_X1 U4919 ( .B1(n4268), .B2(n4267), .A(n4266), .ZN(n4504) );
  NOR2_X1 U4920 ( .A1(n4504), .A2(n4368), .ZN(n4272) );
  INV_X1 U4921 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4270) );
  OAI22_X1 U4922 ( .A1(n4544), .A2(n4270), .B1(n4269), .B2(n4300), .ZN(n4271)
         );
  AOI211_X1 U4923 ( .C1(n4426), .C2(n4544), .A(n4272), .B(n4271), .ZN(n4273)
         );
  OAI21_X1 U4924 ( .B1(n4274), .B2(n4391), .A(n4273), .ZN(U3266) );
  XNOR2_X1 U4925 ( .A(n4275), .B(n4282), .ZN(n4430) );
  INV_X1 U4926 ( .A(n4430), .ZN(n4295) );
  OR2_X1 U4927 ( .A1(n4276), .A2(n4277), .ZN(n4279) );
  NAND2_X1 U4928 ( .A1(n4279), .A2(n4278), .ZN(n4306) );
  INV_X1 U4929 ( .A(n4280), .ZN(n4281) );
  AOI21_X1 U4930 ( .B1(n4306), .B2(n4305), .A(n4281), .ZN(n4283) );
  XNOR2_X1 U4931 ( .A(n4283), .B(n4282), .ZN(n4284) );
  NAND2_X1 U4932 ( .A1(n4284), .A2(n3121), .ZN(n4287) );
  AOI22_X1 U4933 ( .A1(n4438), .A2(n4471), .B1(n4463), .B2(n4285), .ZN(n4286)
         );
  OAI211_X1 U4934 ( .C1(n4288), .C2(n4458), .A(n4287), .B(n4286), .ZN(n4429)
         );
  OAI21_X1 U4935 ( .B1(n4289), .B2(n4290), .A(n4265), .ZN(n4508) );
  AOI22_X1 U4936 ( .A1(n2160), .A2(REG2_REG_23__SCAN_IN), .B1(n4291), .B2(
        n4645), .ZN(n4292) );
  OAI21_X1 U4937 ( .B1(n4508), .B2(n4368), .A(n4292), .ZN(n4293) );
  AOI21_X1 U4938 ( .B1(n4429), .B2(n4544), .A(n4293), .ZN(n4294) );
  OAI21_X1 U4939 ( .B1(n4295), .B2(n4391), .A(n4294), .ZN(U3267) );
  AND2_X1 U4940 ( .A1(n4296), .A2(n4305), .ZN(n4297) );
  OR2_X1 U4941 ( .A1(n4297), .A2(n2183), .ZN(n4434) );
  NOR2_X1 U4942 ( .A1(n4320), .A2(n4298), .ZN(n4299) );
  OR2_X1 U4943 ( .A1(n4289), .A2(n4299), .ZN(n4512) );
  INV_X1 U4944 ( .A(n4512), .ZN(n4304) );
  INV_X1 U4945 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4302) );
  OAI22_X1 U4946 ( .A1(n4544), .A2(n4302), .B1(n4301), .B2(n4300), .ZN(n4303)
         );
  AOI21_X1 U4947 ( .B1(n4304), .B2(n4647), .A(n4303), .ZN(n4314) );
  XNOR2_X1 U4948 ( .A(n4306), .B(n4305), .ZN(n4312) );
  NAND2_X1 U4949 ( .A1(n4307), .A2(n4474), .ZN(n4310) );
  AOI22_X1 U4950 ( .A1(n4334), .A2(n4471), .B1(n4308), .B2(n4463), .ZN(n4309)
         );
  NAND2_X1 U4951 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  AOI21_X1 U4952 ( .B1(n4312), .B2(n3121), .A(n4311), .ZN(n4433) );
  OR2_X1 U4953 ( .A1(n4433), .A2(n2160), .ZN(n4313) );
  OAI211_X1 U4954 ( .C1(n4434), .C2(n4391), .A(n4314), .B(n4313), .ZN(U3268)
         );
  XNOR2_X1 U4955 ( .A(n4276), .B(n4317), .ZN(n4315) );
  NAND2_X1 U4956 ( .A1(n4315), .A2(n3121), .ZN(n4440) );
  XOR2_X1 U4957 ( .A(n4317), .B(n4316), .Z(n4443) );
  NAND2_X1 U4958 ( .A1(n4443), .A2(n4318), .ZN(n4330) );
  INV_X1 U4959 ( .A(n4319), .ZN(n4323) );
  INV_X1 U4960 ( .A(n4320), .ZN(n4321) );
  OAI21_X1 U4961 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4516) );
  INV_X1 U4962 ( .A(n4516), .ZN(n4328) );
  AOI22_X1 U4963 ( .A1(n4379), .A2(n4437), .B1(n4378), .B2(n4438), .ZN(n4326)
         );
  AOI22_X1 U4964 ( .A1(n2160), .A2(REG2_REG_21__SCAN_IN), .B1(n4324), .B2(
        n4645), .ZN(n4325) );
  OAI211_X1 U4965 ( .C1(n4441), .C2(n4383), .A(n4326), .B(n4325), .ZN(n4327)
         );
  AOI21_X1 U4966 ( .B1(n4328), .B2(n4647), .A(n4327), .ZN(n4329) );
  OAI211_X1 U4967 ( .C1(n2160), .C2(n4440), .A(n4330), .B(n4329), .ZN(U3269)
         );
  NAND2_X1 U4968 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  XNOR2_X1 U4969 ( .A(n4333), .B(n4338), .ZN(n4342) );
  AOI22_X1 U4970 ( .A1(n4334), .A2(n4474), .B1(n4463), .B2(n4344), .ZN(n4335)
         );
  OAI21_X1 U4971 ( .B1(n4336), .B2(n4460), .A(n4335), .ZN(n4341) );
  XNOR2_X1 U4972 ( .A(n4337), .B(n4338), .ZN(n4450) );
  NOR2_X1 U4973 ( .A1(n4450), .A2(n4339), .ZN(n4340) );
  AOI211_X1 U4974 ( .C1(n4342), .C2(n3121), .A(n4341), .B(n4340), .ZN(n4448)
         );
  AOI22_X1 U4975 ( .A1(n2160), .A2(REG2_REG_20__SCAN_IN), .B1(n4343), .B2(
        n4645), .ZN(n4346) );
  NAND2_X1 U4976 ( .A1(n4365), .A2(n4344), .ZN(n4446) );
  NAND3_X1 U4977 ( .A1(n4319), .A2(n4647), .A3(n4446), .ZN(n4345) );
  OAI211_X1 U4978 ( .C1(n4450), .C2(n4347), .A(n4346), .B(n4345), .ZN(n4348)
         );
  INV_X1 U4979 ( .A(n4348), .ZN(n4349) );
  OAI21_X1 U4980 ( .B1(n4448), .B2(n2160), .A(n4349), .ZN(U3270) );
  XNOR2_X1 U4981 ( .A(n4350), .B(n4356), .ZN(n4452) );
  INV_X1 U4982 ( .A(n4452), .ZN(n4371) );
  INV_X1 U4983 ( .A(n4351), .ZN(n4353) );
  OAI21_X1 U4984 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4355) );
  XOR2_X1 U4985 ( .A(n4356), .B(n4355), .Z(n4361) );
  OAI22_X1 U4986 ( .A1(n4441), .A2(n4458), .B1(n4459), .B2(n4460), .ZN(n4357)
         );
  AOI21_X1 U4987 ( .B1(n4358), .B2(n4463), .A(n4357), .ZN(n4359) );
  OAI21_X1 U4988 ( .B1(n4361), .B2(n4360), .A(n4359), .ZN(n4451) );
  OR2_X1 U4989 ( .A1(n4363), .A2(n4362), .ZN(n4364) );
  NAND2_X1 U4990 ( .A1(n4365), .A2(n4364), .ZN(n4521) );
  AOI22_X1 U4991 ( .A1(n2160), .A2(REG2_REG_19__SCAN_IN), .B1(n4366), .B2(
        n4645), .ZN(n4367) );
  OAI21_X1 U4992 ( .B1(n4521), .B2(n4368), .A(n4367), .ZN(n4369) );
  AOI21_X1 U4993 ( .B1(n4451), .B2(n4544), .A(n4369), .ZN(n4370) );
  OAI21_X1 U4994 ( .B1(n4371), .B2(n4391), .A(n4370), .ZN(U3271) );
  XOR2_X1 U4995 ( .A(n4384), .B(n4372), .Z(n4467) );
  INV_X1 U4996 ( .A(n4373), .ZN(n4374) );
  OAI21_X1 U4997 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n4527) );
  INV_X1 U4998 ( .A(n4527), .ZN(n4389) );
  AOI22_X1 U4999 ( .A1(n4379), .A2(n4464), .B1(n4378), .B2(n4377), .ZN(n4382)
         );
  AOI22_X1 U5000 ( .A1(n2160), .A2(REG2_REG_17__SCAN_IN), .B1(n4380), .B2(
        n4645), .ZN(n4381) );
  OAI211_X1 U5001 ( .C1(n4461), .C2(n4383), .A(n4382), .B(n4381), .ZN(n4388)
         );
  INV_X1 U5002 ( .A(n4384), .ZN(n4385) );
  XNOR2_X1 U5003 ( .A(n3857), .B(n4385), .ZN(n4386) );
  NAND2_X1 U5004 ( .A1(n4386), .A2(n3121), .ZN(n4465) );
  NOR2_X1 U5005 ( .A1(n4465), .A2(n2160), .ZN(n4387) );
  AOI211_X1 U5006 ( .C1(n4389), .C2(n4647), .A(n4388), .B(n4387), .ZN(n4390)
         );
  OAI21_X1 U5007 ( .B1(n4467), .B2(n4391), .A(n4390), .ZN(U3273) );
  INV_X1 U5008 ( .A(n4542), .ZN(n4488) );
  NAND2_X1 U5009 ( .A1(n4393), .A2(n4392), .ZN(n4401) );
  OAI21_X1 U5010 ( .B1(n4394), .B2(n4476), .A(n4401), .ZN(n4541) );
  NAND2_X1 U5011 ( .A1(n4688), .A2(n4541), .ZN(n4396) );
  NAND2_X1 U5012 ( .A1(n4686), .A2(REG1_REG_31__SCAN_IN), .ZN(n4395) );
  OAI211_X1 U5013 ( .C1(n4488), .C2(n4470), .A(n4396), .B(n4395), .ZN(U3549)
         );
  AOI21_X1 U5014 ( .B1(n4399), .B2(n4398), .A(n4397), .ZN(n4545) );
  INV_X1 U5015 ( .A(n4545), .ZN(n4490) );
  NAND2_X1 U5016 ( .A1(n4399), .A2(n4463), .ZN(n4400) );
  AND2_X1 U5017 ( .A1(n4401), .A2(n4400), .ZN(n4547) );
  INV_X1 U5018 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4402) );
  MUX2_X1 U5019 ( .A(n4547), .B(n4402), .S(n4686), .Z(n4403) );
  OAI21_X1 U5020 ( .B1(n4490), .B2(n4470), .A(n4403), .ZN(U3548) );
  INV_X1 U5021 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5022 ( .A1(n4405), .A2(n4471), .B1(n4404), .B2(n4463), .ZN(n4406)
         );
  OAI211_X1 U5023 ( .C1(n4408), .C2(n4458), .A(n4407), .B(n4406), .ZN(n4409)
         );
  AOI21_X1 U5024 ( .B1(n4410), .B2(n4676), .A(n4409), .ZN(n4491) );
  MUX2_X1 U5025 ( .A(n4411), .B(n4491), .S(n4688), .Z(n4412) );
  OAI21_X1 U5026 ( .B1(n4470), .B2(n4494), .A(n4412), .ZN(U3545) );
  INV_X1 U5027 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4415) );
  AOI21_X1 U5028 ( .B1(n4414), .B2(n4676), .A(n4413), .ZN(n4495) );
  MUX2_X1 U5029 ( .A(n4415), .B(n4495), .S(n4688), .Z(n4416) );
  OAI21_X1 U5030 ( .B1(n4470), .B2(n4497), .A(n4416), .ZN(U3544) );
  INV_X1 U5031 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U5032 ( .A1(n4418), .A2(n4471), .B1(n4417), .B2(n4463), .ZN(n4419)
         );
  OAI211_X1 U5033 ( .C1(n4421), .C2(n4458), .A(n4420), .B(n4419), .ZN(n4422)
         );
  AOI21_X1 U5034 ( .B1(n4423), .B2(n4676), .A(n4422), .ZN(n4498) );
  MUX2_X1 U5035 ( .A(n4424), .B(n4498), .S(n4688), .Z(n4425) );
  OAI21_X1 U5036 ( .B1(n4470), .B2(n4501), .A(n4425), .ZN(U3543) );
  INV_X1 U5037 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4891) );
  AOI21_X1 U5038 ( .B1(n4427), .B2(n4676), .A(n4426), .ZN(n4502) );
  MUX2_X1 U5039 ( .A(n4891), .B(n4502), .S(n4688), .Z(n4428) );
  OAI21_X1 U5040 ( .B1(n4470), .B2(n4504), .A(n4428), .ZN(U3542) );
  INV_X1 U5041 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4431) );
  AOI21_X1 U5042 ( .B1(n4430), .B2(n4676), .A(n4429), .ZN(n4505) );
  MUX2_X1 U5043 ( .A(n4431), .B(n4505), .S(n4688), .Z(n4432) );
  OAI21_X1 U5044 ( .B1(n4470), .B2(n4508), .A(n4432), .ZN(U3541) );
  OAI21_X1 U5045 ( .B1(n4434), .B2(n4483), .A(n4433), .ZN(n4509) );
  MUX2_X1 U5046 ( .A(n4509), .B(REG1_REG_22__SCAN_IN), .S(n4686), .Z(n4435) );
  INV_X1 U5047 ( .A(n4435), .ZN(n4436) );
  OAI21_X1 U5048 ( .B1(n4470), .B2(n4512), .A(n4436), .ZN(U3540) );
  INV_X1 U5049 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U5050 ( .A1(n4438), .A2(n4474), .B1(n4463), .B2(n4437), .ZN(n4439)
         );
  OAI211_X1 U5051 ( .C1(n4441), .C2(n4460), .A(n4440), .B(n4439), .ZN(n4442)
         );
  AOI21_X1 U5052 ( .B1(n4443), .B2(n4676), .A(n4442), .ZN(n4513) );
  MUX2_X1 U5053 ( .A(n4444), .B(n4513), .S(n4688), .Z(n4445) );
  OAI21_X1 U5054 ( .B1(n4470), .B2(n4516), .A(n4445), .ZN(U3539) );
  NAND3_X1 U5055 ( .A1(n4319), .A2(n4479), .A3(n4446), .ZN(n4447) );
  OAI211_X1 U5056 ( .C1(n4450), .C2(n4449), .A(n4448), .B(n4447), .ZN(n4517)
         );
  MUX2_X1 U5057 ( .A(REG1_REG_20__SCAN_IN), .B(n4517), .S(n4688), .Z(U3538) );
  AOI21_X1 U5058 ( .B1(n4452), .B2(n4676), .A(n4451), .ZN(n4518) );
  MUX2_X1 U5059 ( .A(n4181), .B(n4518), .S(n4688), .Z(n4453) );
  OAI21_X1 U5060 ( .B1(n4470), .B2(n4521), .A(n4453), .ZN(U3537) );
  INV_X1 U5061 ( .A(n4454), .ZN(n4457) );
  OAI211_X1 U5062 ( .C1(n4457), .C2(n4483), .A(n4456), .B(n4455), .ZN(n4522)
         );
  MUX2_X1 U5063 ( .A(REG1_REG_18__SCAN_IN), .B(n4522), .S(n4688), .Z(U3536) );
  OAI22_X1 U5064 ( .A1(n4461), .A2(n4460), .B1(n4459), .B2(n4458), .ZN(n4462)
         );
  AOI21_X1 U5065 ( .B1(n4464), .B2(n4463), .A(n4462), .ZN(n4466) );
  OAI211_X1 U5066 ( .C1(n4467), .C2(n4483), .A(n4466), .B(n4465), .ZN(n4468)
         );
  INV_X1 U5067 ( .A(n4468), .ZN(n4523) );
  MUX2_X1 U5068 ( .A(n4700), .B(n4523), .S(n4688), .Z(n4469) );
  OAI21_X1 U5069 ( .B1(n4470), .B2(n4527), .A(n4469), .ZN(U3535) );
  AOI22_X1 U5070 ( .A1(n4474), .A2(n4473), .B1(n4472), .B2(n4471), .ZN(n4475)
         );
  OAI21_X1 U5071 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4478) );
  AOI21_X1 U5072 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4482) );
  OAI211_X1 U5073 ( .C1(n4484), .C2(n4483), .A(n4482), .B(n4481), .ZN(n4528)
         );
  MUX2_X1 U5074 ( .A(REG1_REG_16__SCAN_IN), .B(n4528), .S(n4688), .Z(U3534) );
  NOR2_X1 U5075 ( .A1(n4683), .A2(n4485), .ZN(n4486) );
  AOI21_X1 U5076 ( .B1(n4683), .B2(n4541), .A(n4486), .ZN(n4487) );
  OAI21_X1 U5077 ( .B1(n4488), .B2(n4526), .A(n4487), .ZN(U3517) );
  MUX2_X1 U5078 ( .A(n4547), .B(n2810), .S(n4682), .Z(n4489) );
  OAI21_X1 U5079 ( .B1(n4490), .B2(n4526), .A(n4489), .ZN(U3516) );
  MUX2_X1 U5080 ( .A(n4492), .B(n4491), .S(n4683), .Z(n4493) );
  OAI21_X1 U5081 ( .B1(n4494), .B2(n4526), .A(n4493), .ZN(U3513) );
  MUX2_X1 U5082 ( .A(n4901), .B(n4495), .S(n4683), .Z(n4496) );
  OAI21_X1 U5083 ( .B1(n4497), .B2(n4526), .A(n4496), .ZN(U3512) );
  MUX2_X1 U5084 ( .A(n4499), .B(n4498), .S(n4683), .Z(n4500) );
  OAI21_X1 U5085 ( .B1(n4501), .B2(n4526), .A(n4500), .ZN(U3511) );
  INV_X1 U5086 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4898) );
  MUX2_X1 U5087 ( .A(n4898), .B(n4502), .S(n4683), .Z(n4503) );
  OAI21_X1 U5088 ( .B1(n4504), .B2(n4526), .A(n4503), .ZN(U3510) );
  MUX2_X1 U5089 ( .A(n4506), .B(n4505), .S(n4683), .Z(n4507) );
  OAI21_X1 U5090 ( .B1(n4508), .B2(n4526), .A(n4507), .ZN(U3509) );
  MUX2_X1 U5091 ( .A(n4509), .B(REG0_REG_22__SCAN_IN), .S(n4682), .Z(n4510) );
  INV_X1 U5092 ( .A(n4510), .ZN(n4511) );
  OAI21_X1 U5093 ( .B1(n4512), .B2(n4526), .A(n4511), .ZN(U3508) );
  MUX2_X1 U5094 ( .A(n4514), .B(n4513), .S(n4683), .Z(n4515) );
  OAI21_X1 U5095 ( .B1(n4516), .B2(n4526), .A(n4515), .ZN(U3507) );
  MUX2_X1 U5096 ( .A(REG0_REG_20__SCAN_IN), .B(n4517), .S(n4683), .Z(U3506) );
  MUX2_X1 U5097 ( .A(n4519), .B(n4518), .S(n4683), .Z(n4520) );
  OAI21_X1 U5098 ( .B1(n4521), .B2(n4526), .A(n4520), .ZN(U3505) );
  MUX2_X1 U5099 ( .A(REG0_REG_18__SCAN_IN), .B(n4522), .S(n4683), .Z(U3503) );
  MUX2_X1 U5100 ( .A(n4524), .B(n4523), .S(n4683), .Z(n4525) );
  OAI21_X1 U5101 ( .B1(n4527), .B2(n4526), .A(n4525), .ZN(U3501) );
  MUX2_X1 U5102 ( .A(REG0_REG_16__SCAN_IN), .B(n4528), .S(n4683), .Z(U3499) );
  MUX2_X1 U5103 ( .A(n2522), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5104 ( .A(n4529), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5105 ( .A(n4530), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5106 ( .A(DATAI_25_), .B(n4531), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5107 ( .A(n2815), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5108 ( .A(DATAI_21_), .B(n4532), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5109 ( .A(DATAI_19_), .B(n4533), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5110 ( .A(DATAI_14_), .B(n4534), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5111 ( .A(n4535), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5112 ( .A(n4536), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5113 ( .A(n4537), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5114 ( .A(DATAI_4_), .B(n4538), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5115 ( .A(n4539), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5116 ( .A(n4540), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5117 ( .A(n2482), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5118 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5119 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5120 ( .A1(n4542), .A2(n4647), .B1(n4544), .B2(n4541), .ZN(n4543)
         );
  OAI21_X1 U5121 ( .B1(n4544), .B2(n4736), .A(n4543), .ZN(U3260) );
  AOI22_X1 U5122 ( .A1(n4545), .A2(n4647), .B1(REG2_REG_30__SCAN_IN), .B2(
        n2160), .ZN(n4546) );
  OAI21_X1 U5123 ( .B1(n2160), .B2(n4547), .A(n4546), .ZN(U3261) );
  OAI211_X1 U5124 ( .C1(n4550), .C2(n4549), .A(n4631), .B(n4548), .ZN(n4555)
         );
  OAI211_X1 U5125 ( .C1(n4553), .C2(n4552), .A(n4592), .B(n4551), .ZN(n4554)
         );
  OAI211_X1 U5126 ( .C1(n4637), .C2(n4669), .A(n4555), .B(n4554), .ZN(n4556)
         );
  AOI211_X1 U5127 ( .C1(n4630), .C2(ADDR_REG_9__SCAN_IN), .A(n4557), .B(n4556), 
        .ZN(n4558) );
  INV_X1 U5128 ( .A(n4558), .ZN(U3249) );
  OAI211_X1 U5129 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4560), .A(n4592), .B(n4559), .ZN(n4562) );
  NAND2_X1 U5130 ( .A1(n4562), .A2(n4561), .ZN(n4563) );
  AOI21_X1 U5131 ( .B1(n4630), .B2(ADDR_REG_10__SCAN_IN), .A(n4563), .ZN(n4567) );
  OAI211_X1 U5132 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4565), .A(n4631), .B(n4564), .ZN(n4566) );
  OAI211_X1 U5133 ( .C1(n4637), .C2(n4568), .A(n4567), .B(n4566), .ZN(U3250)
         );
  OAI211_X1 U5134 ( .C1(n4571), .C2(n4570), .A(n4631), .B(n4569), .ZN(n4576)
         );
  OAI211_X1 U5135 ( .C1(n4574), .C2(n4573), .A(n4592), .B(n4572), .ZN(n4575)
         );
  OAI211_X1 U5136 ( .C1(n4637), .C2(n4665), .A(n4576), .B(n4575), .ZN(n4577)
         );
  AOI211_X1 U5137 ( .C1(n4630), .C2(ADDR_REG_11__SCAN_IN), .A(n4578), .B(n4577), .ZN(n4579) );
  INV_X1 U5138 ( .A(n4579), .ZN(U3251) );
  OAI211_X1 U5139 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4581), .A(n4592), .B(n4580), .ZN(n4583) );
  NAND2_X1 U5140 ( .A1(n4583), .A2(n4582), .ZN(n4584) );
  AOI21_X1 U5141 ( .B1(n4630), .B2(ADDR_REG_12__SCAN_IN), .A(n4584), .ZN(n4588) );
  OAI211_X1 U5142 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4586), .A(n4631), .B(n4585), .ZN(n4587) );
  OAI211_X1 U5143 ( .C1(n4637), .C2(n4589), .A(n4588), .B(n4587), .ZN(U3252)
         );
  AOI21_X1 U5144 ( .B1(n4591), .B2(n4603), .A(n4590), .ZN(n4595) );
  OAI21_X1 U5145 ( .B1(n4595), .B2(n4594), .A(n4592), .ZN(n4593) );
  AOI21_X1 U5146 ( .B1(n4595), .B2(n4594), .A(n4593), .ZN(n4597) );
  AOI211_X1 U5147 ( .C1(n4630), .C2(ADDR_REG_13__SCAN_IN), .A(n4597), .B(n4596), .ZN(n4602) );
  OAI211_X1 U5148 ( .C1(n4600), .C2(n4599), .A(n4631), .B(n4598), .ZN(n4601)
         );
  OAI211_X1 U5149 ( .C1(n4637), .C2(n4603), .A(n4602), .B(n4601), .ZN(U3253)
         );
  AOI211_X1 U5150 ( .C1(n4606), .C2(n4605), .A(n4604), .B(n4624), .ZN(n4607)
         );
  AOI211_X1 U5151 ( .C1(n4630), .C2(ADDR_REG_15__SCAN_IN), .A(n4608), .B(n4607), .ZN(n4613) );
  OAI211_X1 U5152 ( .C1(n4611), .C2(n4610), .A(n4631), .B(n4609), .ZN(n4612)
         );
  OAI211_X1 U5153 ( .C1(n4637), .C2(n4614), .A(n4613), .B(n4612), .ZN(U3255)
         );
  AOI221_X1 U5154 ( .B1(n4617), .B2(n4616), .C1(n4615), .C2(n4616), .A(n4624), 
        .ZN(n4618) );
  AOI211_X1 U5155 ( .C1(n4630), .C2(ADDR_REG_16__SCAN_IN), .A(n4619), .B(n4618), .ZN(n4623) );
  OAI221_X1 U5156 ( .B1(n4621), .B2(REG1_REG_16__SCAN_IN), .C1(n4621), .C2(
        n4620), .A(n4631), .ZN(n4622) );
  OAI211_X1 U5157 ( .C1(n4637), .C2(n4660), .A(n4623), .B(n4622), .ZN(U3256)
         );
  AOI221_X1 U5158 ( .B1(n4627), .B2(n4626), .C1(n4625), .C2(n4626), .A(n4624), 
        .ZN(n4628) );
  AOI211_X1 U5159 ( .C1(n4630), .C2(ADDR_REG_17__SCAN_IN), .A(n4629), .B(n4628), .ZN(n4635) );
  OAI221_X1 U5160 ( .B1(n4633), .B2(n2173), .C1(n4633), .C2(n4632), .A(n4631), 
        .ZN(n4634) );
  OAI211_X1 U5161 ( .C1(n4637), .C2(n4636), .A(n4635), .B(n4634), .ZN(U3257)
         );
  AOI22_X1 U5162 ( .A1(n2160), .A2(REG2_REG_8__SCAN_IN), .B1(n4638), .B2(n4645), .ZN(n4643) );
  INV_X1 U5163 ( .A(n4639), .ZN(n4640) );
  AOI22_X1 U5164 ( .A1(n4641), .A2(n4648), .B1(n4647), .B2(n4640), .ZN(n4642)
         );
  OAI211_X1 U5165 ( .C1(n2160), .C2(n4644), .A(n4643), .B(n4642), .ZN(U3282)
         );
  AOI22_X1 U5166 ( .A1(n2160), .A2(REG2_REG_3__SCAN_IN), .B1(n4645), .B2(n2523), .ZN(n4651) );
  AOI22_X1 U5167 ( .A1(n4649), .A2(n4648), .B1(n4647), .B2(n4646), .ZN(n4650)
         );
  OAI211_X1 U5168 ( .C1(n2160), .C2(n4652), .A(n4651), .B(n4650), .ZN(U3287)
         );
  AND2_X1 U5169 ( .A1(D_REG_31__SCAN_IN), .A2(n4654), .ZN(U3291) );
  INV_X1 U5170 ( .A(D_REG_30__SCAN_IN), .ZN(n4879) );
  NOR2_X1 U5171 ( .A1(n4653), .A2(n4879), .ZN(U3292) );
  INV_X1 U5172 ( .A(D_REG_29__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5173 ( .A1(n4653), .A2(n4776), .ZN(U3293) );
  INV_X1 U5174 ( .A(D_REG_28__SCAN_IN), .ZN(n4871) );
  NOR2_X1 U5175 ( .A1(n4653), .A2(n4871), .ZN(U3294) );
  INV_X1 U5176 ( .A(D_REG_27__SCAN_IN), .ZN(n4770) );
  NOR2_X1 U5177 ( .A1(n4653), .A2(n4770), .ZN(U3295) );
  INV_X1 U5178 ( .A(D_REG_26__SCAN_IN), .ZN(n4880) );
  NOR2_X1 U5179 ( .A1(n4653), .A2(n4880), .ZN(U3296) );
  AND2_X1 U5180 ( .A1(D_REG_25__SCAN_IN), .A2(n4654), .ZN(U3297) );
  INV_X1 U5181 ( .A(D_REG_24__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U5182 ( .A1(n4653), .A2(n4877), .ZN(U3298) );
  INV_X1 U5183 ( .A(D_REG_23__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U5184 ( .A1(n4653), .A2(n4771), .ZN(U3299) );
  AND2_X1 U5185 ( .A1(D_REG_22__SCAN_IN), .A2(n4654), .ZN(U3300) );
  AND2_X1 U5186 ( .A1(D_REG_21__SCAN_IN), .A2(n4654), .ZN(U3301) );
  INV_X1 U5187 ( .A(D_REG_20__SCAN_IN), .ZN(n4873) );
  NOR2_X1 U5188 ( .A1(n4653), .A2(n4873), .ZN(U3302) );
  INV_X1 U5189 ( .A(D_REG_19__SCAN_IN), .ZN(n4773) );
  NOR2_X1 U5190 ( .A1(n4653), .A2(n4773), .ZN(U3303) );
  AND2_X1 U5191 ( .A1(D_REG_18__SCAN_IN), .A2(n4654), .ZN(U3304) );
  AND2_X1 U5192 ( .A1(D_REG_17__SCAN_IN), .A2(n4654), .ZN(U3305) );
  INV_X1 U5193 ( .A(D_REG_16__SCAN_IN), .ZN(n4774) );
  NOR2_X1 U5194 ( .A1(n4653), .A2(n4774), .ZN(U3306) );
  AND2_X1 U5195 ( .A1(D_REG_15__SCAN_IN), .A2(n4654), .ZN(U3307) );
  INV_X1 U5196 ( .A(D_REG_14__SCAN_IN), .ZN(n4874) );
  NOR2_X1 U5197 ( .A1(n4653), .A2(n4874), .ZN(U3308) );
  AND2_X1 U5198 ( .A1(D_REG_13__SCAN_IN), .A2(n4654), .ZN(U3309) );
  AND2_X1 U5199 ( .A1(D_REG_12__SCAN_IN), .A2(n4654), .ZN(U3310) );
  AND2_X1 U5200 ( .A1(D_REG_11__SCAN_IN), .A2(n4654), .ZN(U3311) );
  INV_X1 U5201 ( .A(D_REG_10__SCAN_IN), .ZN(n4876) );
  NOR2_X1 U5202 ( .A1(n4653), .A2(n4876), .ZN(U3312) );
  AND2_X1 U5203 ( .A1(D_REG_9__SCAN_IN), .A2(n4654), .ZN(U3313) );
  AND2_X1 U5204 ( .A1(D_REG_8__SCAN_IN), .A2(n4654), .ZN(U3314) );
  AND2_X1 U5205 ( .A1(D_REG_7__SCAN_IN), .A2(n4654), .ZN(U3315) );
  INV_X1 U5206 ( .A(D_REG_6__SCAN_IN), .ZN(n4870) );
  NOR2_X1 U5207 ( .A1(n4653), .A2(n4870), .ZN(U3316) );
  AND2_X1 U5208 ( .A1(D_REG_5__SCAN_IN), .A2(n4654), .ZN(U3317) );
  AND2_X1 U5209 ( .A1(D_REG_4__SCAN_IN), .A2(n4654), .ZN(U3318) );
  AND2_X1 U5210 ( .A1(D_REG_3__SCAN_IN), .A2(n4654), .ZN(U3319) );
  AND2_X1 U5211 ( .A1(D_REG_2__SCAN_IN), .A2(n4654), .ZN(U3320) );
  OAI21_X1 U5212 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4655), .ZN(
        n4656) );
  INV_X1 U5213 ( .A(n4656), .ZN(U3329) );
  OAI22_X1 U5214 ( .A1(U3149), .A2(n4657), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4658) );
  INV_X1 U5215 ( .A(n4658), .ZN(U3335) );
  INV_X1 U5216 ( .A(DATAI_16_), .ZN(n4659) );
  AOI22_X1 U5217 ( .A1(STATE_REG_SCAN_IN), .A2(n4660), .B1(n4659), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5218 ( .A1(U3149), .A2(n4661), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4662) );
  INV_X1 U5219 ( .A(n4662), .ZN(U3337) );
  OAI22_X1 U5220 ( .A1(U3149), .A2(n4663), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4664) );
  INV_X1 U5221 ( .A(n4664), .ZN(U3340) );
  INV_X1 U5222 ( .A(DATAI_11_), .ZN(n4934) );
  AOI22_X1 U5223 ( .A1(STATE_REG_SCAN_IN), .A2(n4665), .B1(n4934), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5224 ( .A1(U3149), .A2(n4666), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4667) );
  INV_X1 U5225 ( .A(n4667), .ZN(U3342) );
  INV_X1 U5226 ( .A(DATAI_9_), .ZN(n4668) );
  AOI22_X1 U5227 ( .A1(STATE_REG_SCAN_IN), .A2(n4669), .B1(n4668), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5228 ( .A1(n4683), .A2(n4670), .B1(n2548), .B2(n4682), .ZN(U3467)
         );
  INV_X1 U5229 ( .A(n4671), .ZN(n4672) );
  AOI211_X1 U5230 ( .C1(n4675), .C2(n4674), .A(n4673), .B(n4672), .ZN(n4685)
         );
  AOI22_X1 U5231 ( .A1(n4683), .A2(n4685), .B1(n2537), .B2(n4682), .ZN(U3475)
         );
  NAND3_X1 U5232 ( .A1(n4678), .A2(n4677), .A3(n4676), .ZN(n4679) );
  AND3_X1 U5233 ( .A1(n4681), .A2(n4680), .A3(n4679), .ZN(n4687) );
  AOI22_X1 U5234 ( .A1(n4683), .A2(n4687), .B1(n2577), .B2(n4682), .ZN(U3481)
         );
  INV_X1 U5235 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5236 ( .A1(n4688), .A2(n4685), .B1(n4684), .B2(n4686), .ZN(U3522)
         );
  INV_X1 U5237 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5238 ( .A1(n4688), .A2(n4687), .B1(n4696), .B2(n4686), .ZN(U3525)
         );
  AOI22_X1 U5239 ( .A1(STATE_REG_SCAN_IN), .A2(n4689), .B1(DATAI_13_), .B2(
        U3149), .ZN(n5005) );
  INV_X1 U5240 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4692) );
  INV_X1 U5241 ( .A(keyinput60), .ZN(n4691) );
  AOI22_X1 U5242 ( .A1(n4692), .A2(keyinput81), .B1(ADDR_REG_15__SCAN_IN), 
        .B2(n4691), .ZN(n4690) );
  OAI221_X1 U5243 ( .B1(n4692), .B2(keyinput81), .C1(n4691), .C2(
        ADDR_REG_15__SCAN_IN), .A(n4690), .ZN(n4704) );
  AOI22_X1 U5244 ( .A1(n3710), .A2(keyinput111), .B1(n4694), .B2(keyinput108), 
        .ZN(n4693) );
  OAI221_X1 U5245 ( .B1(n3710), .B2(keyinput111), .C1(n4694), .C2(keyinput108), 
        .A(n4693), .ZN(n4703) );
  AOI22_X1 U5246 ( .A1(n4697), .A2(keyinput79), .B1(keyinput50), .B2(n4696), 
        .ZN(n4695) );
  OAI221_X1 U5247 ( .B1(n4697), .B2(keyinput79), .C1(n4696), .C2(keyinput50), 
        .A(n4695), .ZN(n4702) );
  AOI22_X1 U5248 ( .A1(n4700), .A2(keyinput37), .B1(keyinput64), .B2(n4699), 
        .ZN(n4698) );
  OAI221_X1 U5249 ( .B1(n4700), .B2(keyinput37), .C1(n4699), .C2(keyinput64), 
        .A(n4698), .ZN(n4701) );
  NOR4_X1 U5250 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n5003)
         );
  AOI22_X1 U5251 ( .A1(n2523), .A2(keyinput84), .B1(keyinput97), .B2(n3437), 
        .ZN(n4705) );
  OAI221_X1 U5252 ( .B1(n2523), .B2(keyinput84), .C1(n3437), .C2(keyinput97), 
        .A(n4705), .ZN(n4714) );
  INV_X1 U5253 ( .A(keyinput36), .ZN(n4707) );
  AOI22_X1 U5254 ( .A1(n2417), .A2(keyinput70), .B1(ADDR_REG_7__SCAN_IN), .B2(
        n4707), .ZN(n4706) );
  OAI221_X1 U5255 ( .B1(n2417), .B2(keyinput70), .C1(n4707), .C2(
        ADDR_REG_7__SCAN_IN), .A(n4706), .ZN(n4713) );
  XOR2_X1 U5256 ( .A(n3188), .B(keyinput94), .Z(n4711) );
  XNOR2_X1 U5257 ( .A(keyinput19), .B(REG2_REG_0__SCAN_IN), .ZN(n4710) );
  XNOR2_X1 U5258 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput62), .ZN(n4709) );
  XNOR2_X1 U5259 ( .A(IR_REG_0__SCAN_IN), .B(keyinput14), .ZN(n4708) );
  NAND4_X1 U5260 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4712)
         );
  NOR3_X1 U5261 ( .A1(n4714), .A2(n4713), .A3(n4712), .ZN(n5002) );
  INV_X1 U5262 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5263 ( .A1(n4717), .A2(keyinput34), .B1(n4716), .B2(keyinput110), 
        .ZN(n4715) );
  OAI221_X1 U5264 ( .B1(n4717), .B2(keyinput34), .C1(n4716), .C2(keyinput110), 
        .A(n4715), .ZN(n4801) );
  INV_X1 U5265 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5266 ( .A1(n4720), .A2(keyinput24), .B1(keyinput74), .B2(n4719), 
        .ZN(n4718) );
  OAI221_X1 U5267 ( .B1(n4720), .B2(keyinput24), .C1(n4719), .C2(keyinput74), 
        .A(n4718), .ZN(n4800) );
  INV_X1 U5268 ( .A(keyinput127), .ZN(n4743) );
  INV_X1 U5269 ( .A(keyinput107), .ZN(n4725) );
  INV_X1 U5270 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4724) );
  INV_X1 U5271 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5272 ( .A1(n4722), .A2(keyinput71), .B1(n4210), .B2(keyinput23), 
        .ZN(n4721) );
  OAI221_X1 U5273 ( .B1(n4722), .B2(keyinput71), .C1(n4210), .C2(keyinput23), 
        .A(n4721), .ZN(n4723) );
  AOI221_X1 U5274 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4725), .C1(n4724), .C2(
        keyinput107), .A(n4723), .ZN(n4742) );
  AOI22_X1 U5275 ( .A1(n4728), .A2(keyinput13), .B1(n4727), .B2(keyinput10), 
        .ZN(n4726) );
  OAI221_X1 U5276 ( .B1(n4728), .B2(keyinput13), .C1(n4727), .C2(keyinput10), 
        .A(n4726), .ZN(n4740) );
  INV_X1 U5277 ( .A(keyinput80), .ZN(n4730) );
  AOI22_X1 U5278 ( .A1(n3352), .A2(keyinput66), .B1(ADDR_REG_3__SCAN_IN), .B2(
        n4730), .ZN(n4729) );
  OAI221_X1 U5279 ( .B1(n3352), .B2(keyinput66), .C1(n4730), .C2(
        ADDR_REG_3__SCAN_IN), .A(n4729), .ZN(n4739) );
  AOI22_X1 U5280 ( .A1(n4733), .A2(keyinput96), .B1(keyinput105), .B2(n4732), 
        .ZN(n4731) );
  OAI221_X1 U5281 ( .B1(n4733), .B2(keyinput96), .C1(n4732), .C2(keyinput105), 
        .A(n4731), .ZN(n4738) );
  INV_X1 U5282 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5283 ( .A1(n4736), .A2(keyinput17), .B1(n4735), .B2(keyinput40), 
        .ZN(n4734) );
  OAI221_X1 U5284 ( .B1(n4736), .B2(keyinput17), .C1(n4735), .C2(keyinput40), 
        .A(n4734), .ZN(n4737) );
  NOR4_X1 U5285 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4741)
         );
  OAI211_X1 U5286 ( .C1(IR_REG_19__SCAN_IN), .C2(n4743), .A(n4742), .B(n4741), 
        .ZN(n4799) );
  AOI22_X1 U5287 ( .A1(n4746), .A2(keyinput48), .B1(n4745), .B2(keyinput58), 
        .ZN(n4744) );
  OAI221_X1 U5288 ( .B1(n4746), .B2(keyinput48), .C1(n4745), .C2(keyinput58), 
        .A(n4744), .ZN(n4756) );
  AOI22_X1 U5289 ( .A1(n4748), .A2(keyinput33), .B1(keyinput52), .B2(n3787), 
        .ZN(n4747) );
  OAI221_X1 U5290 ( .B1(n4748), .B2(keyinput33), .C1(n3787), .C2(keyinput52), 
        .A(n4747), .ZN(n4755) );
  AOI22_X1 U5291 ( .A1(n2614), .A2(keyinput45), .B1(n4750), .B2(keyinput69), 
        .ZN(n4749) );
  OAI221_X1 U5292 ( .B1(n2614), .B2(keyinput45), .C1(n4750), .C2(keyinput69), 
        .A(n4749), .ZN(n4754) );
  INV_X1 U5293 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4752) );
  AOI22_X1 U5294 ( .A1(n4752), .A2(keyinput116), .B1(n2643), .B2(keyinput100), 
        .ZN(n4751) );
  OAI221_X1 U5295 ( .B1(n4752), .B2(keyinput116), .C1(n2643), .C2(keyinput100), 
        .A(n4751), .ZN(n4753) );
  NOR4_X1 U5296 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4797)
         );
  AOI22_X1 U5297 ( .A1(n2204), .A2(keyinput88), .B1(keyinput53), .B2(n2510), 
        .ZN(n4757) );
  OAI221_X1 U5298 ( .B1(n2204), .B2(keyinput88), .C1(n2510), .C2(keyinput53), 
        .A(n4757), .ZN(n4768) );
  INV_X1 U5299 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4758) );
  XNOR2_X1 U5300 ( .A(keyinput31), .B(n4758), .ZN(n4767) );
  XOR2_X1 U5301 ( .A(n4759), .B(keyinput113), .Z(n4763) );
  XNOR2_X1 U5302 ( .A(IR_REG_31__SCAN_IN), .B(keyinput43), .ZN(n4762) );
  XNOR2_X1 U5303 ( .A(IR_REG_27__SCAN_IN), .B(keyinput30), .ZN(n4761) );
  XNOR2_X1 U5304 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput75), .ZN(n4760) );
  NAND4_X1 U5305 ( .A1(n4763), .A2(n4762), .A3(n4761), .A4(n4760), .ZN(n4766)
         );
  XNOR2_X1 U5306 ( .A(keyinput59), .B(n4764), .ZN(n4765) );
  NOR4_X1 U5307 ( .A1(n4768), .A2(n4767), .A3(n4766), .A4(n4765), .ZN(n4796)
         );
  AOI22_X1 U5308 ( .A1(n4771), .A2(keyinput101), .B1(keyinput42), .B2(n4770), 
        .ZN(n4769) );
  OAI221_X1 U5309 ( .B1(n4771), .B2(keyinput101), .C1(n4770), .C2(keyinput42), 
        .A(n4769), .ZN(n4782) );
  AOI22_X1 U5310 ( .A1(n4774), .A2(keyinput87), .B1(keyinput98), .B2(n4773), 
        .ZN(n4772) );
  OAI221_X1 U5311 ( .B1(n4774), .B2(keyinput87), .C1(n4773), .C2(keyinput98), 
        .A(n4772), .ZN(n4781) );
  AOI22_X1 U5312 ( .A1(n3695), .A2(keyinput77), .B1(n4776), .B2(keyinput117), 
        .ZN(n4775) );
  OAI221_X1 U5313 ( .B1(n3695), .B2(keyinput77), .C1(n4776), .C2(keyinput117), 
        .A(n4775), .ZN(n4780) );
  XOR2_X1 U5314 ( .A(n2603), .B(keyinput57), .Z(n4778) );
  XNOR2_X1 U5315 ( .A(IR_REG_7__SCAN_IN), .B(keyinput51), .ZN(n4777) );
  NAND2_X1 U5316 ( .A1(n4778), .A2(n4777), .ZN(n4779) );
  NOR4_X1 U5317 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), .ZN(n4795)
         );
  INV_X1 U5318 ( .A(DATAI_4_), .ZN(n4784) );
  AOI22_X1 U5319 ( .A1(n4784), .A2(keyinput72), .B1(keyinput102), .B2(n2537), 
        .ZN(n4783) );
  OAI221_X1 U5320 ( .B1(n4784), .B2(keyinput72), .C1(n2537), .C2(keyinput102), 
        .A(n4783), .ZN(n4793) );
  AOI22_X1 U5321 ( .A1(n4786), .A2(keyinput22), .B1(keyinput114), .B2(n2201), 
        .ZN(n4785) );
  OAI221_X1 U5322 ( .B1(n4786), .B2(keyinput22), .C1(n2201), .C2(keyinput114), 
        .A(n4785), .ZN(n4792) );
  AOI22_X1 U5323 ( .A1(n2577), .A2(keyinput46), .B1(n2574), .B2(keyinput120), 
        .ZN(n4787) );
  OAI221_X1 U5324 ( .B1(n2577), .B2(keyinput46), .C1(n2574), .C2(keyinput120), 
        .A(n4787), .ZN(n4791) );
  XOR2_X1 U5325 ( .A(n2521), .B(keyinput21), .Z(n4789) );
  XNOR2_X1 U5326 ( .A(IR_REG_1__SCAN_IN), .B(keyinput55), .ZN(n4788) );
  NAND2_X1 U5327 ( .A1(n4789), .A2(n4788), .ZN(n4790) );
  NOR4_X1 U5328 ( .A1(n4793), .A2(n4792), .A3(n4791), .A4(n4790), .ZN(n4794)
         );
  NAND4_X1 U5329 ( .A1(n4797), .A2(n4796), .A3(n4795), .A4(n4794), .ZN(n4798)
         );
  NOR4_X1 U5330 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n5001)
         );
  NAND2_X1 U5331 ( .A1(keyinput59), .A2(keyinput31), .ZN(n4802) );
  NOR3_X1 U5332 ( .A1(keyinput113), .A2(keyinput75), .A3(n4802), .ZN(n4834) );
  INV_X1 U5333 ( .A(keyinput50), .ZN(n4803) );
  NOR4_X1 U5334 ( .A1(keyinput53), .A2(keyinput88), .A3(keyinput30), .A4(n4803), .ZN(n4833) );
  NAND2_X1 U5335 ( .A1(keyinput102), .A2(keyinput72), .ZN(n4804) );
  NOR3_X1 U5336 ( .A1(keyinput21), .A2(keyinput22), .A3(n4804), .ZN(n4805) );
  NAND3_X1 U5337 ( .A1(keyinput69), .A2(keyinput46), .A3(n4805), .ZN(n4814) );
  NAND2_X1 U5338 ( .A1(keyinput100), .A2(keyinput58), .ZN(n4806) );
  NOR3_X1 U5339 ( .A1(keyinput116), .A2(keyinput45), .A3(n4806), .ZN(n4812) );
  NAND2_X1 U5340 ( .A1(keyinput48), .A2(keyinput43), .ZN(n4807) );
  NOR3_X1 U5341 ( .A1(keyinput52), .A2(keyinput33), .A3(n4807), .ZN(n4811) );
  INV_X1 U5342 ( .A(keyinput87), .ZN(n4808) );
  NOR4_X1 U5343 ( .A1(keyinput117), .A2(keyinput101), .A3(keyinput42), .A4(
        n4808), .ZN(n4810) );
  NOR4_X1 U5344 ( .A1(keyinput114), .A2(keyinput51), .A3(keyinput57), .A4(
        keyinput77), .ZN(n4809) );
  NAND4_X1 U5345 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(n4813)
         );
  NOR4_X1 U5346 ( .A1(keyinput120), .A2(keyinput55), .A3(n4814), .A4(n4813), 
        .ZN(n4832) );
  INV_X1 U5347 ( .A(keyinput92), .ZN(n4815) );
  NAND4_X1 U5348 ( .A1(keyinput49), .A2(keyinput1), .A3(keyinput41), .A4(n4815), .ZN(n4816) );
  NOR3_X1 U5349 ( .A1(keyinput104), .A2(keyinput28), .A3(n4816), .ZN(n4817) );
  NAND3_X1 U5350 ( .A1(keyinput29), .A2(keyinput5), .A3(n4817), .ZN(n4830) );
  NOR2_X1 U5351 ( .A1(keyinput8), .A2(keyinput26), .ZN(n4818) );
  NAND3_X1 U5352 ( .A1(keyinput56), .A2(keyinput18), .A3(n4818), .ZN(n4829) );
  NAND4_X1 U5353 ( .A1(keyinput16), .A2(keyinput12), .A3(keyinput32), .A4(
        keyinput68), .ZN(n4828) );
  INV_X1 U5354 ( .A(keyinput82), .ZN(n4819) );
  NOR4_X1 U5355 ( .A1(keyinput54), .A2(keyinput63), .A3(keyinput78), .A4(n4819), .ZN(n4826) );
  NAND2_X1 U5356 ( .A1(keyinput47), .A2(keyinput35), .ZN(n4820) );
  NOR3_X1 U5357 ( .A1(keyinput39), .A2(keyinput38), .A3(n4820), .ZN(n4825) );
  NAND2_X1 U5358 ( .A1(keyinput122), .A2(keyinput106), .ZN(n4821) );
  NOR3_X1 U5359 ( .A1(keyinput99), .A2(keyinput118), .A3(n4821), .ZN(n4824) );
  INV_X1 U5360 ( .A(keyinput83), .ZN(n4822) );
  NOR4_X1 U5361 ( .A1(keyinput90), .A2(keyinput86), .A3(keyinput95), .A4(n4822), .ZN(n4823) );
  NAND4_X1 U5362 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4827)
         );
  NOR4_X1 U5363 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4827), .ZN(n4831)
         );
  NAND4_X1 U5364 ( .A1(n4834), .A2(n4833), .A3(n4832), .A4(n4831), .ZN(n4868)
         );
  NOR2_X1 U5365 ( .A1(keyinput19), .A2(keyinput14), .ZN(n4835) );
  NAND3_X1 U5366 ( .A1(keyinput94), .A2(keyinput36), .A3(n4835), .ZN(n4842) );
  INV_X1 U5367 ( .A(keyinput97), .ZN(n4836) );
  NAND4_X1 U5368 ( .A1(keyinput84), .A2(keyinput105), .A3(keyinput62), .A4(
        n4836), .ZN(n4841) );
  NOR2_X1 U5369 ( .A1(keyinput64), .A2(keyinput37), .ZN(n4837) );
  NAND3_X1 U5370 ( .A1(keyinput81), .A2(keyinput79), .A3(n4837), .ZN(n4840) );
  NOR2_X1 U5371 ( .A1(keyinput70), .A2(keyinput108), .ZN(n4838) );
  NAND3_X1 U5372 ( .A1(keyinput111), .A2(keyinput60), .A3(n4838), .ZN(n4839)
         );
  NOR4_X1 U5373 ( .A1(n4842), .A2(n4841), .A3(n4840), .A4(n4839), .ZN(n4866)
         );
  NOR4_X1 U5374 ( .A1(keyinput107), .A2(keyinput71), .A3(keyinput23), .A4(
        keyinput24), .ZN(n4844) );
  INV_X1 U5375 ( .A(keyinput74), .ZN(n4843) );
  NAND4_X1 U5376 ( .A1(keyinput126), .A2(keyinput34), .A3(n4844), .A4(n4843), 
        .ZN(n4848) );
  NAND2_X1 U5377 ( .A1(keyinput40), .A2(keyinput13), .ZN(n4845) );
  NOR3_X1 U5378 ( .A1(keyinput66), .A2(keyinput96), .A3(n4845), .ZN(n4846) );
  NAND3_X1 U5379 ( .A1(keyinput110), .A2(keyinput80), .A3(n4846), .ZN(n4847)
         );
  NOR4_X1 U5380 ( .A1(keyinput17), .A2(keyinput10), .A3(n4848), .A4(n4847), 
        .ZN(n4865) );
  INV_X1 U5381 ( .A(keyinput7), .ZN(n4849) );
  NAND4_X1 U5382 ( .A1(keyinput119), .A2(keyinput27), .A3(keyinput11), .A4(
        n4849), .ZN(n4855) );
  OR4_X1 U5383 ( .A1(keyinput44), .A2(keyinput112), .A3(keyinput67), .A4(
        keyinput76), .ZN(n4854) );
  INV_X1 U5384 ( .A(keyinput25), .ZN(n4850) );
  NAND4_X1 U5385 ( .A1(keyinput125), .A2(keyinput73), .A3(keyinput109), .A4(
        n4850), .ZN(n4853) );
  NOR2_X1 U5386 ( .A1(keyinput91), .A2(keyinput89), .ZN(n4851) );
  NAND3_X1 U5387 ( .A1(keyinput85), .A2(keyinput65), .A3(n4851), .ZN(n4852) );
  NOR4_X1 U5388 ( .A1(n4855), .A2(n4854), .A3(n4853), .A4(n4852), .ZN(n4864)
         );
  INV_X1 U5389 ( .A(keyinput3), .ZN(n4856) );
  NAND4_X1 U5390 ( .A1(keyinput0), .A2(keyinput123), .A3(keyinput2), .A4(n4856), .ZN(n4862) );
  OR4_X1 U5391 ( .A1(keyinput98), .A2(keyinput103), .A3(keyinput124), .A4(
        keyinput61), .ZN(n4861) );
  INV_X1 U5392 ( .A(keyinput15), .ZN(n4857) );
  NAND4_X1 U5393 ( .A1(keyinput93), .A2(keyinput4), .A3(keyinput9), .A4(n4857), 
        .ZN(n4860) );
  NOR2_X1 U5394 ( .A1(keyinput6), .A2(keyinput115), .ZN(n4858) );
  NAND3_X1 U5395 ( .A1(keyinput121), .A2(keyinput20), .A3(n4858), .ZN(n4859)
         );
  NOR4_X1 U5396 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4863)
         );
  NAND4_X1 U5397 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4867)
         );
  OAI21_X1 U5398 ( .B1(n4868), .B2(n4867), .A(keyinput127), .ZN(n4999) );
  AOI22_X1 U5399 ( .A1(n4871), .A2(keyinput103), .B1(keyinput123), .B2(n4870), 
        .ZN(n4869) );
  OAI221_X1 U5400 ( .B1(n4871), .B2(keyinput103), .C1(n4870), .C2(keyinput123), 
        .A(n4869), .ZN(n4884) );
  AOI22_X1 U5401 ( .A1(n4874), .A2(keyinput0), .B1(keyinput124), .B2(n4873), 
        .ZN(n4872) );
  OAI221_X1 U5402 ( .B1(n4874), .B2(keyinput0), .C1(n4873), .C2(keyinput124), 
        .A(n4872), .ZN(n4883) );
  AOI22_X1 U5403 ( .A1(n4877), .A2(keyinput61), .B1(keyinput3), .B2(n4876), 
        .ZN(n4875) );
  OAI221_X1 U5404 ( .B1(n4877), .B2(keyinput61), .C1(n4876), .C2(keyinput3), 
        .A(n4875), .ZN(n4882) );
  AOI22_X1 U5405 ( .A1(n4880), .A2(keyinput2), .B1(keyinput6), .B2(n4879), 
        .ZN(n4878) );
  OAI221_X1 U5406 ( .B1(n4880), .B2(keyinput2), .C1(n4879), .C2(keyinput6), 
        .A(n4878), .ZN(n4881) );
  NOR4_X1 U5407 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .ZN(n4931)
         );
  AOI22_X1 U5408 ( .A1(n2675), .A2(keyinput121), .B1(keyinput115), .B2(n4886), 
        .ZN(n4885) );
  OAI221_X1 U5409 ( .B1(n2675), .B2(keyinput121), .C1(n4886), .C2(keyinput115), 
        .A(n4885), .ZN(n4895) );
  AOI22_X1 U5410 ( .A1(n4514), .A2(keyinput20), .B1(n4444), .B2(keyinput93), 
        .ZN(n4887) );
  OAI221_X1 U5411 ( .B1(n4514), .B2(keyinput20), .C1(n4444), .C2(keyinput93), 
        .A(n4887), .ZN(n4894) );
  INV_X1 U5412 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U5413 ( .A1(n3938), .A2(keyinput15), .B1(keyinput4), .B2(n4889), 
        .ZN(n4888) );
  OAI221_X1 U5414 ( .B1(n3938), .B2(keyinput15), .C1(n4889), .C2(keyinput4), 
        .A(n4888), .ZN(n4893) );
  AOI22_X1 U5415 ( .A1(n4506), .A2(keyinput9), .B1(keyinput44), .B2(n4891), 
        .ZN(n4890) );
  OAI221_X1 U5416 ( .B1(n4506), .B2(keyinput9), .C1(n4891), .C2(keyinput44), 
        .A(n4890), .ZN(n4892) );
  NOR4_X1 U5417 ( .A1(n4895), .A2(n4894), .A3(n4893), .A4(n4892), .ZN(n4930)
         );
  AOI22_X1 U5418 ( .A1(n2836), .A2(keyinput76), .B1(keyinput7), .B2(n2810), 
        .ZN(n4896) );
  OAI221_X1 U5419 ( .B1(n2836), .B2(keyinput76), .C1(n2810), .C2(keyinput7), 
        .A(n4896), .ZN(n4908) );
  AOI22_X1 U5420 ( .A1(n4898), .A2(keyinput112), .B1(n4424), .B2(keyinput27), 
        .ZN(n4897) );
  OAI221_X1 U5421 ( .B1(n4898), .B2(keyinput112), .C1(n4424), .C2(keyinput27), 
        .A(n4897), .ZN(n4907) );
  AOI22_X1 U5422 ( .A1(n4901), .A2(keyinput119), .B1(n4900), .B2(keyinput67), 
        .ZN(n4899) );
  OAI221_X1 U5423 ( .B1(n4901), .B2(keyinput119), .C1(n4900), .C2(keyinput67), 
        .A(n4899), .ZN(n4906) );
  INV_X1 U5424 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4902) );
  XOR2_X1 U5425 ( .A(n4902), .B(keyinput11), .Z(n4904) );
  XNOR2_X1 U5426 ( .A(IR_REG_28__SCAN_IN), .B(keyinput91), .ZN(n4903) );
  NAND2_X1 U5427 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  NOR4_X1 U5428 ( .A1(n4908), .A2(n4907), .A3(n4906), .A4(n4905), .ZN(n4929)
         );
  INV_X1 U5429 ( .A(DATAI_7_), .ZN(n4911) );
  INV_X1 U5430 ( .A(DATAI_2_), .ZN(n4910) );
  AOI22_X1 U5431 ( .A1(n4911), .A2(keyinput125), .B1(keyinput109), .B2(n4910), 
        .ZN(n4909) );
  OAI221_X1 U5432 ( .B1(n4911), .B2(keyinput125), .C1(n4910), .C2(keyinput109), 
        .A(n4909), .ZN(n4912) );
  INV_X1 U5433 ( .A(n4912), .ZN(n4927) );
  AOI22_X1 U5434 ( .A1(n4915), .A2(keyinput25), .B1(n4914), .B2(keyinput29), 
        .ZN(n4913) );
  OAI221_X1 U5435 ( .B1(n4915), .B2(keyinput25), .C1(n4914), .C2(keyinput29), 
        .A(n4913), .ZN(n4916) );
  INV_X1 U5436 ( .A(n4916), .ZN(n4926) );
  INV_X1 U5437 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4919) );
  AOI22_X1 U5438 ( .A1(n4919), .A2(keyinput85), .B1(n4918), .B2(keyinput89), 
        .ZN(n4917) );
  OAI221_X1 U5439 ( .B1(n4919), .B2(keyinput85), .C1(n4918), .C2(keyinput89), 
        .A(n4917), .ZN(n4921) );
  XNOR2_X1 U5440 ( .A(n2449), .B(keyinput65), .ZN(n4920) );
  NOR2_X1 U5441 ( .A1(n4921), .A2(n4920), .ZN(n4925) );
  INV_X1 U5442 ( .A(keyinput73), .ZN(n4922) );
  XNOR2_X1 U5443 ( .A(n4923), .B(n4922), .ZN(n4924) );
  AND4_X1 U5444 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n4928)
         );
  NAND4_X1 U5445 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(n4998)
         );
  AOI22_X1 U5446 ( .A1(n4934), .A2(keyinput92), .B1(keyinput104), .B2(n4933), 
        .ZN(n4932) );
  OAI221_X1 U5447 ( .B1(n4934), .B2(keyinput92), .C1(n4933), .C2(keyinput104), 
        .A(n4932), .ZN(n4946) );
  AOI22_X1 U5448 ( .A1(n4937), .A2(keyinput5), .B1(n4936), .B2(keyinput1), 
        .ZN(n4935) );
  OAI221_X1 U5449 ( .B1(n4937), .B2(keyinput5), .C1(n4936), .C2(keyinput1), 
        .A(n4935), .ZN(n4945) );
  XOR2_X1 U5450 ( .A(n4938), .B(keyinput49), .Z(n4941) );
  XNOR2_X1 U5451 ( .A(IR_REG_14__SCAN_IN), .B(keyinput41), .ZN(n4940) );
  XNOR2_X1 U5452 ( .A(IR_REG_24__SCAN_IN), .B(keyinput28), .ZN(n4939) );
  NAND3_X1 U5453 ( .A1(n4941), .A2(n4940), .A3(n4939), .ZN(n4944) );
  XNOR2_X1 U5454 ( .A(n4942), .B(keyinput16), .ZN(n4943) );
  NOR4_X1 U5455 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4996)
         );
  AOI22_X1 U5456 ( .A1(n4949), .A2(keyinput68), .B1(keyinput18), .B2(n4948), 
        .ZN(n4947) );
  OAI221_X1 U5457 ( .B1(n4949), .B2(keyinput68), .C1(n4948), .C2(keyinput18), 
        .A(n4947), .ZN(n4961) );
  INV_X1 U5458 ( .A(DATAI_21_), .ZN(n4952) );
  AOI22_X1 U5459 ( .A1(n4952), .A2(keyinput56), .B1(keyinput32), .B2(n4951), 
        .ZN(n4950) );
  OAI221_X1 U5460 ( .B1(n4952), .B2(keyinput56), .C1(n4951), .C2(keyinput32), 
        .A(n4950), .ZN(n4960) );
  INV_X1 U5461 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5462 ( .A1(n4955), .A2(keyinput12), .B1(n4954), .B2(keyinput8), 
        .ZN(n4953) );
  OAI221_X1 U5463 ( .B1(n4955), .B2(keyinput12), .C1(n4954), .C2(keyinput8), 
        .A(n4953), .ZN(n4959) );
  XNOR2_X1 U5464 ( .A(IR_REG_8__SCAN_IN), .B(keyinput35), .ZN(n4957) );
  XNOR2_X1 U5465 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput26), .ZN(n4956) );
  NAND2_X1 U5466 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  NOR4_X1 U5467 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4995)
         );
  AOI22_X1 U5468 ( .A1(n4964), .A2(keyinput82), .B1(n4963), .B2(keyinput83), 
        .ZN(n4962) );
  OAI221_X1 U5469 ( .B1(n4964), .B2(keyinput82), .C1(n4963), .C2(keyinput83), 
        .A(n4962), .ZN(n4969) );
  XNOR2_X1 U5470 ( .A(n4965), .B(keyinput78), .ZN(n4968) );
  XNOR2_X1 U5471 ( .A(n4966), .B(keyinput63), .ZN(n4967) );
  OR3_X1 U5472 ( .A1(n4969), .A2(n4968), .A3(n4967), .ZN(n4978) );
  AOI22_X1 U5473 ( .A1(n4972), .A2(keyinput38), .B1(keyinput39), .B2(n4971), 
        .ZN(n4970) );
  OAI221_X1 U5474 ( .B1(n4972), .B2(keyinput38), .C1(n4971), .C2(keyinput39), 
        .A(n4970), .ZN(n4977) );
  AOI22_X1 U5475 ( .A1(n4975), .A2(keyinput47), .B1(n4974), .B2(keyinput54), 
        .ZN(n4973) );
  OAI221_X1 U5476 ( .B1(n4975), .B2(keyinput47), .C1(n4974), .C2(keyinput54), 
        .A(n4973), .ZN(n4976) );
  NOR3_X1 U5477 ( .A1(n4978), .A2(n4977), .A3(n4976), .ZN(n4994) );
  INV_X1 U5478 ( .A(DATAI_25_), .ZN(n4980) );
  AOI22_X1 U5479 ( .A1(n4981), .A2(keyinput106), .B1(n4980), .B2(keyinput118), 
        .ZN(n4979) );
  OAI221_X1 U5480 ( .B1(n4981), .B2(keyinput106), .C1(n4980), .C2(keyinput118), 
        .A(n4979), .ZN(n4985) );
  XOR2_X1 U5481 ( .A(IR_REG_5__SCAN_IN), .B(keyinput126), .Z(n4984) );
  XOR2_X1 U5482 ( .A(DATAI_1_), .B(keyinput99), .Z(n4983) );
  XOR2_X1 U5483 ( .A(IR_REG_18__SCAN_IN), .B(keyinput86), .Z(n4982) );
  OR4_X1 U5484 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n4992) );
  XNOR2_X1 U5485 ( .A(n4986), .B(keyinput122), .ZN(n4991) );
  XNOR2_X1 U5486 ( .A(n4987), .B(keyinput90), .ZN(n4990) );
  XNOR2_X1 U5487 ( .A(n4988), .B(keyinput95), .ZN(n4989) );
  NOR4_X1 U5488 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n4993)
         );
  NAND4_X1 U5489 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n4997)
         );
  AOI211_X1 U5490 ( .C1(IR_REG_19__SCAN_IN), .C2(n4999), .A(n4998), .B(n4997), 
        .ZN(n5000) );
  NAND4_X1 U5491 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5004)
         );
  XOR2_X1 U5492 ( .A(n5005), .B(n5004), .Z(U3339) );
  CLKBUF_X1 U2403 ( .A(n2857), .Z(n2162) );
  CLKBUF_X1 U2404 ( .A(n2857), .Z(n2161) );
endmodule

