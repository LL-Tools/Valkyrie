

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173;

  INV_X2 U4780 ( .A(n5556), .ZN(n5624) );
  INV_X1 U4781 ( .A(n5558), .ZN(n5627) );
  INV_X2 U4782 ( .A(n5262), .ZN(n5556) );
  INV_X1 U4783 ( .A(n6159), .ZN(n5930) );
  INV_X1 U4784 ( .A(n5893), .ZN(n5884) );
  OAI21_X1 U4785 ( .B1(n6110), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  CLKBUF_X1 U4786 ( .A(n5899), .Z(n6065) );
  INV_X4 U4787 ( .A(n8295), .ZN(n6361) );
  OR2_X1 U4788 ( .A1(n5852), .A2(n5849), .ZN(n5850) );
  OAI21_X1 U4789 ( .B1(n6807), .B2(n4817), .A(n4815), .ZN(n4818) );
  AND2_X1 U4790 ( .A1(n6219), .A2(n5811), .ZN(n5820) );
  NAND2_X1 U4791 ( .A1(n4803), .A2(n4799), .ZN(n8726) );
  AND2_X2 U4792 ( .A1(n5861), .A2(n5950), .ZN(n6222) );
  INV_X1 U4793 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U4794 ( .A1(n9037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U4796 ( .A1(n5854), .A2(n9040), .ZN(n8305) );
  CLKBUF_X3 U4797 ( .A(n8305), .Z(n4275) );
  NAND2_X2 U4798 ( .A1(n8613), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8646) );
  XNOR2_X1 U4799 ( .A(n5865), .B(n5864), .ZN(n8672) );
  NAND2_X2 U4800 ( .A1(n8080), .A2(n9681), .ZN(n6568) );
  XNOR2_X2 U4801 ( .A(n4677), .B(n6649), .ZN(n6664) );
  NAND2_X2 U4802 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  XNOR2_X2 U4803 ( .A(n5823), .B(n5848), .ZN(n6257) );
  OAI22_X2 U4804 ( .A1(n6664), .A2(n6663), .B1(n4676), .B2(n6665), .ZN(n8548)
         );
  AOI21_X2 U4805 ( .B1(n5941), .B2(n4857), .A(n4856), .ZN(n6807) );
  NOR2_X1 U4806 ( .A1(n5480), .A2(n5479), .ZN(n9129) );
  OAI22_X1 U4807 ( .A1(n9071), .A2(n9072), .B1(n5459), .B2(n5458), .ZN(n5480)
         );
  XNOR2_X1 U4808 ( .A(n8581), .B(n8577), .ZN(n8559) );
  NAND3_X1 U4809 ( .A1(n4524), .A2(n7607), .A3(n4523), .ZN(n7606) );
  INV_X1 U4810 ( .A(n6751), .ZN(n9882) );
  INV_X4 U4811 ( .A(n8126), .ZN(n8131) );
  INV_X1 U4812 ( .A(n8528), .ZN(n5927) );
  CLKBUF_X2 U4813 ( .A(n5427), .Z(n7890) );
  INV_X2 U4814 ( .A(n5556), .ZN(n5604) );
  CLKBUF_X2 U4815 ( .A(n4992), .Z(n5427) );
  CLKBUF_X3 U4816 ( .A(n4896), .Z(n5558) );
  NOR2_X1 U4817 ( .A1(n6433), .A2(n6434), .ZN(n6528) );
  CLKBUF_X2 U4818 ( .A(n5905), .Z(n8299) );
  NAND2_X1 U4819 ( .A1(n7989), .A2(n8046), .ZN(n7048) );
  INV_X1 U4820 ( .A(n6520), .ZN(n6430) );
  AND2_X1 U4821 ( .A1(n4416), .A2(n4415), .ZN(n6338) );
  AOI21_X1 U4822 ( .B1(n4474), .B2(n4472), .A(n4471), .ZN(n4470) );
  NOR2_X1 U4823 ( .A1(n4474), .A2(n8454), .ZN(n4469) );
  NAND2_X1 U4824 ( .A1(n4526), .A2(n4343), .ZN(n5653) );
  OAI21_X1 U4825 ( .B1(n4766), .B2(n5792), .A(n4763), .ZN(n5793) );
  AND2_X1 U4826 ( .A1(n5480), .A2(n5479), .ZN(n9131) );
  NAND2_X1 U4827 ( .A1(n4586), .A2(n4585), .ZN(n9381) );
  AND2_X1 U4828 ( .A1(n8838), .A2(n6109), .ZN(n8825) );
  NAND2_X1 U4829 ( .A1(n8559), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U4830 ( .A1(n7545), .A2(n4673), .ZN(n7635) );
  NAND2_X1 U4831 ( .A1(n7153), .A2(n4671), .ZN(n7394) );
  AOI21_X1 U4832 ( .B1(n8481), .B2(n5994), .A(n4283), .ZN(n4825) );
  NAND2_X1 U4833 ( .A1(n6995), .A2(n6994), .ZN(n7153) );
  OAI21_X1 U4834 ( .B1(n4297), .B2(n4510), .A(n4506), .ZN(n4505) );
  INV_X1 U4835 ( .A(n9802), .ZN(n7373) );
  NAND2_X1 U4836 ( .A1(n6713), .A2(n6714), .ZN(n6717) );
  INV_X1 U4837 ( .A(n6679), .ZN(n8126) );
  NAND2_X1 U4838 ( .A1(n4575), .A2(n4930), .ZN(n5683) );
  INV_X1 U4839 ( .A(n4998), .ZN(n5557) );
  INV_X2 U4840 ( .A(n5060), .ZN(n5581) );
  NAND3_X1 U4841 ( .A1(n4965), .A2(n4964), .A3(n4963), .ZN(n6834) );
  NAND3_X1 U4842 ( .A1(n4299), .A2(n5917), .A3(n5916), .ZN(n8528) );
  AND4_X1 U4843 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n9918)
         );
  BUF_X2 U4844 ( .A(n5008), .Z(n5666) );
  NAND2_X1 U4845 ( .A1(n5891), .A2(n4296), .ZN(n6415) );
  INV_X1 U4846 ( .A(n7029), .ZN(n7008) );
  NAND4_X1 U4847 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n5910)
         );
  INV_X2 U4848 ( .A(n6568), .ZN(n5402) );
  NAND4_X1 U4849 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n5893)
         );
  NAND2_X1 U4850 ( .A1(n6304), .A2(n8504), .ZN(n9902) );
  INV_X2 U4851 ( .A(n5913), .ZN(n6159) );
  INV_X2 U4852 ( .A(n5904), .ZN(n8298) );
  NAND2_X1 U4853 ( .A1(n4536), .A2(n4539), .ZN(n8080) );
  XNOR2_X1 U4854 ( .A(n4925), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4928) );
  NAND2_X2 U4855 ( .A1(n6258), .A2(n6257), .ZN(n8296) );
  XNOR2_X1 U4856 ( .A(n4891), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7989) );
  XNOR2_X1 U4857 ( .A(n4895), .B(n4894), .ZN(n8046) );
  OR2_X1 U4858 ( .A1(n4899), .A2(n4540), .ZN(n4539) );
  NAND2_X1 U4859 ( .A1(n4893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U4860 ( .A1(n4887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U4861 ( .A(n4535), .B(n4902), .ZN(n9681) );
  NAND2_X1 U4862 ( .A1(n5863), .A2(n5862), .ZN(n6110) );
  AND2_X1 U4863 ( .A1(n4885), .A2(n4871), .ZN(n4892) );
  INV_X1 U4864 ( .A(n6097), .ZN(n5863) );
  AND2_X1 U4865 ( .A1(n5326), .A2(n4870), .ZN(n4885) );
  AND2_X2 U4866 ( .A1(n4701), .A2(n4702), .ZN(n4913) );
  AND2_X1 U4867 ( .A1(n4778), .A2(n5878), .ZN(n5950) );
  AND2_X1 U4868 ( .A1(n6226), .A2(n4836), .ZN(n6219) );
  AND2_X1 U4869 ( .A1(n5808), .A2(n5807), .ZN(n6226) );
  BUF_X1 U4870 ( .A(n5878), .Z(n5879) );
  AND2_X1 U4871 ( .A1(n5906), .A2(n5812), .ZN(n4778) );
  INV_X1 U4872 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4886) );
  INV_X4 U4873 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X2 U4874 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5906) );
  INV_X1 U4875 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5949) );
  INV_X1 U4876 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5951) );
  INV_X1 U4877 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5853) );
  NOR2_X1 U4878 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4762) );
  NOR2_X1 U4879 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5808) );
  NOR2_X1 U4880 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5807) );
  INV_X1 U4881 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4907) );
  INV_X4 U4882 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4883 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5813) );
  NOR2_X1 U4884 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5814) );
  NOR2_X1 U4885 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4904) );
  INV_X1 U4886 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10073) );
  AOI21_X2 U4887 ( .B1(n5708), .B2(n4862), .A(n4845), .ZN(n9434) );
  OAI22_X2 U4888 ( .A1(n9381), .A2(n5711), .B1(n9112), .B2(n9542), .ZN(n9372)
         );
  INV_X4 U4889 ( .A(n5897), .ZN(n4734) );
  NOR2_X1 U4890 ( .A1(n8725), .A2(n8445), .ZN(n4498) );
  INV_X1 U4891 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5817) );
  INV_X1 U4892 ( .A(n8083), .ZN(n5854) );
  OR2_X1 U4893 ( .A1(n9023), .A2(n8095), .ZN(n8402) );
  NAND3_X1 U4894 ( .A1(n4934), .A2(n5717), .A3(n7048), .ZN(n4896) );
  NAND2_X1 U4895 ( .A1(n4716), .A2(n4719), .ZN(n5612) );
  INV_X1 U4896 ( .A(n4720), .ZN(n4719) );
  OAI21_X1 U4897 ( .B1(n5543), .B2(n4721), .A(n5587), .ZN(n4720) );
  OAI21_X1 U4898 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(n5443) );
  OAI21_X1 U4899 ( .B1(n4913), .B2(n4393), .A(n4940), .ZN(n4958) );
  NAND2_X1 U4900 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U4901 ( .A1(n4331), .A2(n4624), .ZN(n7390) );
  AOI21_X1 U4902 ( .B1(n4801), .B2(n4805), .A(n4800), .ZN(n4799) );
  INV_X1 U4903 ( .A(n8440), .ZN(n4800) );
  INV_X1 U4904 ( .A(n6065), .ZN(n6211) );
  AND2_X1 U4905 ( .A1(n5855), .A2(n8083), .ZN(n5913) );
  INV_X2 U4906 ( .A(n5040), .ZN(n6587) );
  MUX2_X1 U4907 ( .A(n8324), .B(n8878), .S(n8323), .Z(n8329) );
  NAND2_X1 U4908 ( .A1(n4490), .A2(n8418), .ZN(n4489) );
  OAI21_X1 U4909 ( .B1(n8417), .B2(n8416), .A(n4491), .ZN(n4490) );
  AND2_X1 U4910 ( .A1(n8415), .A2(n8414), .ZN(n4491) );
  NAND2_X1 U4911 ( .A1(n8451), .A2(n4317), .ZN(n4474) );
  INV_X1 U4912 ( .A(n9897), .ZN(n6237) );
  OAI21_X1 U4913 ( .B1(n8476), .B2(n4817), .A(n5970), .ZN(n4816) );
  INV_X1 U4914 ( .A(n5346), .ZN(n5347) );
  AOI21_X1 U4915 ( .B1(n4787), .B2(n8195), .A(n4309), .ZN(n4785) );
  INV_X1 U4916 ( .A(n4468), .ZN(n4365) );
  INV_X1 U4917 ( .A(n4829), .ZN(n4828) );
  INV_X1 U4918 ( .A(n8414), .ZN(n4742) );
  INV_X1 U4919 ( .A(n8462), .ZN(n6327) );
  OR2_X1 U4920 ( .A1(n8732), .A2(n8715), .ZN(n8448) );
  NOR2_X1 U4921 ( .A1(n4814), .A2(n6165), .ZN(n4810) );
  INV_X1 U4922 ( .A(n4812), .ZN(n4807) );
  AND2_X1 U4923 ( .A1(n8123), .A2(n8759), .ZN(n6165) );
  AND2_X1 U4924 ( .A1(n8978), .A2(n8516), .ZN(n8439) );
  OR2_X1 U4925 ( .A1(n9018), .A2(n8831), .ZN(n8406) );
  NAND2_X1 U4926 ( .A1(n8296), .A2(n6361), .ZN(n5905) );
  AND2_X1 U4927 ( .A1(n8508), .A2(n6547), .ZN(n8459) );
  OR2_X1 U4928 ( .A1(n6024), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6047) );
  NOR2_X2 U4929 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5878) );
  AND2_X1 U4930 ( .A1(n5527), .A2(n5526), .ZN(n5529) );
  NOR2_X1 U4931 ( .A1(n5159), .A2(n4759), .ZN(n4758) );
  INV_X1 U4932 ( .A(n6351), .ZN(n4759) );
  INV_X1 U4933 ( .A(n7898), .ZN(n8042) );
  INV_X1 U4934 ( .A(n8085), .ZN(n4927) );
  OR2_X1 U4935 ( .A1(n9531), .A2(n9367), .ZN(n7973) );
  AOI21_X1 U4936 ( .B1(n4590), .B2(n4589), .A(n4318), .ZN(n4588) );
  INV_X1 U4937 ( .A(n4295), .ZN(n4589) );
  NOR2_X1 U4938 ( .A1(n4594), .A2(n4311), .ZN(n4592) );
  INV_X1 U4939 ( .A(n4601), .ZN(n4599) );
  INV_X1 U4940 ( .A(n7533), .ZN(n5732) );
  OR2_X1 U4941 ( .A1(n5748), .A2(n5797), .ZN(n7974) );
  INV_X1 U4942 ( .A(n9608), .ZN(n9405) );
  AND2_X1 U4943 ( .A1(n4770), .A2(n5276), .ZN(n4900) );
  NOR3_X1 U4944 ( .A1(n4773), .A2(n4771), .A3(P1_IR_REG_25__SCAN_IN), .ZN(
        n4770) );
  AND2_X1 U4945 ( .A1(n5608), .A2(n5567), .ZN(n5587) );
  OR2_X1 U4946 ( .A1(n5441), .A2(n5442), .ZN(n4715) );
  NOR2_X1 U4947 ( .A1(n5463), .A2(n4712), .ZN(n4711) );
  INV_X1 U4948 ( .A(n4713), .ZN(n4712) );
  NAND2_X1 U4949 ( .A1(n5377), .A2(n5376), .ZN(n5400) );
  OAI21_X1 U4950 ( .B1(n5324), .B2(n4724), .A(n4722), .ZN(n5377) );
  INV_X1 U4951 ( .A(n4728), .ZN(n4724) );
  AND2_X1 U4952 ( .A1(n4723), .A2(n4725), .ZN(n4722) );
  OAI21_X1 U4953 ( .B1(n5297), .B2(n5296), .A(n5295), .ZN(n5324) );
  NOR2_X1 U4954 ( .A1(n5244), .A2(n4693), .ZN(n4692) );
  INV_X1 U4955 ( .A(n5217), .ZN(n4693) );
  INV_X1 U4956 ( .A(n5173), .ZN(n5171) );
  OAI21_X1 U4957 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4907), .ZN(n4702) );
  AOI21_X1 U4958 ( .B1(n4840), .B2(n8316), .A(n4846), .ZN(n8505) );
  NAND2_X1 U4959 ( .A1(n8314), .A2(n8317), .ZN(n8316) );
  NAND2_X1 U4960 ( .A1(n5822), .A2(n4293), .ZN(n6258) );
  MUX2_X1 U4961 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5821), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5822) );
  NAND2_X1 U4962 ( .A1(n4838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  AND2_X1 U4963 ( .A1(n5809), .A2(n5810), .ZN(n4836) );
  XNOR2_X1 U4964 ( .A(n7394), .B(n7387), .ZN(n7155) );
  NAND2_X1 U4965 ( .A1(n7390), .A2(n7389), .ZN(n7543) );
  NAND2_X1 U4966 ( .A1(n8607), .A2(n8643), .ZN(n8631) );
  INV_X1 U4967 ( .A(n8631), .ZN(n4635) );
  OR2_X1 U4968 ( .A1(n6201), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8689) );
  XNOR2_X1 U4969 ( .A(n6336), .B(n8716), .ZN(n8469) );
  OR2_X1 U4970 ( .A1(n6180), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6191) );
  NOR2_X1 U4971 ( .A1(n8792), .A2(n8798), .ZN(n6141) );
  INV_X1 U4972 ( .A(n8820), .ZN(n6247) );
  AND2_X1 U4973 ( .A1(n6034), .A2(n4301), .ZN(n4821) );
  AND2_X1 U4974 ( .A1(n6197), .A2(n6196), .ZN(n8902) );
  OR2_X1 U4975 ( .A1(n8833), .A2(n8842), .ZN(n8414) );
  NAND2_X1 U4976 ( .A1(n7699), .A2(n8405), .ZN(n4745) );
  AND4_X1 U4977 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n8095)
         );
  INV_X1 U4978 ( .A(n8299), .ZN(n6113) );
  INV_X1 U4979 ( .A(n8296), .ZN(n6112) );
  NOR2_X1 U4980 ( .A1(n6493), .A2(n6308), .ZN(n6486) );
  NAND2_X1 U4981 ( .A1(n6285), .A2(n6286), .ZN(n6369) );
  INV_X1 U4982 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U4983 ( .A1(n7244), .A2(n5079), .ZN(n5081) );
  AND2_X2 U4984 ( .A1(n5385), .A2(n8046), .ZN(n7984) );
  OR2_X1 U4985 ( .A1(n5038), .A2(n5037), .ZN(n5039) );
  AND2_X1 U4986 ( .A1(n5422), .A2(n4519), .ZN(n4518) );
  NAND2_X1 U4987 ( .A1(n5417), .A2(n4520), .ZN(n4519) );
  AOI21_X1 U4988 ( .B1(n5741), .B2(n5604), .A(n5437), .ZN(n9117) );
  AOI21_X1 U4989 ( .B1(n4442), .B2(n4444), .A(n8046), .ZN(n4441) );
  OR2_X1 U4990 ( .A1(n9330), .A2(n8030), .ZN(n7898) );
  AND4_X1 U4991 ( .A1(n5046), .A2(n5045), .A3(n5044), .A4(n5043), .ZN(n7021)
         );
  CLKBUF_X3 U4992 ( .A(n4979), .Z(n5518) );
  INV_X1 U4993 ( .A(n5007), .ZN(n5040) );
  AND2_X1 U4994 ( .A1(n4927), .A2(n4926), .ZN(n4979) );
  AND2_X1 U4995 ( .A1(n4927), .A2(n4928), .ZN(n5008) );
  AND2_X1 U4996 ( .A1(n8085), .A2(n4926), .ZN(n5007) );
  NOR2_X1 U4997 ( .A1(n9374), .A2(n9389), .ZN(n9373) );
  NOR2_X1 U4998 ( .A1(n4380), .A2(n9385), .ZN(n4378) );
  AOI21_X1 U4999 ( .B1(n7312), .B2(n4611), .A(n4320), .ZN(n4610) );
  AND2_X1 U5000 ( .A1(n4900), .A2(n4898), .ZN(n4922) );
  NOR2_X1 U5001 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4919) );
  OR2_X1 U5002 ( .A1(n4883), .A2(n4882), .ZN(n4884) );
  XNOR2_X1 U5003 ( .A(n5443), .B(n5426), .ZN(n7325) );
  INV_X1 U5004 ( .A(n8738), .ZN(n8715) );
  INV_X1 U5005 ( .A(n8775), .ZN(n8916) );
  XNOR2_X1 U5006 ( .A(n5650), .B(n5649), .ZN(n6567) );
  NAND2_X1 U5007 ( .A1(n5648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5650) );
  AND2_X1 U5008 ( .A1(n5786), .A2(n5785), .ZN(n4864) );
  AOI21_X1 U5009 ( .B1(n8329), .B2(n8325), .A(n8459), .ZN(n8326) );
  INV_X1 U5010 ( .A(n8362), .ZN(n4483) );
  OAI211_X1 U5011 ( .C1(n8369), .C2(n8368), .A(n8483), .B(n8367), .ZN(n8381)
         );
  NAND2_X1 U5012 ( .A1(n4484), .A2(n4480), .ZN(n8367) );
  MUX2_X1 U5013 ( .A(n8353), .B(n8352), .S(n8459), .Z(n8369) );
  NAND2_X1 U5014 ( .A1(n8403), .A2(n8404), .ZN(n4359) );
  AOI21_X1 U5015 ( .B1(n4448), .B2(n4306), .A(n7178), .ZN(n4447) );
  OAI21_X1 U5016 ( .B1(n7783), .B2(n7778), .A(n4305), .ZN(n4448) );
  AOI21_X1 U5017 ( .B1(n4450), .B2(n7919), .A(n7784), .ZN(n4449) );
  OAI21_X1 U5018 ( .B1(n7783), .B2(n7782), .A(n7917), .ZN(n4450) );
  NAND2_X1 U5019 ( .A1(n4494), .A2(n4488), .ZN(n8425) );
  NAND2_X1 U5020 ( .A1(n4489), .A2(n8459), .ZN(n4488) );
  NAND2_X1 U5021 ( .A1(n4502), .A2(n8442), .ZN(n4501) );
  NAND2_X1 U5022 ( .A1(n4456), .A2(n4453), .ZN(n7857) );
  NAND2_X1 U5023 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  AOI21_X1 U5024 ( .B1(n4460), .B2(n4458), .A(n4457), .ZN(n4456) );
  AND2_X1 U5025 ( .A1(n7851), .A2(n7905), .ZN(n4454) );
  INV_X1 U5026 ( .A(n8454), .ZN(n4473) );
  OAI21_X1 U5027 ( .B1(n7874), .B2(n7863), .A(n7862), .ZN(n7864) );
  NAND2_X1 U5028 ( .A1(n4546), .A2(n4545), .ZN(n4544) );
  NAND2_X1 U5029 ( .A1(n5772), .A2(n5771), .ZN(n7750) );
  NAND2_X1 U5030 ( .A1(n4728), .A2(n4733), .ZN(n4723) );
  INV_X1 U5031 ( .A(SI_15_), .ZN(n5323) );
  INV_X1 U5032 ( .A(n4690), .ZN(n4689) );
  OAI21_X1 U5033 ( .B1(n4692), .B2(n4691), .A(n5268), .ZN(n4690) );
  INV_X1 U5034 ( .A(n5243), .ZN(n4691) );
  INV_X1 U5035 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5271) );
  AND2_X1 U5036 ( .A1(n4683), .A2(n4478), .ZN(n4476) );
  NAND2_X1 U5037 ( .A1(n6285), .A2(n4796), .ZN(n4795) );
  AND2_X1 U5038 ( .A1(n6286), .A2(n4797), .ZN(n4796) );
  AOI21_X1 U5039 ( .B1(n4794), .B2(n6920), .A(n4323), .ZN(n4792) );
  INV_X1 U5040 ( .A(n4794), .ZN(n4793) );
  NAND2_X1 U5041 ( .A1(n4367), .A2(n4366), .ZN(n4468) );
  NOR2_X1 U5042 ( .A1(n4469), .A2(n4325), .ZN(n4367) );
  INV_X1 U5043 ( .A(n4470), .ZN(n4366) );
  NAND2_X1 U5044 ( .A1(n6439), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5045 ( .A1(n6867), .A2(n4672), .ZN(n6989) );
  OR2_X1 U5046 ( .A1(n6868), .A2(n6715), .ZN(n4672) );
  INV_X1 U5047 ( .A(n4849), .ZN(n4830) );
  NOR2_X1 U5048 ( .A1(n8443), .A2(n4423), .ZN(n4422) );
  INV_X1 U5049 ( .A(n4425), .ZN(n4423) );
  OR2_X1 U5050 ( .A1(n8931), .A2(n8924), .ZN(n8420) );
  OR2_X1 U5051 ( .A1(n5957), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U5052 ( .A1(n9897), .A2(n9904), .ZN(n8357) );
  OR2_X1 U5053 ( .A1(n5910), .A2(n6796), .ZN(n8330) );
  NAND2_X1 U5054 ( .A1(n8983), .A2(n6251), .ZN(n4812) );
  OR2_X1 U5055 ( .A1(n8123), .A2(n6251), .ZN(n8435) );
  OR2_X1 U5056 ( .A1(n8921), .A2(n8925), .ZN(n8432) );
  AND2_X1 U5057 ( .A1(n8371), .A2(n4401), .ZN(n4400) );
  NAND2_X1 U5058 ( .A1(n8364), .A2(n4402), .ZN(n4401) );
  AOI21_X1 U5059 ( .B1(n6962), .B2(n8365), .A(n6240), .ZN(n7033) );
  INV_X1 U5060 ( .A(n4816), .ZN(n4815) );
  OR2_X1 U5061 ( .A1(n5995), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U5062 ( .A1(n6352), .A2(n6350), .ZN(n5108) );
  INV_X1 U5063 ( .A(n8044), .ZN(n4444) );
  AOI21_X1 U5064 ( .B1(n4559), .B2(n4561), .A(n4558), .ZN(n4557) );
  INV_X1 U5065 ( .A(n7877), .ZN(n4558) );
  OR2_X1 U5066 ( .A1(n5776), .A2(n6846), .ZN(n7975) );
  NOR2_X1 U5067 ( .A1(n5776), .A2(n4552), .ZN(n4550) );
  NAND2_X1 U5068 ( .A1(n4284), .A2(n9504), .ZN(n4375) );
  AND2_X1 U5069 ( .A1(n4286), .A2(n9504), .ZN(n4372) );
  INV_X1 U5070 ( .A(n4376), .ZN(n4374) );
  AOI21_X1 U5071 ( .B1(n4284), .B2(n4623), .A(n4326), .ZN(n4376) );
  NOR2_X1 U5072 ( .A1(n7669), .A2(n9581), .ZN(n4546) );
  AND2_X1 U5073 ( .A1(n4294), .A2(n7938), .ZN(n4392) );
  AND2_X1 U5074 ( .A1(n7669), .A2(n9178), .ZN(n5700) );
  NAND2_X1 U5075 ( .A1(n5695), .A2(n4530), .ZN(n4529) );
  NOR2_X1 U5076 ( .A1(n7811), .A2(n9838), .ZN(n4530) );
  INV_X1 U5077 ( .A(n4395), .ZN(n8007) );
  OAI21_X1 U5078 ( .B1(n7787), .B2(n7791), .A(n7795), .ZN(n4395) );
  XNOR2_X1 U5079 ( .A(n5683), .B(n4369), .ZN(n6836) );
  INV_X1 U5080 ( .A(n9613), .ZN(n9441) );
  AND2_X1 U5081 ( .A1(n7599), .A2(n4542), .ZN(n9491) );
  NOR2_X1 U5082 ( .A1(n4544), .A2(n9492), .ZN(n4542) );
  INV_X1 U5083 ( .A(n7476), .ZN(n7226) );
  NAND2_X1 U5084 ( .A1(n4303), .A2(n4278), .ZN(n4773) );
  INV_X1 U5085 ( .A(n4302), .ZN(n4771) );
  NAND2_X1 U5086 ( .A1(n5544), .A2(n5543), .ZN(n5563) );
  NOR2_X1 U5087 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4775) );
  AND2_X1 U5088 ( .A1(n5537), .A2(n5515), .ZN(n5535) );
  INV_X1 U5089 ( .A(n5462), .ZN(n4709) );
  INV_X1 U5090 ( .A(n4711), .ZN(n4707) );
  INV_X1 U5091 ( .A(n5481), .ZN(n4706) );
  INV_X1 U5092 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4882) );
  OAI21_X1 U5093 ( .B1(n5400), .B2(n5380), .A(n5379), .ZN(n5425) );
  OAI21_X1 U5094 ( .B1(n4913), .B2(n4911), .A(n4910), .ZN(n4960) );
  OAI21_X1 U5095 ( .B1(n6683), .B2(n4783), .A(n6911), .ZN(n4782) );
  NAND2_X1 U5096 ( .A1(n6438), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5097 ( .A1(n5879), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U5098 ( .A1(n6529), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4678) );
  OAI21_X1 U5099 ( .B1(n6647), .B2(n6646), .A(n8537), .ZN(n8542) );
  NAND2_X1 U5100 ( .A1(n8542), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5101 ( .A1(n8533), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4669) );
  OR2_X1 U5102 ( .A1(n6702), .A2(n6701), .ZN(n6857) );
  NAND2_X1 U5103 ( .A1(n6717), .A2(n6716), .ZN(n6867) );
  XNOR2_X1 U5104 ( .A(n6989), .B(n6974), .ZN(n6869) );
  NAND2_X1 U5105 ( .A1(n7151), .A2(n7150), .ZN(n7385) );
  NAND2_X1 U5106 ( .A1(n7396), .A2(n7397), .ZN(n7399) );
  NAND2_X1 U5107 ( .A1(n7399), .A2(n7398), .ZN(n7545) );
  XNOR2_X1 U5108 ( .A(n7635), .B(n7630), .ZN(n7547) );
  NAND2_X1 U5109 ( .A1(n4655), .A2(n4653), .ZN(n8607) );
  NOR2_X1 U5110 ( .A1(n4654), .A2(n4356), .ZN(n4653) );
  INV_X1 U5111 ( .A(n4656), .ZN(n4654) );
  NAND2_X1 U5112 ( .A1(n4635), .A2(n4355), .ZN(n4626) );
  NOR2_X1 U5113 ( .A1(n8469), .A2(n4754), .ZN(n4753) );
  INV_X1 U5114 ( .A(n8319), .ZN(n4754) );
  OR2_X1 U5115 ( .A1(n8968), .A2(n8902), .ZN(n8319) );
  OR2_X1 U5116 ( .A1(n8151), .A2(n8902), .ZN(n4849) );
  OR2_X1 U5117 ( .A1(n4421), .A2(n8756), .ZN(n4418) );
  INV_X1 U5118 ( .A(n4422), .ZN(n4421) );
  AOI21_X1 U5119 ( .B1(n4422), .B2(n4420), .A(n4334), .ZN(n4419) );
  INV_X1 U5120 ( .A(n4427), .ZN(n4420) );
  OR2_X1 U5121 ( .A1(n8444), .A2(n8446), .ZN(n8725) );
  OR2_X1 U5122 ( .A1(n6144), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6154) );
  AOI21_X1 U5123 ( .B1(n4833), .B2(n8808), .A(n4319), .ZN(n4832) );
  AND2_X1 U5124 ( .A1(n4736), .A2(n8418), .ZN(n4741) );
  NOR2_X1 U5125 ( .A1(n6246), .A2(n4742), .ZN(n4737) );
  NAND2_X1 U5126 ( .A1(n9007), .A2(n8944), .ZN(n4834) );
  AND2_X1 U5127 ( .A1(n8797), .A2(n4834), .ZN(n4833) );
  OR2_X1 U5128 ( .A1(n8807), .A2(n8808), .ZN(n4835) );
  AND2_X1 U5129 ( .A1(n8372), .A2(n7137), .ZN(n8364) );
  AND2_X1 U5130 ( .A1(n8375), .A2(n8374), .ZN(n8483) );
  NAND2_X1 U5131 ( .A1(n7033), .A2(n8356), .ZN(n7138) );
  NAND2_X1 U5132 ( .A1(n4823), .A2(n6022), .ZN(n4822) );
  OR2_X1 U5133 ( .A1(n6950), .A2(n6952), .ZN(n6962) );
  OR2_X1 U5134 ( .A1(n6964), .A2(n8481), .ZN(n6966) );
  NAND2_X1 U5135 ( .A1(n8350), .A2(n8357), .ZN(n8478) );
  NAND2_X1 U5136 ( .A1(n6807), .A2(n8476), .ZN(n6806) );
  INV_X1 U5137 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5138 ( .A1(n5854), .A2(n5855), .ZN(n5899) );
  OR2_X1 U5139 ( .A1(n5904), .A2(n6365), .ZN(n5882) );
  NAND2_X1 U5140 ( .A1(n6210), .A2(n6209), .ZN(n6312) );
  AND2_X1 U5141 ( .A1(n6207), .A2(n6206), .ZN(n8716) );
  NAND2_X1 U5142 ( .A1(n4812), .A2(n4809), .ZN(n4808) );
  INV_X1 U5143 ( .A(n6164), .ZN(n4809) );
  AOI21_X1 U5144 ( .B1(n4427), .B2(n8321), .A(n4426), .ZN(n4425) );
  INV_X1 U5145 ( .A(n8435), .ZN(n4426) );
  NOR2_X1 U5146 ( .A1(n8434), .A2(n4428), .ZN(n4427) );
  AND2_X1 U5147 ( .A1(n8441), .A2(n8440), .ZN(n8737) );
  OR2_X1 U5148 ( .A1(n8758), .A2(n6164), .ZN(n4811) );
  AND2_X1 U5149 ( .A1(n6250), .A2(n8435), .ZN(n8747) );
  AND2_X1 U5150 ( .A1(n8432), .A2(n8430), .ZN(n8767) );
  INV_X1 U5151 ( .A(n4274), .ZN(n6270) );
  AND2_X1 U5152 ( .A1(n8415), .A2(n8418), .ZN(n8808) );
  NOR2_X1 U5153 ( .A1(n4746), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U5154 ( .A1(n6247), .A2(n6246), .ZN(n8822) );
  AND4_X1 U5155 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8841)
         );
  NAND2_X1 U5156 ( .A1(n8854), .A2(n4308), .ZN(n7694) );
  AOI21_X1 U5157 ( .B1(n4408), .B2(n4410), .A(n4405), .ZN(n4404) );
  INV_X1 U5158 ( .A(n8402), .ZN(n4405) );
  AND2_X1 U5159 ( .A1(n8402), .A2(n8400), .ZN(n8853) );
  NOR2_X1 U5160 ( .A1(n4750), .A2(n4412), .ZN(n4411) );
  INV_X1 U5161 ( .A(n6243), .ZN(n4412) );
  INV_X1 U5162 ( .A(n8397), .ZN(n4750) );
  NAND2_X1 U5163 ( .A1(n4820), .A2(n4819), .ZN(n7422) );
  AOI21_X1 U5164 ( .B1(n4821), .B2(n6021), .A(n4281), .ZN(n4819) );
  INV_X1 U5165 ( .A(n8522), .ZN(n9920) );
  INV_X1 U5166 ( .A(n9919), .ZN(n9872) );
  INV_X1 U5167 ( .A(n9874), .ZN(n9917) );
  NAND2_X1 U5168 ( .A1(n6542), .A2(n8459), .ZN(n9919) );
  NAND2_X1 U5169 ( .A1(n6302), .A2(n6301), .ZN(n6491) );
  AND2_X1 U5170 ( .A1(n4752), .A2(n5848), .ZN(n4751) );
  OR2_X1 U5171 ( .A1(n4858), .A2(n6276), .ZN(n6277) );
  AND2_X1 U5172 ( .A1(n6226), .A2(n5809), .ZN(n6221) );
  OR2_X1 U5173 ( .A1(n6224), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6097) );
  XNOR2_X1 U5174 ( .A(n6035), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7546) );
  NOR2_X1 U5175 ( .A1(n6007), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6010) );
  INV_X1 U5176 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5649) );
  AND2_X1 U5177 ( .A1(n5153), .A2(n5152), .ZN(n7474) );
  INV_X1 U5178 ( .A(n5417), .ZN(n4515) );
  AND2_X1 U5179 ( .A1(n5158), .A2(n6350), .ZN(n4522) );
  NAND2_X1 U5180 ( .A1(n5210), .A2(n4756), .ZN(n4521) );
  NOR2_X1 U5181 ( .A1(n5224), .A2(n5223), .ZN(n5252) );
  INV_X1 U5182 ( .A(n5061), .ZN(n5059) );
  INV_X1 U5183 ( .A(n5039), .ZN(n4509) );
  INV_X1 U5184 ( .A(n7130), .ZN(n4510) );
  NOR2_X1 U5185 ( .A1(n4768), .A2(n4282), .ZN(n4765) );
  OR2_X1 U5186 ( .A1(n9147), .A2(n9148), .ZN(n4768) );
  NAND2_X1 U5187 ( .A1(n9110), .A2(n4767), .ZN(n4766) );
  INV_X1 U5188 ( .A(n9078), .ZN(n4767) );
  NOR2_X1 U5189 ( .A1(n5659), .A2(n8051), .ZN(n5664) );
  INV_X1 U5190 ( .A(n5316), .ZN(n5313) );
  AND2_X1 U5191 ( .A1(n7906), .A2(n4335), .ZN(n4445) );
  INV_X1 U5192 ( .A(n4550), .ZN(n4549) );
  NAND2_X1 U5193 ( .A1(n4541), .A2(n9394), .ZN(n9389) );
  NAND2_X1 U5194 ( .A1(n9437), .A2(n4381), .ZN(n4379) );
  NOR2_X1 U5195 ( .A1(n4565), .A2(n4457), .ZN(n4381) );
  INV_X1 U5196 ( .A(n5745), .ZN(n4565) );
  INV_X1 U5197 ( .A(n7950), .ZN(n4563) );
  INV_X1 U5198 ( .A(n5744), .ZN(n4564) );
  AOI21_X1 U5199 ( .B1(n4588), .B2(n4591), .A(n4324), .ZN(n4585) );
  INV_X1 U5200 ( .A(n7860), .ZN(n9399) );
  NAND2_X1 U5201 ( .A1(n9435), .A2(n5744), .ZN(n9423) );
  INV_X1 U5202 ( .A(n4574), .ZN(n9437) );
  OAI21_X1 U5203 ( .B1(n9452), .B2(n9449), .A(n7962), .ZN(n4574) );
  NAND2_X1 U5204 ( .A1(n9437), .A2(n9436), .ZN(n9435) );
  OAI21_X1 U5205 ( .B1(n9471), .B2(n9469), .A(n7839), .ZN(n9452) );
  AND2_X1 U5206 ( .A1(n9492), .A2(n9175), .ZN(n5706) );
  NOR2_X1 U5207 ( .A1(n9581), .A2(n9177), .ZN(n5701) );
  INV_X1 U5208 ( .A(n5737), .ZN(n4391) );
  NAND2_X1 U5209 ( .A1(n5737), .A2(n4392), .ZN(n7711) );
  AOI21_X1 U5210 ( .B1(n4604), .B2(n4602), .A(n4332), .ZN(n4601) );
  INV_X1 U5211 ( .A(n5699), .ZN(n4602) );
  NAND2_X1 U5212 ( .A1(n7530), .A2(n5697), .ZN(n7615) );
  NAND2_X1 U5213 ( .A1(n4382), .A2(n7806), .ZN(n7533) );
  OR2_X1 U5214 ( .A1(n5730), .A2(n4566), .ZN(n4383) );
  NAND2_X1 U5215 ( .A1(n7293), .A2(n5694), .ZN(n7439) );
  NAND2_X1 U5216 ( .A1(n7223), .A2(n5691), .ZN(n7282) );
  NAND2_X1 U5217 ( .A1(n7282), .A2(n7281), .ZN(n7280) );
  OAI21_X1 U5218 ( .B1(n7999), .B2(n4584), .A(n7178), .ZN(n4580) );
  INV_X1 U5219 ( .A(n5690), .ZN(n4584) );
  NAND2_X1 U5220 ( .A1(n7197), .A2(n5689), .ZN(n7018) );
  NAND2_X1 U5221 ( .A1(n7018), .A2(n7999), .ZN(n7017) );
  AND2_X1 U5222 ( .A1(n8041), .A2(n6773), .ZN(n9425) );
  INV_X1 U5223 ( .A(n9458), .ZN(n9427) );
  NOR2_X1 U5224 ( .A1(n6905), .A2(n6909), .ZN(n7199) );
  NAND2_X1 U5225 ( .A1(n4452), .A2(n5721), .ZN(n6830) );
  INV_X1 U5226 ( .A(n9425), .ZN(n9456) );
  AOI21_X1 U5227 ( .B1(n9815), .B2(n5755), .A(n5754), .ZN(n7004) );
  NAND2_X1 U5228 ( .A1(n8046), .A2(n5749), .ZN(n9509) );
  NAND2_X1 U5229 ( .A1(n7767), .A2(n7766), .ZN(n9330) );
  OAI21_X1 U5230 ( .B1(n9354), .B2(n4620), .A(n5714), .ZN(n4619) );
  NAND2_X1 U5231 ( .A1(n5713), .A2(n5712), .ZN(n4620) );
  NOR2_X1 U5232 ( .A1(n9354), .A2(n4622), .ZN(n4621) );
  INV_X1 U5233 ( .A(n5712), .ZN(n4622) );
  NAND2_X1 U5234 ( .A1(n5569), .A2(n5568), .ZN(n9374) );
  NAND2_X1 U5235 ( .A1(n5493), .A2(n5492), .ZN(n9550) );
  INV_X1 U5236 ( .A(n7203), .ZN(n9817) );
  OR2_X1 U5237 ( .A1(n7030), .A2(n7984), .ZN(n9831) );
  AND2_X1 U5238 ( .A1(n6568), .A2(n6361), .ZN(n4984) );
  OAI21_X1 U5239 ( .B1(n4901), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4899) );
  INV_X1 U5240 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4540) );
  INV_X1 U5241 ( .A(n4917), .ZN(n4538) );
  XNOR2_X1 U5242 ( .A(n5593), .B(n5592), .ZN(n7734) );
  XNOR2_X1 U5243 ( .A(n5588), .B(n5587), .ZN(n7729) );
  NAND2_X1 U5244 ( .A1(n5563), .A2(n5562), .ZN(n5588) );
  NAND2_X1 U5245 ( .A1(n4710), .A2(n5462), .ZN(n5483) );
  NAND2_X1 U5246 ( .A1(n4714), .A2(n4711), .ZN(n4710) );
  INV_X1 U5247 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5248 ( .A1(n4727), .A2(n5348), .ZN(n5375) );
  NAND2_X1 U5249 ( .A1(n4731), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U5250 ( .A1(n4688), .A2(n5243), .ZN(n5269) );
  NAND2_X1 U5251 ( .A1(n5218), .A2(n4692), .ZN(n4688) );
  NAND2_X1 U5252 ( .A1(n5218), .A2(n5217), .ZN(n5245) );
  XNOR2_X1 U5253 ( .A(n4497), .B(n5192), .ZN(n6409) );
  NAND2_X1 U5254 ( .A1(n5162), .A2(n5161), .ZN(n4497) );
  NAND2_X1 U5255 ( .A1(n5071), .A2(n5070), .ZN(n5075) );
  NAND2_X1 U5256 ( .A1(n4986), .A2(n4985), .ZN(n4990) );
  OR2_X1 U5257 ( .A1(n8878), .A2(n6551), .ZN(n6579) );
  AND4_X1 U5258 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8842)
         );
  NOR2_X1 U5259 ( .A1(n8087), .A2(n8520), .ZN(n4791) );
  AND2_X1 U5260 ( .A1(n6485), .A2(n6484), .ZN(n8280) );
  NAND2_X1 U5261 ( .A1(n8503), .A2(n4363), .ZN(n4362) );
  INV_X1 U5262 ( .A(n4364), .ZN(n4363) );
  OAI21_X1 U5263 ( .B1(n8505), .B2(n8504), .A(n8502), .ZN(n4364) );
  NAND2_X1 U5264 ( .A1(n4293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U5265 ( .A(n6220), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U5266 ( .A1(n6186), .A2(n6185), .ZN(n8738) );
  NAND2_X1 U5267 ( .A1(n6177), .A2(n6176), .ZN(n8516) );
  NAND2_X1 U5268 ( .A1(n5860), .A2(n5859), .ZN(n8759) );
  NAND2_X1 U5269 ( .A1(n6162), .A2(n6161), .ZN(n8775) );
  INV_X1 U5270 ( .A(n6438), .ZN(n6461) );
  XNOR2_X1 U5271 ( .A(n4668), .B(n4667), .ZN(n6648) );
  NOR2_X1 U5272 ( .A1(n6648), .A2(n6955), .ZN(n6698) );
  OR2_X1 U5273 ( .A1(n7152), .A2(n7160), .ZN(n4624) );
  XNOR2_X1 U5274 ( .A(n7385), .B(n7395), .ZN(n7152) );
  NAND2_X1 U5275 ( .A1(n7636), .A2(n4665), .ZN(n4663) );
  NOR2_X1 U5276 ( .A1(n7636), .A2(n4665), .ZN(n4664) );
  INV_X1 U5277 ( .A(n8678), .ZN(n8624) );
  INV_X1 U5278 ( .A(n6267), .ZN(n6268) );
  OAI21_X1 U5279 ( .B1(n8701), .B2(n9866), .A(n6266), .ZN(n6267) );
  INV_X1 U5280 ( .A(n8516), .ZN(n8901) );
  NAND2_X1 U5281 ( .A1(n6115), .A2(n6114), .ZN(n8833) );
  NAND2_X1 U5282 ( .A1(n6089), .A2(n6088), .ZN(n8098) );
  INV_X1 U5283 ( .A(n6312), .ZN(n8695) );
  NAND2_X1 U5284 ( .A1(n4417), .A2(n9884), .ZN(n4416) );
  AOI21_X1 U5285 ( .B1(n8702), .B2(n9902), .A(n6323), .ZN(n4415) );
  INV_X1 U5286 ( .A(n8709), .ZN(n4417) );
  AND2_X1 U5287 ( .A1(n6299), .A2(n6298), .ZN(n6727) );
  INV_X1 U5288 ( .A(n7387), .ZN(n7395) );
  NOR2_X1 U5289 ( .A1(n7731), .A2(n7692), .ZN(n4880) );
  AND2_X1 U5290 ( .A1(n5094), .A2(n5093), .ZN(n9825) );
  AND4_X1 U5291 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9457)
         );
  NAND2_X1 U5292 ( .A1(n5614), .A2(n5613), .ZN(n5748) );
  NAND2_X1 U5293 ( .A1(n5446), .A2(n5445), .ZN(n9562) );
  AND4_X1 U5294 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n7131)
         );
  NAND2_X1 U5295 ( .A1(n4516), .A2(n4518), .ZN(n9120) );
  NAND2_X1 U5296 ( .A1(n4517), .A2(n5417), .ZN(n4516) );
  NAND2_X1 U5297 ( .A1(n5429), .A2(n5428), .ZN(n5741) );
  INV_X1 U5298 ( .A(n9151), .ZN(n9671) );
  INV_X1 U5299 ( .A(n4441), .ZN(n4440) );
  AND2_X1 U5300 ( .A1(n4445), .A2(n4434), .ZN(n4432) );
  AOI21_X1 U5301 ( .B1(n4435), .B2(n4434), .A(n4357), .ZN(n4433) );
  NAND2_X1 U5302 ( .A1(n4438), .A2(n4436), .ZN(n4435) );
  INV_X1 U5303 ( .A(n9457), .ZN(n9426) );
  INV_X1 U5304 ( .A(n7585), .ZN(n9185) );
  NAND4_X1 U5305 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n9191)
         );
  OR2_X1 U5306 ( .A1(n5040), .A2(n4978), .ZN(n4982) );
  NAND2_X1 U5307 ( .A1(n4864), .A2(n4572), .ZN(n4571) );
  AND2_X1 U5308 ( .A1(n5787), .A2(n4573), .ZN(n4572) );
  INV_X1 U5309 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5310 ( .A1(n8339), .A2(n8338), .ZN(n8347) );
  NAND2_X1 U5311 ( .A1(n4487), .A2(n4486), .ZN(n4485) );
  INV_X1 U5312 ( .A(n8365), .ZN(n4486) );
  OAI21_X1 U5313 ( .B1(n8366), .B2(n8363), .A(n4481), .ZN(n4480) );
  NOR2_X1 U5314 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U5315 ( .A1(n8361), .A2(n8459), .ZN(n4482) );
  NAND2_X1 U5316 ( .A1(n4493), .A2(n4492), .ZN(n8417) );
  NAND2_X1 U5317 ( .A1(n8410), .A2(n8459), .ZN(n4492) );
  OAI21_X1 U5318 ( .B1(n4449), .B2(n7905), .A(n4447), .ZN(n7794) );
  NAND2_X1 U5319 ( .A1(n7840), .A2(n7954), .ZN(n4460) );
  NOR2_X1 U5320 ( .A1(n7905), .A2(n4459), .ZN(n4458) );
  INV_X1 U5321 ( .A(n7841), .ZN(n4459) );
  NAND2_X1 U5322 ( .A1(n7850), .A2(n7849), .ZN(n4455) );
  INV_X1 U5323 ( .A(n8737), .ZN(n4500) );
  OAI21_X1 U5324 ( .B1(n4462), .B2(n4461), .A(n7861), .ZN(n7874) );
  NOR2_X1 U5325 ( .A1(n7858), .A2(n7897), .ZN(n4461) );
  OAI21_X1 U5326 ( .B1(n7859), .B2(n7905), .A(n9399), .ZN(n4462) );
  NAND2_X1 U5327 ( .A1(n4696), .A2(n8513), .ZN(n8318) );
  NAND2_X1 U5328 ( .A1(n8458), .A2(n8310), .ZN(n8470) );
  NAND2_X1 U5329 ( .A1(n8470), .A2(n4495), .ZN(n4694) );
  INV_X1 U5330 ( .A(n8456), .ZN(n4471) );
  NAND2_X1 U5331 ( .A1(n6217), .A2(n4473), .ZN(n4472) );
  INV_X1 U5332 ( .A(n8759), .ZN(n6251) );
  INV_X1 U5333 ( .A(n5956), .ZN(n4817) );
  NOR2_X1 U5334 ( .A1(n7870), .A2(n7897), .ZN(n7871) );
  AND2_X1 U5335 ( .A1(n7789), .A2(n7229), .ZN(n7787) );
  INV_X1 U5336 ( .A(n5562), .ZN(n4721) );
  NOR2_X1 U5337 ( .A1(n4718), .A2(n4721), .ZN(n4717) );
  INV_X1 U5338 ( .A(n5537), .ZN(n4718) );
  NOR2_X1 U5339 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4873) );
  NOR2_X1 U5340 ( .A1(n5374), .A2(n4726), .ZN(n4725) );
  INV_X1 U5341 ( .A(n5348), .ZN(n4726) );
  NAND2_X1 U5342 ( .A1(n5351), .A2(n10088), .ZN(n5376) );
  INV_X1 U5343 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U5344 ( .A1(n5273), .A2(n5272), .ZN(n5295) );
  INV_X1 U5345 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5219) );
  NOR2_X1 U5346 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  INV_X1 U5347 ( .A(n5161), .ZN(n4699) );
  INV_X1 U5348 ( .A(n5192), .ZN(n4700) );
  INV_X1 U5349 ( .A(n5113), .ZN(n4684) );
  AOI21_X1 U5350 ( .B1(n5083), .B2(n4479), .A(n4327), .ZN(n4478) );
  INV_X1 U5351 ( .A(n5074), .ZN(n4479) );
  NAND2_X1 U5352 ( .A1(n8467), .A2(n8311), .ZN(n8312) );
  INV_X1 U5353 ( .A(n8470), .ZN(n8311) );
  INV_X1 U5354 ( .A(SI_17_), .ZN(n10088) );
  AOI21_X1 U5355 ( .B1(n6511), .B2(n6512), .A(n4368), .ZN(n6431) );
  OR2_X1 U5356 ( .A1(n7154), .A2(n6993), .ZN(n4671) );
  INV_X1 U5357 ( .A(n8580), .ZN(n4658) );
  NAND2_X1 U5358 ( .A1(n8556), .A2(n4670), .ZN(n8581) );
  OR2_X1 U5359 ( .A1(n8558), .A2(n8557), .ZN(n4670) );
  OR2_X1 U5360 ( .A1(n6312), .A2(n9990), .ZN(n8317) );
  NOR2_X1 U5361 ( .A1(n4806), .A2(n8439), .ZN(n4804) );
  NOR2_X1 U5362 ( .A1(n8439), .A2(n4802), .ZN(n4801) );
  INV_X1 U5363 ( .A(n4808), .ZN(n4802) );
  NAND2_X1 U5364 ( .A1(n5844), .A2(n5843), .ZN(n6144) );
  OR2_X1 U5365 ( .A1(n6127), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6134) );
  INV_X1 U5366 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U5367 ( .A1(n4734), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5874) );
  OR2_X1 U5368 ( .A1(n6369), .A2(n6297), .ZN(n6324) );
  AND2_X1 U5369 ( .A1(n4795), .A2(n6379), .ZN(n6728) );
  OR2_X1 U5370 ( .A1(n8792), .A2(n8934), .ZN(n8427) );
  INV_X1 U5371 ( .A(n8396), .ZN(n4410) );
  INV_X1 U5372 ( .A(n4409), .ZN(n4408) );
  OAI21_X1 U5373 ( .B1(n4411), .B2(n4410), .A(n8400), .ZN(n4409) );
  NOR2_X1 U5374 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4752) );
  INV_X1 U5375 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6275) );
  INV_X1 U5376 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5809) );
  OR2_X1 U5377 ( .A1(n5983), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5995) );
  INV_X1 U5378 ( .A(n4758), .ZN(n4757) );
  INV_X1 U5379 ( .A(n9094), .ZN(n4520) );
  AND2_X1 U5380 ( .A1(n5289), .A2(n5293), .ZN(n4525) );
  NOR2_X1 U5381 ( .A1(n8047), .A2(n4443), .ZN(n4442) );
  NOR2_X1 U5382 ( .A1(n4444), .A2(n8027), .ZN(n4443) );
  OR2_X1 U5383 ( .A1(n5741), .A2(n9455), .ZN(n7839) );
  NOR2_X1 U5384 ( .A1(n4612), .A2(n4609), .ZN(n4608) );
  INV_X1 U5385 ( .A(n7281), .ZN(n4609) );
  INV_X1 U5386 ( .A(n5692), .ZN(n4611) );
  NOR2_X1 U5387 ( .A1(n7226), .A2(n4532), .ZN(n4531) );
  INV_X1 U5388 ( .A(n4533), .ZN(n4532) );
  AND2_X1 U5389 ( .A1(n7921), .A2(n4612), .ZN(n4384) );
  NAND2_X1 U5390 ( .A1(n7226), .A2(n7524), .ZN(n7789) );
  NOR2_X1 U5391 ( .A1(n7188), .A2(n9802), .ZN(n4533) );
  INV_X1 U5392 ( .A(n6836), .ZN(n7992) );
  INV_X1 U5393 ( .A(n5671), .ZN(n8041) );
  OR2_X1 U5394 ( .A1(n9562), .A2(n9475), .ZN(n9459) );
  INV_X1 U5395 ( .A(n4544), .ZN(n4543) );
  NAND2_X1 U5396 ( .A1(n6839), .A2(n7910), .ZN(n6879) );
  AND2_X1 U5397 ( .A1(n7564), .A2(n7993), .ZN(n5749) );
  XNOR2_X1 U5398 ( .A(n7750), .B(n7751), .ZN(n7748) );
  AOI21_X1 U5399 ( .B1(n5612), .B2(n5611), .A(n5610), .ZN(n5768) );
  INV_X1 U5400 ( .A(n5609), .ZN(n5610) );
  AND2_X1 U5401 ( .A1(n5562), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U5402 ( .A1(n4881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U5403 ( .A1(n5441), .A2(n5442), .ZN(n4713) );
  INV_X1 U5404 ( .A(SI_20_), .ZN(n5442) );
  NOR2_X1 U5405 ( .A1(n4729), .A2(n5349), .ZN(n4728) );
  INV_X1 U5406 ( .A(n4730), .ZN(n4729) );
  NAND2_X1 U5407 ( .A1(n5322), .A2(n5323), .ZN(n4730) );
  AOI21_X1 U5408 ( .B1(n4689), .B2(n4691), .A(n4328), .ZN(n4687) );
  INV_X1 U5409 ( .A(SI_11_), .ZN(n5167) );
  NAND2_X1 U5410 ( .A1(n4682), .A2(n4680), .ZN(n5160) );
  AOI21_X1 U5411 ( .B1(n5109), .B2(n4683), .A(n4681), .ZN(n4680) );
  NAND2_X1 U5412 ( .A1(n4476), .A2(n4477), .ZN(n4682) );
  INV_X1 U5413 ( .A(n5119), .ZN(n4681) );
  OAI21_X1 U5414 ( .B1(n8295), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4396), .ZN(
        n5017) );
  NAND2_X1 U5415 ( .A1(n8295), .A2(n4397), .ZN(n4396) );
  INV_X1 U5416 ( .A(n8262), .ZN(n8107) );
  INV_X1 U5417 ( .A(n4788), .ZN(n4787) );
  OAI21_X1 U5418 ( .B1(n8225), .B2(n8195), .A(n8194), .ZN(n4788) );
  NAND2_X1 U5419 ( .A1(n8224), .A2(n8225), .ZN(n8223) );
  NAND2_X1 U5420 ( .A1(n5846), .A2(n5845), .ZN(n6171) );
  INV_X1 U5421 ( .A(n6156), .ZN(n5846) );
  NAND2_X1 U5422 ( .A1(n6683), .A2(n6684), .ZN(n6767) );
  CLKBUF_X1 U5423 ( .A(n8183), .Z(n8232) );
  XNOR2_X1 U5424 ( .A(n6679), .B(n8884), .ZN(n6552) );
  NAND2_X1 U5425 ( .A1(n4468), .A2(n4466), .ZN(n4465) );
  NAND2_X1 U5426 ( .A1(n4365), .A2(n4495), .ZN(n4467) );
  INV_X1 U5427 ( .A(n8460), .ZN(n4466) );
  AND4_X1 U5428 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n7488)
         );
  OAI211_X1 U5429 ( .C1(n4652), .C2(n4645), .A(n6516), .B(n4641), .ZN(n6514)
         );
  INV_X1 U5430 ( .A(n4651), .ZN(n4650) );
  OAI22_X1 U5431 ( .A1(n4277), .A2(n6429), .B1(n5886), .B2(n4639), .ZN(n6512)
         );
  XNOR2_X1 U5432 ( .A(n6431), .B(n6478), .ZN(n6468) );
  OR2_X1 U5433 ( .A1(n6469), .A2(n6852), .ZN(n6471) );
  NAND2_X1 U5434 ( .A1(n4659), .A2(n8538), .ZN(n4660) );
  INV_X1 U5435 ( .A(n4677), .ZN(n4676) );
  XNOR2_X1 U5436 ( .A(n6712), .B(n6697), .ZN(n6667) );
  NAND2_X1 U5437 ( .A1(n6667), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U5438 ( .A1(n6857), .A2(n6856), .ZN(n4666) );
  OR2_X1 U5439 ( .A1(n6979), .A2(n6978), .ZN(n7151) );
  NAND2_X1 U5440 ( .A1(n6991), .A2(n6992), .ZN(n6995) );
  INV_X1 U5441 ( .A(n7542), .ZN(n4665) );
  OR2_X1 U5442 ( .A1(n7546), .A2(n7407), .ZN(n4673) );
  AOI21_X1 U5443 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8554), .A(n8553), .ZN(
        n8576) );
  NAND2_X1 U5444 ( .A1(n8579), .A2(n4658), .ZN(n4656) );
  OR2_X1 U5445 ( .A1(n8555), .A2(n4657), .ZN(n4655) );
  NAND2_X1 U5446 ( .A1(n4658), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4657) );
  OR2_X1 U5447 ( .A1(n8609), .A2(n10130), .ZN(n8632) );
  NAND2_X1 U5448 ( .A1(n4636), .A2(n4633), .ZN(n4631) );
  OAI21_X1 U5449 ( .B1(n8666), .B2(n4629), .A(n4628), .ZN(n4627) );
  NOR2_X1 U5450 ( .A1(n4638), .A2(n8660), .ZN(n4629) );
  NAND2_X1 U5451 ( .A1(n8666), .A2(n8659), .ZN(n4628) );
  NAND2_X1 U5452 ( .A1(n6319), .A2(n6254), .ZN(n8314) );
  AOI21_X1 U5453 ( .B1(n4828), .B2(n4830), .A(n4329), .ZN(n4826) );
  NAND2_X1 U5454 ( .A1(n6190), .A2(n9993), .ZN(n6201) );
  NAND2_X1 U5455 ( .A1(n4740), .A2(n4738), .ZN(n8783) );
  AOI21_X1 U5456 ( .B1(n4298), .B2(n4741), .A(n4739), .ZN(n4738) );
  INV_X1 U5457 ( .A(n8420), .ZN(n4739) );
  NAND2_X1 U5458 ( .A1(n5842), .A2(n5841), .ZN(n6127) );
  INV_X1 U5459 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5841) );
  INV_X1 U5460 ( .A(n6118), .ZN(n5842) );
  NAND2_X1 U5461 ( .A1(n5840), .A2(n5839), .ZN(n6116) );
  INV_X1 U5462 ( .A(n6102), .ZN(n5840) );
  NAND2_X1 U5463 ( .A1(n5838), .A2(n5837), .ZN(n6090) );
  INV_X1 U5464 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5837) );
  INV_X1 U5465 ( .A(n6079), .ZN(n5838) );
  OR2_X1 U5466 ( .A1(n6063), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U5467 ( .A1(n5834), .A2(n7400), .ZN(n6051) );
  INV_X1 U5468 ( .A(n6038), .ZN(n5834) );
  NAND2_X1 U5469 ( .A1(n5836), .A2(n5835), .ZN(n6063) );
  INV_X1 U5470 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5835) );
  INV_X1 U5471 ( .A(n6051), .ZN(n5836) );
  INV_X1 U5472 ( .A(n5999), .ZN(n5833) );
  OR2_X1 U5473 ( .A1(n6015), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U5474 ( .A1(n5831), .A2(n5830), .ZN(n5988) );
  INV_X1 U5475 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5830) );
  INV_X1 U5476 ( .A(n5972), .ZN(n5831) );
  OR2_X1 U5477 ( .A1(n5988), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5999) );
  AND2_X1 U5478 ( .A1(n5980), .A2(n5979), .ZN(n6937) );
  NAND2_X1 U5479 ( .A1(n4749), .A2(n4747), .ZN(n6892) );
  AOI21_X1 U5480 ( .B1(n8341), .B2(n8345), .A(n4748), .ZN(n4747) );
  INV_X1 U5481 ( .A(n8348), .ZN(n4748) );
  INV_X1 U5482 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5828) );
  OR2_X1 U5483 ( .A1(n6159), .A2(n6852), .ZN(n5915) );
  AND3_X1 U5484 ( .A1(n5909), .A2(n5908), .A3(n5907), .ZN(n6796) );
  NAND2_X1 U5485 ( .A1(n8330), .A2(n8331), .ZN(n6793) );
  NAND2_X1 U5486 ( .A1(n8877), .A2(n6232), .ZN(n6791) );
  NAND2_X1 U5487 ( .A1(n5898), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U5488 ( .A1(n8879), .A2(n8878), .ZN(n8877) );
  AND2_X1 U5489 ( .A1(n8688), .A2(n8687), .ZN(n8962) );
  NAND2_X1 U5490 ( .A1(n5825), .A2(n5824), .ZN(n8123) );
  AND2_X1 U5491 ( .A1(n8854), .A2(n6086), .ZN(n7695) );
  AND2_X1 U5492 ( .A1(n8385), .A2(n8384), .ZN(n8382) );
  AOI21_X1 U5493 ( .B1(n4400), .B2(n4403), .A(n8370), .ZN(n4399) );
  INV_X1 U5494 ( .A(n8364), .ZN(n4403) );
  OR2_X1 U5495 ( .A1(n6305), .A2(n8508), .ZN(n9930) );
  AND2_X1 U5496 ( .A1(n6500), .A2(n6499), .ZN(n6481) );
  XNOR2_X1 U5497 ( .A(n6303), .B(n10073), .ZN(n6490) );
  INV_X1 U5498 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U5499 ( .A(n6284), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6286) );
  XNOR2_X1 U5500 ( .A(n6223), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6547) );
  INV_X1 U5501 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U5502 ( .A(n6073), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8558) );
  AND2_X1 U5503 ( .A1(n6025), .A2(n6047), .ZN(n7387) );
  NOR2_X1 U5504 ( .A1(n5963), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5966) );
  INV_X1 U5505 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5812) );
  AND2_X1 U5506 ( .A1(n5878), .A2(n5906), .ZN(n5918) );
  NAND2_X1 U5507 ( .A1(n4640), .A2(n4639), .ZN(n4646) );
  NOR2_X1 U5508 ( .A1(n5906), .A2(n5849), .ZN(n4640) );
  AND2_X1 U5509 ( .A1(n5849), .A2(n5906), .ZN(n4648) );
  AND2_X1 U5510 ( .A1(n5879), .A2(n5906), .ZN(n4649) );
  NAND2_X1 U5511 ( .A1(n4883), .A2(n4882), .ZN(n5648) );
  OR2_X1 U5512 ( .A1(n5290), .A2(n5289), .ZN(n4777) );
  NAND2_X1 U5513 ( .A1(n5290), .A2(n5289), .ZN(n5294) );
  INV_X1 U5514 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U5515 ( .A1(n4761), .A2(n5321), .ZN(n9086) );
  OR2_X1 U5516 ( .A1(n5304), .A2(n5303), .ZN(n5332) );
  NOR2_X1 U5517 ( .A1(n5358), .A2(n5357), .ZN(n5405) );
  OR2_X1 U5518 ( .A1(n5406), .A2(n5388), .ZN(n5430) );
  NAND2_X1 U5519 ( .A1(n5251), .A2(n5250), .ZN(n7811) );
  AND2_X1 U5520 ( .A1(n5252), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5280) );
  NOR2_X1 U5521 ( .A1(n9129), .A2(n9128), .ZN(n9127) );
  NOR2_X1 U5522 ( .A1(n10115), .A2(n5471), .ZN(n5494) );
  INV_X1 U5523 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5181) );
  OR2_X1 U5524 ( .A1(n5199), .A2(n5181), .ZN(n5224) );
  NAND2_X1 U5525 ( .A1(n5108), .A2(n4758), .ZN(n4755) );
  INV_X1 U5526 ( .A(n5753), .ZN(n8051) );
  NAND2_X1 U5527 ( .A1(n5373), .A2(n9094), .ZN(n9058) );
  AND2_X1 U5528 ( .A1(n7896), .A2(n9326), .ZN(n7901) );
  NAND2_X1 U5529 ( .A1(n4441), .A2(n4439), .ZN(n4438) );
  INV_X1 U5530 ( .A(n4442), .ZN(n4439) );
  AND2_X1 U5531 ( .A1(n8048), .A2(n4437), .ZN(n4436) );
  NAND2_X1 U5532 ( .A1(n4445), .A2(n4446), .ZN(n4437) );
  INV_X1 U5533 ( .A(n8054), .ZN(n4434) );
  AND3_X1 U5534 ( .A1(n6590), .A2(n6589), .A3(n6588), .ZN(n8030) );
  INV_X1 U5535 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4869) );
  OAI21_X1 U5536 ( .B1(n8024), .B2(n4280), .A(n4555), .ZN(n4554) );
  NAND2_X1 U5537 ( .A1(n8024), .A2(n4557), .ZN(n4555) );
  NAND2_X1 U5538 ( .A1(n5778), .A2(n4557), .ZN(n4556) );
  AND2_X1 U5539 ( .A1(n5665), .A2(n5619), .ZN(n8056) );
  AND3_X1 U5540 ( .A1(n4371), .A2(n4370), .A3(n4373), .ZN(n8059) );
  AOI21_X1 U5541 ( .B1(n4374), .B2(n9504), .A(n5747), .ZN(n4373) );
  NAND2_X1 U5542 ( .A1(n9374), .A2(n9387), .ZN(n9355) );
  AND4_X1 U5543 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n9367)
         );
  NOR2_X1 U5544 ( .A1(n9459), .A2(n9441), .ZN(n9440) );
  NAND2_X1 U5545 ( .A1(n9440), .A2(n9419), .ZN(n9414) );
  NAND2_X1 U5546 ( .A1(n5740), .A2(n7909), .ZN(n9471) );
  OAI21_X1 U5547 ( .B1(n5737), .B2(n4389), .A(n4387), .ZN(n9487) );
  AND2_X1 U5548 ( .A1(n4388), .A2(n7844), .ZN(n4387) );
  OR2_X1 U5549 ( .A1(n4392), .A2(n4389), .ZN(n4388) );
  NAND2_X1 U5550 ( .A1(n4390), .A2(n7940), .ZN(n4389) );
  NAND2_X1 U5551 ( .A1(n7599), .A2(n4546), .ZN(n9510) );
  NAND2_X1 U5552 ( .A1(n7599), .A2(n9632), .ZN(n7715) );
  AOI21_X1 U5553 ( .B1(n8015), .B2(n4599), .A(n5700), .ZN(n4598) );
  NAND2_X1 U5554 ( .A1(n8015), .A2(n4604), .ZN(n4600) );
  INV_X1 U5555 ( .A(n5736), .ZN(n4569) );
  AOI21_X1 U5556 ( .B1(n5736), .B2(n4568), .A(n7828), .ZN(n4567) );
  NAND2_X1 U5557 ( .A1(n7532), .A2(n5733), .ZN(n7618) );
  AND2_X1 U5558 ( .A1(n4528), .A2(n4527), .ZN(n7623) );
  NOR2_X1 U5559 ( .A1(n4529), .A2(n7624), .ZN(n4528) );
  NAND2_X1 U5560 ( .A1(n7295), .A2(n7802), .ZN(n7441) );
  NAND2_X1 U5561 ( .A1(n7313), .A2(n5730), .ZN(n7295) );
  NOR2_X1 U5562 ( .A1(n4534), .A2(n7527), .ZN(n7315) );
  OR2_X1 U5563 ( .A1(n7924), .A2(n5728), .ZN(n4386) );
  NAND2_X1 U5564 ( .A1(n4384), .A2(n4386), .ZN(n7313) );
  NAND2_X1 U5565 ( .A1(n4582), .A2(n4581), .ZN(n7224) );
  AOI21_X1 U5566 ( .B1(n4583), .B2(n4584), .A(n4321), .ZN(n4581) );
  NAND2_X1 U5567 ( .A1(n7200), .A2(n4533), .ZN(n7225) );
  AND2_X1 U5568 ( .A1(n5041), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U5569 ( .A1(n7200), .A2(n7373), .ZN(n7185) );
  AND2_X1 U5570 ( .A1(n7775), .A2(n7780), .ZN(n7776) );
  NAND2_X1 U5571 ( .A1(n4451), .A2(n4576), .ZN(n6906) );
  OAI21_X1 U5572 ( .B1(n4577), .B2(n5724), .A(n7914), .ZN(n4576) );
  INV_X1 U5573 ( .A(n5723), .ZN(n4577) );
  OR2_X1 U5574 ( .A1(n6879), .A2(n6899), .ZN(n6905) );
  NAND2_X1 U5575 ( .A1(n6828), .A2(n5685), .ZN(n6877) );
  NAND2_X1 U5576 ( .A1(n6837), .A2(n5684), .ZN(n4579) );
  XNOR2_X1 U5577 ( .A(n9192), .B(n7910), .ZN(n7991) );
  NOR2_X1 U5578 ( .A1(n6843), .A2(n7008), .ZN(n6839) );
  NAND2_X1 U5579 ( .A1(n5656), .A2(n5753), .ZN(n7103) );
  AND2_X1 U5580 ( .A1(n5647), .A2(n9634), .ZN(n5761) );
  AND2_X1 U5581 ( .A1(n8059), .A2(n8055), .ZN(n5750) );
  NAND2_X1 U5582 ( .A1(n5595), .A2(n5594), .ZN(n9531) );
  AOI211_X1 U5583 ( .C1(n5741), .C2(n9477), .A(n9509), .B(n9476), .ZN(n9566)
         );
  INV_X1 U5584 ( .A(n9831), .ZN(n9837) );
  INV_X1 U5585 ( .A(n9835), .ZN(n9583) );
  NAND3_X1 U5586 ( .A1(n4916), .A2(n4915), .A3(n4914), .ZN(n5682) );
  OR2_X1 U5587 ( .A1(n6568), .A2(n6617), .ZN(n4916) );
  NAND2_X1 U5588 ( .A1(n4984), .A2(n6365), .ZN(n4914) );
  INV_X1 U5589 ( .A(n5761), .ZN(n7005) );
  AND2_X1 U5590 ( .A1(n7004), .A2(n5758), .ZN(n5762) );
  INV_X1 U5591 ( .A(n9642), .ZN(n4463) );
  AND3_X1 U5592 ( .A1(n4934), .A2(P1_STATE_REG_SCAN_IN), .A3(n6567), .ZN(n5753) );
  XNOR2_X1 U5593 ( .A(n7765), .B(n7764), .ZN(n9036) );
  NAND2_X1 U5594 ( .A1(n7888), .A2(n7887), .ZN(n9041) );
  XNOR2_X1 U5595 ( .A(n7748), .B(SI_29_), .ZN(n8081) );
  XNOR2_X1 U5596 ( .A(n5768), .B(n5767), .ZN(n8078) );
  XNOR2_X1 U5597 ( .A(n4876), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U5598 ( .A1(n4776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4872) );
  AND2_X1 U5599 ( .A1(n4775), .A2(n4338), .ZN(n4774) );
  OAI21_X1 U5600 ( .B1(n4704), .B2(n4703), .A(n4705), .ZN(n5490) );
  AOI21_X1 U5601 ( .B1(n4707), .B2(n4708), .A(n4706), .ZN(n4705) );
  NAND2_X1 U5602 ( .A1(n4708), .A2(n4715), .ZN(n4703) );
  OR2_X1 U5603 ( .A1(n5193), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5220) );
  CLKBUF_X1 U5604 ( .A(n5087), .Z(n5088) );
  NAND2_X1 U5605 ( .A1(n5052), .A2(n5051), .ZN(n5071) );
  NAND2_X1 U5606 ( .A1(n4475), .A2(n4961), .ZN(n4986) );
  NAND2_X1 U5607 ( .A1(n4394), .A2(n4958), .ZN(n4475) );
  INV_X1 U5608 ( .A(n4959), .ZN(n4394) );
  CLKBUF_X1 U5609 ( .A(n4904), .Z(n4954) );
  AND2_X1 U5610 ( .A1(n6933), .A2(n6932), .ZN(n6935) );
  NAND2_X1 U5611 ( .A1(n8270), .A2(n4312), .ZN(n8145) );
  NAND2_X1 U5612 ( .A1(n8270), .A2(n8130), .ZN(n8144) );
  AND2_X1 U5613 ( .A1(n6150), .A2(n6149), .ZN(n8925) );
  INV_X1 U5614 ( .A(n9877), .ZN(n5926) );
  XNOR2_X1 U5615 ( .A(n6552), .B(n5884), .ZN(n6580) );
  CLKBUF_X1 U5616 ( .A(n8153), .Z(n8240) );
  OR2_X1 U5617 ( .A1(n6543), .A2(n6542), .ZN(n8257) );
  NAND2_X1 U5618 ( .A1(n6143), .A2(n6142), .ZN(n8921) );
  NAND2_X1 U5619 ( .A1(n6502), .A2(n6501), .ZN(n8267) );
  NAND2_X1 U5620 ( .A1(n5969), .A2(n4430), .ZN(n9897) );
  AND2_X1 U5621 ( .A1(n5968), .A2(n4333), .ZN(n4430) );
  NAND2_X1 U5622 ( .A1(n6488), .A2(n8882), .ZN(n8259) );
  NAND2_X1 U5623 ( .A1(n4784), .A2(n6915), .ZN(n6919) );
  INV_X1 U5624 ( .A(n8286), .ZN(n8277) );
  INV_X1 U5625 ( .A(n8280), .ZN(n8272) );
  NOR2_X1 U5626 ( .A1(n8281), .A2(n4780), .ZN(n4779) );
  INV_X1 U5627 ( .A(n8094), .ZN(n4780) );
  NAND2_X1 U5628 ( .A1(n8152), .A2(n8094), .ZN(n8282) );
  INV_X1 U5629 ( .A(n8925), .ZN(n8787) );
  NAND2_X1 U5630 ( .A1(n4652), .A2(n6439), .ZN(n6456) );
  INV_X1 U5631 ( .A(n8683), .ZN(n8617) );
  INV_X1 U5632 ( .A(n4668), .ZN(n6696) );
  XNOR2_X1 U5633 ( .A(n4666), .B(n6990), .ZN(n6858) );
  NOR2_X1 U5634 ( .A1(n6858), .A2(n7036), .ZN(n6975) );
  NOR2_X1 U5635 ( .A1(n7631), .A2(n7632), .ZN(n7634) );
  NOR2_X1 U5636 ( .A1(n8555), .A2(n8563), .ZN(n8578) );
  NAND2_X1 U5637 ( .A1(n4655), .A2(n4656), .ZN(n8606) );
  NAND2_X1 U5638 ( .A1(n4635), .A2(n4638), .ZN(n4634) );
  OR2_X1 U5639 ( .A1(n6491), .A2(n6347), .ZN(n8641) );
  OAI211_X1 U5640 ( .C1(n4635), .C2(n4630), .A(n4627), .B(n4626), .ZN(n4632)
         );
  OR2_X1 U5641 ( .A1(n8666), .A2(n8660), .ZN(n4630) );
  XNOR2_X1 U5642 ( .A(n8314), .B(n8453), .ZN(n8701) );
  NOR2_X1 U5643 ( .A1(n6322), .A2(n6321), .ZN(n8709) );
  AND2_X1 U5644 ( .A1(n6320), .A2(n8469), .ZN(n6321) );
  NAND2_X1 U5645 ( .A1(n8718), .A2(n4849), .ZN(n6318) );
  NAND2_X1 U5646 ( .A1(n4418), .A2(n4419), .ZN(n8724) );
  NAND2_X1 U5647 ( .A1(n6179), .A2(n6178), .ZN(n8732) );
  OAI21_X1 U5648 ( .B1(n6247), .B2(n4298), .A(n4741), .ZN(n8795) );
  NAND2_X1 U5649 ( .A1(n4835), .A2(n4833), .ZN(n8796) );
  NAND2_X1 U5650 ( .A1(n6126), .A2(n6125), .ZN(n8931) );
  AND4_X1 U5651 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n8831)
         );
  OR2_X1 U5652 ( .A1(n6306), .A2(n9886), .ZN(n8752) );
  NAND2_X1 U5653 ( .A1(n7138), .A2(n8364), .ZN(n7236) );
  NAND2_X1 U5654 ( .A1(n4822), .A2(n4821), .ZN(n7238) );
  NAND2_X1 U5655 ( .A1(n4496), .A2(n6013), .ZN(n9934) );
  NAND2_X1 U5656 ( .A1(n6409), .A2(n8298), .ZN(n4496) );
  NAND2_X1 U5657 ( .A1(n6966), .A2(n5994), .ZN(n7040) );
  NAND2_X1 U5658 ( .A1(n6806), .A2(n5956), .ZN(n6887) );
  NAND2_X1 U5659 ( .A1(n6499), .A2(n6487), .ZN(n8882) );
  OR2_X1 U5660 ( .A1(n6745), .A2(n8341), .ZN(n6804) );
  CLKBUF_X1 U5661 ( .A(n5893), .Z(n9863) );
  OR2_X1 U5662 ( .A1(n5897), .A2(n5885), .ZN(n5891) );
  CLKBUF_X1 U5663 ( .A(n5884), .Z(n6739) );
  INV_X1 U5664 ( .A(n8882), .ZN(n8848) );
  INV_X1 U5665 ( .A(n8691), .ZN(n8961) );
  NAND2_X1 U5666 ( .A1(n6189), .A2(n6188), .ZN(n8968) );
  INV_X1 U5667 ( .A(n8732), .ZN(n8975) );
  NAND2_X1 U5668 ( .A1(n6168), .A2(n6167), .ZN(n8978) );
  NAND2_X1 U5669 ( .A1(n4798), .A2(n4805), .ZN(n8736) );
  OR2_X1 U5670 ( .A1(n8758), .A2(n4808), .ZN(n4798) );
  NAND2_X1 U5671 ( .A1(n4424), .A2(n4425), .ZN(n8735) );
  NAND2_X1 U5672 ( .A1(n8756), .A2(n4427), .ZN(n4424) );
  INV_X1 U5673 ( .A(n8123), .ZN(n8983) );
  NAND2_X1 U5674 ( .A1(n4811), .A2(n4813), .ZN(n8748) );
  NAND2_X1 U5675 ( .A1(n4429), .A2(n8471), .ZN(n8746) );
  OR2_X1 U5676 ( .A1(n8756), .A2(n8321), .ZN(n4429) );
  NAND2_X1 U5677 ( .A1(n6153), .A2(n6152), .ZN(n8989) );
  NAND2_X1 U5678 ( .A1(n5867), .A2(n5866), .ZN(n9007) );
  NAND2_X1 U5679 ( .A1(n8822), .A2(n8414), .ZN(n8806) );
  NAND2_X1 U5680 ( .A1(n6101), .A2(n6100), .ZN(n9018) );
  NAND2_X1 U5681 ( .A1(n4745), .A2(n8404), .ZN(n8837) );
  NAND2_X1 U5682 ( .A1(n6078), .A2(n6077), .ZN(n9023) );
  NAND2_X1 U5683 ( .A1(n4407), .A2(n8396), .ZN(n8851) );
  NAND2_X1 U5684 ( .A1(n6244), .A2(n4411), .ZN(n4407) );
  NAND2_X1 U5685 ( .A1(n6244), .A2(n6243), .ZN(n7507) );
  NAND2_X1 U5686 ( .A1(n6050), .A2(n6049), .ZN(n8870) );
  NAND2_X1 U5687 ( .A1(n6037), .A2(n6036), .ZN(n7494) );
  AND2_X1 U5688 ( .A1(n6491), .A2(n6381), .ZN(n6499) );
  INV_X1 U5689 ( .A(n6286), .ZN(n7738) );
  XNOR2_X1 U5690 ( .A(n6281), .B(n6280), .ZN(n7733) );
  INV_X1 U5691 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7658) );
  INV_X1 U5692 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10005) );
  INV_X1 U5693 ( .A(n6547), .ZN(n8323) );
  INV_X1 U5694 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7430) );
  NAND2_X1 U5695 ( .A1(n6229), .A2(n6228), .ZN(n8462) );
  INV_X1 U5696 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7264) );
  INV_X1 U5697 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7045) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6947) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6761) );
  INV_X1 U5700 ( .A(n8558), .ZN(n8554) );
  INV_X1 U5701 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10132) );
  INV_X1 U5702 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6506) );
  INV_X1 U5703 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6413) );
  OR2_X1 U5704 ( .A1(n6012), .A2(n6011), .ZN(n7149) );
  INV_X1 U5705 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U5706 ( .A1(n5880), .A2(n4639), .ZN(n6438) );
  INV_X1 U5707 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5708 ( .B1(n4765), .B2(n5792), .A(n5791), .ZN(n4764) );
  INV_X1 U5709 ( .A(n5653), .ZN(n5795) );
  AND4_X1 U5710 ( .A1(n5135), .A2(n5134), .A3(n5133), .A4(n5132), .ZN(n7585)
         );
  AND2_X1 U5711 ( .A1(n5664), .A2(n7984), .ZN(n9066) );
  AOI21_X1 U5712 ( .B1(n4276), .B2(n4515), .A(n4330), .ZN(n4514) );
  AND4_X1 U5713 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n7610)
         );
  NOR2_X1 U5714 ( .A1(n9110), .A2(n5534), .ZN(n9079) );
  NOR2_X1 U5715 ( .A1(n9079), .A2(n9078), .ZN(n9149) );
  NAND2_X1 U5716 ( .A1(n4507), .A2(n5061), .ZN(n7128) );
  NAND2_X1 U5717 ( .A1(n7094), .A2(n5039), .ZN(n4507) );
  INV_X1 U5718 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10115) );
  AND4_X1 U5719 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n9663)
         );
  AND4_X1 U5720 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9660)
         );
  XNOR2_X1 U5721 ( .A(n4973), .B(n4974), .ZN(n6822) );
  NOR2_X1 U5722 ( .A1(n5061), .A2(n7130), .ZN(n4511) );
  AND4_X1 U5723 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n9366)
         );
  AND2_X1 U5724 ( .A1(n5664), .A2(n5652), .ZN(n9151) );
  AND2_X1 U5725 ( .A1(n5618), .A2(n5573), .ZN(n9375) );
  INV_X1 U5726 ( .A(n9678), .ZN(n9161) );
  INV_X1 U5727 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U5728 ( .A1(n5302), .A2(n5301), .ZN(n9167) );
  AND4_X1 U5729 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n6846)
         );
  INV_X1 U5730 ( .A(n9388), .ZN(n9428) );
  INV_X1 U5731 ( .A(n7610), .ZN(n9183) );
  NAND4_X1 U5732 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n7009)
         );
  INV_X1 U5733 ( .A(n9758), .ZN(n9784) );
  INV_X1 U5734 ( .A(n9764), .ZN(n9788) );
  NOR2_X1 U5735 ( .A1(n9326), .A2(n4549), .ZN(n4548) );
  NOR2_X1 U5736 ( .A1(n9334), .A2(n9509), .ZN(n9527) );
  XNOR2_X1 U5737 ( .A(n5775), .B(n8024), .ZN(n9339) );
  NAND2_X1 U5738 ( .A1(n4379), .A2(n4562), .ZN(n9384) );
  NAND2_X1 U5739 ( .A1(n4587), .A2(n4590), .ZN(n9397) );
  NAND2_X1 U5740 ( .A1(n9434), .A2(n4295), .ZN(n4587) );
  NAND2_X1 U5741 ( .A1(n9423), .A2(n5745), .ZN(n9398) );
  AND2_X1 U5742 ( .A1(n4593), .A2(n4596), .ZN(n9413) );
  NAND2_X1 U5743 ( .A1(n9434), .A2(n5709), .ZN(n4593) );
  CLKBUF_X1 U5744 ( .A(n9448), .Z(n9450) );
  NAND2_X1 U5745 ( .A1(n7711), .A2(n7940), .ZN(n9503) );
  NOR2_X1 U5746 ( .A1(n4391), .A2(n7941), .ZN(n4859) );
  OAI21_X1 U5747 ( .B1(n7615), .B2(n4603), .A(n4601), .ZN(n7660) );
  NAND2_X1 U5748 ( .A1(n7615), .A2(n5699), .ZN(n4605) );
  NAND2_X1 U5749 ( .A1(n5180), .A2(n5179), .ZN(n9838) );
  NAND2_X1 U5750 ( .A1(n7310), .A2(n7312), .ZN(n7309) );
  NAND2_X1 U5751 ( .A1(n7280), .A2(n5692), .ZN(n7310) );
  OAI21_X1 U5752 ( .B1(n7018), .B2(n4584), .A(n4583), .ZN(n7176) );
  NAND2_X1 U5753 ( .A1(n7017), .A2(n5690), .ZN(n7174) );
  NAND2_X1 U5754 ( .A1(n4578), .A2(n5723), .ZN(n6880) );
  INV_X1 U5755 ( .A(n9518), .ZN(n9494) );
  INV_X1 U5756 ( .A(n9806), .ZN(n9512) );
  OAI21_X1 U5757 ( .B1(n9813), .B2(n7622), .A(n7629), .ZN(n9809) );
  OR2_X1 U5758 ( .A1(n5750), .A2(n5802), .ZN(n4613) );
  NAND2_X1 U5759 ( .A1(n5031), .A2(n4855), .ZN(n6909) );
  CLKBUF_X1 U5760 ( .A(n5682), .Z(n6843) );
  AND2_X1 U5761 ( .A1(n9854), .A2(n9837), .ZN(n7450) );
  INV_X1 U5762 ( .A(n9330), .ZN(n9595) );
  AND2_X1 U5763 ( .A1(n9522), .A2(n9525), .ZN(n9592) );
  INV_X1 U5764 ( .A(n5748), .ZN(n8058) );
  OR2_X1 U5765 ( .A1(n5750), .A2(n9846), .ZN(n4615) );
  OAI21_X1 U5766 ( .B1(n9372), .B2(n4619), .A(n4616), .ZN(n5715) );
  INV_X1 U5767 ( .A(n4617), .ZN(n4616) );
  OAI21_X1 U5768 ( .B1(n4619), .B2(n4621), .A(n8023), .ZN(n4617) );
  INV_X1 U5769 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4614) );
  INV_X1 U5770 ( .A(n9374), .ZN(n9603) );
  AND2_X1 U5771 ( .A1(n5517), .A2(n5516), .ZN(n9608) );
  AND2_X1 U5772 ( .A1(n5470), .A2(n5469), .ZN(n9613) );
  INV_X1 U5773 ( .A(n5741), .ZN(n9618) );
  INV_X1 U5774 ( .A(n9167), .ZN(n7690) );
  AND2_X1 U5775 ( .A1(n9627), .A2(n9837), .ZN(n7448) );
  AND2_X1 U5776 ( .A1(n5145), .A2(n5144), .ZN(n7476) );
  INV_X1 U5777 ( .A(n6909), .ZN(n7329) );
  INV_X1 U5778 ( .A(n7448), .ZN(n9631) );
  NAND2_X1 U5779 ( .A1(n5751), .A2(n5753), .ZN(n9815) );
  NAND2_X1 U5780 ( .A1(n4924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U5781 ( .A1(n4923), .A2(n4924), .ZN(n8085) );
  NOR2_X1 U5782 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  NOR2_X1 U5783 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4537) );
  INV_X1 U5784 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U5785 ( .A1(n4901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4535) );
  INV_X1 U5786 ( .A(n5645), .ZN(n7731) );
  XNOR2_X1 U5787 ( .A(n4879), .B(n4878), .ZN(n7692) );
  INV_X1 U5788 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4878) );
  INV_X1 U5789 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7565) );
  INV_X1 U5790 ( .A(n5651), .ZN(n7564) );
  INV_X1 U5791 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7421) );
  INV_X1 U5792 ( .A(n7989), .ZN(n7993) );
  AOI21_X1 U5793 ( .B1(n5401), .B2(n4888), .A(n4875), .ZN(n4512) );
  INV_X1 U5794 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10018) );
  INV_X1 U5795 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7047) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10114) );
  INV_X1 U5797 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10071) );
  XNOR2_X1 U5798 ( .A(n4362), .B(n4274), .ZN(n8512) );
  INV_X1 U5799 ( .A(n4624), .ZN(n7388) );
  INV_X1 U5800 ( .A(n6343), .ZN(n6344) );
  OAI22_X1 U5801 ( .A1(n8695), .A2(n8957), .B1(n9956), .B2(n6342), .ZN(n6343)
         );
  OAI21_X1 U5802 ( .B1(n6338), .B2(n4414), .A(n4347), .ZN(P2_U3487) );
  NAND2_X1 U5803 ( .A1(n4414), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4413) );
  AOI211_X1 U5804 ( .C1(n5741), .C2(n9675), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI211_X1 U5805 ( .C1(n8028), .C2(n4285), .A(n4433), .B(n4431), .ZN(P1_U3242) );
  OAI21_X1 U5806 ( .B1(n7988), .B2(n4446), .A(n7987), .ZN(n8028) );
  NOR2_X1 U5807 ( .A1(n4842), .A2(n5805), .ZN(n5806) );
  NAND2_X1 U5808 ( .A1(n4571), .A2(n9854), .ZN(n4570) );
  NOR2_X1 U5809 ( .A1(n4853), .A2(n5789), .ZN(n5790) );
  NOR2_X1 U5810 ( .A1(n9627), .A2(n5788), .ZN(n5789) );
  AND2_X2 U5811 ( .A1(n4934), .A2(n4933), .ZN(n5262) );
  INV_X1 U5812 ( .A(n8666), .ZN(n4633) );
  NAND2_X1 U5813 ( .A1(n5774), .A2(n5773), .ZN(n5776) );
  AND2_X1 U5814 ( .A1(n4518), .A2(n4314), .ZN(n4276) );
  OR3_X1 U5815 ( .A1(n8042), .A2(n8026), .A3(n8025), .ZN(n8044) );
  AOI21_X1 U5816 ( .B1(n5745), .B2(n4564), .A(n4563), .ZN(n4562) );
  NAND2_X1 U5817 ( .A1(n8301), .A2(n8300), .ZN(n8895) );
  INV_X1 U5818 ( .A(n7312), .ZN(n4612) );
  AND2_X1 U5819 ( .A1(n4674), .A2(n4300), .ZN(n4277) );
  INV_X1 U5820 ( .A(n8023), .ZN(n4377) );
  INV_X1 U5821 ( .A(n8471), .ZN(n4428) );
  INV_X1 U5822 ( .A(n7876), .ZN(n4561) );
  NAND2_X1 U5823 ( .A1(n5404), .A2(n5403), .ZN(n9511) );
  INV_X1 U5824 ( .A(n9511), .ZN(n4545) );
  AND4_X1 U5825 ( .A1(n5649), .A2(n4874), .A3(n4886), .A4(n4889), .ZN(n4278)
         );
  OR2_X1 U5826 ( .A1(n8609), .A2(n4358), .ZN(n4279) );
  NAND2_X1 U5827 ( .A1(n4790), .A2(n4345), .ZN(n8166) );
  AND2_X1 U5828 ( .A1(n7973), .A2(n7876), .ZN(n9354) );
  INV_X1 U5829 ( .A(n9354), .ZN(n4623) );
  AND2_X1 U5830 ( .A1(n4557), .A2(n4560), .ZN(n4280) );
  INV_X1 U5831 ( .A(n4591), .ZN(n4590) );
  NOR2_X1 U5832 ( .A1(n4592), .A2(n5710), .ZN(n4591) );
  AND2_X1 U5833 ( .A1(n9939), .A2(n8521), .ZN(n4281) );
  NOR2_X1 U5834 ( .A1(n9078), .A2(n5533), .ZN(n4282) );
  NOR2_X1 U5835 ( .A1(n9922), .A2(n8523), .ZN(n4283) );
  AND2_X1 U5836 ( .A1(n4377), .A2(n7876), .ZN(n4284) );
  INV_X1 U5837 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4837) );
  INV_X2 U5838 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4894) );
  OR2_X1 U5839 ( .A1(n4440), .A2(n8054), .ZN(n4285) );
  AND2_X1 U5840 ( .A1(n8023), .A2(n9354), .ZN(n4286) );
  AND2_X1 U5841 ( .A1(n6085), .A2(n6071), .ZN(n4287) );
  INV_X1 U5842 ( .A(n6697), .ZN(n4667) );
  AND2_X1 U5843 ( .A1(n6200), .A2(n6199), .ZN(n8455) );
  INV_X1 U5844 ( .A(n8455), .ZN(n6336) );
  OR2_X1 U5845 ( .A1(n8105), .A2(n8517), .ZN(n4288) );
  AND2_X1 U5846 ( .A1(n4605), .A2(n4606), .ZN(n7593) );
  AND2_X1 U5847 ( .A1(n4760), .A2(n5321), .ZN(n4289) );
  AND2_X1 U5848 ( .A1(n7508), .A2(n6071), .ZN(n8852) );
  NAND2_X1 U5849 ( .A1(n4777), .A2(n5294), .ZN(n7739) );
  NOR3_X1 U5850 ( .A1(n7316), .A2(n9838), .A3(n7454), .ZN(n4290) );
  OR2_X1 U5851 ( .A1(n9627), .A2(n4614), .ZN(n4291) );
  OR2_X1 U5852 ( .A1(n9854), .A2(n10010), .ZN(n4292) );
  INV_X1 U5853 ( .A(n8630), .ZN(n4638) );
  INV_X1 U5854 ( .A(n5010), .ZN(n5783) );
  AND2_X2 U5855 ( .A1(n6568), .A2(n8295), .ZN(n4992) );
  NAND3_X1 U5856 ( .A1(n6222), .A2(n5820), .A3(n4752), .ZN(n4293) );
  AND2_X1 U5857 ( .A1(n7940), .A2(n7835), .ZN(n4294) );
  AND3_X1 U5858 ( .A1(n4997), .A2(n4996), .A3(n4995), .ZN(n5686) );
  XNOR2_X1 U5859 ( .A(n9441), .B(n9426), .ZN(n9436) );
  INV_X1 U5860 ( .A(n9436), .ZN(n4457) );
  AND2_X1 U5861 ( .A1(n4595), .A2(n5709), .ZN(n4295) );
  AND3_X1 U5862 ( .A1(n5890), .A2(n5889), .A3(n5888), .ZN(n4296) );
  NAND2_X1 U5863 ( .A1(n6133), .A2(n6132), .ZN(n8792) );
  NAND2_X1 U5864 ( .A1(n5356), .A2(n5355), .ZN(n9581) );
  NAND2_X1 U5865 ( .A1(n5330), .A2(n5329), .ZN(n7669) );
  AND2_X1 U5866 ( .A1(n5059), .A2(n5039), .ZN(n4297) );
  OR2_X1 U5867 ( .A1(n6248), .A2(n4742), .ZN(n4298) );
  AND2_X1 U5868 ( .A1(n5915), .A2(n4854), .ZN(n4299) );
  OR3_X1 U5869 ( .A1(n5879), .A2(P2_IR_REG_0__SCAN_IN), .A3(n5886), .ZN(n4300)
         );
  OR2_X1 U5870 ( .A1(n9934), .A2(n8522), .ZN(n4301) );
  NAND2_X1 U5871 ( .A1(n4731), .A2(n4730), .ZN(n5350) );
  AND2_X1 U5872 ( .A1(n4869), .A2(n4772), .ZN(n4302) );
  NAND2_X1 U5873 ( .A1(n8355), .A2(n8356), .ZN(n8366) );
  INV_X1 U5874 ( .A(n8366), .ZN(n4487) );
  NAND2_X1 U5875 ( .A1(n4922), .A2(n4921), .ZN(n4924) );
  AND4_X1 U5876 ( .A1(n4873), .A2(n4882), .A3(n4894), .A4(n4888), .ZN(n4303)
         );
  OR2_X1 U5877 ( .A1(n8609), .A2(n4631), .ZN(n4304) );
  AND2_X1 U5878 ( .A1(n7919), .A2(n7781), .ZN(n4305) );
  NAND2_X1 U5879 ( .A1(n7892), .A2(n7891), .ZN(n9326) );
  AND2_X1 U5880 ( .A1(n7779), .A2(n7905), .ZN(n4306) );
  INV_X1 U5881 ( .A(n9502), .ZN(n4390) );
  INV_X1 U5882 ( .A(n5879), .ZN(n4639) );
  OR2_X1 U5883 ( .A1(n8098), .A2(n8841), .ZN(n8404) );
  INV_X1 U5884 ( .A(n8404), .ZN(n4744) );
  AND3_X1 U5885 ( .A1(n8399), .A2(n8853), .A3(n8398), .ZN(n4307) );
  AND2_X1 U5886 ( .A1(n8491), .A2(n6086), .ZN(n4308) );
  AND2_X1 U5887 ( .A1(n8125), .A2(n8901), .ZN(n4309) );
  NOR2_X1 U5888 ( .A1(n5141), .A2(n4684), .ZN(n4683) );
  NOR2_X1 U5889 ( .A1(n8578), .A2(n8579), .ZN(n4310) );
  AND2_X1 U5890 ( .A1(n9550), .A2(n9173), .ZN(n4311) );
  INV_X1 U5891 ( .A(n4541), .ZN(n9404) );
  NOR2_X1 U5892 ( .A1(n9414), .A2(n9405), .ZN(n4541) );
  INV_X1 U5893 ( .A(n4604), .ZN(n4603) );
  NOR2_X1 U5894 ( .A1(n5698), .A2(n4315), .ZN(n4604) );
  AND2_X1 U5895 ( .A1(n8130), .A2(n8132), .ZN(n4312) );
  INV_X1 U5896 ( .A(n4814), .ZN(n4813) );
  INV_X1 U5897 ( .A(n4560), .ZN(n4559) );
  OAI21_X1 U5898 ( .B1(n9354), .B2(n4561), .A(n7974), .ZN(n4560) );
  INV_X1 U5899 ( .A(n9492), .ZN(n9622) );
  NAND2_X1 U5900 ( .A1(n5387), .A2(n5386), .ZN(n9492) );
  AND2_X1 U5901 ( .A1(n4646), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4313) );
  INV_X1 U5902 ( .A(n7624), .ZN(n7742) );
  NAND2_X1 U5903 ( .A1(n5279), .A2(n5278), .ZN(n7624) );
  NAND2_X1 U5904 ( .A1(n9118), .A2(n9117), .ZN(n4314) );
  NOR2_X1 U5905 ( .A1(n9167), .A2(n9179), .ZN(n4315) );
  INV_X1 U5906 ( .A(n4806), .ZN(n4805) );
  NOR2_X1 U5907 ( .A1(n4810), .A2(n4807), .ZN(n4806) );
  AND2_X1 U5908 ( .A1(n7543), .A2(n7542), .ZN(n4316) );
  INV_X1 U5909 ( .A(n5710), .ZN(n4595) );
  INV_X1 U5910 ( .A(n4733), .ZN(n4732) );
  NOR2_X1 U5911 ( .A1(n5322), .A2(n5323), .ZN(n4733) );
  AND2_X1 U5912 ( .A1(n6217), .A2(n8452), .ZN(n4317) );
  AND2_X1 U5913 ( .A1(n8123), .A2(n6251), .ZN(n8434) );
  AND2_X1 U5914 ( .A1(n9608), .A2(n9388), .ZN(n4318) );
  AND2_X1 U5915 ( .A1(n9004), .A2(n8924), .ZN(n4319) );
  OR2_X1 U5916 ( .A1(n9939), .A2(n7488), .ZN(n8375) );
  NOR2_X1 U5917 ( .A1(n7318), .A2(n9184), .ZN(n4320) );
  NAND2_X1 U5918 ( .A1(n8317), .A2(n8310), .ZN(n8453) );
  INV_X1 U5919 ( .A(n8453), .ZN(n6217) );
  AND2_X1 U5920 ( .A1(n7477), .A2(n9825), .ZN(n4321) );
  INV_X1 U5921 ( .A(n4562), .ZN(n4380) );
  XNOR2_X1 U5922 ( .A(n4960), .B(SI_1_), .ZN(n4959) );
  NAND2_X1 U5923 ( .A1(n6226), .A2(n6225), .ZN(n4322) );
  AND2_X1 U5924 ( .A1(n7113), .A2(n9895), .ZN(n4323) );
  XNOR2_X1 U5925 ( .A(n4937), .B(n5558), .ZN(n4950) );
  INV_X1 U5926 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4874) );
  AND2_X1 U5927 ( .A1(n9405), .A2(n9428), .ZN(n4324) );
  NAND2_X1 U5928 ( .A1(n4695), .A2(n4694), .ZN(n4325) );
  AND2_X1 U5929 ( .A1(n8023), .A2(n4561), .ZN(n4326) );
  AND2_X1 U5930 ( .A1(n5085), .A2(SI_6_), .ZN(n4327) );
  AND2_X1 U5931 ( .A1(n5270), .A2(SI_13_), .ZN(n4328) );
  AND2_X1 U5932 ( .A1(n6336), .A2(n8514), .ZN(n4329) );
  INV_X1 U5933 ( .A(n4552), .ZN(n4551) );
  NAND2_X1 U5934 ( .A1(n8058), .A2(n9352), .ZN(n4552) );
  AND2_X1 U5935 ( .A1(n5439), .A2(n5438), .ZN(n4330) );
  OR2_X1 U5936 ( .A1(n7387), .A2(n7386), .ZN(n4331) );
  NAND2_X1 U5937 ( .A1(n4766), .A2(n4765), .ZN(n4526) );
  NOR2_X1 U5938 ( .A1(n7690), .A2(n5734), .ZN(n4332) );
  OR2_X1 U5939 ( .A1(n8296), .A2(n8533), .ZN(n4333) );
  AND2_X1 U5940 ( .A1(n8978), .A2(n8901), .ZN(n4334) );
  OR2_X1 U5941 ( .A1(n8040), .A2(n7905), .ZN(n4335) );
  AND2_X1 U5942 ( .A1(n5083), .A2(n5070), .ZN(n4336) );
  AND2_X1 U5943 ( .A1(n8354), .A2(n8359), .ZN(n8481) );
  INV_X1 U5944 ( .A(n7802), .ZN(n4566) );
  OR2_X1 U5945 ( .A1(n8088), .A2(n8244), .ZN(n4337) );
  AND2_X1 U5946 ( .A1(n4882), .A2(n5649), .ZN(n4338) );
  AND2_X1 U5947 ( .A1(n8024), .A2(n4559), .ZN(n4339) );
  AND2_X1 U5948 ( .A1(n4835), .A2(n4834), .ZN(n4340) );
  OR2_X1 U5949 ( .A1(n9007), .A2(n8933), .ZN(n8415) );
  AND2_X1 U5950 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4341) );
  INV_X1 U5951 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6273) );
  INV_X1 U5952 ( .A(n8356), .ZN(n4402) );
  NAND2_X1 U5953 ( .A1(n4755), .A2(n5158), .ZN(n7580) );
  NAND2_X1 U5954 ( .A1(n5108), .A2(n6351), .ZN(n7471) );
  AND2_X1 U5955 ( .A1(n5648), .A2(n4884), .ZN(n5651) );
  NAND2_X1 U5956 ( .A1(n9330), .A2(n8030), .ZN(n8040) );
  INV_X1 U5957 ( .A(n8040), .ZN(n4446) );
  AND2_X1 U5958 ( .A1(n7974), .A2(n7877), .ZN(n8023) );
  INV_X1 U5959 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4397) );
  OAI21_X1 U5960 ( .B1(n8216), .B2(n8217), .A(n8103), .ZN(n8262) );
  NAND2_X1 U5961 ( .A1(n4406), .A2(n4404), .ZN(n7699) );
  NAND2_X1 U5962 ( .A1(n8101), .A2(n8206), .ZN(n8216) );
  INV_X1 U5963 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4889) );
  AND2_X1 U5964 ( .A1(n7623), .A2(n7690), .ZN(n7599) );
  NAND2_X1 U5965 ( .A1(n5317), .A2(n5321), .ZN(n9158) );
  AND3_X1 U5966 ( .A1(n4777), .A2(n5293), .A3(n5294), .ZN(n4342) );
  NOR2_X1 U5967 ( .A1(n5792), .A2(n5791), .ZN(n4343) );
  NAND2_X1 U5968 ( .A1(n5276), .A2(n4869), .ZN(n5299) );
  XOR2_X1 U5969 ( .A(n8989), .B(n8131), .Z(n4344) );
  INV_X1 U5970 ( .A(n9394), .ZN(n9542) );
  AND2_X1 U5971 ( .A1(n5547), .A2(n5546), .ZN(n9394) );
  NAND2_X1 U5972 ( .A1(n7599), .A2(n4543), .ZN(n4547) );
  AND2_X1 U5973 ( .A1(n4344), .A2(n8252), .ZN(n4345) );
  NOR2_X1 U5974 ( .A1(n5741), .A2(n9065), .ZN(n4346) );
  AND2_X1 U5975 ( .A1(n5276), .A2(n4302), .ZN(n5326) );
  AND2_X1 U5976 ( .A1(n6337), .A2(n4413), .ZN(n4347) );
  NOR2_X1 U5977 ( .A1(n5482), .A2(n4709), .ZN(n4708) );
  AND2_X1 U5978 ( .A1(n4822), .A2(n4301), .ZN(n4348) );
  INV_X1 U5979 ( .A(n4596), .ZN(n4594) );
  NAND2_X1 U5980 ( .A1(n9441), .A2(n9426), .ZN(n4596) );
  INV_X1 U5981 ( .A(n9956), .ZN(n4414) );
  NAND2_X1 U5982 ( .A1(n4789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6303) );
  OR2_X1 U5983 ( .A1(n7316), .A2(n9838), .ZN(n4349) );
  AND2_X1 U5984 ( .A1(n7564), .A2(n9321), .ZN(n7905) );
  OR2_X1 U5985 ( .A1(n4529), .A2(n7316), .ZN(n4350) );
  NAND2_X1 U5986 ( .A1(n6767), .A2(n6766), .ZN(n6912) );
  OAI21_X1 U5987 ( .B1(n7094), .B2(n4511), .A(n4508), .ZN(n7244) );
  NAND2_X1 U5988 ( .A1(n5222), .A2(n5221), .ZN(n7454) );
  NAND2_X1 U5989 ( .A1(n6933), .A2(n4794), .ZN(n7114) );
  NAND2_X1 U5990 ( .A1(n7094), .A2(n4297), .ZN(n7127) );
  AND2_X1 U5991 ( .A1(n4524), .A2(n4523), .ZN(n4351) );
  AND2_X1 U5992 ( .A1(n4386), .A2(n7921), .ZN(n4352) );
  NAND2_X1 U5993 ( .A1(n6917), .A2(n6916), .ZN(n6933) );
  NAND2_X1 U5994 ( .A1(n5036), .A2(n5035), .ZN(n7094) );
  OR2_X1 U5995 ( .A1(n9583), .A2(n5802), .ZN(n4353) );
  OR2_X1 U5996 ( .A1(n9583), .A2(n9846), .ZN(n4354) );
  INV_X1 U5997 ( .A(n5698), .ZN(n4606) );
  INV_X1 U5998 ( .A(n9030), .ZN(n9024) );
  INV_X1 U5999 ( .A(n8459), .ZN(n4495) );
  NAND2_X1 U6000 ( .A1(n4638), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U6001 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  AND2_X1 U6002 ( .A1(n9866), .A2(n9930), .ZN(n9935) );
  AND2_X1 U6003 ( .A1(n8666), .A2(n4638), .ZN(n4355) );
  NOR2_X1 U6004 ( .A1(n8612), .A2(n8605), .ZN(n4356) );
  NOR2_X1 U6005 ( .A1(n8053), .A2(n8052), .ZN(n4357) );
  NAND2_X1 U6006 ( .A1(n4636), .A2(n8666), .ZN(n4358) );
  INV_X1 U6007 ( .A(n4637), .ZN(n4636) );
  OR2_X1 U6008 ( .A1(n6438), .A2(n6437), .ZN(n4652) );
  INV_X1 U6009 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7087) );
  INV_X1 U6010 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4464) );
  NAND3_X1 U6011 ( .A1(n8349), .A2(n8348), .A3(n8357), .ZN(n8351) );
  NAND2_X1 U6012 ( .A1(n8419), .A2(n4495), .ZN(n4494) );
  OAI21_X1 U6013 ( .B1(n4307), .B2(n4359), .A(n8836), .ZN(n8408) );
  NAND2_X1 U6014 ( .A1(n4360), .A2(n8489), .ZN(n8399) );
  NAND2_X1 U6015 ( .A1(n8392), .A2(n4361), .ZN(n4360) );
  OR2_X1 U6016 ( .A1(n8394), .A2(n8393), .ZN(n4361) );
  NAND2_X1 U6017 ( .A1(n4501), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U6018 ( .A1(n4499), .A2(n4498), .ZN(n8450) );
  NAND2_X1 U6019 ( .A1(n8409), .A2(n4495), .ZN(n4493) );
  OAI21_X2 U6020 ( .B1(n6917), .B2(n4793), .A(n4792), .ZN(n7348) );
  AOI21_X2 U6021 ( .B1(n7358), .B2(n7351), .A(n7357), .ZN(n7359) );
  OAI21_X2 U6022 ( .B1(n7486), .B2(n7485), .A(n7484), .ZN(n7502) );
  OAI21_X2 U6023 ( .B1(n8107), .B2(n8106), .A(n4288), .ZN(n8174) );
  NAND2_X1 U6024 ( .A1(n8250), .A2(n8251), .ZN(n4790) );
  NAND2_X1 U6025 ( .A1(n8121), .A2(n8120), .ZN(n8167) );
  OAI21_X1 U6026 ( .B1(n6684), .B2(n4783), .A(n4781), .ZN(n4784) );
  INV_X4 U6027 ( .A(n4913), .ZN(n8295) );
  OAI21_X1 U6028 ( .B1(n8089), .B2(n4791), .A(n4337), .ZN(n8241) );
  NAND2_X1 U6029 ( .A1(n4900), .A2(n4898), .ZN(n4901) );
  NAND2_X1 U6030 ( .A1(n7198), .A2(n7996), .ZN(n7197) );
  NAND2_X1 U6031 ( .A1(n7531), .A2(n8010), .ZN(n7530) );
  NAND2_X1 U6032 ( .A1(n4570), .A2(n5806), .ZN(P1_U3551) );
  NAND2_X1 U6033 ( .A1(n4786), .A2(n4785), .ZN(n8129) );
  AOI21_X1 U6034 ( .B1(n7710), .B2(n5702), .A(n5701), .ZN(n9500) );
  NOR2_X1 U6035 ( .A1(n8241), .A2(n8242), .ZN(n8153) );
  OAI22_X1 U6036 ( .A1(n5704), .A2(n5703), .B1(n5739), .B2(n4545), .ZN(n9485)
         );
  AOI21_X1 U6037 ( .B1(n9372), .B2(n4621), .A(n4619), .ZN(n4618) );
  AOI21_X1 U6038 ( .B1(n8521), .B2(n7503), .A(n7501), .ZN(n8089) );
  AOI211_X2 U6039 ( .C1(n8683), .C2(n8682), .A(n8681), .B(n8680), .ZN(n8684)
         );
  AND2_X1 U6040 ( .A1(n6520), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U6041 ( .A1(n7639), .A2(n7640), .ZN(n8556) );
  NOR2_X1 U6042 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  INV_X1 U6043 ( .A(n6528), .ZN(n4679) );
  INV_X1 U6044 ( .A(n4571), .ZN(n5803) );
  NAND2_X1 U6045 ( .A1(n4607), .A2(n4610), .ZN(n7291) );
  AND3_X1 U6046 ( .A1(n4932), .A2(n4929), .A3(n4931), .ZN(n4575) );
  NAND2_X1 U6047 ( .A1(n9339), .A2(n9835), .ZN(n4573) );
  NAND2_X1 U6048 ( .A1(n6836), .A2(n6838), .ZN(n6837) );
  INV_X1 U6049 ( .A(n5682), .ZN(n4369) );
  INV_X1 U6050 ( .A(n4597), .ZN(n7710) );
  OR2_X1 U6051 ( .A1(n5746), .A2(n4375), .ZN(n4371) );
  NAND2_X1 U6052 ( .A1(n5746), .A2(n4372), .ZN(n4370) );
  NAND2_X1 U6053 ( .A1(n5746), .A2(n9354), .ZN(n9357) );
  NAND2_X1 U6054 ( .A1(n4379), .A2(n4378), .ZN(n9382) );
  NAND3_X1 U6055 ( .A1(n4385), .A2(n4383), .A3(n8008), .ZN(n4382) );
  NAND3_X1 U6056 ( .A1(n4384), .A2(n4386), .A3(n7802), .ZN(n4385) );
  NAND2_X1 U6057 ( .A1(n5071), .A2(n4336), .ZN(n4477) );
  NAND2_X2 U6058 ( .A1(n6361), .A2(P1_U3086), .ZN(n9640) );
  MUX2_X1 U6059 ( .A(n6372), .B(n6385), .S(n8295), .Z(n5049) );
  MUX2_X1 U6060 ( .A(n5114), .B(n10020), .S(n8295), .Z(n5116) );
  MUX2_X1 U6061 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8295), .Z(n5085) );
  MUX2_X1 U6062 ( .A(n5053), .B(n6386), .S(n8295), .Z(n5072) );
  MUX2_X1 U6063 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8295), .Z(n5112) );
  MUX2_X1 U6064 ( .A(n10071), .B(n6411), .S(n8295), .Z(n5121) );
  MUX2_X1 U6065 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n8295), .Z(n5270) );
  MUX2_X1 U6066 ( .A(n5271), .B(n6761), .S(n8295), .Z(n5273) );
  MUX2_X1 U6067 ( .A(n8079), .B(n6198), .S(n8295), .Z(n5770) );
  NAND2_X1 U6068 ( .A1(n4398), .A2(n4399), .ZN(n7424) );
  NAND2_X1 U6069 ( .A1(n7033), .A2(n4400), .ZN(n4398) );
  NAND2_X1 U6070 ( .A1(n6244), .A2(n4408), .ZN(n4406) );
  NAND3_X1 U6071 ( .A1(n4418), .A2(n4419), .A3(n8447), .ZN(n6252) );
  NAND2_X1 U6072 ( .A1(n7904), .A2(n4432), .ZN(n4431) );
  NAND3_X1 U6073 ( .A1(n5722), .A2(n7914), .A3(n6830), .ZN(n4451) );
  NAND2_X1 U6074 ( .A1(n7992), .A2(n7010), .ZN(n4452) );
  MUX2_X1 U6075 ( .A(n4464), .B(n4463), .S(n6568), .Z(n7029) );
  NAND3_X1 U6076 ( .A1(n4467), .A2(n4465), .A3(n8461), .ZN(n8466) );
  NAND2_X1 U6077 ( .A1(n4477), .A2(n4478), .ZN(n5111) );
  NAND2_X1 U6078 ( .A1(n5075), .A2(n5074), .ZN(n5084) );
  NAND3_X1 U6079 ( .A1(n8364), .A2(n4485), .A3(n4495), .ZN(n4484) );
  NAND4_X1 U6080 ( .A1(n4503), .A2(n8747), .A3(n8433), .A4(n8472), .ZN(n4502)
         );
  NAND3_X1 U6081 ( .A1(n8429), .A2(n8428), .A3(n8767), .ZN(n4503) );
  NOR2_X2 U6082 ( .A1(n5087), .A2(n4504), .ZN(n5276) );
  NAND4_X1 U6083 ( .A1(n4866), .A2(n4868), .A3(n4867), .A4(n5089), .ZN(n4504)
         );
  NAND4_X1 U6084 ( .A1(n4762), .A2(n5022), .A3(n4904), .A4(n4865), .ZN(n5087)
         );
  INV_X1 U6085 ( .A(n4505), .ZN(n4508) );
  NAND2_X1 U6086 ( .A1(n4509), .A2(n5061), .ZN(n4506) );
  XNOR2_X2 U6087 ( .A(n4512), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6088 ( .A1(n5373), .A2(n4276), .ZN(n4513) );
  NAND2_X1 U6089 ( .A1(n4513), .A2(n4514), .ZN(n9071) );
  INV_X1 U6090 ( .A(n5373), .ZN(n4517) );
  NAND2_X1 U6091 ( .A1(n4521), .A2(n5216), .ZN(n4523) );
  NAND3_X1 U6092 ( .A1(n6352), .A2(n5216), .A3(n4522), .ZN(n4524) );
  OAI22_X1 U6093 ( .A1(n5290), .A2(n4525), .B1(n5289), .B2(n5293), .ZN(n5316)
         );
  INV_X1 U6094 ( .A(n7316), .ZN(n4527) );
  NAND2_X1 U6095 ( .A1(n4531), .A2(n7200), .ZN(n4534) );
  INV_X1 U6096 ( .A(n4534), .ZN(n7283) );
  INV_X1 U6097 ( .A(n4547), .ZN(n9508) );
  AND2_X1 U6098 ( .A1(n9373), .A2(n4550), .ZN(n9333) );
  NAND2_X1 U6099 ( .A1(n9373), .A2(n4548), .ZN(n9327) );
  NAND2_X1 U6100 ( .A1(n9373), .A2(n4551), .ZN(n5777) );
  AND2_X1 U6101 ( .A1(n9373), .A2(n9352), .ZN(n9348) );
  NAND2_X1 U6102 ( .A1(n5746), .A2(n4339), .ZN(n4553) );
  OAI211_X1 U6103 ( .C1(n5746), .C2(n4556), .A(n4554), .B(n4553), .ZN(n5779)
         );
  INV_X1 U6104 ( .A(n5733), .ZN(n4568) );
  OAI21_X1 U6105 ( .B1(n7532), .B2(n4569), .A(n4567), .ZN(n7662) );
  NAND2_X1 U6106 ( .A1(n7662), .A2(n7661), .ZN(n5737) );
  NAND2_X1 U6107 ( .A1(n6830), .A2(n5722), .ZN(n4578) );
  NAND2_X1 U6108 ( .A1(n4579), .A2(n7991), .ZN(n6828) );
  OAI21_X1 U6109 ( .B1(n7991), .B2(n4579), .A(n6828), .ZN(n7109) );
  NAND2_X1 U6110 ( .A1(n7018), .A2(n4583), .ZN(n4582) );
  INV_X1 U6111 ( .A(n4580), .ZN(n4583) );
  NAND2_X1 U6112 ( .A1(n9434), .A2(n4588), .ZN(n4586) );
  OAI21_X1 U6113 ( .B1(n7615), .B2(n4600), .A(n4598), .ZN(n4597) );
  NAND2_X1 U6114 ( .A1(n7282), .A2(n4608), .ZN(n4607) );
  OAI211_X1 U6115 ( .C1(n8064), .C2(n4353), .A(n4292), .B(n4613), .ZN(n5759)
         );
  OAI211_X1 U6116 ( .C1(n8064), .C2(n4354), .A(n4615), .B(n4291), .ZN(n5763)
         );
  OAI21_X1 U6117 ( .B1(n9372), .B2(n5713), .A(n5712), .ZN(n9347) );
  INV_X1 U6118 ( .A(n5707), .ZN(n9468) );
  INV_X1 U6119 ( .A(n9448), .ZN(n5708) );
  OAI21_X1 U6120 ( .B1(n5707), .B2(n4346), .A(n4847), .ZN(n9448) );
  NAND2_X1 U6121 ( .A1(n4909), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U6122 ( .A1(n5732), .A2(n5731), .ZN(n7532) );
  NAND2_X1 U6123 ( .A1(n5111), .A2(n5110), .ZN(n4685) );
  NAND2_X1 U6124 ( .A1(n4685), .A2(n5113), .ZN(n5142) );
  NAND2_X1 U6125 ( .A1(n4625), .A2(n4279), .ZN(n8686) );
  NAND2_X1 U6126 ( .A1(n4304), .A2(n4632), .ZN(n4625) );
  OAI21_X1 U6127 ( .B1(n4637), .B2(n8609), .A(n4634), .ZN(n8661) );
  NAND2_X1 U6128 ( .A1(n4647), .A2(n4646), .ZN(n6520) );
  NAND2_X1 U6129 ( .A1(n6454), .A2(n6439), .ZN(n6515) );
  NAND2_X1 U6130 ( .A1(n4652), .A2(n4650), .ZN(n6454) );
  NAND2_X1 U6131 ( .A1(n4651), .A2(n6439), .ZN(n4641) );
  NAND2_X1 U6132 ( .A1(n4643), .A2(n4642), .ZN(n6516) );
  NAND2_X1 U6133 ( .A1(n4647), .A2(n4313), .ZN(n4642) );
  INV_X1 U6134 ( .A(n4644), .ZN(n4643) );
  AOI21_X1 U6135 ( .B1(n4647), .B2(n4646), .A(P2_REG2_REG_2__SCAN_IN), .ZN(
        n4644) );
  INV_X1 U6136 ( .A(n6439), .ZN(n4645) );
  NAND3_X1 U6137 ( .A1(n4659), .A2(n8538), .A3(P2_REG2_REG_5__SCAN_IN), .ZN(
        n8540) );
  NAND2_X1 U6138 ( .A1(n4661), .A2(n6665), .ZN(n4659) );
  NAND2_X1 U6139 ( .A1(n4660), .A2(n5942), .ZN(n6533) );
  INV_X1 U6140 ( .A(n6532), .ZN(n4661) );
  NAND2_X1 U6141 ( .A1(n7543), .A2(n4664), .ZN(n4662) );
  OAI211_X1 U6142 ( .C1(n7543), .C2(n7630), .A(n4662), .B(n4663), .ZN(n7544)
         );
  NOR2_X1 U6143 ( .A1(n7544), .A2(n7551), .ZN(n7631) );
  INV_X1 U6144 ( .A(n4666), .ZN(n6973) );
  NAND2_X1 U6145 ( .A1(n5218), .A2(n4689), .ZN(n4686) );
  NAND2_X1 U6146 ( .A1(n4686), .A2(n4687), .ZN(n5297) );
  NAND2_X1 U6147 ( .A1(n8895), .A2(n8315), .ZN(n8458) );
  NAND2_X1 U6148 ( .A1(n8468), .A2(n8459), .ZN(n4695) );
  NAND2_X1 U6149 ( .A1(n8318), .A2(n8317), .ZN(n8468) );
  INV_X1 U6150 ( .A(n8895), .ZN(n4696) );
  NAND2_X1 U6151 ( .A1(n4697), .A2(n5166), .ZN(n5174) );
  NAND2_X1 U6152 ( .A1(n5162), .A2(n4698), .ZN(n4697) );
  MUX2_X1 U6153 ( .A(n6367), .B(n4957), .S(n4913), .Z(n4987) );
  NAND2_X1 U6154 ( .A1(n5443), .A2(n4715), .ZN(n4714) );
  INV_X1 U6155 ( .A(n5443), .ZN(n4704) );
  NAND2_X1 U6156 ( .A1(n4714), .A2(n4713), .ZN(n5464) );
  NAND2_X1 U6157 ( .A1(n5538), .A2(n5537), .ZN(n5544) );
  NAND2_X1 U6158 ( .A1(n5538), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U6159 ( .A1(n5324), .A2(n4732), .ZN(n4731) );
  NAND2_X2 U6160 ( .A1(n8083), .A2(n9040), .ZN(n5897) );
  XNOR2_X2 U6161 ( .A(n4735), .B(n5853), .ZN(n9040) );
  XNOR2_X2 U6162 ( .A(n5850), .B(n5851), .ZN(n8083) );
  INV_X1 U6163 ( .A(n8879), .ZN(n6231) );
  AND2_X2 U6164 ( .A1(n6232), .A2(n8325), .ZN(n8879) );
  NAND2_X1 U6165 ( .A1(n6247), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U6166 ( .A1(n8415), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U6167 ( .A1(n4745), .A2(n4743), .ZN(n6245) );
  INV_X1 U6168 ( .A(n8406), .ZN(n4746) );
  NAND2_X1 U6169 ( .A1(n6745), .A2(n8345), .ZN(n4749) );
  AND3_X2 U6170 ( .A1(n6222), .A2(n5820), .A3(n4751), .ZN(n5852) );
  NAND3_X1 U6171 ( .A1(n6222), .A2(n5820), .A3(n4837), .ZN(n4838) );
  NAND2_X1 U6172 ( .A1(n6253), .A2(n8319), .ZN(n6320) );
  NAND2_X1 U6173 ( .A1(n6253), .A2(n4753), .ZN(n6319) );
  NAND2_X1 U6174 ( .A1(n4757), .A2(n5158), .ZN(n4756) );
  NAND2_X1 U6175 ( .A1(n5317), .A2(n5320), .ZN(n4761) );
  NAND3_X1 U6176 ( .A1(n5022), .A2(n4762), .A3(n4954), .ZN(n5068) );
  NOR2_X2 U6177 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5022) );
  NAND2_X1 U6178 ( .A1(n5276), .A2(n4769), .ZN(n4877) );
  NOR2_X1 U6179 ( .A1(n4773), .A2(n4771), .ZN(n4769) );
  NAND2_X1 U6180 ( .A1(n4892), .A2(n4775), .ZN(n4881) );
  NAND2_X1 U6181 ( .A1(n4892), .A2(n4774), .ZN(n4776) );
  NAND2_X1 U6182 ( .A1(n4892), .A2(n4894), .ZN(n4890) );
  NAND2_X1 U6183 ( .A1(n8152), .A2(n4779), .ZN(n8283) );
  NAND2_X1 U6184 ( .A1(n8283), .A2(n8097), .ZN(n8207) );
  INV_X1 U6185 ( .A(n4782), .ZN(n4781) );
  INV_X1 U6186 ( .A(n6766), .ZN(n4783) );
  OAI21_X1 U6187 ( .B1(n8224), .B2(n8195), .A(n4787), .ZN(n8197) );
  NAND2_X1 U6188 ( .A1(n8224), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U6189 ( .A1(n6222), .A2(n6219), .ZN(n6272) );
  NAND3_X1 U6190 ( .A1(n6222), .A2(n6219), .A3(n6273), .ZN(n4789) );
  NAND2_X1 U6191 ( .A1(n4790), .A2(n8252), .ZN(n8121) );
  NAND2_X1 U6192 ( .A1(n8145), .A2(n8135), .ZN(n8137) );
  NAND3_X1 U6193 ( .A1(n6560), .A2(n6559), .A3(n6563), .ZN(n6682) );
  NAND2_X1 U6194 ( .A1(n6682), .A2(n6681), .ZN(n6686) );
  AND2_X1 U6195 ( .A1(n6934), .A2(n6932), .ZN(n4794) );
  NAND3_X1 U6196 ( .A1(n4795), .A2(n6379), .A3(n8499), .ZN(n6550) );
  INV_X1 U6197 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U6198 ( .A1(n8758), .A2(n4804), .ZN(n4803) );
  NOR2_X1 U6199 ( .A1(n6163), .A2(n8916), .ZN(n4814) );
  NAND2_X1 U6200 ( .A1(n4818), .A2(n5971), .ZN(n6951) );
  NAND2_X1 U6201 ( .A1(n7140), .A2(n4821), .ZN(n4820) );
  INV_X1 U6202 ( .A(n7140), .ZN(n4823) );
  NAND2_X1 U6203 ( .A1(n4824), .A2(n4825), .ZN(n6006) );
  NAND2_X1 U6204 ( .A1(n6964), .A2(n5994), .ZN(n4824) );
  NAND2_X1 U6205 ( .A1(n8712), .A2(n8710), .ZN(n8718) );
  NAND2_X1 U6206 ( .A1(n4827), .A2(n4826), .ZN(n6218) );
  NAND2_X1 U6207 ( .A1(n8712), .A2(n4828), .ZN(n4827) );
  OAI21_X1 U6208 ( .B1(n8710), .B2(n4830), .A(n6208), .ZN(n4829) );
  NAND2_X1 U6209 ( .A1(n8807), .A2(n4833), .ZN(n4831) );
  NAND2_X1 U6210 ( .A1(n4831), .A2(n4832), .ZN(n8786) );
  INV_X1 U6211 ( .A(n4835), .ZN(n8811) );
  NAND2_X1 U6212 ( .A1(n7508), .A2(n4287), .ZN(n8854) );
  NAND2_X1 U6213 ( .A1(n5820), .A2(n6222), .ZN(n6283) );
  NAND2_X1 U6214 ( .A1(n7884), .A2(n7883), .ZN(n7896) );
  NAND2_X1 U6215 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  NAND2_X1 U6216 ( .A1(n7872), .A2(n7871), .ZN(n7884) );
  NAND2_X1 U6217 ( .A1(n4841), .A2(n9551), .ZN(n9522) );
  INV_X1 U6218 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U6219 ( .A1(n7760), .A2(n7759), .ZN(n7888) );
  NAND2_X1 U6220 ( .A1(n7888), .A2(n7761), .ZN(n7765) );
  NAND2_X1 U6221 ( .A1(n5766), .A2(n5715), .ZN(n8064) );
  OR2_X1 U6222 ( .A1(n4900), .A2(n4875), .ZN(n4876) );
  OR2_X1 U6223 ( .A1(n4885), .A2(n4875), .ZN(n5354) );
  XNOR2_X1 U6224 ( .A(n6318), .B(n6317), .ZN(n8702) );
  NAND2_X1 U6225 ( .A1(n5927), .A2(n5926), .ZN(n6234) );
  AOI22_X1 U6226 ( .A1(n4998), .A2(n7008), .B1(n5604), .B2(n7009), .ZN(n4949)
         );
  NAND2_X1 U6227 ( .A1(n5913), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5875) );
  INV_X1 U6228 ( .A(n6258), .ZN(n8506) );
  CLKBUF_X1 U6229 ( .A(n9500), .Z(n9501) );
  NAND2_X4 U6230 ( .A1(n5558), .A2(n5060), .ZN(n4998) );
  CLKBUF_X1 U6231 ( .A(n7348), .Z(n7209) );
  CLKBUF_X1 U6232 ( .A(n8250), .Z(n8254) );
  AOI22_X2 U6233 ( .A1(n8726), .A2(n6187), .B1(n8715), .B2(n8975), .ZN(n8712)
         );
  AOI21_X2 U6234 ( .B1(n8786), .B2(n8785), .A(n6141), .ZN(n8766) );
  AOI21_X2 U6235 ( .B1(n8183), .B2(n8117), .A(n4848), .ZN(n8250) );
  OAI21_X2 U6236 ( .B1(n8766), .B2(n8767), .A(n6151), .ZN(n8758) );
  INV_X1 U6237 ( .A(n9040), .ZN(n5855) );
  NAND2_X2 U6238 ( .A1(n6735), .A2(n8882), .ZN(n8859) );
  AND2_X2 U6239 ( .A1(n6729), .A2(n6334), .ZN(n9956) );
  INV_X2 U6240 ( .A(n9943), .ZN(n9941) );
  NOR2_X1 U6241 ( .A1(n8695), .A2(n9030), .ZN(n6313) );
  INV_X1 U6242 ( .A(n6378), .ZN(n6375) );
  AND2_X1 U6243 ( .A1(n6140), .A2(n6139), .ZN(n8934) );
  INV_X1 U6244 ( .A(P1_U3973), .ZN(n9170) );
  AND4_X1 U6245 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n5797)
         );
  AND2_X1 U6246 ( .A1(n5161), .A2(n5123), .ZN(n4839) );
  INV_X1 U6247 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4865) );
  NOR2_X1 U6248 ( .A1(n8313), .A2(n8312), .ZN(n4840) );
  XOR2_X1 U6249 ( .A(n9330), .B(n9327), .Z(n4841) );
  AND2_X1 U6250 ( .A1(n5776), .A2(n7450), .ZN(n4842) );
  OR2_X1 U6251 ( .A1(n8058), .A2(n9590), .ZN(n4843) );
  OR2_X1 U6252 ( .A1(n9352), .A2(n9157), .ZN(n4844) );
  AND2_X1 U6253 ( .A1(n9465), .A2(n5742), .ZN(n4845) );
  AND2_X1 U6254 ( .A1(n8961), .A2(n8457), .ZN(n4846) );
  OR2_X1 U6255 ( .A1(n9618), .A2(n9455), .ZN(n4847) );
  NOR2_X1 U6256 ( .A1(n8116), .A2(n8115), .ZN(n4848) );
  AND4_X1 U6257 ( .A1(n8713), .A2(n8747), .A3(n8497), .A4(n8496), .ZN(n4850)
         );
  OR2_X1 U6258 ( .A1(n8058), .A2(n9631), .ZN(n4851) );
  AND3_X1 U6259 ( .A1(n5676), .A2(n9151), .A3(n5675), .ZN(n4852) );
  AND2_X1 U6260 ( .A1(n5776), .A2(n7448), .ZN(n4853) );
  OR2_X1 U6261 ( .A1(n4275), .A2(n5914), .ZN(n4854) );
  INV_X1 U6262 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n6166) );
  INV_X1 U6263 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4898) );
  AND2_X1 U6264 ( .A1(n5030), .A2(n5029), .ZN(n4855) );
  AND2_X1 U6265 ( .A1(n9873), .A2(n6751), .ZN(n4856) );
  OR2_X1 U6266 ( .A1(n9873), .A2(n6751), .ZN(n4857) );
  INV_X1 U6267 ( .A(n8884), .ZN(n5883) );
  INV_X1 U6268 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4911) );
  INV_X1 U6269 ( .A(n7454), .ZN(n5695) );
  INV_X1 U6270 ( .A(n8924), .ZN(n8177) );
  AND3_X1 U6271 ( .A1(n6131), .A2(n6130), .A3(n6129), .ZN(n8924) );
  NOR2_X1 U6272 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4858) );
  AND2_X1 U6273 ( .A1(n7974), .A2(n7973), .ZN(n4860) );
  INV_X1 U6274 ( .A(n6070), .ZN(n8855) );
  AND4_X1 U6275 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6070)
         );
  NOR2_X1 U6276 ( .A1(n5280), .A2(n5253), .ZN(n4861) );
  NAND2_X1 U6277 ( .A1(n9562), .A2(n9174), .ZN(n4862) );
  OR2_X1 U6278 ( .A1(n8870), .A2(n8161), .ZN(n4863) );
  INV_X1 U6279 ( .A(n8853), .ZN(n6085) );
  INV_X1 U6280 ( .A(n4984), .ZN(n5086) );
  AND2_X1 U6281 ( .A1(n7006), .A2(n7103), .ZN(n9813) );
  AND2_X2 U6282 ( .A1(n5762), .A2(n7005), .ZN(n9627) );
  AND2_X2 U6283 ( .A1(n5762), .A2(n5761), .ZN(n9854) );
  INV_X1 U6284 ( .A(n9854), .ZN(n5802) );
  NOR2_X1 U6285 ( .A1(n7880), .A2(n7905), .ZN(n7881) );
  AND2_X1 U6286 ( .A1(n7352), .A2(n9918), .ZN(n7349) );
  INV_X1 U6287 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U6288 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  AND4_X1 U6289 ( .A1(n6273), .A2(n6275), .A3(n10073), .A4(n6280), .ZN(n5811)
         );
  AOI21_X1 U6290 ( .B1(n7355), .B2(n7354), .A(n7353), .ZN(n7356) );
  NOR2_X1 U6291 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  INV_X1 U6292 ( .A(n7356), .ZN(n7357) );
  INV_X1 U6293 ( .A(n6134), .ZN(n5844) );
  NAND2_X1 U6294 ( .A1(n7895), .A2(n7894), .ZN(n7903) );
  INV_X1 U6295 ( .A(n8010), .ZN(n5731) );
  AND3_X1 U6296 ( .A1(n4888), .A2(n4886), .A3(n4889), .ZN(n4871) );
  INV_X1 U6297 ( .A(n6920), .ZN(n6916) );
  OR2_X1 U6298 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  INV_X1 U6299 ( .A(n8175), .ZN(n8108) );
  OAI21_X1 U6300 ( .B1(n8463), .B2(n8462), .A(n8467), .ZN(n8464) );
  INV_X1 U6301 ( .A(n6171), .ZN(n6170) );
  INV_X1 U6302 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5832) );
  OR2_X1 U6303 ( .A1(n8305), .A2(n5886), .ZN(n5890) );
  INV_X1 U6304 ( .A(n7385), .ZN(n7386) );
  INV_X1 U6305 ( .A(n8341), .ZN(n6236) );
  OR2_X1 U6306 ( .A1(n8921), .A2(n8787), .ZN(n6151) );
  INV_X1 U6307 ( .A(n8483), .ZN(n6034) );
  NOR2_X1 U6308 ( .A1(n7624), .A2(n9180), .ZN(n5698) );
  OR2_X1 U6309 ( .A1(n7750), .A2(n7751), .ZN(n7752) );
  INV_X1 U6310 ( .A(n5460), .ZN(n5461) );
  INV_X1 U6311 ( .A(SI_19_), .ZN(n5381) );
  INV_X1 U6312 ( .A(SI_14_), .ZN(n5272) );
  NAND2_X1 U6313 ( .A1(n4913), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4910) );
  INV_X1 U6314 ( .A(n4344), .ZN(n8120) );
  INV_X1 U6315 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6316 ( .A1(n8093), .A2(n6070), .ZN(n8094) );
  NAND2_X1 U6317 ( .A1(n6170), .A2(n6169), .ZN(n6180) );
  NAND2_X1 U6318 ( .A1(n5833), .A2(n5832), .ZN(n6015) );
  INV_X1 U6319 ( .A(n7392), .ZN(n7389) );
  INV_X1 U6320 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5848) );
  INV_X1 U6321 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5839) );
  OR2_X1 U6322 ( .A1(n6028), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6038) );
  INV_X1 U6323 ( .A(n6727), .ZN(n6331) );
  INV_X1 U6324 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10082) );
  OR2_X1 U6325 ( .A1(n6047), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6048) );
  AND2_X1 U6326 ( .A1(n5586), .A2(n5585), .ZN(n5792) );
  NAND2_X1 U6327 ( .A1(n5313), .A2(n5314), .ZN(n5321) );
  NOR2_X1 U6328 ( .A1(n5430), .A2(n9122), .ZN(n5447) );
  AND2_X1 U6329 ( .A1(n9772), .A2(n9296), .ZN(n9787) );
  NAND2_X1 U6330 ( .A1(n5695), .A2(n9660), .ZN(n5696) );
  AND2_X1 U6331 ( .A1(n5510), .A2(n5488), .ZN(n5489) );
  NAND2_X1 U6332 ( .A1(n5382), .A2(n5381), .ZN(n5423) );
  INV_X1 U6333 ( .A(n5240), .ZN(n5244) );
  OR2_X1 U6334 ( .A1(n6090), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6102) );
  OR2_X1 U6335 ( .A1(n6116), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6118) );
  XNOR2_X1 U6336 ( .A(n8129), .B(n8127), .ZN(n8271) );
  INV_X1 U6337 ( .A(n8469), .ZN(n6317) );
  OR2_X1 U6338 ( .A1(n6154), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6156) );
  INV_X1 U6339 ( .A(n8824), .ZN(n6246) );
  OR2_X1 U6340 ( .A1(n7462), .A2(n8388), .ZN(n8487) );
  INV_X1 U6341 ( .A(n9902), .ZN(n8917) );
  OR2_X1 U6342 ( .A1(n6369), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6299) );
  INV_X1 U6343 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5965) );
  AND2_X1 U6344 ( .A1(n5062), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5095) );
  INV_X1 U6345 ( .A(n5520), .ZN(n5519) );
  OR2_X1 U6346 ( .A1(n5332), .A2(n5331), .ZN(n5358) );
  OAI21_X1 U6347 ( .B1(n9127), .B2(n9131), .A(n9051), .ZN(n9108) );
  AND2_X1 U6348 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5041) );
  NAND2_X1 U6349 ( .A1(n5447), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5471) );
  OR2_X1 U6350 ( .A1(n9685), .A2(n8049), .ZN(n9758) );
  INV_X1 U6351 ( .A(n9531), .ZN(n9352) );
  AND2_X1 U6352 ( .A1(n7836), .A2(n7909), .ZN(n9486) );
  INV_X1 U6353 ( .A(n8015), .ZN(n7661) );
  OR2_X1 U6354 ( .A1(n7811), .A2(n9181), .ZN(n5697) );
  OR2_X1 U6355 ( .A1(n5751), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5647) );
  INV_X1 U6356 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5089) );
  INV_X1 U6357 ( .A(n8174), .ZN(n8176) );
  INV_X1 U6358 ( .A(n8257), .ZN(n8290) );
  AND2_X1 U6359 ( .A1(n8309), .A2(n6216), .ZN(n9990) );
  AND3_X1 U6360 ( .A1(n5871), .A2(n5870), .A3(n5869), .ZN(n8933) );
  INV_X1 U6361 ( .A(n8673), .ZN(n8587) );
  AND2_X1 U6362 ( .A1(n6479), .A2(n8459), .ZN(n9874) );
  NOR2_X1 U6363 ( .A1(n8890), .A2(n8917), .ZN(n8826) );
  INV_X1 U6364 ( .A(n8885), .ZN(n8861) );
  INV_X1 U6365 ( .A(n8957), .ZN(n8953) );
  AND2_X1 U6366 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  INV_X1 U6367 ( .A(n9886), .ZN(n9940) );
  INV_X1 U6368 ( .A(n9935), .ZN(n9884) );
  INV_X1 U6369 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5864) );
  INV_X1 U6370 ( .A(n9661), .ZN(n9152) );
  INV_X1 U6371 ( .A(n9157), .ZN(n9675) );
  AND4_X1 U6372 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n9388)
         );
  AND4_X1 U6373 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n9099)
         );
  AND4_X1 U6374 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n7810)
         );
  INV_X1 U6375 ( .A(n9795), .ZN(n9777) );
  INV_X1 U6376 ( .A(n5385), .ZN(n9321) );
  NOR2_X1 U6377 ( .A1(n9854), .A2(n5804), .ZN(n5805) );
  NAND2_X1 U6378 ( .A1(n7622), .A2(n5720), .ZN(n9835) );
  NAND2_X1 U6379 ( .A1(n5643), .A2(n5645), .ZN(n5751) );
  INV_X1 U6380 ( .A(n8267), .ZN(n8287) );
  OR2_X1 U6381 ( .A1(n6543), .A2(n6479), .ZN(n8286) );
  INV_X1 U6382 ( .A(n8259), .ZN(n8293) );
  INV_X1 U6383 ( .A(n8716), .ZN(n8514) );
  INV_X1 U6384 ( .A(n8841), .ZN(n8856) );
  INV_X1 U6385 ( .A(n7488), .ZN(n8521) );
  OR2_X1 U6386 ( .A1(P2_U3150), .A2(n6395), .ZN(n8653) );
  OR2_X1 U6387 ( .A1(n6446), .A2(n8665), .ZN(n8685) );
  INV_X1 U6388 ( .A(n8859), .ZN(n8890) );
  NAND2_X1 U6389 ( .A1(n9956), .A2(n9940), .ZN(n8957) );
  NOR2_X1 U6390 ( .A1(n6313), .A2(n6315), .ZN(n6316) );
  OR2_X1 U6391 ( .A1(n9943), .A2(n9886), .ZN(n9030) );
  OR2_X1 U6392 ( .A1(n9943), .A2(n9935), .ZN(n9032) );
  AND2_X1 U6393 ( .A1(n6311), .A2(n6310), .ZN(n9943) );
  AND2_X1 U6394 ( .A1(n6499), .A2(n6369), .ZN(n6378) );
  AND2_X1 U6395 ( .A1(n6490), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6381) );
  INV_X1 U6396 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10120) );
  INV_X1 U6397 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10006) );
  INV_X1 U6398 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10020) );
  AND2_X1 U6399 ( .A1(n5663), .A2(n8054), .ZN(n9678) );
  AND2_X1 U6400 ( .A1(n5657), .A2(n7103), .ZN(n9157) );
  INV_X1 U6401 ( .A(n5797), .ZN(n9359) );
  INV_X1 U6402 ( .A(n9099), .ZN(n9178) );
  INV_X1 U6403 ( .A(n7810), .ZN(n9181) );
  OR2_X1 U6404 ( .A1(n9685), .A2(n6636), .ZN(n9764) );
  INV_X1 U6405 ( .A(n9683), .ZN(n9799) );
  OR2_X1 U6406 ( .A1(n9813), .A2(n9321), .ZN(n9806) );
  OR2_X1 U6407 ( .A1(n9813), .A2(n7049), .ZN(n7629) );
  INV_X1 U6408 ( .A(n9809), .ZN(n9520) );
  INV_X1 U6409 ( .A(n7450), .ZN(n9590) );
  INV_X1 U6410 ( .A(n9326), .ZN(n9598) );
  INV_X1 U6411 ( .A(n7669), .ZN(n9632) );
  INV_X1 U6412 ( .A(n9627), .ZN(n9846) );
  INV_X1 U6413 ( .A(n9815), .ZN(n9814) );
  INV_X1 U6414 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7693) );
  INV_X1 U6415 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10128) );
  INV_X1 U6416 ( .A(n8641), .ZN(P2_U3893) );
  AND2_X2 U6417 ( .A1(n6346), .A2(n6567), .ZN(P1_U3973) );
  OAI21_X1 U6418 ( .B1(n5803), .B2(n9846), .A(n5790), .ZN(P1_U3519) );
  NOR2_X1 U6419 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4868) );
  NOR2_X1 U6420 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4867) );
  NOR2_X1 U6421 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4866) );
  INV_X1 U6422 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4870) );
  XNOR2_X1 U6423 ( .A(n4872), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5641) );
  INV_X1 U6424 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6425 ( .A1(n4877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6426 ( .A1(n5641), .A2(n4880), .ZN(n4934) );
  NAND2_X1 U6427 ( .A1(n5354), .A2(n4886), .ZN(n4887) );
  NAND2_X1 U6428 ( .A1(n5651), .A2(n5385), .ZN(n5717) );
  NAND2_X1 U6429 ( .A1(n4890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4891) );
  INV_X1 U6430 ( .A(n4892), .ZN(n4893) );
  INV_X1 U6431 ( .A(n7048), .ZN(n4933) );
  OAI21_X1 U6432 ( .B1(n7984), .B2(n4933), .A(n5717), .ZN(n4897) );
  NAND2_X2 U6433 ( .A1(n4897), .A2(n4934), .ZN(n5060) );
  NAND2_X1 U6434 ( .A1(n4922), .A2(n4919), .ZN(n4917) );
  NAND2_X1 U6435 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4903) );
  MUX2_X1 U6436 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4903), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n4906) );
  INV_X1 U6437 ( .A(n4954), .ZN(n4905) );
  NAND2_X1 U6438 ( .A1(n4906), .A2(n4905), .ZN(n6617) );
  INV_X1 U6439 ( .A(n6617), .ZN(n9199) );
  INV_X1 U6440 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4908) );
  NAND2_X1 U6441 ( .A1(n4908), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U6442 ( .A1(n4992), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4915) );
  AND2_X1 U6443 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U6444 ( .A1(n4913), .A2(n4912), .ZN(n4940) );
  XNOR2_X1 U6445 ( .A(n4959), .B(n4958), .ZN(n6365) );
  NAND2_X1 U6446 ( .A1(n4998), .A2(n5682), .ZN(n4936) );
  NAND2_X1 U6447 ( .A1(n4917), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4918) );
  MUX2_X1 U6448 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4918), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4923) );
  AND2_X1 U6449 ( .A1(n4920), .A2(n4919), .ZN(n4921) );
  NAND2_X1 U6450 ( .A1(n5008), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4932) );
  INV_X1 U6451 ( .A(n4928), .ZN(n4926) );
  NAND2_X1 U6452 ( .A1(n5007), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U6453 ( .A1(n4979), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4930) );
  AND2_X2 U6454 ( .A1(n8085), .A2(n4928), .ZN(n5010) );
  NAND2_X1 U6455 ( .A1(n5010), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6456 ( .A1(n5683), .A2(n5262), .ZN(n4935) );
  NAND2_X1 U6457 ( .A1(n4936), .A2(n4935), .ZN(n4937) );
  AOI22_X1 U6458 ( .A1(n5683), .A2(n5581), .B1(n6843), .B2(n5604), .ZN(n4951)
         );
  XNOR2_X1 U6459 ( .A(n4950), .B(n4951), .ZN(n8070) );
  INV_X1 U6460 ( .A(SI_0_), .ZN(n4939) );
  INV_X1 U6461 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U6462 ( .B1(n8295), .B2(n4939), .A(n4938), .ZN(n4941) );
  AND2_X1 U6463 ( .A1(n4941), .A2(n4940), .ZN(n9642) );
  NAND2_X1 U6464 ( .A1(n4979), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U6465 ( .A1(n5007), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U6466 ( .A1(n5008), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6467 ( .A1(n5010), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4942) );
  INV_X1 U6468 ( .A(n4934), .ZN(n5662) );
  NAND2_X1 U6469 ( .A1(n5662), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U6470 ( .A1(n4949), .A2(n4946), .ZN(n6756) );
  NAND2_X1 U6471 ( .A1(n7009), .A2(n5581), .ZN(n4948) );
  AOI22_X1 U6472 ( .A1(n7008), .A2(n5262), .B1(n5662), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6473 ( .A1(n4948), .A2(n4947), .ZN(n6757) );
  AOI22_X1 U6474 ( .A1(n6756), .A2(n6757), .B1(n4949), .B2(n5627), .ZN(n8072)
         );
  NAND2_X1 U6475 ( .A1(n8070), .A2(n8072), .ZN(n8071) );
  INV_X1 U6476 ( .A(n4950), .ZN(n4952) );
  NAND2_X1 U6477 ( .A1(n4952), .A2(n4951), .ZN(n4953) );
  NAND2_X1 U6478 ( .A1(n8071), .A2(n4953), .ZN(n6821) );
  OR2_X1 U6479 ( .A1(n4954), .A2(n4875), .ZN(n5024) );
  INV_X1 U6480 ( .A(n5024), .ZN(n4955) );
  NAND2_X1 U6481 ( .A1(n4955), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4956) );
  INV_X1 U6482 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10106) );
  NAND2_X1 U6483 ( .A1(n5024), .A2(n10106), .ZN(n4993) );
  AND2_X1 U6484 ( .A1(n4956), .A2(n4993), .ZN(n6784) );
  NAND2_X1 U6485 ( .A1(n5402), .A2(n6784), .ZN(n4965) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4957) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6367) );
  XNOR2_X1 U6488 ( .A(n4987), .B(SI_2_), .ZN(n4985) );
  NAND2_X1 U6489 ( .A1(n4960), .A2(SI_1_), .ZN(n4961) );
  XNOR2_X1 U6490 ( .A(n4986), .B(n4985), .ZN(n6368) );
  INV_X1 U6491 ( .A(n6368), .ZN(n4962) );
  NAND2_X1 U6492 ( .A1(n4984), .A2(n4962), .ZN(n4964) );
  NAND2_X1 U6493 ( .A1(n4992), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6494 ( .A1(n6834), .A2(n4998), .ZN(n4971) );
  NAND2_X1 U6495 ( .A1(n5007), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6496 ( .A1(n5008), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6497 ( .A1(n4979), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6498 ( .A1(n5010), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4966) );
  NAND4_X1 U6499 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n9192)
         );
  NAND2_X1 U6500 ( .A1(n9192), .A2(n5262), .ZN(n4970) );
  NAND2_X1 U6501 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  XNOR2_X1 U6502 ( .A(n4972), .B(n5558), .ZN(n4973) );
  AOI22_X1 U6503 ( .A1(n9192), .A2(n5581), .B1(n6834), .B2(n5624), .ZN(n4974)
         );
  NAND2_X1 U6504 ( .A1(n6821), .A2(n6822), .ZN(n4977) );
  INV_X1 U6505 ( .A(n4973), .ZN(n4975) );
  NAND2_X1 U6506 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NAND2_X1 U6507 ( .A1(n4977), .A2(n4976), .ZN(n6896) );
  INV_X1 U6508 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U6509 ( .A1(n5008), .A2(n7268), .ZN(n4983) );
  INV_X1 U6510 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6511 ( .A1(n5518), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6512 ( .A1(n5010), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6513 ( .A1(n9191), .A2(n5624), .ZN(n5000) );
  INV_X1 U6514 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6515 ( .A1(n4988), .A2(SI_2_), .ZN(n4989) );
  NAND2_X1 U6516 ( .A1(n4990), .A2(n4989), .ZN(n5016) );
  XNOR2_X1 U6517 ( .A(n5017), .B(SI_3_), .ZN(n5015) );
  XNOR2_X1 U6518 ( .A(n5016), .B(n5015), .ZN(n6366) );
  INV_X1 U6519 ( .A(n6366), .ZN(n4991) );
  NAND2_X1 U6520 ( .A1(n4984), .A2(n4991), .ZN(n4997) );
  NAND2_X1 U6521 ( .A1(n5427), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6522 ( .A1(n4993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4994) );
  XNOR2_X1 U6523 ( .A(n4994), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U6524 ( .A1(n5402), .A2(n9207), .ZN(n4995) );
  INV_X1 U6525 ( .A(n5686), .ZN(n6899) );
  NAND2_X1 U6526 ( .A1(n6899), .A2(n4998), .ZN(n4999) );
  NAND2_X1 U6527 ( .A1(n5000), .A2(n4999), .ZN(n5001) );
  XNOR2_X1 U6528 ( .A(n5001), .B(n5558), .ZN(n5002) );
  AOI22_X1 U6529 ( .A1(n9191), .A2(n5581), .B1(n6899), .B2(n5624), .ZN(n5003)
         );
  XNOR2_X1 U6530 ( .A(n5002), .B(n5003), .ZN(n6897) );
  NAND2_X1 U6531 ( .A1(n6896), .A2(n6897), .ZN(n5006) );
  INV_X1 U6532 ( .A(n5002), .ZN(n5004) );
  NAND2_X1 U6533 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NAND2_X1 U6534 ( .A1(n5006), .A2(n5005), .ZN(n7093) );
  INV_X1 U6535 ( .A(n7093), .ZN(n5036) );
  NAND2_X1 U6536 ( .A1(n5518), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U6537 ( .A1(n5007), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U6538 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5009) );
  NOR2_X1 U6539 ( .A1(n5041), .A2(n5009), .ZN(n7099) );
  NAND2_X1 U6540 ( .A1(n5666), .A2(n7099), .ZN(n5012) );
  INV_X2 U6541 ( .A(n5783), .ZN(n6586) );
  NAND2_X1 U6542 ( .A1(n6586), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5011) );
  NAND4_X1 U6543 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n9190)
         );
  NAND2_X1 U6544 ( .A1(n9190), .A2(n5262), .ZN(n5033) );
  NAND2_X1 U6545 ( .A1(n5427), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6546 ( .A1(n5016), .A2(n5015), .ZN(n5020) );
  INV_X1 U6547 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6548 ( .A1(n5018), .A2(SI_3_), .ZN(n5019) );
  NAND2_X1 U6549 ( .A1(n5020), .A2(n5019), .ZN(n5048) );
  INV_X1 U6550 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6385) );
  INV_X1 U6551 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6372) );
  XNOR2_X1 U6552 ( .A(n5049), .B(SI_4_), .ZN(n5047) );
  XNOR2_X1 U6553 ( .A(n5048), .B(n5047), .ZN(n6384) );
  INV_X1 U6554 ( .A(n6384), .ZN(n5021) );
  NAND2_X1 U6555 ( .A1(n4984), .A2(n5021), .ZN(n5030) );
  OR2_X1 U6556 ( .A1(n5022), .A2(n4875), .ZN(n5023) );
  AND2_X1 U6557 ( .A1(n5024), .A2(n5023), .ZN(n5026) );
  INV_X1 U6558 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6559 ( .A1(n5026), .A2(n5025), .ZN(n5054) );
  INV_X1 U6560 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6561 ( .A1(n5027), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5028) );
  AND2_X1 U6562 ( .A1(n5054), .A2(n5028), .ZN(n6623) );
  NAND2_X1 U6563 ( .A1(n5402), .A2(n6623), .ZN(n5029) );
  NAND2_X1 U6564 ( .A1(n6909), .A2(n4998), .ZN(n5032) );
  NAND2_X1 U6565 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  XNOR2_X1 U6566 ( .A(n5034), .B(n5627), .ZN(n5038) );
  AOI22_X1 U6567 ( .A1(n9190), .A2(n5581), .B1(n6909), .B2(n5624), .ZN(n5037)
         );
  XNOR2_X1 U6568 ( .A(n5038), .B(n5037), .ZN(n7096) );
  INV_X1 U6569 ( .A(n7096), .ZN(n5035) );
  NAND2_X1 U6570 ( .A1(n5518), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6571 ( .A1(n6587), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U6572 ( .A1(n5041), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5042) );
  NOR2_X1 U6573 ( .A1(n5062), .A2(n5042), .ZN(n7202) );
  NAND2_X1 U6574 ( .A1(n5666), .A2(n7202), .ZN(n5044) );
  NAND2_X1 U6575 ( .A1(n6586), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6576 ( .A1(n5048), .A2(n5047), .ZN(n5052) );
  INV_X1 U6577 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6578 ( .A1(n5050), .A2(SI_4_), .ZN(n5051) );
  INV_X1 U6579 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6386) );
  INV_X1 U6580 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5053) );
  XNOR2_X1 U6581 ( .A(n5072), .B(SI_5_), .ZN(n5070) );
  XNOR2_X1 U6582 ( .A(n5071), .B(n5070), .ZN(n6387) );
  NAND2_X1 U6583 ( .A1(n7890), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6584 ( .A1(n5054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U6585 ( .A(n5055), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U6586 ( .A1(n5402), .A2(n9234), .ZN(n5056) );
  OAI211_X1 U6587 ( .C1(n5086), .C2(n6387), .A(n5057), .B(n5056), .ZN(n7203)
         );
  OAI22_X1 U6588 ( .A1(n7021), .A2(n5556), .B1(n9817), .B2(n5557), .ZN(n5058)
         );
  XNOR2_X1 U6589 ( .A(n5058), .B(n5558), .ZN(n5061) );
  OAI22_X1 U6590 ( .A1(n7021), .A2(n5060), .B1(n9817), .B2(n5556), .ZN(n7130)
         );
  NAND2_X1 U6591 ( .A1(n5518), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6592 ( .A1(n6587), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5066) );
  NOR2_X1 U6593 ( .A1(n5062), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5063) );
  NOR2_X1 U6594 ( .A1(n5095), .A2(n5063), .ZN(n9801) );
  NAND2_X1 U6595 ( .A1(n5666), .A2(n9801), .ZN(n5065) );
  NAND2_X1 U6596 ( .A1(n6586), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6597 ( .A1(n5068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5069) );
  XNOR2_X1 U6598 ( .A(n5069), .B(n4865), .ZN(n9244) );
  INV_X1 U6599 ( .A(n5072), .ZN(n5073) );
  NAND2_X1 U6600 ( .A1(n5073), .A2(SI_5_), .ZN(n5074) );
  XNOR2_X1 U6601 ( .A(n5085), .B(SI_6_), .ZN(n5082) );
  XNOR2_X1 U6602 ( .A(n5084), .B(n5082), .ZN(n6376) );
  INV_X4 U6603 ( .A(n5086), .ZN(n7889) );
  NAND2_X1 U6604 ( .A1(n6376), .A2(n7889), .ZN(n5077) );
  NAND2_X1 U6605 ( .A1(n5427), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5076) );
  OAI211_X1 U6606 ( .C1(n6568), .C2(n9244), .A(n5077), .B(n5076), .ZN(n9802)
         );
  OAI22_X1 U6607 ( .A1(n7131), .A2(n5556), .B1(n7373), .B2(n5557), .ZN(n5078)
         );
  XNOR2_X1 U6608 ( .A(n5078), .B(n5558), .ZN(n7246) );
  OAI22_X1 U6609 ( .A1(n7131), .A2(n5060), .B1(n7373), .B2(n5556), .ZN(n7245)
         );
  OR2_X1 U6610 ( .A1(n7246), .A2(n7245), .ZN(n5079) );
  NAND2_X1 U6611 ( .A1(n7246), .A2(n7245), .ZN(n5080) );
  NAND2_X1 U6612 ( .A1(n5081), .A2(n5080), .ZN(n6352) );
  INV_X1 U6613 ( .A(n5082), .ZN(n5083) );
  XNOR2_X1 U6614 ( .A(n5112), .B(SI_7_), .ZN(n5109) );
  XNOR2_X1 U6615 ( .A(n5111), .B(n5109), .ZN(n6388) );
  NAND2_X1 U6616 ( .A1(n6388), .A2(n7889), .ZN(n5094) );
  NAND2_X1 U6617 ( .A1(n5088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  MUX2_X1 U6618 ( .A(n5090), .B(P1_IR_REG_31__SCAN_IN), .S(n5089), .Z(n5092)
         );
  NOR2_X1 U6619 ( .A1(n5088), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5177) );
  INV_X1 U6620 ( .A(n5177), .ZN(n5091) );
  NAND2_X1 U6621 ( .A1(n5092), .A2(n5091), .ZN(n6629) );
  INV_X1 U6622 ( .A(n6629), .ZN(n9261) );
  AOI22_X1 U6623 ( .A1(n7890), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5402), .B2(
        n9261), .ZN(n5093) );
  NAND2_X1 U6624 ( .A1(n5518), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6625 ( .A1(n6587), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6626 ( .A1(n5095), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5146) );
  OAI21_X1 U6627 ( .B1(n5095), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5146), .ZN(
        n6356) );
  INV_X1 U6628 ( .A(n6356), .ZN(n7187) );
  NAND2_X1 U6629 ( .A1(n5666), .A2(n7187), .ZN(n5097) );
  NAND2_X1 U6630 ( .A1(n6586), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5096) );
  NAND4_X1 U6631 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n9187)
         );
  NAND2_X1 U6632 ( .A1(n9187), .A2(n5262), .ZN(n5100) );
  OAI21_X1 U6633 ( .B1(n9825), .B2(n5557), .A(n5100), .ZN(n5101) );
  XNOR2_X1 U6634 ( .A(n5101), .B(n5627), .ZN(n5104) );
  OR2_X1 U6635 ( .A1(n9825), .A2(n5556), .ZN(n5103) );
  NAND2_X1 U6636 ( .A1(n9187), .A2(n5581), .ZN(n5102) );
  AND2_X1 U6637 ( .A1(n5103), .A2(n5102), .ZN(n5105) );
  NAND2_X1 U6638 ( .A1(n5104), .A2(n5105), .ZN(n6350) );
  INV_X1 U6639 ( .A(n5104), .ZN(n5107) );
  INV_X1 U6640 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6641 ( .A1(n5107), .A2(n5106), .ZN(n6351) );
  INV_X1 U6642 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6643 ( .A1(n5112), .A2(SI_7_), .ZN(n5113) );
  INV_X1 U6644 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5114) );
  INV_X1 U6645 ( .A(SI_8_), .ZN(n5115) );
  NAND2_X1 U6646 ( .A1(n5116), .A2(n5115), .ZN(n5119) );
  INV_X1 U6647 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6648 ( .A1(n5117), .A2(SI_8_), .ZN(n5118) );
  NAND2_X1 U6649 ( .A1(n5119), .A2(n5118), .ZN(n5141) );
  INV_X1 U6650 ( .A(SI_9_), .ZN(n5120) );
  NAND2_X1 U6651 ( .A1(n5121), .A2(n5120), .ZN(n5161) );
  INV_X1 U6652 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6653 ( .A1(n5122), .A2(SI_9_), .ZN(n5123) );
  XNOR2_X1 U6654 ( .A(n5160), .B(n4839), .ZN(n6407) );
  NAND2_X1 U6655 ( .A1(n6407), .A2(n7889), .ZN(n5128) );
  OR2_X1 U6656 ( .A1(n5177), .A2(n4875), .ZN(n5143) );
  INV_X1 U6657 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6658 ( .A1(n5143), .A2(n5124), .ZN(n5125) );
  NAND2_X1 U6659 ( .A1(n5125), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6660 ( .A(n5126), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9300) );
  AOI22_X1 U6661 ( .A1(n5427), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5402), .B2(
        n9300), .ZN(n5127) );
  NAND2_X1 U6662 ( .A1(n5128), .A2(n5127), .ZN(n7527) );
  NAND2_X1 U6663 ( .A1(n7527), .A2(n4998), .ZN(n5137) );
  NAND2_X1 U6664 ( .A1(n5518), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6665 ( .A1(n6587), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5134) );
  INV_X1 U6666 ( .A(n5146), .ZN(n5129) );
  AOI21_X1 U6667 ( .B1(n5129), .B2(P1_REG3_REG_8__SCAN_IN), .A(
        P1_REG3_REG_9__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6668 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n5130) );
  NOR2_X1 U6669 ( .A1(n5146), .A2(n5130), .ZN(n5197) );
  OR2_X1 U6670 ( .A1(n5131), .A2(n5197), .ZN(n7521) );
  INV_X1 U6671 ( .A(n7521), .ZN(n7279) );
  NAND2_X1 U6672 ( .A1(n5666), .A2(n7279), .ZN(n5133) );
  NAND2_X1 U6673 ( .A1(n6586), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6674 ( .A1(n9185), .A2(n5262), .ZN(n5136) );
  NAND2_X1 U6675 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  XNOR2_X1 U6676 ( .A(n5138), .B(n5627), .ZN(n7518) );
  NAND2_X1 U6677 ( .A1(n7527), .A2(n5624), .ZN(n5140) );
  NAND2_X1 U6678 ( .A1(n9185), .A2(n5581), .ZN(n5139) );
  AND2_X1 U6679 ( .A1(n5140), .A2(n5139), .ZN(n7517) );
  XNOR2_X1 U6680 ( .A(n5142), .B(n5141), .ZN(n6392) );
  NAND2_X1 U6681 ( .A1(n6392), .A2(n7889), .ZN(n5145) );
  XNOR2_X1 U6682 ( .A(n5143), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9274) );
  AOI22_X1 U6683 ( .A1(n5427), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5402), .B2(
        n9274), .ZN(n5144) );
  NAND2_X1 U6684 ( .A1(n6587), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6685 ( .A1(n5518), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5149) );
  XNOR2_X1 U6686 ( .A(n5146), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U6687 ( .A1(n5666), .A2(n7481), .ZN(n5148) );
  NAND2_X1 U6688 ( .A1(n6586), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5147) );
  NAND4_X1 U6689 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n9186)
         );
  INV_X1 U6690 ( .A(n9186), .ZN(n7524) );
  OAI22_X1 U6691 ( .A1(n7476), .A2(n5557), .B1(n7524), .B2(n5556), .ZN(n5151)
         );
  XNOR2_X1 U6692 ( .A(n5151), .B(n5627), .ZN(n7472) );
  OR2_X1 U6693 ( .A1(n7476), .A2(n5556), .ZN(n5153) );
  NAND2_X1 U6694 ( .A1(n9186), .A2(n5581), .ZN(n5152) );
  OAI22_X1 U6695 ( .A1(n7518), .A2(n7517), .B1(n7472), .B2(n7474), .ZN(n5159)
         );
  INV_X1 U6696 ( .A(n7472), .ZN(n7516) );
  INV_X1 U6697 ( .A(n7474), .ZN(n5154) );
  INV_X1 U6698 ( .A(n7517), .ZN(n5155) );
  OAI21_X1 U6699 ( .B1(n7516), .B2(n5154), .A(n5155), .ZN(n5157) );
  NOR2_X1 U6700 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  AOI22_X1 U6701 ( .A1(n5157), .A2(n7518), .B1(n7472), .B2(n5156), .ZN(n5158)
         );
  NAND2_X1 U6702 ( .A1(n5160), .A2(n4839), .ZN(n5162) );
  INV_X1 U6703 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5163) );
  MUX2_X1 U6704 ( .A(n6413), .B(n5163), .S(n6361), .Z(n5164) );
  XNOR2_X1 U6705 ( .A(n5164), .B(SI_10_), .ZN(n5192) );
  INV_X1 U6706 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6707 ( .A1(n5165), .A2(SI_10_), .ZN(n5166) );
  INV_X1 U6708 ( .A(n5174), .ZN(n5172) );
  MUX2_X1 U6709 ( .A(n6506), .B(n10128), .S(n6361), .Z(n5168) );
  NAND2_X1 U6710 ( .A1(n5168), .A2(n5167), .ZN(n5217) );
  INV_X1 U6711 ( .A(n5168), .ZN(n5169) );
  NAND2_X1 U6712 ( .A1(n5169), .A2(SI_11_), .ZN(n5170) );
  NAND2_X1 U6713 ( .A1(n5217), .A2(n5170), .ZN(n5173) );
  NAND2_X1 U6714 ( .A1(n5172), .A2(n5171), .ZN(n5218) );
  NAND2_X1 U6715 ( .A1(n5174), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6716 ( .A1(n5218), .A2(n5175), .ZN(n6505) );
  NAND2_X1 U6717 ( .A1(n6505), .A2(n7889), .ZN(n5180) );
  NOR2_X1 U6718 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5176) );
  NAND2_X1 U6719 ( .A1(n5177), .A2(n5176), .ZN(n5193) );
  NAND2_X1 U6720 ( .A1(n5220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5178) );
  XNOR2_X1 U6721 ( .A(n5178), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U6722 ( .A1(n5427), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5402), .B2(
        n9695), .ZN(n5179) );
  NAND2_X1 U6723 ( .A1(n9838), .A2(n4998), .ZN(n5188) );
  NAND2_X1 U6724 ( .A1(n6587), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6725 ( .A1(n5518), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6726 ( .A1(n6586), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6727 ( .A1(n5197), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6728 ( .A1(n5199), .A2(n5181), .ZN(n5182) );
  NAND2_X1 U6729 ( .A1(n5224), .A2(n5182), .ZN(n9677) );
  INV_X1 U6730 ( .A(n9677), .ZN(n7303) );
  NAND2_X1 U6731 ( .A1(n5666), .A2(n7303), .ZN(n5183) );
  NAND2_X1 U6732 ( .A1(n9183), .A2(n5262), .ZN(n5187) );
  NAND2_X1 U6733 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  XNOR2_X1 U6734 ( .A(n5189), .B(n5558), .ZN(n9665) );
  NAND2_X1 U6735 ( .A1(n9838), .A2(n5624), .ZN(n5191) );
  NAND2_X1 U6736 ( .A1(n9183), .A2(n5581), .ZN(n5190) );
  NAND2_X1 U6737 ( .A1(n5191), .A2(n5190), .ZN(n9666) );
  NAND2_X1 U6738 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  INV_X1 U6739 ( .A(n9664), .ZN(n5209) );
  NAND2_X1 U6740 ( .A1(n6409), .A2(n7889), .ZN(n5196) );
  NAND2_X1 U6741 ( .A1(n5193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6742 ( .A(n5194), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9651) );
  AOI22_X1 U6743 ( .A1(n5427), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5402), .B2(
        n9651), .ZN(n5195) );
  NAND2_X1 U6744 ( .A1(n5196), .A2(n5195), .ZN(n7318) );
  NAND2_X1 U6745 ( .A1(n7318), .A2(n4998), .ZN(n5205) );
  OR2_X1 U6746 ( .A1(n5197), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5198) );
  AND2_X1 U6747 ( .A1(n5199), .A2(n5198), .ZN(n7583) );
  NAND2_X1 U6748 ( .A1(n5666), .A2(n7583), .ZN(n5203) );
  NAND2_X1 U6749 ( .A1(n6587), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6750 ( .A1(n6586), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6751 ( .A1(n5518), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5200) );
  INV_X1 U6752 ( .A(n9663), .ZN(n9184) );
  NAND2_X1 U6753 ( .A1(n9184), .A2(n5262), .ZN(n5204) );
  NAND2_X1 U6754 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  XNOR2_X1 U6755 ( .A(n5206), .B(n5627), .ZN(n9668) );
  NOR2_X1 U6756 ( .A1(n9663), .A2(n5060), .ZN(n5207) );
  AOI21_X1 U6757 ( .B1(n7318), .B2(n5604), .A(n5207), .ZN(n5211) );
  NOR2_X1 U6758 ( .A1(n9668), .A2(n5211), .ZN(n5208) );
  INV_X1 U6759 ( .A(n9668), .ZN(n5212) );
  INV_X1 U6760 ( .A(n5211), .ZN(n7581) );
  OAI21_X1 U6761 ( .B1(n5212), .B2(n7581), .A(n9666), .ZN(n5215) );
  INV_X1 U6762 ( .A(n9665), .ZN(n5214) );
  NOR2_X1 U6763 ( .A1(n9666), .A2(n7581), .ZN(n5213) );
  AOI22_X1 U6764 ( .A1(n5215), .A2(n5214), .B1(n9668), .B2(n5213), .ZN(n5216)
         );
  MUX2_X1 U6765 ( .A(n10132), .B(n5219), .S(n6361), .Z(n5241) );
  XNOR2_X1 U6766 ( .A(n5241), .B(SI_12_), .ZN(n5240) );
  XNOR2_X1 U6767 ( .A(n5245), .B(n5240), .ZN(n6642) );
  NAND2_X1 U6768 ( .A1(n6642), .A2(n7889), .ZN(n5222) );
  OAI21_X1 U6769 ( .B1(n5220), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6770 ( .A(n5247), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U6771 ( .A1(n5427), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5402), .B2(
        n9699), .ZN(n5221) );
  NAND2_X1 U6772 ( .A1(n7454), .A2(n4998), .ZN(n5231) );
  NAND2_X1 U6773 ( .A1(n6587), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6774 ( .A1(n6586), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5228) );
  AND2_X1 U6775 ( .A1(n5224), .A2(n5223), .ZN(n5225) );
  NOR2_X1 U6776 ( .A1(n5252), .A2(n5225), .ZN(n7612) );
  NAND2_X1 U6777 ( .A1(n5666), .A2(n7612), .ZN(n5227) );
  NAND2_X1 U6778 ( .A1(n5518), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5226) );
  INV_X1 U6779 ( .A(n9660), .ZN(n9182) );
  NAND2_X1 U6780 ( .A1(n9182), .A2(n5624), .ZN(n5230) );
  NAND2_X1 U6781 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  XNOR2_X1 U6782 ( .A(n5232), .B(n5627), .ZN(n5234) );
  NOR2_X1 U6783 ( .A1(n9660), .A2(n5060), .ZN(n5233) );
  AOI21_X1 U6784 ( .B1(n7454), .B2(n5604), .A(n5233), .ZN(n5235) );
  NAND2_X1 U6785 ( .A1(n5234), .A2(n5235), .ZN(n5239) );
  INV_X1 U6786 ( .A(n5234), .ZN(n5237) );
  INV_X1 U6787 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6788 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  AND2_X1 U6789 ( .A1(n5239), .A2(n5238), .ZN(n7607) );
  NAND2_X1 U6790 ( .A1(n7606), .A2(n5239), .ZN(n7676) );
  INV_X1 U6791 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6792 ( .A1(n5242), .A2(SI_12_), .ZN(n5243) );
  XNOR2_X1 U6793 ( .A(n5270), .B(SI_13_), .ZN(n5267) );
  XNOR2_X1 U6794 ( .A(n5269), .B(n5267), .ZN(n6677) );
  NAND2_X1 U6795 ( .A1(n6677), .A2(n7889), .ZN(n5251) );
  INV_X1 U6796 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6797 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  NAND2_X1 U6798 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6799 ( .A(n5249), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U6800 ( .A1(n5427), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5402), .B2(
        n9715), .ZN(n5250) );
  NAND2_X1 U6801 ( .A1(n7811), .A2(n4998), .ZN(n5259) );
  NAND2_X1 U6802 ( .A1(n5518), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6803 ( .A1(n6587), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5256) );
  NOR2_X1 U6804 ( .A1(n5252), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6805 ( .A1(n5666), .A2(n4861), .ZN(n5255) );
  NAND2_X1 U6806 ( .A1(n6586), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6807 ( .A1(n9181), .A2(n5624), .ZN(n5258) );
  NAND2_X1 U6808 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  XNOR2_X1 U6809 ( .A(n5260), .B(n5558), .ZN(n5263) );
  NOR2_X1 U6810 ( .A1(n7810), .A2(n5060), .ZN(n5261) );
  AOI21_X1 U6811 ( .B1(n7811), .B2(n5262), .A(n5261), .ZN(n5264) );
  XNOR2_X1 U6812 ( .A(n5263), .B(n5264), .ZN(n7677) );
  NAND2_X1 U6813 ( .A1(n7676), .A2(n7677), .ZN(n7675) );
  INV_X1 U6814 ( .A(n5263), .ZN(n5265) );
  NAND2_X1 U6815 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6816 ( .A1(n7675), .A2(n5266), .ZN(n5290) );
  INV_X1 U6817 ( .A(n5267), .ZN(n5268) );
  INV_X1 U6818 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6819 ( .A1(n5274), .A2(SI_14_), .ZN(n5275) );
  NAND2_X1 U6820 ( .A1(n5295), .A2(n5275), .ZN(n5296) );
  XNOR2_X1 U6821 ( .A(n5297), .B(n5296), .ZN(n6740) );
  NAND2_X1 U6822 ( .A1(n6740), .A2(n7889), .ZN(n5279) );
  OR2_X1 U6823 ( .A1(n5276), .A2(n4875), .ZN(n5277) );
  XNOR2_X1 U6824 ( .A(n5277), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U6825 ( .A1(n5427), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5402), .B2(
        n9731), .ZN(n5278) );
  NAND2_X1 U6826 ( .A1(n7624), .A2(n4998), .ZN(n5287) );
  NAND2_X1 U6827 ( .A1(n6587), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6828 ( .A1(n5280), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6829 ( .A1(n5280), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5281) );
  AND2_X1 U6830 ( .A1(n5304), .A2(n5281), .ZN(n7745) );
  NAND2_X1 U6831 ( .A1(n5666), .A2(n7745), .ZN(n5284) );
  NAND2_X1 U6832 ( .A1(n5518), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6833 ( .A1(n6586), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5282) );
  NAND4_X1 U6834 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n9180)
         );
  NAND2_X1 U6835 ( .A1(n9180), .A2(n5624), .ZN(n5286) );
  NAND2_X1 U6836 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  XNOR2_X1 U6837 ( .A(n5288), .B(n5627), .ZN(n5289) );
  NAND2_X1 U6838 ( .A1(n7624), .A2(n5624), .ZN(n5292) );
  NAND2_X1 U6839 ( .A1(n9180), .A2(n5581), .ZN(n5291) );
  NAND2_X1 U6840 ( .A1(n5292), .A2(n5291), .ZN(n7740) );
  INV_X1 U6841 ( .A(n7740), .ZN(n5293) );
  INV_X1 U6842 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6820) );
  MUX2_X1 U6843 ( .A(n10006), .B(n6820), .S(n6361), .Z(n5322) );
  XNOR2_X1 U6844 ( .A(n5322), .B(SI_15_), .ZN(n5298) );
  XNOR2_X1 U6845 ( .A(n5324), .B(n5298), .ZN(n6819) );
  NAND2_X1 U6846 ( .A1(n6819), .A2(n7889), .ZN(n5302) );
  NAND2_X1 U6847 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  XNOR2_X1 U6848 ( .A(n5300), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U6849 ( .A1(n4992), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5402), .B2(
        n9754), .ZN(n5301) );
  NAND2_X1 U6850 ( .A1(n9167), .A2(n4998), .ZN(n5311) );
  NAND2_X1 U6851 ( .A1(n5518), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6852 ( .A1(n6587), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5308) );
  INV_X1 U6853 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6854 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  AND2_X1 U6855 ( .A1(n5332), .A2(n5305), .ZN(n9160) );
  NAND2_X1 U6856 ( .A1(n5666), .A2(n9160), .ZN(n5307) );
  NAND2_X1 U6857 ( .A1(n6586), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5306) );
  NAND4_X1 U6858 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n9179)
         );
  NAND2_X1 U6859 ( .A1(n9179), .A2(n5624), .ZN(n5310) );
  NAND2_X1 U6860 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  XNOR2_X1 U6861 ( .A(n5312), .B(n5627), .ZN(n5314) );
  INV_X1 U6862 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6863 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6864 ( .A1(n9167), .A2(n5624), .ZN(n5319) );
  NAND2_X1 U6865 ( .A1(n9179), .A2(n5581), .ZN(n5318) );
  NAND2_X1 U6866 ( .A1(n5319), .A2(n5318), .ZN(n9159) );
  INV_X1 U6867 ( .A(n9159), .ZN(n5320) );
  MUX2_X1 U6868 ( .A(n6947), .B(n10114), .S(n6361), .Z(n5346) );
  XNOR2_X1 U6869 ( .A(n5346), .B(SI_16_), .ZN(n5325) );
  XNOR2_X1 U6870 ( .A(n5350), .B(n5325), .ZN(n6946) );
  NAND2_X1 U6871 ( .A1(n6946), .A2(n7889), .ZN(n5330) );
  INV_X1 U6872 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6873 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5328) );
  XNOR2_X1 U6874 ( .A(n5328), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9309) );
  AOI22_X1 U6875 ( .A1(n4992), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5402), .B2(
        n9309), .ZN(n5329) );
  NAND2_X1 U6876 ( .A1(n7669), .A2(n4998), .ZN(n5339) );
  NAND2_X1 U6877 ( .A1(n5518), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6878 ( .A1(n6587), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5336) );
  INV_X1 U6879 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6880 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  AND2_X1 U6881 ( .A1(n5358), .A2(n5333), .ZN(n9091) );
  NAND2_X1 U6882 ( .A1(n5666), .A2(n9091), .ZN(n5335) );
  NAND2_X1 U6883 ( .A1(n6586), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6884 ( .A1(n9178), .A2(n5262), .ZN(n5338) );
  NAND2_X1 U6885 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  XNOR2_X1 U6886 ( .A(n5340), .B(n5558), .ZN(n5342) );
  NOR2_X1 U6887 ( .A1(n9099), .A2(n5060), .ZN(n5341) );
  AOI21_X1 U6888 ( .B1(n7669), .B2(n5604), .A(n5341), .ZN(n5343) );
  XNOR2_X1 U6889 ( .A(n5342), .B(n5343), .ZN(n9087) );
  NAND2_X1 U6890 ( .A1(n9086), .A2(n9087), .ZN(n9085) );
  INV_X1 U6891 ( .A(n5342), .ZN(n5344) );
  NAND2_X1 U6892 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U6893 ( .A1(n9085), .A2(n5345), .ZN(n9097) );
  NOR2_X1 U6894 ( .A1(n5347), .A2(SI_16_), .ZN(n5349) );
  NAND2_X1 U6895 ( .A1(n5347), .A2(SI_16_), .ZN(n5348) );
  MUX2_X1 U6896 ( .A(n7045), .B(n7047), .S(n6361), .Z(n5351) );
  INV_X1 U6897 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6898 ( .A1(n5352), .A2(SI_17_), .ZN(n5353) );
  NAND2_X1 U6899 ( .A1(n5376), .A2(n5353), .ZN(n5374) );
  XNOR2_X1 U6900 ( .A(n5375), .B(n5374), .ZN(n7044) );
  NAND2_X1 U6901 ( .A1(n7044), .A2(n7889), .ZN(n5356) );
  XNOR2_X1 U6902 ( .A(n5354), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U6903 ( .A1(n4992), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5402), .B2(
        n9778), .ZN(n5355) );
  NAND2_X1 U6904 ( .A1(n9581), .A2(n4998), .ZN(n5365) );
  NAND2_X1 U6905 ( .A1(n6587), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5363) );
  INV_X1 U6906 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5357) );
  AND2_X1 U6907 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  NOR2_X1 U6908 ( .A1(n5405), .A2(n5359), .ZN(n9103) );
  NAND2_X1 U6909 ( .A1(n5666), .A2(n9103), .ZN(n5362) );
  NAND2_X1 U6910 ( .A1(n5518), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6911 ( .A1(n6586), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5360) );
  NAND4_X1 U6912 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n9177)
         );
  NAND2_X1 U6913 ( .A1(n9177), .A2(n5604), .ZN(n5364) );
  NAND2_X1 U6914 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  XNOR2_X1 U6915 ( .A(n5366), .B(n5558), .ZN(n5369) );
  NAND2_X1 U6916 ( .A1(n9581), .A2(n5624), .ZN(n5368) );
  NAND2_X1 U6917 ( .A1(n9177), .A2(n5581), .ZN(n5367) );
  NAND2_X1 U6918 ( .A1(n5368), .A2(n5367), .ZN(n5370) );
  NAND2_X1 U6919 ( .A1(n5369), .A2(n5370), .ZN(n9095) );
  NAND2_X1 U6920 ( .A1(n9097), .A2(n9095), .ZN(n5373) );
  INV_X1 U6921 ( .A(n5369), .ZN(n5372) );
  INV_X1 U6922 ( .A(n5370), .ZN(n5371) );
  NAND2_X1 U6923 ( .A1(n5372), .A2(n5371), .ZN(n9094) );
  MUX2_X1 U6924 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6361), .Z(n5378) );
  XNOR2_X1 U6925 ( .A(n5378), .B(n10061), .ZN(n5399) );
  INV_X1 U6926 ( .A(n5399), .ZN(n5380) );
  NAND2_X1 U6927 ( .A1(n5378), .A2(SI_18_), .ZN(n5379) );
  MUX2_X1 U6928 ( .A(n7264), .B(n10018), .S(n6361), .Z(n5382) );
  INV_X1 U6929 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6930 ( .A1(n5383), .A2(SI_19_), .ZN(n5384) );
  NAND2_X1 U6931 ( .A1(n5423), .A2(n5384), .ZN(n5424) );
  XNOR2_X1 U6932 ( .A(n5425), .B(n5424), .ZN(n7263) );
  NAND2_X1 U6933 ( .A1(n7263), .A2(n7889), .ZN(n5387) );
  AOI22_X1 U6934 ( .A1(n4992), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9321), .B2(
        n5402), .ZN(n5386) );
  NAND2_X1 U6935 ( .A1(n9492), .A2(n4998), .ZN(n5395) );
  NAND2_X1 U6936 ( .A1(n5405), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5406) );
  INV_X1 U6937 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6938 ( .A1(n5406), .A2(n5388), .ZN(n5389) );
  AND2_X1 U6939 ( .A1(n5430), .A2(n5389), .ZN(n9493) );
  NAND2_X1 U6940 ( .A1(n9493), .A2(n5666), .ZN(n5393) );
  NAND2_X1 U6941 ( .A1(n6587), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6942 ( .A1(n6586), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6943 ( .A1(n5518), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5390) );
  NAND4_X1 U6944 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n9175)
         );
  NAND2_X1 U6945 ( .A1(n9175), .A2(n5624), .ZN(n5394) );
  NAND2_X1 U6946 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  XNOR2_X1 U6947 ( .A(n5396), .B(n5558), .ZN(n5418) );
  NAND2_X1 U6948 ( .A1(n9492), .A2(n5624), .ZN(n5398) );
  NAND2_X1 U6949 ( .A1(n9175), .A2(n5581), .ZN(n5397) );
  NAND2_X1 U6950 ( .A1(n5398), .A2(n5397), .ZN(n9060) );
  XNOR2_X1 U6951 ( .A(n5400), .B(n5399), .ZN(n7101) );
  NAND2_X1 U6952 ( .A1(n7101), .A2(n7889), .ZN(n5404) );
  XNOR2_X1 U6953 ( .A(n5401), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9313) );
  AOI22_X1 U6954 ( .A1(n7890), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5402), .B2(
        n9313), .ZN(n5403) );
  NAND2_X1 U6955 ( .A1(n9511), .A2(n5624), .ZN(n5413) );
  NAND2_X1 U6956 ( .A1(n6587), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6957 ( .A1(n5518), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6958 ( .A1(n5405), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5407) );
  AND2_X1 U6959 ( .A1(n5407), .A2(n5406), .ZN(n9513) );
  NAND2_X1 U6960 ( .A1(n5666), .A2(n9513), .ZN(n5409) );
  NAND2_X1 U6961 ( .A1(n6586), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5408) );
  NAND4_X1 U6962 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n9176)
         );
  NAND2_X1 U6963 ( .A1(n9176), .A2(n5581), .ZN(n5412) );
  NAND2_X1 U6964 ( .A1(n5413), .A2(n5412), .ZN(n9139) );
  NAND2_X1 U6965 ( .A1(n9511), .A2(n4998), .ZN(n5415) );
  NAND2_X1 U6966 ( .A1(n9176), .A2(n5624), .ZN(n5414) );
  NAND2_X1 U6967 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  XNOR2_X1 U6968 ( .A(n5416), .B(n5558), .ZN(n5419) );
  AOI22_X1 U6969 ( .A1(n5418), .A2(n9060), .B1(n9139), .B2(n5419), .ZN(n5417)
         );
  INV_X1 U6970 ( .A(n5418), .ZN(n9061) );
  OAI21_X1 U6971 ( .B1(n5419), .B2(n9139), .A(n9060), .ZN(n5421) );
  NOR2_X1 U6972 ( .A1(n9060), .A2(n9139), .ZN(n5420) );
  INV_X1 U6973 ( .A(n5419), .ZN(n9059) );
  AOI22_X1 U6974 ( .A1(n9061), .A2(n5421), .B1(n5420), .B2(n9059), .ZN(n5422)
         );
  MUX2_X1 U6975 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6361), .Z(n5440) );
  XNOR2_X1 U6976 ( .A(n5440), .B(n5442), .ZN(n5426) );
  NAND2_X1 U6977 ( .A1(n7325), .A2(n7889), .ZN(n5429) );
  NAND2_X1 U6978 ( .A1(n5427), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6979 ( .A1(n5741), .A2(n4998), .ZN(n5435) );
  INV_X1 U6980 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9122) );
  AND2_X1 U6981 ( .A1(n5430), .A2(n9122), .ZN(n5431) );
  OR2_X1 U6982 ( .A1(n5431), .A2(n5447), .ZN(n9478) );
  INV_X1 U6983 ( .A(n5666), .ZN(n5451) );
  AOI22_X1 U6984 ( .A1(n6586), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6587), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6985 ( .A1(n5518), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5432) );
  OAI211_X1 U6986 ( .C1(n9478), .C2(n5451), .A(n5433), .B(n5432), .ZN(n9065)
         );
  NAND2_X1 U6987 ( .A1(n9065), .A2(n5262), .ZN(n5434) );
  NAND2_X1 U6988 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  XNOR2_X1 U6989 ( .A(n5436), .B(n5627), .ZN(n9118) );
  AND2_X1 U6990 ( .A1(n9065), .A2(n5581), .ZN(n5437) );
  INV_X1 U6991 ( .A(n9118), .ZN(n5439) );
  INV_X1 U6992 ( .A(n9117), .ZN(n5438) );
  INV_X1 U6993 ( .A(n5440), .ZN(n5441) );
  MUX2_X1 U6994 ( .A(n7430), .B(n7421), .S(n6361), .Z(n5460) );
  XNOR2_X1 U6995 ( .A(n5460), .B(SI_21_), .ZN(n5444) );
  XNOR2_X1 U6996 ( .A(n5464), .B(n5444), .ZN(n7420) );
  NAND2_X1 U6997 ( .A1(n7420), .A2(n7889), .ZN(n5446) );
  NAND2_X1 U6998 ( .A1(n7890), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6999 ( .A1(n9562), .A2(n4998), .ZN(n5453) );
  OR2_X1 U7000 ( .A1(n5447), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7001 ( .A1(n5448), .A2(n5471), .ZN(n9461) );
  AOI22_X1 U7002 ( .A1(n6586), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n6587), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7003 ( .A1(n5518), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U7004 ( .C1(n9461), .C2(n5451), .A(n5450), .B(n5449), .ZN(n9174)
         );
  NAND2_X1 U7005 ( .A1(n9174), .A2(n5624), .ZN(n5452) );
  NAND2_X1 U7006 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  XNOR2_X1 U7007 ( .A(n5454), .B(n5627), .ZN(n5457) );
  AND2_X1 U7008 ( .A1(n9174), .A2(n5581), .ZN(n5455) );
  AOI21_X1 U7009 ( .B1(n9562), .B2(n5604), .A(n5455), .ZN(n5456) );
  XNOR2_X1 U7010 ( .A(n5457), .B(n5456), .ZN(n9072) );
  INV_X1 U7011 ( .A(n5456), .ZN(n5459) );
  INV_X1 U7012 ( .A(n5457), .ZN(n5458) );
  NOR2_X1 U7013 ( .A1(n5461), .A2(SI_21_), .ZN(n5463) );
  NAND2_X1 U7014 ( .A1(n5461), .A2(SI_21_), .ZN(n5462) );
  MUX2_X1 U7015 ( .A(n10005), .B(n7565), .S(n6361), .Z(n5466) );
  INV_X1 U7016 ( .A(SI_22_), .ZN(n5465) );
  NAND2_X1 U7017 ( .A1(n5466), .A2(n5465), .ZN(n5481) );
  INV_X1 U7018 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U7019 ( .A1(n5467), .A2(SI_22_), .ZN(n5468) );
  NAND2_X1 U7020 ( .A1(n5481), .A2(n5468), .ZN(n5482) );
  XNOR2_X1 U7021 ( .A(n5483), .B(n5482), .ZN(n7563) );
  NAND2_X1 U7022 ( .A1(n7563), .A2(n7889), .ZN(n5470) );
  NAND2_X1 U7023 ( .A1(n7890), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7024 ( .A1(n5518), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7025 ( .A1(n6587), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5474) );
  AOI21_X1 U7026 ( .B1(n10115), .B2(n5471), .A(n5494), .ZN(n9442) );
  NAND2_X1 U7027 ( .A1(n5666), .A2(n9442), .ZN(n5473) );
  NAND2_X1 U7028 ( .A1(n6586), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5472) );
  OAI22_X1 U7029 ( .A1(n9613), .A2(n5557), .B1(n9457), .B2(n5556), .ZN(n5476)
         );
  XNOR2_X1 U7030 ( .A(n5476), .B(n5627), .ZN(n5479) );
  OR2_X1 U7031 ( .A1(n9613), .A2(n5556), .ZN(n5478) );
  NAND2_X1 U7032 ( .A1(n9426), .A2(n5581), .ZN(n5477) );
  NAND2_X1 U7033 ( .A1(n5478), .A2(n5477), .ZN(n9128) );
  INV_X1 U7034 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5484) );
  MUX2_X1 U7035 ( .A(n10120), .B(n5484), .S(n6361), .Z(n5486) );
  INV_X1 U7036 ( .A(SI_23_), .ZN(n5485) );
  NAND2_X1 U7037 ( .A1(n5486), .A2(n5485), .ZN(n5510) );
  INV_X1 U7038 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U7039 ( .A1(n5487), .A2(SI_23_), .ZN(n5488) );
  NAND2_X1 U7040 ( .A1(n5490), .A2(n5489), .ZN(n5511) );
  OR2_X1 U7041 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U7042 ( .A1(n5511), .A2(n5491), .ZN(n7577) );
  NAND2_X1 U7043 ( .A1(n7577), .A2(n7889), .ZN(n5493) );
  NAND2_X1 U7044 ( .A1(n7890), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7045 ( .A1(n9550), .A2(n4998), .ZN(n5502) );
  NAND2_X1 U7046 ( .A1(n5518), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7047 ( .A1(n6587), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5499) );
  INV_X1 U7048 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5496) );
  INV_X1 U7049 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U7050 ( .A1(n5494), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5520) );
  AOI21_X1 U7051 ( .B1(n5496), .B2(n5495), .A(n5519), .ZN(n9417) );
  NAND2_X1 U7052 ( .A1(n5666), .A2(n9417), .ZN(n5498) );
  NAND2_X1 U7053 ( .A1(n6586), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U7054 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n9173)
         );
  NAND2_X1 U7055 ( .A1(n9173), .A2(n5624), .ZN(n5501) );
  NAND2_X1 U7056 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  XNOR2_X1 U7057 ( .A(n5503), .B(n5627), .ZN(n5505) );
  AND2_X1 U7058 ( .A1(n9173), .A2(n5581), .ZN(n5504) );
  AOI21_X1 U7059 ( .B1(n9550), .B2(n5604), .A(n5504), .ZN(n5506) );
  NAND2_X1 U7060 ( .A1(n5505), .A2(n5506), .ZN(n9107) );
  INV_X1 U7061 ( .A(n5505), .ZN(n5508) );
  INV_X1 U7062 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U7063 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  AND2_X1 U7064 ( .A1(n9107), .A2(n5509), .ZN(n9051) );
  NAND2_X1 U7065 ( .A1(n5511), .A2(n5510), .ZN(n5536) );
  INV_X1 U7066 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8067) );
  MUX2_X1 U7067 ( .A(n7658), .B(n8067), .S(n6361), .Z(n5513) );
  INV_X1 U7068 ( .A(SI_24_), .ZN(n5512) );
  NAND2_X1 U7069 ( .A1(n5513), .A2(n5512), .ZN(n5537) );
  INV_X1 U7070 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7071 ( .A1(n5514), .A2(SI_24_), .ZN(n5515) );
  XNOR2_X1 U7072 ( .A(n5536), .B(n5535), .ZN(n7657) );
  NAND2_X1 U7073 ( .A1(n7657), .A2(n7889), .ZN(n5517) );
  NAND2_X1 U7074 ( .A1(n7890), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7075 ( .A1(n5518), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7076 ( .A1(n6587), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5523) );
  INV_X1 U7077 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U7078 ( .A1(n5519), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5548) );
  INV_X1 U7079 ( .A(n5548), .ZN(n5550) );
  AOI21_X1 U7080 ( .B1(n9113), .B2(n5520), .A(n5550), .ZN(n9406) );
  NAND2_X1 U7081 ( .A1(n5666), .A2(n9406), .ZN(n5522) );
  NAND2_X1 U7082 ( .A1(n6586), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5521) );
  OAI22_X1 U7083 ( .A1(n9608), .A2(n5557), .B1(n9388), .B2(n5556), .ZN(n5525)
         );
  XNOR2_X1 U7084 ( .A(n5525), .B(n5627), .ZN(n5528) );
  OR2_X1 U7085 ( .A1(n9608), .A2(n5556), .ZN(n5527) );
  NAND2_X1 U7086 ( .A1(n9428), .A2(n5581), .ZN(n5526) );
  NAND2_X1 U7087 ( .A1(n5528), .A2(n5529), .ZN(n5533) );
  INV_X1 U7088 ( .A(n5528), .ZN(n5531) );
  INV_X1 U7089 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7090 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  NAND2_X1 U7091 ( .A1(n5533), .A2(n5532), .ZN(n9106) );
  AOI21_X1 U7092 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9110) );
  INV_X1 U7093 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7094 ( .A1(n5536), .A2(n5535), .ZN(n5538) );
  MUX2_X1 U7095 ( .A(n6166), .B(n7693), .S(n6361), .Z(n5540) );
  INV_X1 U7096 ( .A(SI_25_), .ZN(n5539) );
  NAND2_X1 U7097 ( .A1(n5540), .A2(n5539), .ZN(n5562) );
  INV_X1 U7098 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7099 ( .A1(n5541), .A2(SI_25_), .ZN(n5542) );
  OR2_X1 U7100 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  NAND2_X1 U7101 ( .A1(n5563), .A2(n5545), .ZN(n7691) );
  NAND2_X1 U7102 ( .A1(n7691), .A2(n7889), .ZN(n5547) );
  NAND2_X1 U7103 ( .A1(n7890), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7104 ( .A1(n6587), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7105 ( .A1(n5518), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5554) );
  INV_X1 U7106 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7107 ( .A1(n5549), .A2(n5548), .ZN(n5551) );
  NAND2_X1 U7108 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5550), .ZN(n5572) );
  AND2_X1 U7109 ( .A1(n5551), .A2(n5572), .ZN(n9391) );
  NAND2_X1 U7110 ( .A1(n5666), .A2(n9391), .ZN(n5553) );
  NAND2_X1 U7111 ( .A1(n5010), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5552) );
  OAI22_X1 U7112 ( .A1(n9394), .A2(n5557), .B1(n9366), .B2(n5556), .ZN(n5559)
         );
  XNOR2_X1 U7113 ( .A(n5559), .B(n5558), .ZN(n5561) );
  OAI22_X1 U7114 ( .A1(n9394), .A2(n5556), .B1(n9366), .B2(n5060), .ZN(n5560)
         );
  XNOR2_X1 U7115 ( .A(n5561), .B(n5560), .ZN(n9078) );
  NOR2_X1 U7116 ( .A1(n5561), .A2(n5560), .ZN(n9148) );
  INV_X1 U7117 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10076) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7730) );
  MUX2_X1 U7119 ( .A(n10076), .B(n7730), .S(n6361), .Z(n5565) );
  INV_X1 U7120 ( .A(SI_26_), .ZN(n5564) );
  NAND2_X1 U7121 ( .A1(n5565), .A2(n5564), .ZN(n5608) );
  INV_X1 U7122 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7123 ( .A1(n5566), .A2(SI_26_), .ZN(n5567) );
  NAND2_X1 U7124 ( .A1(n7729), .A2(n7889), .ZN(n5569) );
  NAND2_X1 U7125 ( .A1(n7890), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7126 ( .A1(n9374), .A2(n4998), .ZN(n5579) );
  NAND2_X1 U7127 ( .A1(n5518), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7128 ( .A1(n6587), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5576) );
  INV_X1 U7129 ( .A(n5572), .ZN(n5570) );
  NAND2_X1 U7130 ( .A1(n5570), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5618) );
  INV_X1 U7131 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7132 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  NAND2_X1 U7133 ( .A1(n5666), .A2(n9375), .ZN(n5575) );
  NAND2_X1 U7134 ( .A1(n6586), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5574) );
  NAND4_X1 U7135 ( .A1(n5577), .A2(n5576), .A3(n5575), .A4(n5574), .ZN(n9358)
         );
  NAND2_X1 U7136 ( .A1(n9358), .A2(n5624), .ZN(n5578) );
  NAND2_X1 U7137 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  XNOR2_X1 U7138 ( .A(n5580), .B(n5627), .ZN(n5583) );
  AND2_X1 U7139 ( .A1(n9358), .A2(n5581), .ZN(n5582) );
  AOI21_X1 U7140 ( .B1(n9374), .B2(n5604), .A(n5582), .ZN(n5584) );
  XNOR2_X1 U7141 ( .A(n5583), .B(n5584), .ZN(n9147) );
  INV_X1 U7142 ( .A(n5583), .ZN(n5586) );
  INV_X1 U7143 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7144 ( .A1(n5612), .A2(n5608), .ZN(n5593) );
  INV_X1 U7145 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8065) );
  MUX2_X1 U7146 ( .A(n10082), .B(n8065), .S(n6361), .Z(n5590) );
  INV_X1 U7147 ( .A(SI_27_), .ZN(n5589) );
  NAND2_X1 U7148 ( .A1(n5590), .A2(n5589), .ZN(n5607) );
  INV_X1 U7149 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7150 ( .A1(n5591), .A2(SI_27_), .ZN(n5609) );
  AND2_X1 U7151 ( .A1(n5607), .A2(n5609), .ZN(n5592) );
  NAND2_X1 U7152 ( .A1(n7734), .A2(n7889), .ZN(n5595) );
  NAND2_X1 U7153 ( .A1(n7890), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7154 ( .A1(n9531), .A2(n4998), .ZN(n5601) );
  NAND2_X1 U7155 ( .A1(n6587), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7156 ( .A1(n5518), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5598) );
  XNOR2_X1 U7157 ( .A(n5618), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U7158 ( .A1(n5666), .A2(n9350), .ZN(n5597) );
  NAND2_X1 U7159 ( .A1(n5010), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5596) );
  INV_X1 U7160 ( .A(n9367), .ZN(n9172) );
  NAND2_X1 U7161 ( .A1(n9172), .A2(n5624), .ZN(n5600) );
  NAND2_X1 U7162 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  XNOR2_X1 U7163 ( .A(n5602), .B(n5627), .ZN(n5606) );
  NOR2_X1 U7164 ( .A1(n9367), .A2(n5060), .ZN(n5603) );
  AOI21_X1 U7165 ( .B1(n9531), .B2(n5604), .A(n5603), .ZN(n5605) );
  NAND2_X1 U7166 ( .A1(n5606), .A2(n5605), .ZN(n5675) );
  OAI21_X1 U7167 ( .B1(n5606), .B2(n5605), .A(n5675), .ZN(n5791) );
  AND2_X1 U7168 ( .A1(n5608), .A2(n5607), .ZN(n5611) );
  INV_X1 U7169 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6198) );
  INV_X1 U7170 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U7171 ( .A(n5770), .B(SI_28_), .ZN(n5767) );
  NAND2_X1 U7172 ( .A1(n8078), .A2(n7889), .ZN(n5614) );
  NAND2_X1 U7173 ( .A1(n7890), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7174 ( .A1(n5748), .A2(n4998), .ZN(n5626) );
  NAND2_X1 U7175 ( .A1(n6587), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7176 ( .A1(n5518), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5622) );
  INV_X1 U7177 ( .A(n5618), .ZN(n5616) );
  AND2_X1 U7178 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n5615) );
  NAND2_X1 U7179 ( .A1(n5616), .A2(n5615), .ZN(n5665) );
  INV_X1 U7180 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5796) );
  INV_X1 U7181 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5617) );
  OAI21_X1 U7182 ( .B1(n5618), .B2(n5796), .A(n5617), .ZN(n5619) );
  NAND2_X1 U7183 ( .A1(n5666), .A2(n8056), .ZN(n5621) );
  NAND2_X1 U7184 ( .A1(n5010), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7185 ( .A1(n9359), .A2(n5624), .ZN(n5625) );
  NAND2_X1 U7186 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  XNOR2_X1 U7187 ( .A(n5628), .B(n5627), .ZN(n5631) );
  NAND2_X1 U7188 ( .A1(n5748), .A2(n5262), .ZN(n5629) );
  OAI21_X1 U7189 ( .B1(n5797), .B2(n5060), .A(n5629), .ZN(n5630) );
  XNOR2_X1 U7190 ( .A(n5631), .B(n5630), .ZN(n5654) );
  INV_X1 U7191 ( .A(n5654), .ZN(n5676) );
  NOR2_X1 U7192 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10125) );
  NOR4_X1 U7193 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5634) );
  NOR4_X1 U7194 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5633) );
  NOR4_X1 U7195 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5632) );
  NAND4_X1 U7196 ( .A1(n10125), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n5640)
         );
  NOR4_X1 U7197 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5638) );
  NOR4_X1 U7198 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5637) );
  NOR4_X1 U7199 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5636) );
  NOR4_X1 U7200 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5635) );
  NAND4_X1 U7201 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n5639)
         );
  NOR2_X1 U7202 ( .A1(n5640), .A2(n5639), .ZN(n5752) );
  NAND2_X1 U7203 ( .A1(n7692), .A2(P1_B_REG_SCAN_IN), .ZN(n5642) );
  MUX2_X1 U7204 ( .A(n5642), .B(P1_B_REG_SCAN_IN), .S(n5641), .Z(n5643) );
  OR2_X1 U7205 ( .A1(n5751), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5646) );
  INV_X1 U7206 ( .A(n7692), .ZN(n5644) );
  OR2_X1 U7207 ( .A1(n5645), .A2(n5644), .ZN(n9633) );
  NAND2_X1 U7208 ( .A1(n5646), .A2(n9633), .ZN(n5757) );
  INV_X1 U7209 ( .A(n5757), .ZN(n7003) );
  INV_X1 U7210 ( .A(n5641), .ZN(n8068) );
  NAND2_X1 U7211 ( .A1(n8068), .A2(n7731), .ZN(n9634) );
  OAI211_X1 U7212 ( .C1(n5752), .C2(n5751), .A(n7003), .B(n5761), .ZN(n5659)
         );
  INV_X1 U7213 ( .A(n5749), .ZN(n7030) );
  NAND2_X1 U7214 ( .A1(n5651), .A2(n7989), .ZN(n5671) );
  AND2_X1 U7215 ( .A1(n9831), .A2(n5671), .ZN(n5652) );
  NAND2_X1 U7216 ( .A1(n5653), .A2(n4852), .ZN(n5681) );
  NAND3_X1 U7217 ( .A1(n5795), .A2(n5654), .A3(n9151), .ZN(n5680) );
  INV_X1 U7218 ( .A(n5664), .ZN(n5655) );
  INV_X1 U7219 ( .A(n8046), .ZN(n7907) );
  NAND2_X1 U7220 ( .A1(n5749), .A2(n7907), .ZN(n7007) );
  OR2_X1 U7221 ( .A1(n5655), .A2(n7007), .ZN(n5657) );
  AND2_X1 U7222 ( .A1(n7905), .A2(n8046), .ZN(n9842) );
  NAND2_X1 U7223 ( .A1(n9842), .A2(n7993), .ZN(n5756) );
  INV_X1 U7224 ( .A(n5756), .ZN(n5656) );
  OR2_X1 U7225 ( .A1(n8046), .A2(P1_U3086), .ZN(n7327) );
  NAND2_X1 U7226 ( .A1(n9837), .A2(n7327), .ZN(n5658) );
  NAND2_X1 U7227 ( .A1(n5659), .A2(n5658), .ZN(n5661) );
  NOR2_X1 U7228 ( .A1(n5671), .A2(n7984), .ZN(n5754) );
  INV_X1 U7229 ( .A(n5754), .ZN(n5660) );
  NAND2_X1 U7230 ( .A1(n5661), .A2(n5660), .ZN(n6758) );
  OAI21_X1 U7231 ( .B1(n6758), .B2(n5662), .A(P1_STATE_REG_SCAN_IN), .ZN(n5663) );
  OR2_X1 U7232 ( .A1(n6567), .A2(P1_U3086), .ZN(n8054) );
  INV_X1 U7233 ( .A(n8056), .ZN(n5674) );
  NAND2_X1 U7234 ( .A1(n6587), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7235 ( .A1(n5518), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5669) );
  INV_X1 U7236 ( .A(n5665), .ZN(n9340) );
  NAND2_X1 U7237 ( .A1(n5666), .A2(n9340), .ZN(n5668) );
  NAND2_X1 U7238 ( .A1(n5010), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7239 ( .A1(n8041), .A2(n8080), .ZN(n9458) );
  INV_X1 U7240 ( .A(n8080), .ZN(n6773) );
  OR2_X1 U7241 ( .A1(n9367), .A2(n9456), .ZN(n5672) );
  OAI21_X1 U7242 ( .B1(n6846), .B2(n9458), .A(n5672), .ZN(n5747) );
  AOI22_X1 U7243 ( .A1(n9066), .A2(n5747), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5673) );
  OAI21_X1 U7244 ( .B1(n9678), .B2(n5674), .A(n5673), .ZN(n5678) );
  NOR3_X1 U7245 ( .A1(n5676), .A2(n9671), .A3(n5675), .ZN(n5677) );
  AOI211_X1 U7246 ( .C1(n5748), .C2(n9675), .A(n5678), .B(n5677), .ZN(n5679)
         );
  NAND3_X1 U7247 ( .A1(n5681), .A2(n5680), .A3(n5679), .ZN(P1_U3220) );
  INV_X1 U7248 ( .A(n9179), .ZN(n5734) );
  NAND2_X1 U7249 ( .A1(n7009), .A2(n7008), .ZN(n6838) );
  INV_X1 U7250 ( .A(n5683), .ZN(n6832) );
  NAND2_X1 U7251 ( .A1(n6832), .A2(n4369), .ZN(n5684) );
  INV_X2 U7252 ( .A(n6834), .ZN(n7910) );
  INV_X1 U7253 ( .A(n9192), .ZN(n6881) );
  NAND2_X1 U7254 ( .A1(n6881), .A2(n7910), .ZN(n5685) );
  XNOR2_X1 U7255 ( .A(n9191), .B(n5686), .ZN(n7990) );
  NAND2_X1 U7256 ( .A1(n6877), .A2(n7990), .ZN(n6876) );
  INV_X1 U7257 ( .A(n9191), .ZN(n6833) );
  NAND2_X1 U7258 ( .A1(n6833), .A2(n5686), .ZN(n5687) );
  NAND2_X1 U7259 ( .A1(n6876), .A2(n5687), .ZN(n6904) );
  XNOR2_X1 U7260 ( .A(n9190), .B(n7329), .ZN(n7997) );
  NAND2_X1 U7261 ( .A1(n6904), .A2(n7997), .ZN(n6903) );
  INV_X1 U7262 ( .A(n9190), .ZN(n7132) );
  NAND2_X1 U7263 ( .A1(n7132), .A2(n7329), .ZN(n5688) );
  NAND2_X1 U7264 ( .A1(n6903), .A2(n5688), .ZN(n7198) );
  NAND2_X1 U7265 ( .A1(n7021), .A2(n7203), .ZN(n7781) );
  INV_X1 U7266 ( .A(n7021), .ZN(n9189) );
  NAND2_X1 U7267 ( .A1(n9189), .A2(n9817), .ZN(n7917) );
  NAND2_X1 U7268 ( .A1(n7781), .A2(n7917), .ZN(n7996) );
  NAND2_X1 U7269 ( .A1(n7021), .A2(n9817), .ZN(n5689) );
  NAND2_X1 U7270 ( .A1(n7131), .A2(n9802), .ZN(n7919) );
  INV_X1 U7271 ( .A(n7131), .ZN(n9188) );
  NAND2_X1 U7272 ( .A1(n9188), .A2(n7373), .ZN(n7779) );
  NAND2_X1 U7273 ( .A1(n7919), .A2(n7779), .ZN(n7999) );
  NAND2_X1 U7274 ( .A1(n7131), .A2(n7373), .ZN(n5690) );
  XNOR2_X1 U7275 ( .A(n9187), .B(n9825), .ZN(n7178) );
  INV_X1 U7276 ( .A(n9187), .ZN(n7477) );
  NAND2_X1 U7277 ( .A1(n7476), .A2(n9186), .ZN(n7786) );
  NAND2_X1 U7278 ( .A1(n7786), .A2(n7789), .ZN(n7227) );
  NAND2_X1 U7279 ( .A1(n7224), .A2(n7227), .ZN(n7223) );
  NAND2_X1 U7280 ( .A1(n7476), .A2(n7524), .ZN(n5691) );
  OR2_X1 U7281 ( .A1(n7527), .A2(n7585), .ZN(n7798) );
  NAND2_X1 U7282 ( .A1(n7527), .A2(n7585), .ZN(n7795) );
  NAND2_X1 U7283 ( .A1(n7798), .A2(n7795), .ZN(n7281) );
  OR2_X1 U7284 ( .A1(n7527), .A2(n9185), .ZN(n5692) );
  OR2_X1 U7285 ( .A1(n7318), .A2(n9663), .ZN(n7922) );
  NAND2_X1 U7286 ( .A1(n7318), .A2(n9663), .ZN(n7799) );
  NAND2_X1 U7287 ( .A1(n7922), .A2(n7799), .ZN(n7312) );
  OR2_X1 U7288 ( .A1(n9838), .A2(n7610), .ZN(n7802) );
  NAND2_X1 U7289 ( .A1(n9838), .A2(n7610), .ZN(n7804) );
  NAND2_X1 U7290 ( .A1(n7802), .A2(n7804), .ZN(n8005) );
  NAND2_X1 U7291 ( .A1(n7291), .A2(n8005), .ZN(n7293) );
  INV_X1 U7292 ( .A(n9838), .ZN(n5693) );
  NAND2_X1 U7293 ( .A1(n5693), .A2(n7610), .ZN(n5694) );
  OR2_X1 U7294 ( .A1(n7454), .A2(n9660), .ZN(n7806) );
  NAND2_X1 U7295 ( .A1(n7454), .A2(n9660), .ZN(n7928) );
  NAND2_X1 U7296 ( .A1(n7806), .A2(n7928), .ZN(n7440) );
  NAND2_X1 U7297 ( .A1(n7439), .A2(n7440), .ZN(n7438) );
  NAND2_X1 U7298 ( .A1(n7438), .A2(n5696), .ZN(n7531) );
  OR2_X1 U7299 ( .A1(n7811), .A2(n7810), .ZN(n7931) );
  NAND2_X1 U7300 ( .A1(n7811), .A2(n7810), .ZN(n7929) );
  NAND2_X1 U7301 ( .A1(n7931), .A2(n7929), .ZN(n8010) );
  NAND2_X1 U7302 ( .A1(n7624), .A2(n9180), .ZN(n5699) );
  INV_X1 U7303 ( .A(n9180), .ZN(n7535) );
  OR2_X1 U7304 ( .A1(n7669), .A2(n9099), .ZN(n7939) );
  NAND2_X1 U7305 ( .A1(n7669), .A2(n9099), .ZN(n7938) );
  NAND2_X1 U7306 ( .A1(n7939), .A2(n7938), .ZN(n8015) );
  NAND2_X1 U7307 ( .A1(n9581), .A2(n9177), .ZN(n5702) );
  INV_X1 U7308 ( .A(n9581), .ZN(n9100) );
  INV_X1 U7309 ( .A(n9177), .ZN(n5738) );
  INV_X1 U7310 ( .A(n9500), .ZN(n5704) );
  NOR2_X1 U7311 ( .A1(n9511), .A2(n9176), .ZN(n5703) );
  INV_X1 U7312 ( .A(n9176), .ZN(n5739) );
  INV_X1 U7313 ( .A(n9175), .ZN(n7770) );
  NAND2_X1 U7314 ( .A1(n9622), .A2(n7770), .ZN(n5705) );
  OAI21_X1 U7315 ( .B1(n9485), .B2(n5706), .A(n5705), .ZN(n5707) );
  INV_X1 U7316 ( .A(n9065), .ZN(n9455) );
  INV_X1 U7317 ( .A(n9562), .ZN(n9465) );
  INV_X1 U7318 ( .A(n9174), .ZN(n5742) );
  NAND2_X1 U7319 ( .A1(n9613), .A2(n9457), .ZN(n5709) );
  NOR2_X1 U7320 ( .A1(n9550), .A2(n9173), .ZN(n5710) );
  NOR2_X1 U7321 ( .A1(n9394), .A2(n9366), .ZN(n5711) );
  INV_X1 U7322 ( .A(n9366), .ZN(n9112) );
  NOR2_X1 U7323 ( .A1(n9374), .A2(n9358), .ZN(n5713) );
  NAND2_X1 U7324 ( .A1(n9374), .A2(n9358), .ZN(n5712) );
  NAND2_X1 U7325 ( .A1(n9531), .A2(n9367), .ZN(n7876) );
  NAND2_X1 U7326 ( .A1(n9352), .A2(n9367), .ZN(n5714) );
  NAND2_X1 U7327 ( .A1(n5748), .A2(n5797), .ZN(n7877) );
  NAND2_X1 U7328 ( .A1(n4618), .A2(n4377), .ZN(n5766) );
  INV_X1 U7329 ( .A(n7984), .ZN(n5716) );
  NAND2_X1 U7330 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  AND2_X1 U7331 ( .A1(n5718), .A2(n7030), .ZN(n5719) );
  NAND2_X1 U7332 ( .A1(n8041), .A2(n7984), .ZN(n8050) );
  NAND2_X1 U7333 ( .A1(n5719), .A2(n8050), .ZN(n7622) );
  INV_X1 U7334 ( .A(n9842), .ZN(n5720) );
  NOR2_X1 U7335 ( .A1(n7009), .A2(n7029), .ZN(n7010) );
  NAND2_X1 U7336 ( .A1(n6832), .A2(n6843), .ZN(n5721) );
  INV_X1 U7337 ( .A(n7991), .ZN(n5722) );
  NAND2_X1 U7338 ( .A1(n6881), .A2(n6834), .ZN(n5723) );
  NOR2_X1 U7339 ( .A1(n9191), .A2(n5686), .ZN(n5724) );
  NAND2_X1 U7340 ( .A1(n9191), .A2(n5686), .ZN(n7914) );
  NAND2_X1 U7341 ( .A1(n9190), .A2(n7329), .ZN(n7916) );
  NAND2_X1 U7342 ( .A1(n6906), .A2(n7916), .ZN(n7775) );
  NAND2_X1 U7343 ( .A1(n7132), .A2(n6909), .ZN(n7780) );
  INV_X1 U7344 ( .A(n7996), .ZN(n5725) );
  NAND2_X1 U7345 ( .A1(n7776), .A2(n5725), .ZN(n5726) );
  NAND2_X1 U7346 ( .A1(n5726), .A2(n7917), .ZN(n7019) );
  NAND2_X1 U7347 ( .A1(n7798), .A2(n7786), .ZN(n7791) );
  INV_X1 U7348 ( .A(n9825), .ZN(n7188) );
  NAND2_X1 U7349 ( .A1(n7477), .A2(n7188), .ZN(n7229) );
  NAND2_X1 U7350 ( .A1(n7019), .A2(n8007), .ZN(n7924) );
  INV_X1 U7351 ( .A(n7919), .ZN(n5728) );
  INV_X1 U7352 ( .A(n7791), .ZN(n8002) );
  NAND2_X1 U7353 ( .A1(n9187), .A2(n9825), .ZN(n8000) );
  NAND3_X1 U7354 ( .A1(n8002), .A2(n8000), .A3(n7779), .ZN(n5727) );
  NAND2_X1 U7355 ( .A1(n8007), .A2(n5727), .ZN(n7921) );
  INV_X1 U7356 ( .A(n7799), .ZN(n5729) );
  NOR2_X1 U7357 ( .A1(n8005), .A2(n5729), .ZN(n5730) );
  INV_X1 U7358 ( .A(n7440), .ZN(n8008) );
  OR2_X1 U7359 ( .A1(n7624), .A2(n7535), .ZN(n7930) );
  NAND2_X1 U7360 ( .A1(n7624), .A2(n7535), .ZN(n7815) );
  NAND2_X1 U7361 ( .A1(n7930), .A2(n7815), .ZN(n7819) );
  INV_X1 U7362 ( .A(n7929), .ZN(n7616) );
  NOR2_X1 U7363 ( .A1(n7819), .A2(n7616), .ZN(n5733) );
  OR2_X1 U7364 ( .A1(n9167), .A2(n5734), .ZN(n7825) );
  NAND2_X1 U7365 ( .A1(n9167), .A2(n5734), .ZN(n7827) );
  NAND2_X1 U7366 ( .A1(n7825), .A2(n7827), .ZN(n7594) );
  INV_X1 U7367 ( .A(n7930), .ZN(n5735) );
  NOR2_X1 U7368 ( .A1(n7594), .A2(n5735), .ZN(n5736) );
  OR2_X1 U7369 ( .A1(n9581), .A2(n5738), .ZN(n7940) );
  NAND2_X1 U7370 ( .A1(n9581), .A2(n5738), .ZN(n7835) );
  OR2_X1 U7371 ( .A1(n9511), .A2(n5739), .ZN(n7842) );
  NAND2_X1 U7372 ( .A1(n9511), .A2(n5739), .ZN(n7844) );
  NAND2_X1 U7373 ( .A1(n7842), .A2(n7844), .ZN(n9502) );
  OR2_X1 U7374 ( .A1(n9492), .A2(n7770), .ZN(n7836) );
  NAND2_X1 U7375 ( .A1(n9492), .A2(n7770), .ZN(n7909) );
  NAND2_X1 U7376 ( .A1(n9487), .A2(n9486), .ZN(n5740) );
  NAND2_X1 U7377 ( .A1(n5741), .A2(n9455), .ZN(n7771) );
  NAND2_X1 U7378 ( .A1(n7839), .A2(n7771), .ZN(n9469) );
  XNOR2_X1 U7379 ( .A(n9562), .B(n5742), .ZN(n9449) );
  NAND2_X1 U7380 ( .A1(n9562), .A2(n5742), .ZN(n7841) );
  NAND2_X1 U7381 ( .A1(n7841), .A2(n7771), .ZN(n7848) );
  OR2_X1 U7382 ( .A1(n9562), .A2(n5742), .ZN(n7851) );
  NAND2_X1 U7383 ( .A1(n7848), .A2(n7851), .ZN(n7962) );
  INV_X1 U7384 ( .A(n9173), .ZN(n5743) );
  OR2_X1 U7385 ( .A1(n9550), .A2(n5743), .ZN(n7854) );
  NAND2_X1 U7386 ( .A1(n9550), .A2(n5743), .ZN(n9400) );
  NAND2_X1 U7387 ( .A1(n7854), .A2(n9400), .ZN(n9420) );
  NOR2_X1 U7388 ( .A1(n9441), .A2(n9457), .ZN(n9421) );
  NOR2_X1 U7389 ( .A1(n9420), .A2(n9421), .ZN(n5744) );
  OR2_X1 U7390 ( .A1(n9405), .A2(n9388), .ZN(n7950) );
  NAND2_X1 U7391 ( .A1(n9405), .A2(n9388), .ZN(n7964) );
  NAND2_X1 U7392 ( .A1(n7950), .A2(n7964), .ZN(n7860) );
  INV_X1 U7393 ( .A(n9400), .ZN(n7856) );
  NOR2_X1 U7394 ( .A1(n7860), .A2(n7856), .ZN(n5745) );
  OR2_X1 U7395 ( .A1(n9542), .A2(n9366), .ZN(n7952) );
  NAND2_X1 U7396 ( .A1(n9542), .A2(n9366), .ZN(n7965) );
  NAND2_X1 U7397 ( .A1(n7952), .A2(n7965), .ZN(n9385) );
  NAND2_X1 U7398 ( .A1(n9382), .A2(n7965), .ZN(n9364) );
  XNOR2_X1 U7399 ( .A(n9374), .B(n9358), .ZN(n9371) );
  NAND2_X1 U7400 ( .A1(n9364), .A2(n9371), .ZN(n9353) );
  INV_X1 U7401 ( .A(n9358), .ZN(n9387) );
  NAND2_X1 U7402 ( .A1(n9353), .A2(n9355), .ZN(n5746) );
  NAND2_X1 U7403 ( .A1(n5651), .A2(n9321), .ZN(n7986) );
  NAND2_X1 U7404 ( .A1(n7989), .A2(n7907), .ZN(n7768) );
  NAND2_X2 U7405 ( .A1(n7986), .A2(n7768), .ZN(n9504) );
  INV_X1 U7406 ( .A(n9550), .ZN(n9419) );
  AND2_X1 U7407 ( .A1(n7199), .A2(n9817), .ZN(n7200) );
  INV_X1 U7408 ( .A(n7527), .ZN(n9832) );
  INV_X1 U7409 ( .A(n7318), .ZN(n7586) );
  NAND2_X1 U7410 ( .A1(n7315), .A2(n7586), .ZN(n7316) );
  NAND2_X1 U7411 ( .A1(n9491), .A2(n9618), .ZN(n9475) );
  INV_X1 U7412 ( .A(n9509), .ZN(n9551) );
  OAI211_X1 U7413 ( .C1(n8058), .C2(n9348), .A(n9551), .B(n5777), .ZN(n8055)
         );
  NAND2_X1 U7414 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  AND2_X1 U7415 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  INV_X1 U7416 ( .A(n5759), .ZN(n5760) );
  NAND2_X1 U7417 ( .A1(n5760), .A2(n4843), .ZN(P1_U3550) );
  INV_X1 U7418 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7419 ( .A1(n5764), .A2(n4851), .ZN(P1_U3518) );
  NAND2_X1 U7420 ( .A1(n5748), .A2(n9359), .ZN(n5765) );
  NAND2_X1 U7421 ( .A1(n5766), .A2(n5765), .ZN(n5775) );
  NAND2_X1 U7422 ( .A1(n5768), .A2(n5767), .ZN(n5772) );
  INV_X1 U7423 ( .A(SI_28_), .ZN(n5769) );
  NAND2_X1 U7424 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  INV_X1 U7425 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8082) );
  INV_X1 U7426 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9991) );
  MUX2_X1 U7427 ( .A(n8082), .B(n9991), .S(n6361), .Z(n7751) );
  NAND2_X1 U7428 ( .A1(n8081), .A2(n7889), .ZN(n5774) );
  NAND2_X1 U7429 ( .A1(n7890), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7430 ( .A1(n5776), .A2(n6846), .ZN(n7869) );
  AND2_X2 U7431 ( .A1(n7975), .A2(n7869), .ZN(n8024) );
  AOI211_X1 U7432 ( .C1(n5776), .C2(n5777), .A(n9509), .B(n9333), .ZN(n9344)
         );
  INV_X1 U7433 ( .A(n9344), .ZN(n5787) );
  INV_X1 U7434 ( .A(n8024), .ZN(n5778) );
  NAND2_X1 U7435 ( .A1(n5779), .A2(n9504), .ZN(n5786) );
  INV_X1 U7436 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7437 ( .A1(n5518), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7438 ( .A1(n6587), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5780) );
  OAI211_X1 U7439 ( .C1(n5783), .C2(n5782), .A(n5781), .B(n5780), .ZN(n9171)
         );
  INV_X1 U7440 ( .A(n9681), .ZN(n6636) );
  AND2_X1 U7441 ( .A1(n6636), .A2(P1_B_REG_SCAN_IN), .ZN(n5784) );
  NOR2_X1 U7442 ( .A1(n9458), .A2(n5784), .ZN(n9328) );
  AOI22_X1 U7443 ( .A1(n9359), .A2(n9425), .B1(n9171), .B2(n9328), .ZN(n5785)
         );
  INV_X1 U7444 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5788) );
  INV_X1 U7445 ( .A(n5793), .ZN(n5794) );
  OAI21_X1 U7446 ( .B1(n5795), .B2(n5794), .A(n9151), .ZN(n5801) );
  NAND2_X1 U7447 ( .A1(n9066), .A2(n9425), .ZN(n9662) );
  NOR2_X1 U7448 ( .A1(n9662), .A2(n9387), .ZN(n5799) );
  NAND2_X1 U7449 ( .A1(n9066), .A2(n9427), .ZN(n9661) );
  OAI22_X1 U7450 ( .A1(n9661), .A2(n5797), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5796), .ZN(n5798) );
  AOI211_X1 U7451 ( .C1(n9350), .C2(n9161), .A(n5799), .B(n5798), .ZN(n5800)
         );
  NAND3_X1 U7452 ( .A1(n5801), .A2(n5800), .A3(n4844), .ZN(P1_U3214) );
  INV_X1 U7453 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5804) );
  NOR2_X1 U7454 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5816) );
  NOR2_X1 U7455 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5815) );
  NAND4_X1 U7456 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n5819)
         );
  NAND4_X1 U7457 ( .A1(n5965), .A2(n5951), .A3(n5817), .A4(n5949), .ZN(n5818)
         );
  NOR2_X2 U7458 ( .A1(n5819), .A2(n5818), .ZN(n5861) );
  NAND2_X2 U7459 ( .A1(n8296), .A2(n8295), .ZN(n5904) );
  NAND2_X1 U7460 ( .A1(n7657), .A2(n8298), .ZN(n5825) );
  OR2_X1 U7461 ( .A1(n8299), .A2(n7658), .ZN(n5824) );
  NAND2_X1 U7462 ( .A1(n5827), .A2(n5826), .ZN(n5943) );
  INV_X1 U7463 ( .A(n5943), .ZN(n5829) );
  NAND2_X1 U7464 ( .A1(n5829), .A2(n5828), .ZN(n5957) );
  INV_X1 U7465 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5843) );
  INV_X1 U7466 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7467 ( .A1(n6156), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7468 ( .A1(n6171), .A2(n5847), .ZN(n8750) );
  NAND2_X1 U7469 ( .A1(n5852), .A2(n5851), .ZN(n9037) );
  NAND2_X1 U7470 ( .A1(n8750), .A2(n6211), .ZN(n5860) );
  INV_X1 U7471 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U7472 ( .A1(n5930), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7473 ( .A1(n4734), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5856) );
  OAI211_X1 U7474 ( .C1(n10131), .C2(n4275), .A(n5857), .B(n5856), .ZN(n5858)
         );
  INV_X1 U7475 ( .A(n5858), .ZN(n5859) );
  NAND2_X1 U7476 ( .A1(n7263), .A2(n8298), .ZN(n5867) );
  NAND2_X1 U7477 ( .A1(n5950), .A2(n5861), .ZN(n6224) );
  AOI22_X1 U7478 ( .A1(n6113), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6270), .B2(
        n6112), .ZN(n5866) );
  NAND2_X1 U7479 ( .A1(n6118), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7480 ( .A1(n6127), .A2(n5868), .ZN(n8816) );
  NAND2_X1 U7481 ( .A1(n8816), .A2(n6211), .ZN(n5871) );
  AOI22_X1 U7482 ( .A1(n5930), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n4734), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7483 ( .A1(n5898), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5869) );
  INV_X1 U7484 ( .A(n8933), .ZN(n8944) );
  NAND2_X1 U7485 ( .A1(n5898), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5876) );
  INV_X1 U7486 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5872) );
  INV_X1 U7487 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8883) );
  OR2_X1 U7488 ( .A1(n5899), .A2(n8883), .ZN(n5873) );
  NAND2_X1 U7489 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5877) );
  MUX2_X1 U7490 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5877), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5880) );
  OR2_X1 U7491 ( .A1(n5905), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5881) );
  OAI211_X2 U7492 ( .C1(n6461), .C2(n8296), .A(n5882), .B(n5881), .ZN(n8884)
         );
  NAND2_X1 U7493 ( .A1(n5884), .A2(n5883), .ZN(n6232) );
  NAND2_X1 U7494 ( .A1(n5893), .A2(n8884), .ZN(n8325) );
  INV_X1 U7495 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5885) );
  INV_X1 U7496 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5886) );
  INV_X1 U7497 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7498 ( .A1(n5913), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5889) );
  INV_X1 U7499 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7500 ( .A1(n5899), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U7501 ( .A1(n8295), .A2(SI_0_), .ZN(n5892) );
  XNOR2_X1 U7502 ( .A(n5892), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9050) );
  MUX2_X1 U7503 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9050), .S(n8296), .Z(n6736) );
  NAND2_X1 U7504 ( .A1(n6415), .A2(n6736), .ZN(n8888) );
  NAND2_X1 U7505 ( .A1(n6231), .A2(n8888), .ZN(n5895) );
  NAND2_X1 U7506 ( .A1(n5884), .A2(n8884), .ZN(n5894) );
  NAND2_X1 U7507 ( .A1(n5895), .A2(n5894), .ZN(n6792) );
  INV_X1 U7508 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5896) );
  OR2_X1 U7509 ( .A1(n5897), .A2(n5896), .ZN(n5903) );
  INV_X1 U7510 ( .A(n8305), .ZN(n5898) );
  INV_X1 U7511 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6795) );
  OR2_X1 U7512 ( .A1(n5899), .A2(n6795), .ZN(n5901) );
  NAND2_X1 U7513 ( .A1(n5913), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5900) );
  OR2_X1 U7514 ( .A1(n5904), .A2(n6368), .ZN(n5909) );
  OR2_X1 U7515 ( .A1(n5905), .A2(n6367), .ZN(n5908) );
  OR2_X1 U7516 ( .A1(n8296), .A2(n6520), .ZN(n5907) );
  NAND2_X1 U7517 ( .A1(n5910), .A2(n6796), .ZN(n8331) );
  NAND2_X1 U7518 ( .A1(n6792), .A2(n6793), .ZN(n5912) );
  INV_X1 U7519 ( .A(n5910), .ZN(n6556) );
  NAND2_X1 U7520 ( .A1(n6556), .A2(n6796), .ZN(n5911) );
  NAND2_X1 U7521 ( .A1(n5912), .A2(n5911), .ZN(n6848) );
  INV_X1 U7522 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6852) );
  INV_X1 U7523 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7524 ( .A1(n6065), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7525 ( .A1(n4734), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7526 ( .A1(n5904), .A2(n6366), .ZN(n5925) );
  OR2_X1 U7527 ( .A1(n8299), .A2(n4397), .ZN(n5924) );
  NOR2_X1 U7528 ( .A1(n5918), .A2(n5849), .ZN(n5919) );
  MUX2_X1 U7529 ( .A(n5849), .B(n5919), .S(P2_IR_REG_3__SCAN_IN), .Z(n5920) );
  INV_X1 U7530 ( .A(n5920), .ZN(n5922) );
  INV_X1 U7531 ( .A(n5950), .ZN(n5921) );
  NAND2_X1 U7532 ( .A1(n5922), .A2(n5921), .ZN(n6478) );
  OR2_X1 U7533 ( .A1(n8296), .A2(n6478), .ZN(n5923) );
  AND3_X2 U7534 ( .A1(n5925), .A2(n5924), .A3(n5923), .ZN(n9877) );
  NAND2_X1 U7535 ( .A1(n8528), .A2(n9877), .ZN(n8340) );
  NAND2_X1 U7536 ( .A1(n6234), .A2(n8340), .ZN(n6849) );
  NAND2_X1 U7537 ( .A1(n6848), .A2(n6849), .ZN(n5929) );
  NAND2_X1 U7538 ( .A1(n5927), .A2(n9877), .ZN(n5928) );
  NAND2_X1 U7539 ( .A1(n5929), .A2(n5928), .ZN(n6742) );
  INV_X1 U7540 ( .A(n6742), .ZN(n5941) );
  NAND2_X1 U7541 ( .A1(n5930), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5937) );
  INV_X1 U7542 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7543 ( .A1(n5897), .A2(n5931), .ZN(n5936) );
  NAND2_X1 U7544 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5932) );
  AND2_X1 U7545 ( .A1(n5943), .A2(n5932), .ZN(n6690) );
  OR2_X1 U7546 ( .A1(n6065), .A2(n6690), .ZN(n5935) );
  INV_X1 U7547 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5933) );
  OR2_X1 U7548 ( .A1(n4275), .A2(n5933), .ZN(n5934) );
  NAND4_X1 U7549 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n9873)
         );
  OR2_X1 U7550 ( .A1(n5950), .A2(n5849), .ZN(n5938) );
  XNOR2_X1 U7551 ( .A(n5938), .B(n5949), .ZN(n6529) );
  OR2_X1 U7552 ( .A1(n8299), .A2(n6385), .ZN(n5940) );
  OR2_X1 U7553 ( .A1(n5904), .A2(n6384), .ZN(n5939) );
  OAI211_X1 U7554 ( .C1(n8296), .C2(n6529), .A(n5940), .B(n5939), .ZN(n6751)
         );
  NAND2_X1 U7555 ( .A1(n4734), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5948) );
  INV_X1 U7556 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7557 ( .A1(n6159), .A2(n5942), .ZN(n5947) );
  NAND2_X1 U7558 ( .A1(n5943), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5944) );
  AND2_X1 U7559 ( .A1(n5957), .A2(n5944), .ZN(n6814) );
  OR2_X1 U7560 ( .A1(n6065), .A2(n6814), .ZN(n5946) );
  INV_X1 U7561 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6663) );
  OR2_X1 U7562 ( .A1(n4275), .A2(n6663), .ZN(n5945) );
  NAND4_X1 U7563 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8527)
         );
  OR2_X1 U7564 ( .A1(n5904), .A2(n6387), .ZN(n5955) );
  OR2_X1 U7565 ( .A1(n8299), .A2(n6386), .ZN(n5954) );
  NAND2_X1 U7566 ( .A1(n5950), .A2(n5949), .ZN(n5963) );
  NAND2_X1 U7567 ( .A1(n5963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7568 ( .A(n5952), .B(n5951), .ZN(n6649) );
  OR2_X1 U7569 ( .A1(n8296), .A2(n6649), .ZN(n5953) );
  AND3_X2 U7570 ( .A1(n5955), .A2(n5954), .A3(n5953), .ZN(n9887) );
  OR2_X1 U7571 ( .A1(n8527), .A2(n9887), .ZN(n8348) );
  NAND2_X1 U7572 ( .A1(n8527), .A2(n9887), .ZN(n8343) );
  NAND2_X1 U7573 ( .A1(n8348), .A2(n8343), .ZN(n8476) );
  INV_X1 U7574 ( .A(n8527), .ZN(n9894) );
  NAND2_X1 U7575 ( .A1(n9894), .A2(n9887), .ZN(n5956) );
  NAND2_X1 U7576 ( .A1(n4734), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5962) );
  INV_X1 U7577 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6888) );
  OR2_X1 U7578 ( .A1(n6159), .A2(n6888), .ZN(n5961) );
  NAND2_X1 U7579 ( .A1(n5957), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5958) );
  AND2_X1 U7580 ( .A1(n5972), .A2(n5958), .ZN(n6922) );
  OR2_X1 U7581 ( .A1(n6065), .A2(n6922), .ZN(n5960) );
  INV_X1 U7582 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7583 ( .A1(n4275), .A2(n6662), .ZN(n5959) );
  NAND4_X1 U7584 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8526)
         );
  OR2_X1 U7585 ( .A1(n5966), .A2(n5849), .ZN(n5964) );
  MUX2_X1 U7586 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5964), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5967) );
  NAND2_X1 U7587 ( .A1(n5966), .A2(n5965), .ZN(n5983) );
  NAND2_X1 U7588 ( .A1(n5967), .A2(n5983), .ZN(n8533) );
  NAND2_X1 U7589 ( .A1(n6376), .A2(n8298), .ZN(n5969) );
  INV_X1 U7590 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6382) );
  OR2_X1 U7591 ( .A1(n8299), .A2(n6382), .ZN(n5968) );
  NAND2_X1 U7592 ( .A1(n8526), .A2(n9897), .ZN(n5970) );
  INV_X1 U7593 ( .A(n8526), .ZN(n9904) );
  NAND2_X1 U7594 ( .A1(n9904), .A2(n6237), .ZN(n5971) );
  NAND2_X1 U7595 ( .A1(n4734), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5977) );
  INV_X1 U7596 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6955) );
  OR2_X1 U7597 ( .A1(n6159), .A2(n6955), .ZN(n5976) );
  NAND2_X1 U7598 ( .A1(n5972), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5973) );
  AND2_X1 U7599 ( .A1(n5988), .A2(n5973), .ZN(n6938) );
  OR2_X1 U7600 ( .A1(n6065), .A2(n6938), .ZN(n5975) );
  INV_X1 U7601 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6655) );
  OR2_X1 U7602 ( .A1(n4275), .A2(n6655), .ZN(n5974) );
  NAND4_X1 U7603 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8525)
         );
  NAND2_X1 U7604 ( .A1(n6388), .A2(n8298), .ZN(n5980) );
  NAND2_X1 U7605 ( .A1(n5983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7606 ( .A(n5978), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6697) );
  AOI22_X1 U7607 ( .A1(n6113), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6112), .B2(
        n6697), .ZN(n5979) );
  OR2_X1 U7608 ( .A1(n8525), .A2(n6937), .ZN(n8358) );
  NAND2_X1 U7609 ( .A1(n6937), .A2(n8525), .ZN(n6961) );
  NAND2_X1 U7610 ( .A1(n8358), .A2(n6961), .ZN(n6952) );
  NAND2_X1 U7611 ( .A1(n6951), .A2(n6952), .ZN(n5982) );
  INV_X1 U7612 ( .A(n8525), .ZN(n9895) );
  NAND2_X1 U7613 ( .A1(n9895), .A2(n6937), .ZN(n5981) );
  NAND2_X1 U7614 ( .A1(n5982), .A2(n5981), .ZN(n6964) );
  NAND2_X1 U7615 ( .A1(n6392), .A2(n8298), .ZN(n5986) );
  NAND2_X1 U7616 ( .A1(n5995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U7617 ( .A(n5984), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6868) );
  AOI22_X1 U7618 ( .A1(n6113), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6112), .B2(
        n6868), .ZN(n5985) );
  NAND2_X1 U7619 ( .A1(n5986), .A2(n5985), .ZN(n9916) );
  NAND2_X1 U7620 ( .A1(n5930), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5993) );
  INV_X1 U7621 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5987) );
  OR2_X1 U7622 ( .A1(n5897), .A2(n5987), .ZN(n5992) );
  NAND2_X1 U7623 ( .A1(n5988), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5989) );
  AND2_X1 U7624 ( .A1(n5999), .A2(n5989), .ZN(n7116) );
  OR2_X1 U7625 ( .A1(n6065), .A2(n7116), .ZN(n5991) );
  INV_X1 U7626 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6715) );
  OR2_X1 U7627 ( .A1(n4275), .A2(n6715), .ZN(n5990) );
  OR2_X1 U7628 ( .A1(n9916), .A2(n9918), .ZN(n8354) );
  NAND2_X1 U7629 ( .A1(n9916), .A2(n9918), .ZN(n8359) );
  INV_X1 U7630 ( .A(n9918), .ZN(n8524) );
  NAND2_X1 U7631 ( .A1(n9916), .A2(n8524), .ZN(n5994) );
  NAND2_X1 U7632 ( .A1(n6407), .A2(n8298), .ZN(n5998) );
  NAND2_X1 U7633 ( .A1(n6007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7634 ( .A(n5996), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U7635 ( .A1(n6113), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6112), .B2(
        n6974), .ZN(n5997) );
  NAND2_X1 U7636 ( .A1(n5998), .A2(n5997), .ZN(n9922) );
  NAND2_X1 U7637 ( .A1(n4734), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6004) );
  INV_X1 U7638 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7036) );
  OR2_X1 U7639 ( .A1(n6159), .A2(n7036), .ZN(n6003) );
  NAND2_X1 U7640 ( .A1(n5999), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6000) );
  AND2_X1 U7641 ( .A1(n6015), .A2(n6000), .ZN(n7214) );
  OR2_X1 U7642 ( .A1(n6065), .A2(n7214), .ZN(n6002) );
  INV_X1 U7643 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6859) );
  OR2_X1 U7644 ( .A1(n4275), .A2(n6859), .ZN(n6001) );
  NAND4_X1 U7645 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n8523)
         );
  NAND2_X1 U7646 ( .A1(n9922), .A2(n8523), .ZN(n6005) );
  NAND2_X1 U7647 ( .A1(n6006), .A2(n6005), .ZN(n7140) );
  NOR2_X1 U7648 ( .A1(n6010), .A2(n5849), .ZN(n6008) );
  MUX2_X1 U7649 ( .A(n5849), .B(n6008), .S(P2_IR_REG_10__SCAN_IN), .Z(n6012)
         );
  INV_X1 U7650 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7651 ( .A1(n6010), .A2(n6009), .ZN(n6024) );
  INV_X1 U7652 ( .A(n6024), .ZN(n6011) );
  INV_X1 U7653 ( .A(n7149), .ZN(n7154) );
  AOI22_X1 U7654 ( .A1(n6113), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6112), .B2(
        n7154), .ZN(n6013) );
  NAND2_X1 U7655 ( .A1(n5930), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6020) );
  INV_X1 U7656 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7657 ( .A1(n5897), .A2(n6014), .ZN(n6019) );
  NAND2_X1 U7658 ( .A1(n6015), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6016) );
  AND2_X1 U7659 ( .A1(n6028), .A2(n6016), .ZN(n7363) );
  OR2_X1 U7660 ( .A1(n6065), .A2(n7363), .ZN(n6018) );
  INV_X1 U7661 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6993) );
  OR2_X1 U7662 ( .A1(n4275), .A2(n6993), .ZN(n6017) );
  NAND4_X1 U7663 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n8522)
         );
  AND2_X1 U7664 ( .A1(n9934), .A2(n8522), .ZN(n6021) );
  INV_X1 U7665 ( .A(n6021), .ZN(n6022) );
  NAND2_X1 U7666 ( .A1(n6505), .A2(n8298), .ZN(n6027) );
  NAND2_X1 U7667 ( .A1(n6024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6023) );
  MUX2_X1 U7668 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6023), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n6025) );
  AOI22_X1 U7669 ( .A1(n6113), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6112), .B2(
        n7387), .ZN(n6026) );
  NAND2_X1 U7670 ( .A1(n6027), .A2(n6026), .ZN(n9939) );
  NAND2_X1 U7671 ( .A1(n4734), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6033) );
  INV_X1 U7672 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7160) );
  OR2_X1 U7673 ( .A1(n6159), .A2(n7160), .ZN(n6032) );
  NAND2_X1 U7674 ( .A1(n6028), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6029) );
  AND2_X1 U7675 ( .A1(n6038), .A2(n6029), .ZN(n7500) );
  OR2_X1 U7676 ( .A1(n6065), .A2(n7500), .ZN(n6031) );
  INV_X1 U7677 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7159) );
  OR2_X1 U7678 ( .A1(n4275), .A2(n7159), .ZN(n6030) );
  NAND2_X1 U7679 ( .A1(n9939), .A2(n7488), .ZN(n8374) );
  NAND2_X1 U7680 ( .A1(n6642), .A2(n8298), .ZN(n6037) );
  NAND2_X1 U7681 ( .A1(n6047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6035) );
  AOI22_X1 U7682 ( .A1(n6113), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6112), .B2(
        n7546), .ZN(n6036) );
  NAND2_X1 U7683 ( .A1(n5930), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6043) );
  INV_X1 U7684 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7427) );
  OR2_X1 U7685 ( .A1(n5897), .A2(n7427), .ZN(n6042) );
  NAND2_X1 U7686 ( .A1(n6038), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6039) );
  AND2_X1 U7687 ( .A1(n6051), .A2(n6039), .ZN(n7492) );
  OR2_X1 U7688 ( .A1(n6065), .A2(n7492), .ZN(n6041) );
  INV_X1 U7689 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7407) );
  OR2_X1 U7690 ( .A1(n4275), .A2(n7407), .ZN(n6040) );
  NAND4_X1 U7691 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8520)
         );
  OR2_X1 U7692 ( .A1(n7494), .A2(n8520), .ZN(n6044) );
  NAND2_X1 U7693 ( .A1(n7422), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7694 ( .A1(n7494), .A2(n8520), .ZN(n6045) );
  NAND2_X1 U7695 ( .A1(n6046), .A2(n6045), .ZN(n7463) );
  NAND2_X1 U7696 ( .A1(n6677), .A2(n8298), .ZN(n6050) );
  NAND2_X1 U7697 ( .A1(n6048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6059) );
  XNOR2_X1 U7698 ( .A(n6059), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7630) );
  AOI22_X1 U7699 ( .A1(n6112), .A2(n7630), .B1(n6113), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7700 ( .A1(n4734), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6056) );
  INV_X1 U7701 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7551) );
  OR2_X1 U7702 ( .A1(n6159), .A2(n7551), .ZN(n6055) );
  NAND2_X1 U7703 ( .A1(n6051), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6052) );
  AND2_X1 U7704 ( .A1(n6063), .A2(n6052), .ZN(n8866) );
  OR2_X1 U7705 ( .A1(n6065), .A2(n8866), .ZN(n6054) );
  INV_X1 U7706 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7550) );
  OR2_X1 U7707 ( .A1(n4275), .A2(n7550), .ZN(n6053) );
  NAND4_X1 U7708 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n8519)
         );
  AND2_X1 U7709 ( .A1(n8870), .A2(n8519), .ZN(n8388) );
  OR2_X1 U7710 ( .A1(n8870), .A2(n8519), .ZN(n8393) );
  OAI21_X1 U7711 ( .B1(n7463), .B2(n8388), .A(n8393), .ZN(n6057) );
  INV_X1 U7712 ( .A(n6057), .ZN(n7509) );
  NAND2_X1 U7713 ( .A1(n6740), .A2(n8298), .ZN(n6062) );
  INV_X1 U7714 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7715 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7716 ( .A1(n6060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  AOI22_X1 U7717 ( .A1(n8558), .A2(n6112), .B1(n6113), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7718 ( .A1(n6062), .A2(n6061), .ZN(n8092) );
  NAND2_X1 U7719 ( .A1(n4734), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6069) );
  INV_X1 U7720 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7642) );
  OR2_X1 U7721 ( .A1(n6159), .A2(n7642), .ZN(n6068) );
  NAND2_X1 U7722 ( .A1(n6063), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6064) );
  AND2_X1 U7723 ( .A1(n6079), .A2(n6064), .ZN(n8158) );
  OR2_X1 U7724 ( .A1(n6065), .A2(n8158), .ZN(n6067) );
  INV_X1 U7725 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8557) );
  OR2_X1 U7726 ( .A1(n4275), .A2(n8557), .ZN(n6066) );
  OR2_X1 U7727 ( .A1(n8092), .A2(n6070), .ZN(n8396) );
  NAND2_X1 U7728 ( .A1(n8092), .A2(n6070), .ZN(n8397) );
  NAND2_X1 U7729 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  NAND2_X1 U7730 ( .A1(n7509), .A2(n8395), .ZN(n7508) );
  NAND2_X1 U7731 ( .A1(n8092), .A2(n8855), .ZN(n6071) );
  NAND2_X1 U7732 ( .A1(n6819), .A2(n8298), .ZN(n6078) );
  INV_X1 U7733 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7734 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U7735 ( .A1(n6074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6075) );
  XNOR2_X1 U7736 ( .A(n6075), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8577) );
  NOR2_X1 U7737 ( .A1(n8299), .A2(n10006), .ZN(n6076) );
  AOI21_X1 U7738 ( .B1(n8577), .B2(n6112), .A(n6076), .ZN(n6077) );
  INV_X1 U7739 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8563) );
  OR2_X1 U7740 ( .A1(n6159), .A2(n8563), .ZN(n6084) );
  INV_X1 U7741 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10119) );
  OR2_X1 U7742 ( .A1(n5897), .A2(n10119), .ZN(n6083) );
  NAND2_X1 U7743 ( .A1(n6079), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6080) );
  AND2_X1 U7744 ( .A1(n6090), .A2(n6080), .ZN(n8858) );
  OR2_X1 U7745 ( .A1(n6065), .A2(n8858), .ZN(n6082) );
  INV_X1 U7746 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10113) );
  OR2_X1 U7747 ( .A1(n4275), .A2(n10113), .ZN(n6081) );
  NAND2_X1 U7748 ( .A1(n9023), .A2(n8095), .ZN(n8400) );
  INV_X1 U7749 ( .A(n8095), .ZN(n8518) );
  OR2_X1 U7750 ( .A1(n9023), .A2(n8518), .ZN(n6086) );
  NAND2_X1 U7751 ( .A1(n6946), .A2(n8298), .ZN(n6089) );
  NAND2_X1 U7752 ( .A1(n6224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U7753 ( .A(n6087), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8612) );
  AOI22_X1 U7754 ( .A1(n6113), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6112), .B2(
        n8612), .ZN(n6088) );
  NAND2_X1 U7755 ( .A1(n6090), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7756 ( .A1(n6102), .A2(n6091), .ZN(n8213) );
  NAND2_X1 U7757 ( .A1(n6211), .A2(n8213), .ZN(n6095) );
  INV_X1 U7758 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8605) );
  OR2_X1 U7759 ( .A1(n6159), .A2(n8605), .ZN(n6094) );
  INV_X1 U7760 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10074) );
  OR2_X1 U7761 ( .A1(n5897), .A2(n10074), .ZN(n6093) );
  INV_X1 U7762 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8611) );
  OR2_X1 U7763 ( .A1(n4275), .A2(n8611), .ZN(n6092) );
  NAND2_X1 U7764 ( .A1(n8098), .A2(n8841), .ZN(n8405) );
  NAND2_X1 U7765 ( .A1(n8404), .A2(n8405), .ZN(n8491) );
  NAND2_X1 U7766 ( .A1(n8098), .A2(n8856), .ZN(n6096) );
  NAND2_X1 U7767 ( .A1(n7694), .A2(n6096), .ZN(n8840) );
  NAND2_X1 U7768 ( .A1(n7044), .A2(n8298), .ZN(n6101) );
  NAND2_X1 U7769 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6098) );
  MUX2_X1 U7770 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6098), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6099) );
  NAND2_X1 U7771 ( .A1(n6099), .A2(n6110), .ZN(n8643) );
  INV_X1 U7772 ( .A(n8643), .ZN(n8637) );
  AOI22_X1 U7773 ( .A1(n6113), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6112), .B2(
        n8637), .ZN(n6100) );
  NAND2_X1 U7774 ( .A1(n6102), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7775 ( .A1(n6116), .A2(n6103), .ZN(n8847) );
  NAND2_X1 U7776 ( .A1(n6211), .A2(n8847), .ZN(n6108) );
  INV_X1 U7777 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10130) );
  OR2_X1 U7778 ( .A1(n6159), .A2(n10130), .ZN(n6107) );
  INV_X1 U7779 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9016) );
  OR2_X1 U7780 ( .A1(n5897), .A2(n9016), .ZN(n6106) );
  INV_X1 U7781 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7782 ( .A1(n4275), .A2(n6104), .ZN(n6105) );
  NAND2_X1 U7783 ( .A1(n9018), .A2(n8831), .ZN(n8412) );
  NAND2_X1 U7784 ( .A1(n8406), .A2(n8412), .ZN(n8839) );
  NAND2_X1 U7785 ( .A1(n8840), .A2(n8839), .ZN(n8838) );
  INV_X1 U7786 ( .A(n8831), .ZN(n8943) );
  NAND2_X1 U7787 ( .A1(n9018), .A2(n8943), .ZN(n6109) );
  NAND2_X1 U7788 ( .A1(n7101), .A2(n8298), .ZN(n6115) );
  NAND2_X1 U7789 ( .A1(n6110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6111) );
  XNOR2_X1 U7790 ( .A(n6111), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8663) );
  AOI22_X1 U7791 ( .A1(n6113), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6112), .B2(
        n8663), .ZN(n6114) );
  NAND2_X1 U7792 ( .A1(n6116), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7793 ( .A1(n6118), .A2(n6117), .ZN(n8827) );
  NAND2_X1 U7794 ( .A1(n8827), .A2(n6211), .ZN(n6122) );
  NAND2_X1 U7795 ( .A1(n5930), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7796 ( .A1(n4734), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6120) );
  INV_X1 U7797 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9997) );
  OR2_X1 U7798 ( .A1(n4275), .A2(n9997), .ZN(n6119) );
  NAND2_X1 U7799 ( .A1(n8833), .A2(n8842), .ZN(n8413) );
  NAND2_X1 U7800 ( .A1(n8414), .A2(n8413), .ZN(n8824) );
  NAND2_X1 U7801 ( .A1(n8825), .A2(n8824), .ZN(n8823) );
  INV_X1 U7802 ( .A(n8842), .ZN(n8517) );
  OR2_X1 U7803 ( .A1(n8833), .A2(n8517), .ZN(n6123) );
  NAND2_X1 U7804 ( .A1(n8823), .A2(n6123), .ZN(n8807) );
  NAND2_X1 U7805 ( .A1(n9007), .A2(n8933), .ZN(n8418) );
  NAND2_X1 U7806 ( .A1(n7325), .A2(n8298), .ZN(n6126) );
  INV_X1 U7807 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7808 ( .A1(n8299), .A2(n6124), .ZN(n6125) );
  NAND2_X1 U7809 ( .A1(n6127), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7810 ( .A1(n6134), .A2(n6128), .ZN(n8799) );
  NAND2_X1 U7811 ( .A1(n8799), .A2(n6211), .ZN(n6131) );
  AOI22_X1 U7812 ( .A1(n5930), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n4734), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7813 ( .A1(n5898), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7814 ( .A1(n8931), .A2(n8924), .ZN(n8782) );
  NAND2_X1 U7815 ( .A1(n8420), .A2(n8782), .ZN(n8797) );
  NAND2_X1 U7816 ( .A1(n7420), .A2(n8298), .ZN(n6133) );
  OR2_X1 U7817 ( .A1(n8299), .A2(n7430), .ZN(n6132) );
  NAND2_X1 U7818 ( .A1(n6134), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7819 ( .A1(n6144), .A2(n6135), .ZN(n8788) );
  NAND2_X1 U7820 ( .A1(n8788), .A2(n6211), .ZN(n6140) );
  INV_X1 U7821 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U7822 ( .A1(n5930), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7823 ( .A1(n4734), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6136) );
  OAI211_X1 U7824 ( .C1(n8929), .C2(n4275), .A(n6137), .B(n6136), .ZN(n6138)
         );
  INV_X1 U7825 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7826 ( .A1(n8792), .A2(n8934), .ZN(n8426) );
  NAND2_X1 U7827 ( .A1(n8427), .A2(n8426), .ZN(n8785) );
  INV_X1 U7828 ( .A(n8792), .ZN(n9000) );
  NAND2_X1 U7829 ( .A1(n7563), .A2(n8298), .ZN(n6143) );
  OR2_X1 U7830 ( .A1(n8299), .A2(n10005), .ZN(n6142) );
  NAND2_X1 U7831 ( .A1(n6144), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7832 ( .A1(n6154), .A2(n6145), .ZN(n8771) );
  NAND2_X1 U7833 ( .A1(n8771), .A2(n6211), .ZN(n6150) );
  INV_X1 U7834 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U7835 ( .A1(n4734), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7836 ( .A1(n5930), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6146) );
  OAI211_X1 U7837 ( .C1(n4275), .C2(n10104), .A(n6147), .B(n6146), .ZN(n6148)
         );
  INV_X1 U7838 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7839 ( .A1(n8921), .A2(n8925), .ZN(n8430) );
  NAND2_X1 U7840 ( .A1(n7577), .A2(n8298), .ZN(n6153) );
  OR2_X1 U7841 ( .A1(n8299), .A2(n10120), .ZN(n6152) );
  NAND2_X1 U7842 ( .A1(n6154), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7843 ( .A1(n6156), .A2(n6155), .ZN(n8762) );
  NAND2_X1 U7844 ( .A1(n8762), .A2(n6211), .ZN(n6162) );
  INV_X1 U7845 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U7846 ( .A1(n5898), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7847 ( .A1(n4734), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6157) );
  OAI211_X1 U7848 ( .C1(n6159), .C2(n8761), .A(n6158), .B(n6157), .ZN(n6160)
         );
  INV_X1 U7849 ( .A(n6160), .ZN(n6161) );
  NOR2_X1 U7850 ( .A1(n8989), .A2(n8775), .ZN(n6164) );
  INV_X1 U7851 ( .A(n8989), .ZN(n6163) );
  NAND2_X1 U7852 ( .A1(n7691), .A2(n8298), .ZN(n6168) );
  OR2_X1 U7853 ( .A1(n8299), .A2(n6166), .ZN(n6167) );
  INV_X1 U7854 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7855 ( .A1(n6171), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7856 ( .A1(n6180), .A2(n6172), .ZN(n8200) );
  NAND2_X1 U7857 ( .A1(n8200), .A2(n6211), .ZN(n6177) );
  INV_X1 U7858 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U7859 ( .A1(n5930), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7860 ( .A1(n4734), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7861 ( .C1(n8908), .C2(n4275), .A(n6174), .B(n6173), .ZN(n6175)
         );
  INV_X1 U7862 ( .A(n6175), .ZN(n6176) );
  OR2_X1 U7863 ( .A1(n8978), .A2(n8516), .ZN(n8440) );
  NAND2_X1 U7864 ( .A1(n7729), .A2(n8298), .ZN(n6179) );
  OR2_X1 U7865 ( .A1(n8299), .A2(n10076), .ZN(n6178) );
  NAND2_X1 U7866 ( .A1(n6180), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7867 ( .A1(n6191), .A2(n6181), .ZN(n8728) );
  NAND2_X1 U7868 ( .A1(n8728), .A2(n6211), .ZN(n6186) );
  INV_X1 U7869 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U7870 ( .A1(n5930), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7871 ( .A1(n4734), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6182) );
  OAI211_X1 U7872 ( .C1(n8906), .C2(n4275), .A(n6183), .B(n6182), .ZN(n6184)
         );
  INV_X1 U7873 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7874 ( .A1(n8732), .A2(n8738), .ZN(n6187) );
  NAND2_X1 U7875 ( .A1(n7734), .A2(n8298), .ZN(n6189) );
  OR2_X1 U7876 ( .A1(n8299), .A2(n10082), .ZN(n6188) );
  INV_X1 U7877 ( .A(n6191), .ZN(n6190) );
  INV_X1 U7878 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7879 ( .A1(n6191), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7880 ( .A1(n6201), .A2(n6192), .ZN(n8721) );
  NAND2_X1 U7881 ( .A1(n8721), .A2(n6211), .ZN(n6197) );
  INV_X1 U7882 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U7883 ( .A1(n5930), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7884 ( .A1(n4734), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7885 ( .C1(n10058), .C2(n4275), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7886 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U7887 ( .A1(n8968), .A2(n8902), .ZN(n8320) );
  NAND2_X1 U7888 ( .A1(n8319), .A2(n8320), .ZN(n8710) );
  INV_X1 U7889 ( .A(n8968), .ZN(n8151) );
  NAND2_X1 U7890 ( .A1(n8078), .A2(n8298), .ZN(n6200) );
  OR2_X1 U7891 ( .A1(n8299), .A2(n6198), .ZN(n6199) );
  NAND2_X1 U7892 ( .A1(n6201), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7893 ( .A1(n8689), .A2(n6202), .ZN(n8703) );
  NAND2_X1 U7894 ( .A1(n8703), .A2(n6211), .ZN(n6207) );
  INV_X1 U7895 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7896 ( .A1(n5930), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7897 ( .A1(n4734), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6203) );
  OAI211_X1 U7898 ( .C1(n6335), .C2(n4275), .A(n6204), .B(n6203), .ZN(n6205)
         );
  INV_X1 U7899 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7900 ( .A1(n8455), .A2(n8716), .ZN(n6208) );
  NAND2_X1 U7901 ( .A1(n8081), .A2(n8298), .ZN(n6210) );
  OR2_X1 U7902 ( .A1(n8299), .A2(n8082), .ZN(n6209) );
  INV_X1 U7903 ( .A(n8689), .ZN(n6212) );
  NAND2_X1 U7904 ( .A1(n6212), .A2(n6211), .ZN(n8309) );
  INV_X1 U7905 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7906 ( .A1(n4734), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7907 ( .A1(n5930), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6213) );
  OAI211_X1 U7908 ( .C1(n4275), .C2(n6342), .A(n6214), .B(n6213), .ZN(n6215)
         );
  INV_X1 U7909 ( .A(n6215), .ZN(n6216) );
  NAND2_X1 U7910 ( .A1(n6312), .A2(n9990), .ZN(n8310) );
  XNOR2_X1 U7911 ( .A(n6218), .B(n6217), .ZN(n6230) );
  NAND2_X1 U7912 ( .A1(n6272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7913 ( .A1(n8508), .A2(n6270), .ZN(n6304) );
  NAND2_X1 U7914 ( .A1(n6222), .A2(n6221), .ZN(n6228) );
  NAND2_X1 U7915 ( .A1(n6228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6223) );
  INV_X1 U7916 ( .A(n6224), .ZN(n6225) );
  NAND2_X1 U7917 ( .A1(n4322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6227) );
  MUX2_X1 U7918 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6227), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6229) );
  NAND2_X1 U7919 ( .A1(n6547), .A2(n6327), .ZN(n8504) );
  NAND2_X1 U7920 ( .A1(n6230), .A2(n9902), .ZN(n6269) );
  INV_X1 U7921 ( .A(n6736), .ZN(n6418) );
  NOR2_X2 U7922 ( .A1(n6415), .A2(n6418), .ZN(n8878) );
  INV_X1 U7923 ( .A(n6793), .ZN(n8474) );
  NAND2_X1 U7924 ( .A1(n6791), .A2(n8474), .ZN(n6233) );
  NAND2_X1 U7925 ( .A1(n6233), .A2(n8330), .ZN(n6847) );
  INV_X1 U7926 ( .A(n6849), .ZN(n8473) );
  NAND2_X1 U7927 ( .A1(n6847), .A2(n8473), .ZN(n6235) );
  NAND2_X1 U7928 ( .A1(n6235), .A2(n6234), .ZN(n6745) );
  NOR2_X1 U7929 ( .A1(n9873), .A2(n9882), .ZN(n8341) );
  NAND2_X1 U7930 ( .A1(n9873), .A2(n9882), .ZN(n6803) );
  AND2_X1 U7931 ( .A1(n6803), .A2(n8343), .ZN(n8345) );
  NAND2_X1 U7932 ( .A1(n8526), .A2(n6237), .ZN(n8350) );
  INV_X1 U7933 ( .A(n8478), .ZN(n6238) );
  NAND2_X1 U7934 ( .A1(n6892), .A2(n6238), .ZN(n6239) );
  NAND2_X1 U7935 ( .A1(n6239), .A2(n8357), .ZN(n6950) );
  AND2_X1 U7936 ( .A1(n8354), .A2(n6961), .ZN(n8365) );
  INV_X1 U7937 ( .A(n8359), .ZN(n6240) );
  XNOR2_X1 U7938 ( .A(n9922), .B(n8523), .ZN(n8356) );
  OR2_X1 U7939 ( .A1(n9934), .A2(n9920), .ZN(n8372) );
  INV_X1 U7940 ( .A(n8523), .ZN(n8360) );
  OR2_X1 U7941 ( .A1(n9922), .A2(n8360), .ZN(n7137) );
  NAND2_X1 U7942 ( .A1(n9934), .A2(n9920), .ZN(n8362) );
  AND2_X1 U7943 ( .A1(n8374), .A2(n8362), .ZN(n8371) );
  INV_X1 U7944 ( .A(n8520), .ZN(n8244) );
  OR2_X1 U7945 ( .A1(n7494), .A2(n8244), .ZN(n8385) );
  NAND2_X1 U7946 ( .A1(n7494), .A2(n8244), .ZN(n8384) );
  NAND2_X1 U7947 ( .A1(n7424), .A2(n8382), .ZN(n6241) );
  NAND2_X1 U7948 ( .A1(n6241), .A2(n8385), .ZN(n7465) );
  INV_X1 U7949 ( .A(n7465), .ZN(n6242) );
  INV_X1 U7950 ( .A(n8519), .ZN(n8161) );
  NAND2_X1 U7951 ( .A1(n6242), .A2(n4863), .ZN(n6244) );
  NAND2_X1 U7952 ( .A1(n8870), .A2(n8161), .ZN(n6243) );
  NAND2_X1 U7953 ( .A1(n6245), .A2(n8412), .ZN(n8820) );
  INV_X1 U7954 ( .A(n8415), .ZN(n6248) );
  AND2_X1 U7955 ( .A1(n8426), .A2(n8782), .ZN(n8422) );
  NAND2_X1 U7956 ( .A1(n8783), .A2(n8422), .ZN(n6249) );
  NAND2_X1 U7957 ( .A1(n6249), .A2(n8427), .ZN(n8768) );
  NAND2_X1 U7958 ( .A1(n8768), .A2(n8767), .ZN(n8770) );
  NAND2_X1 U7959 ( .A1(n8770), .A2(n8432), .ZN(n8756) );
  NOR2_X1 U7960 ( .A1(n8989), .A2(n8916), .ZN(n8321) );
  NAND2_X1 U7961 ( .A1(n8989), .A2(n8916), .ZN(n8471) );
  INV_X1 U7962 ( .A(n8434), .ZN(n6250) );
  NOR2_X1 U7963 ( .A1(n8978), .A2(n8901), .ZN(n8443) );
  AND2_X1 U7964 ( .A1(n8732), .A2(n8715), .ZN(n8446) );
  NAND2_X1 U7965 ( .A1(n6252), .A2(n8448), .ZN(n8711) );
  NAND2_X1 U7966 ( .A1(n8711), .A2(n8320), .ZN(n6253) );
  NAND2_X1 U7967 ( .A1(n6336), .A2(n8716), .ZN(n6254) );
  INV_X1 U7968 ( .A(n8508), .ZN(n8322) );
  NAND2_X1 U7969 ( .A1(n8322), .A2(n8323), .ZN(n9886) );
  OAI211_X1 U7970 ( .C1(n8508), .C2(n8462), .A(n9886), .B(n4274), .ZN(n6255)
         );
  INV_X1 U7971 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7972 ( .A1(n8672), .A2(n8462), .ZN(n6548) );
  OR2_X1 U7973 ( .A1(n4495), .A2(n6548), .ZN(n6731) );
  NAND2_X1 U7974 ( .A1(n6256), .A2(n6731), .ZN(n9866) );
  INV_X1 U7975 ( .A(n6257), .ZN(n6402) );
  NAND2_X1 U7976 ( .A1(n6402), .A2(n8506), .ZN(n6259) );
  NAND2_X1 U7977 ( .A1(n8296), .A2(n6259), .ZN(n6542) );
  INV_X1 U7978 ( .A(n6542), .ZN(n6479) );
  INV_X1 U7979 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7980 ( .A1(n5930), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7981 ( .A1(n4734), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U7982 ( .C1(n6262), .C2(n4275), .A(n6261), .B(n6260), .ZN(n6263)
         );
  INV_X1 U7983 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7984 ( .A1(n8309), .A2(n6264), .ZN(n8513) );
  AND2_X1 U7985 ( .A1(n8296), .A2(P2_B_REG_SCAN_IN), .ZN(n6265) );
  NOR2_X1 U7986 ( .A1(n9919), .A2(n6265), .ZN(n8687) );
  AOI22_X1 U7987 ( .A1(n9874), .A2(n8514), .B1(n8513), .B2(n8687), .ZN(n6266)
         );
  NAND2_X1 U7988 ( .A1(n6269), .A2(n6268), .ZN(n8694) );
  NAND2_X1 U7989 ( .A1(n6270), .A2(n8462), .ZN(n6305) );
  NOR2_X1 U7990 ( .A1(n8701), .A2(n9930), .ZN(n6271) );
  NOR2_X1 U7991 ( .A1(n8694), .A2(n6271), .ZN(n6345) );
  NAND2_X1 U7992 ( .A1(n6303), .A2(n10073), .ZN(n6274) );
  NAND2_X1 U7993 ( .A1(n6274), .A2(n4341), .ZN(n6278) );
  AND2_X1 U7994 ( .A1(n10073), .A2(n6275), .ZN(n6276) );
  NAND2_X1 U7995 ( .A1(n6303), .A2(n6277), .ZN(n6279) );
  NAND2_X1 U7996 ( .A1(n6278), .A2(n6279), .ZN(n7659) );
  XNOR2_X1 U7997 ( .A(n7659), .B(P2_B_REG_SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7998 ( .A1(n6279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7999 ( .A1(n6282), .A2(n7733), .ZN(n6285) );
  NAND2_X1 U8000 ( .A1(n6283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U8001 ( .A1(n7659), .A2(n7738), .ZN(n6379) );
  NOR2_X1 U8002 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n6290) );
  NOR4_X1 U8003 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6289) );
  NOR4_X1 U8004 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6288) );
  NOR4_X1 U8005 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6287) );
  NAND4_X1 U8006 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n6296)
         );
  NOR4_X1 U8007 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6294) );
  NOR4_X1 U8008 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6293) );
  NOR4_X1 U8009 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6292) );
  NOR4_X1 U8010 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6291) );
  NAND4_X1 U8011 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n6295)
         );
  NOR2_X1 U8012 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  INV_X1 U8013 ( .A(n6324), .ZN(n6307) );
  NOR2_X1 U8014 ( .A1(n6728), .A2(n6307), .ZN(n6300) );
  NAND2_X1 U8015 ( .A1(n7733), .A2(n7738), .ZN(n6298) );
  AND2_X1 U8016 ( .A1(n6300), .A2(n6331), .ZN(n6500) );
  INV_X1 U8017 ( .A(n7733), .ZN(n6302) );
  NOR2_X1 U8018 ( .A1(n7659), .A2(n7738), .ZN(n6301) );
  NAND2_X1 U8019 ( .A1(n8323), .A2(n6327), .ZN(n6546) );
  OR2_X1 U8020 ( .A1(n6546), .A2(n6304), .ZN(n6496) );
  NAND3_X1 U8021 ( .A1(n4495), .A2(n6496), .A3(n9886), .ZN(n6482) );
  INV_X1 U8022 ( .A(n6305), .ZN(n6306) );
  NAND2_X1 U8023 ( .A1(n6482), .A2(n8752), .ZN(n6492) );
  NAND2_X1 U8024 ( .A1(n6481), .A2(n6492), .ZN(n6311) );
  NAND2_X1 U8025 ( .A1(n6727), .A2(n6728), .ZN(n6326) );
  OR2_X1 U8026 ( .A1(n6326), .A2(n6307), .ZN(n6493) );
  INV_X1 U8027 ( .A(n6499), .ZN(n6308) );
  NAND2_X1 U8028 ( .A1(n6496), .A2(n6731), .ZN(n6309) );
  NAND2_X1 U8029 ( .A1(n6486), .A2(n6309), .ZN(n6310) );
  INV_X1 U8030 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6314) );
  NOR2_X1 U8031 ( .A1(n9941), .A2(n6314), .ZN(n6315) );
  OAI21_X1 U8032 ( .B1(n6345), .B2(n9943), .A(n6316), .ZN(P2_U3456) );
  INV_X1 U8033 ( .A(n6319), .ZN(n6322) );
  OAI22_X1 U8034 ( .A1(n9990), .A2(n9919), .B1(n8902), .B2(n9917), .ZN(n6323)
         );
  NAND2_X1 U8035 ( .A1(n8459), .A2(n6548), .ZN(n6489) );
  AND3_X1 U8036 ( .A1(n6324), .A2(n6499), .A3(n6489), .ZN(n6325) );
  AND2_X1 U8037 ( .A1(n6326), .A2(n6325), .ZN(n6729) );
  INV_X1 U8038 ( .A(n6728), .ZN(n6329) );
  NOR2_X1 U8039 ( .A1(n9930), .A2(n6547), .ZN(n6487) );
  NAND3_X1 U8040 ( .A1(n8508), .A2(n4274), .A3(n6327), .ZN(n6328) );
  AND2_X1 U8041 ( .A1(n4495), .A2(n6328), .ZN(n6726) );
  OAI21_X1 U8042 ( .B1(n6329), .B2(n6487), .A(n6726), .ZN(n6333) );
  INV_X1 U8043 ( .A(n6726), .ZN(n6330) );
  NAND2_X1 U8044 ( .A1(n6331), .A2(n6330), .ZN(n6332) );
  NAND2_X1 U8045 ( .A1(n6336), .A2(n8953), .ZN(n6337) );
  INV_X1 U8046 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6339) );
  MUX2_X1 U8047 ( .A(n6339), .B(n6338), .S(n9941), .Z(n6341) );
  NAND2_X1 U8048 ( .A1(n6336), .A2(n9024), .ZN(n6340) );
  NAND2_X1 U8049 ( .A1(n6341), .A2(n6340), .ZN(P2_U3455) );
  OAI21_X1 U8050 ( .B1(n6345), .B2(n4414), .A(n6344), .ZN(P2_U3488) );
  NOR2_X1 U8051 ( .A1(n4934), .A2(P1_U3086), .ZN(n6346) );
  INV_X1 U8052 ( .A(n6381), .ZN(n6347) );
  NAND2_X1 U8053 ( .A1(n6491), .A2(n4495), .ZN(n6348) );
  NAND2_X1 U8054 ( .A1(n6348), .A2(n6490), .ZN(n6401) );
  NAND2_X1 U8055 ( .A1(n6401), .A2(n8296), .ZN(n6349) );
  NAND2_X1 U8056 ( .A1(n6349), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8057 ( .A1(n6351), .A2(n6350), .ZN(n6353) );
  XOR2_X1 U8058 ( .A(n6353), .B(n6352), .Z(n6354) );
  NOR2_X1 U8059 ( .A1(n6354), .A2(n9671), .ZN(n6360) );
  NOR2_X1 U8060 ( .A1(n9662), .A2(n7131), .ZN(n6359) );
  INV_X1 U8061 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6355) );
  OAI22_X1 U8062 ( .A1(n9661), .A2(n7524), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6355), .ZN(n6358) );
  OAI22_X1 U8063 ( .A1(n9678), .A2(n6356), .B1(n9157), .B2(n9825), .ZN(n6357)
         );
  OR4_X1 U8064 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(P1_U3213)
         );
  NOR2_X2 U8065 ( .A1(n6361), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9638) );
  AOI22_X1 U8066 ( .A1(n9638), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6784), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6362) );
  OAI21_X1 U8067 ( .B1(n6368), .B2(n9640), .A(n6362), .ZN(P1_U3353) );
  AOI22_X1 U8068 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9207), .B1(n9638), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8069 ( .B1(n6366), .B2(n9640), .A(n6363), .ZN(P1_U3352) );
  AOI22_X1 U8070 ( .A1(n9234), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9638), .ZN(n6364) );
  OAI21_X1 U8071 ( .B1(n6387), .B2(n9640), .A(n6364), .ZN(P1_U3350) );
  NAND2_X1 U8072 ( .A1(n8295), .A2(P2_U3151), .ZN(n9044) );
  INV_X1 U8073 ( .A(n6365), .ZN(n6373) );
  NOR2_X1 U8074 ( .A1(n8295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9046) );
  INV_X2 U8075 ( .A(n9046), .ZN(n9042) );
  OAI222_X1 U8076 ( .A1(P2_U3151), .A2(n6438), .B1(n9044), .B2(n6373), .C1(
        n4911), .C2(n9042), .ZN(P2_U3294) );
  OAI222_X1 U8077 ( .A1(n6478), .A2(P2_U3151), .B1(n9044), .B2(n6366), .C1(
        n4397), .C2(n9042), .ZN(P2_U3292) );
  OAI222_X1 U8078 ( .A1(n6520), .A2(P2_U3151), .B1(n9044), .B2(n6368), .C1(
        n6367), .C2(n9042), .ZN(P2_U3293) );
  INV_X1 U8079 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U8080 ( .A1(n6378), .A2(n9996), .ZN(P2_U3240) );
  INV_X1 U8081 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U8082 ( .A1(n6378), .A2(n10109), .ZN(P2_U3258) );
  INV_X1 U8083 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8084 ( .A1(n6727), .A2(n6499), .ZN(n6370) );
  OAI21_X1 U8085 ( .B1(n6499), .B2(n6371), .A(n6370), .ZN(P2_U3377) );
  INV_X1 U8086 ( .A(n9638), .ZN(n8084) );
  INV_X1 U8087 ( .A(n6623), .ZN(n9219) );
  OAI222_X1 U8088 ( .A1(n8084), .A2(n6372), .B1(n9640), .B2(n6384), .C1(
        P1_U3086), .C2(n9219), .ZN(P1_U3351) );
  INV_X1 U8089 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6374) );
  OAI222_X1 U8090 ( .A1(n8084), .A2(n6374), .B1(n9640), .B2(n6373), .C1(
        P1_U3086), .C2(n6617), .ZN(P1_U3354) );
  AND2_X1 U8091 ( .A1(n6375), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8092 ( .A1(n6375), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8093 ( .A1(n6375), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8094 ( .A1(n6375), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8095 ( .A1(n6375), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8096 ( .A1(n6375), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8097 ( .A1(n6375), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8098 ( .A1(n6375), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8099 ( .A1(n6375), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8100 ( .A1(n6375), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8101 ( .A1(n6375), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8102 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6377) );
  INV_X1 U8103 ( .A(n6376), .ZN(n6383) );
  OAI222_X1 U8104 ( .A1(n8084), .A2(n6377), .B1(n9640), .B2(n6383), .C1(
        P1_U3086), .C2(n9244), .ZN(P1_U3349) );
  INV_X1 U8105 ( .A(n6379), .ZN(n6380) );
  AOI22_X1 U8106 ( .A1(n6375), .A2(n4797), .B1(n6381), .B2(n6380), .ZN(
        P2_U3376) );
  INV_X1 U8107 ( .A(n9044), .ZN(n7576) );
  INV_X1 U8108 ( .A(n7576), .ZN(n9048) );
  OAI222_X1 U8109 ( .A1(n8533), .A2(P2_U3151), .B1(n9048), .B2(n6383), .C1(
        n6382), .C2(n9042), .ZN(P2_U3289) );
  OAI222_X1 U8110 ( .A1(n9042), .A2(n6385), .B1(n9048), .B2(n6384), .C1(n6529), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  OAI222_X1 U8111 ( .A1(n6649), .A2(P2_U3151), .B1(n9048), .B2(n6387), .C1(
        n6386), .C2(n9042), .ZN(P2_U3290) );
  INV_X1 U8112 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6389) );
  INV_X1 U8113 ( .A(n6388), .ZN(n6390) );
  OAI222_X1 U8114 ( .A1(n8084), .A2(n6389), .B1(n9640), .B2(n6390), .C1(
        P1_U3086), .C2(n6629), .ZN(P1_U3348) );
  INV_X1 U8115 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6391) );
  OAI222_X1 U8116 ( .A1(n9042), .A2(n6391), .B1(n9048), .B2(n6390), .C1(n4667), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  AND2_X1 U8117 ( .A1(n6375), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8118 ( .A1(n6375), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8119 ( .A1(n6375), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8120 ( .A1(n6375), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8121 ( .A1(n6375), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8122 ( .A1(n6375), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8123 ( .A1(n6375), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8124 ( .A1(n6375), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8125 ( .A1(n6375), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8126 ( .A1(n6375), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8127 ( .A1(n6375), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8128 ( .A1(n6375), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8129 ( .A1(n6375), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8130 ( .A1(n6375), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8131 ( .A1(n6375), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8132 ( .A1(n6375), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8133 ( .A1(n6375), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  INV_X1 U8134 ( .A(n6392), .ZN(n6394) );
  AOI22_X1 U8135 ( .A1(n9274), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9638), .ZN(n6393) );
  OAI21_X1 U8136 ( .B1(n6394), .B2(n9640), .A(n6393), .ZN(P1_U3347) );
  INV_X1 U8137 ( .A(n6868), .ZN(n6720) );
  OAI222_X1 U8138 ( .A1(n6720), .A2(P2_U3151), .B1(n9048), .B2(n6394), .C1(
        n10020), .C2(n9042), .ZN(P2_U3287) );
  INV_X1 U8139 ( .A(n6490), .ZN(n7578) );
  NOR2_X1 U8140 ( .A1(n6491), .A2(n7578), .ZN(n6395) );
  INV_X1 U8141 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6406) );
  NOR2_X1 U8142 ( .A1(n6257), .A2(P2_U3151), .ZN(n9045) );
  NAND2_X1 U8143 ( .A1(n6401), .A2(n9045), .ZN(n6446) );
  NOR2_X2 U8144 ( .A1(n8641), .A2(n6402), .ZN(n8683) );
  INV_X1 U8145 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6398) );
  INV_X2 U8146 ( .A(n8506), .ZN(n8665) );
  MUX2_X1 U8147 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8665), .Z(n6397) );
  MUX2_X1 U8148 ( .A(n6734), .B(n5886), .S(n8665), .Z(n6396) );
  AND2_X1 U8149 ( .A1(n6396), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6452) );
  AOI21_X1 U8150 ( .B1(n6398), .B2(n6397), .A(n6452), .ZN(n6399) );
  AOI21_X1 U8151 ( .B1(n6446), .B2(n8617), .A(n6399), .ZN(n6400) );
  AOI21_X1 U8152 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6400), .ZN(
        n6405) );
  NOR2_X1 U8153 ( .A1(n8665), .A2(P2_U3151), .ZN(n7735) );
  NAND2_X1 U8154 ( .A1(n6401), .A2(n7735), .ZN(n6403) );
  MUX2_X1 U8155 ( .A(n6403), .B(n8641), .S(n6402), .Z(n8673) );
  NAND2_X1 U8156 ( .A1(n8587), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6404) );
  OAI211_X1 U8157 ( .C1(n8653), .C2(n6406), .A(n6405), .B(n6404), .ZN(P2_U3182) );
  INV_X1 U8158 ( .A(n6407), .ZN(n6412) );
  INV_X1 U8159 ( .A(n9300), .ZN(n6408) );
  OAI222_X1 U8160 ( .A1(n9640), .A2(n6412), .B1(n6408), .B2(P1_U3086), .C1(
        n10071), .C2(n8084), .ZN(P1_U3346) );
  INV_X1 U8161 ( .A(n6409), .ZN(n6414) );
  AOI22_X1 U8162 ( .A1(n9651), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9638), .ZN(n6410) );
  OAI21_X1 U8163 ( .B1(n6414), .B2(n9640), .A(n6410), .ZN(P1_U3345) );
  INV_X1 U8164 ( .A(n6974), .ZN(n6990) );
  OAI222_X1 U8165 ( .A1(P2_U3151), .A2(n6990), .B1(n9048), .B2(n6412), .C1(
        n6411), .C2(n9042), .ZN(P2_U3286) );
  OAI222_X1 U8166 ( .A1(P2_U3151), .A2(n7149), .B1(n9048), .B2(n6414), .C1(
        n6413), .C2(n9042), .ZN(P2_U3285) );
  NAND2_X1 U8167 ( .A1(n6415), .A2(n6418), .ZN(n8327) );
  INV_X1 U8168 ( .A(n8327), .ZN(n6416) );
  NOR2_X1 U8169 ( .A1(n8878), .A2(n6416), .ZN(n8475) );
  NOR2_X1 U8170 ( .A1(n9884), .A2(n9902), .ZN(n6417) );
  OAI222_X1 U8171 ( .A1(n6418), .A2(n9886), .B1(n8475), .B2(n6417), .C1(n9919), 
        .C2(n6739), .ZN(n6571) );
  NAND2_X1 U8172 ( .A1(n6571), .A2(n9956), .ZN(n6419) );
  OAI21_X1 U8173 ( .B1(n9956), .B2(n5886), .A(n6419), .ZN(P2_U3459) );
  MUX2_X1 U8174 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8665), .Z(n6420) );
  XNOR2_X1 U8175 ( .A(n6420), .B(n6438), .ZN(n6453) );
  INV_X1 U8176 ( .A(n6420), .ZN(n6421) );
  OAI22_X1 U8177 ( .A1(n6453), .A2(n6452), .B1(n6461), .B2(n6421), .ZN(n6509)
         );
  MUX2_X1 U8178 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8665), .Z(n6422) );
  XNOR2_X1 U8179 ( .A(n6422), .B(n6430), .ZN(n6510) );
  AOI22_X1 U8180 ( .A1(n6509), .A2(n6510), .B1(n6422), .B2(n6520), .ZN(n6466)
         );
  MUX2_X1 U8181 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8665), .Z(n6423) );
  XOR2_X1 U8182 ( .A(n6478), .B(n6423), .Z(n6465) );
  NAND2_X1 U8183 ( .A1(n6466), .A2(n6465), .ZN(n6464) );
  INV_X1 U8184 ( .A(n6423), .ZN(n6425) );
  INV_X1 U8185 ( .A(n6478), .ZN(n6424) );
  NAND2_X1 U8186 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  AND2_X1 U8187 ( .A1(n6464), .A2(n6426), .ZN(n6428) );
  MUX2_X1 U8188 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8665), .Z(n6524) );
  INV_X1 U8189 ( .A(n6529), .ZN(n6527) );
  XNOR2_X1 U8190 ( .A(n6524), .B(n6527), .ZN(n6427) );
  NAND3_X1 U8191 ( .A1(n6464), .A2(n6426), .A3(n6427), .ZN(n6525) );
  OAI211_X1 U8192 ( .C1(n6428), .C2(n6427), .A(n8683), .B(n6525), .ZN(n6451)
         );
  MUX2_X1 U8193 ( .A(n5933), .B(P2_REG1_REG_4__SCAN_IN), .S(n6529), .Z(n6434)
         );
  INV_X1 U8194 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U8195 ( .A(n6430), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6511) );
  INV_X1 U8196 ( .A(n6431), .ZN(n6432) );
  AOI22_X1 U8197 ( .A1(n6468), .A2(P2_REG1_REG_3__SCAN_IN), .B1(n6478), .B2(
        n6432), .ZN(n6433) );
  AOI21_X1 U8198 ( .B1(n6434), .B2(n6433), .A(n6528), .ZN(n6436) );
  OR2_X1 U8199 ( .A1(n6446), .A2(n8506), .ZN(n8678) );
  INV_X1 U8200 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6435) );
  OAI22_X1 U8201 ( .A1(n6436), .A2(n8678), .B1(n8653), .B2(n6435), .ZN(n6449)
         );
  NOR2_X1 U8202 ( .A1(n6734), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8203 ( .A1(n5879), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6439) );
  INV_X1 U8204 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U8205 ( .A1(n6520), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8206 ( .A1(n6514), .A2(n6440), .ZN(n6441) );
  NAND2_X1 U8207 ( .A1(n6441), .A2(n6478), .ZN(n6444) );
  OAI21_X1 U8208 ( .B1(n6441), .B2(n6478), .A(n6444), .ZN(n6469) );
  NAND2_X1 U8209 ( .A1(n6471), .A2(n6444), .ZN(n6442) );
  INV_X1 U8210 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6753) );
  MUX2_X1 U8211 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6753), .S(n6529), .Z(n6443)
         );
  NAND2_X1 U8212 ( .A1(n6442), .A2(n6443), .ZN(n6531) );
  INV_X1 U8213 ( .A(n6443), .ZN(n6445) );
  NAND3_X1 U8214 ( .A1(n6471), .A2(n6445), .A3(n6444), .ZN(n6447) );
  AOI21_X1 U8215 ( .B1(n6531), .B2(n6447), .A(n8685), .ZN(n6448) );
  AND2_X1 U8216 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6689) );
  NOR3_X1 U8217 ( .A1(n6449), .A2(n6448), .A3(n6689), .ZN(n6450) );
  OAI211_X1 U8218 ( .C1(n8673), .C2(n6529), .A(n6451), .B(n6450), .ZN(P2_U3186) );
  XNOR2_X1 U8219 ( .A(n6453), .B(n6452), .ZN(n6463) );
  INV_X1 U8220 ( .A(n6454), .ZN(n6455) );
  AOI21_X1 U8221 ( .B1(n10102), .B2(n6456), .A(n6455), .ZN(n6457) );
  OAI22_X1 U8222 ( .A1(n8685), .A2(n6457), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8883), .ZN(n6460) );
  INV_X1 U8223 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9961) );
  XNOR2_X1 U8224 ( .A(n4277), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6458) );
  OAI22_X1 U8225 ( .A1(n8653), .A2(n9961), .B1(n8678), .B2(n6458), .ZN(n6459)
         );
  AOI211_X1 U8226 ( .C1(n6461), .C2(n8587), .A(n6460), .B(n6459), .ZN(n6462)
         );
  OAI21_X1 U8227 ( .B1(n8617), .B2(n6463), .A(n6462), .ZN(P2_U3183) );
  OAI21_X1 U8228 ( .B1(n6466), .B2(n6465), .A(n6464), .ZN(n6467) );
  NAND2_X1 U8229 ( .A1(n6467), .A2(n8683), .ZN(n6477) );
  XNOR2_X1 U8230 ( .A(n6468), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6475) );
  NOR2_X1 U8231 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5827), .ZN(n6545) );
  INV_X1 U8232 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8233 ( .A1(n6469), .A2(n6852), .ZN(n6470) );
  AND2_X1 U8234 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  OAI22_X1 U8235 ( .A1(n8653), .A2(n6473), .B1(n8685), .B2(n6472), .ZN(n6474)
         );
  AOI211_X1 U8236 ( .C1(n8624), .C2(n6475), .A(n6545), .B(n6474), .ZN(n6476)
         );
  OAI211_X1 U8237 ( .C1(n8673), .C2(n6478), .A(n6477), .B(n6476), .ZN(P2_U3185) );
  INV_X1 U8238 ( .A(n6731), .ZN(n6498) );
  NAND2_X1 U8239 ( .A1(n6481), .A2(n6498), .ZN(n6543) );
  INV_X1 U8240 ( .A(n6496), .ZN(n6480) );
  NAND2_X1 U8241 ( .A1(n6481), .A2(n6480), .ZN(n6485) );
  INV_X1 U8242 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8243 ( .A1(n6486), .A2(n6483), .ZN(n6484) );
  INV_X1 U8244 ( .A(n8475), .ZN(n6732) );
  NAND2_X1 U8245 ( .A1(n6486), .A2(n9940), .ZN(n6488) );
  AOI22_X1 U8246 ( .A1(n8272), .A2(n6732), .B1(n6736), .B2(n8259), .ZN(n6504)
         );
  AND3_X1 U8247 ( .A1(n6491), .A2(n6490), .A3(n6489), .ZN(n6495) );
  NAND2_X1 U8248 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  OAI211_X1 U8249 ( .C1(n6500), .C2(n6496), .A(n6495), .B(n6494), .ZN(n6497)
         );
  NAND2_X1 U8250 ( .A1(n6497), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8251 ( .A1(n6499), .A2(n6498), .ZN(n8507) );
  OR2_X1 U8252 ( .A1(n6500), .A2(n8507), .ZN(n6501) );
  NAND2_X1 U8253 ( .A1(n8287), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8254 ( .A1(n6583), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6503) );
  OAI211_X1 U8255 ( .C1(n6739), .C2(n8286), .A(n6504), .B(n6503), .ZN(P2_U3172) );
  INV_X1 U8256 ( .A(n6505), .ZN(n6508) );
  OAI222_X1 U8257 ( .A1(n7395), .A2(P2_U3151), .B1(n9048), .B2(n6508), .C1(
        n6506), .C2(n9042), .ZN(P2_U3284) );
  INV_X1 U8258 ( .A(n9695), .ZN(n6507) );
  OAI222_X1 U8259 ( .A1(n8084), .A2(n10128), .B1(n9640), .B2(n6508), .C1(
        P1_U3086), .C2(n6507), .ZN(P1_U3344) );
  XOR2_X1 U8260 ( .A(n6510), .B(n6509), .Z(n6522) );
  INV_X1 U8261 ( .A(n8653), .ZN(n8669) );
  XNOR2_X1 U8262 ( .A(n6512), .B(n6511), .ZN(n6513) );
  AOI22_X1 U8263 ( .A1(n8669), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8624), .B2(
        n6513), .ZN(n6519) );
  INV_X1 U8264 ( .A(n8685), .ZN(n6535) );
  OAI21_X1 U8265 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6517) );
  AOI22_X1 U8266 ( .A1(n6535), .A2(n6517), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6518) );
  OAI211_X1 U8267 ( .C1(n6520), .C2(n8673), .A(n6519), .B(n6518), .ZN(n6521)
         );
  AOI21_X1 U8268 ( .B1(n8683), .B2(n6522), .A(n6521), .ZN(n6523) );
  INV_X1 U8269 ( .A(n6523), .ZN(P2_U3184) );
  INV_X1 U8270 ( .A(n6524), .ZN(n6526) );
  OAI21_X1 U8271 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n6652) );
  MUX2_X1 U8272 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8665), .Z(n6650) );
  XOR2_X1 U8273 ( .A(n6649), .B(n6650), .Z(n6651) );
  XNOR2_X1 U8274 ( .A(n6652), .B(n6651), .ZN(n6541) );
  XOR2_X1 U8275 ( .A(n6664), .B(P2_REG1_REG_5__SCAN_IN), .Z(n6539) );
  INV_X1 U8276 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10124) );
  INV_X1 U8277 ( .A(n6649), .ZN(n6665) );
  NAND2_X1 U8278 ( .A1(n8587), .A2(n6665), .ZN(n6537) );
  NAND2_X1 U8279 ( .A1(n6529), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8280 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  NAND2_X1 U8281 ( .A1(n6532), .A2(n6649), .ZN(n8538) );
  NAND2_X1 U8282 ( .A1(n8540), .A2(n6533), .ZN(n6534) );
  AND2_X1 U8283 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6770) );
  AOI21_X1 U8284 ( .B1(n6535), .B2(n6534), .A(n6770), .ZN(n6536) );
  OAI211_X1 U8285 ( .C1(n10124), .C2(n8653), .A(n6537), .B(n6536), .ZN(n6538)
         );
  AOI21_X1 U8286 ( .B1(n6539), .B2(n8624), .A(n6538), .ZN(n6540) );
  OAI21_X1 U8287 ( .B1(n6541), .B2(n8617), .A(n6540), .ZN(P2_U3187) );
  INV_X1 U8288 ( .A(n9873), .ZN(n6764) );
  OAI22_X1 U8289 ( .A1(n6556), .A2(n8257), .B1(n8286), .B2(n6764), .ZN(n6544)
         );
  AOI211_X1 U8290 ( .C1(n5926), .C2(n8259), .A(n6545), .B(n6544), .ZN(n6566)
         );
  INV_X1 U8291 ( .A(n6546), .ZN(n8499) );
  NAND2_X1 U8292 ( .A1(n6547), .A2(n8462), .ZN(n6746) );
  AND2_X1 U8293 ( .A1(n6548), .A2(n6746), .ZN(n6549) );
  NAND2_X2 U8294 ( .A1(n6550), .A2(n6549), .ZN(n6679) );
  NOR2_X1 U8295 ( .A1(n6679), .A2(n6736), .ZN(n6551) );
  NAND2_X1 U8296 ( .A1(n6580), .A2(n6579), .ZN(n6555) );
  INV_X1 U8297 ( .A(n6552), .ZN(n6553) );
  NAND2_X1 U8298 ( .A1(n6553), .A2(n6739), .ZN(n6554) );
  NAND2_X1 U8299 ( .A1(n6555), .A2(n6554), .ZN(n6573) );
  XNOR2_X1 U8300 ( .A(n6679), .B(n6796), .ZN(n6557) );
  XNOR2_X1 U8301 ( .A(n6557), .B(n6556), .ZN(n6574) );
  NAND2_X1 U8302 ( .A1(n6573), .A2(n6574), .ZN(n6560) );
  INV_X1 U8303 ( .A(n6557), .ZN(n6558) );
  NAND2_X1 U8304 ( .A1(n6558), .A2(n6556), .ZN(n6559) );
  XNOR2_X1 U8305 ( .A(n6679), .B(n9877), .ZN(n6680) );
  XNOR2_X1 U8306 ( .A(n6680), .B(n8528), .ZN(n6562) );
  AOI21_X1 U8307 ( .B1(n6561), .B2(n6562), .A(n8280), .ZN(n6564) );
  INV_X1 U8308 ( .A(n6562), .ZN(n6563) );
  NAND2_X1 U8309 ( .A1(n6564), .A2(n6682), .ZN(n6565) );
  OAI211_X1 U8310 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8287), .A(n6566), .B(
        n6565), .ZN(P2_U3158) );
  NAND2_X1 U8311 ( .A1(n8051), .A2(n8054), .ZN(n6615) );
  NAND2_X1 U8312 ( .A1(n8041), .A2(n6567), .ZN(n6569) );
  AND2_X1 U8313 ( .A1(n6569), .A2(n6568), .ZN(n6614) );
  INV_X1 U8314 ( .A(n6614), .ZN(n6570) );
  AND2_X1 U8315 ( .A1(n6615), .A2(n6570), .ZN(n9683) );
  NOR2_X1 U8316 ( .A1(n9683), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8317 ( .A1(n6571), .A2(n9941), .ZN(n6572) );
  OAI21_X1 U8318 ( .B1(n5885), .B2(n9941), .A(n6572), .ZN(P2_U3390) );
  XOR2_X1 U8319 ( .A(n6573), .B(n6574), .Z(n6578) );
  INV_X1 U8320 ( .A(n6796), .ZN(n9862) );
  AOI22_X1 U8321 ( .A1(n8290), .A2(n9863), .B1(n9862), .B2(n8259), .ZN(n6575)
         );
  OAI21_X1 U8322 ( .B1(n5927), .B2(n8286), .A(n6575), .ZN(n6576) );
  AOI21_X1 U8323 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6583), .A(n6576), .ZN(
        n6577) );
  OAI21_X1 U8324 ( .B1(n8280), .B2(n6578), .A(n6577), .ZN(P2_U3177) );
  XOR2_X1 U8325 ( .A(n6580), .B(n6579), .Z(n6585) );
  AOI22_X1 U8326 ( .A1(n8290), .A2(n6415), .B1(n5883), .B2(n8259), .ZN(n6581)
         );
  OAI21_X1 U8327 ( .B1(n6556), .B2(n8286), .A(n6581), .ZN(n6582) );
  AOI21_X1 U8328 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6583), .A(n6582), .ZN(
        n6584) );
  OAI21_X1 U8329 ( .B1(n8280), .B2(n6585), .A(n6584), .ZN(P2_U3162) );
  INV_X1 U8330 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8331 ( .A1(n5518), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8332 ( .A1(n6586), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U8333 ( .A1(n6587), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6588) );
  INV_X1 U8334 ( .A(n8030), .ZN(n9329) );
  NAND2_X1 U8335 ( .A1(n9329), .A2(P1_U3973), .ZN(n6591) );
  OAI21_X1 U8336 ( .B1(P1_U3973), .B2(n6592), .A(n6591), .ZN(P1_U3585) );
  INV_X1 U8337 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8338 ( .A1(n7009), .A2(P1_U3973), .ZN(n6593) );
  OAI21_X1 U8339 ( .B1(P1_U3973), .B2(n6594), .A(n6593), .ZN(P1_U3554) );
  NAND2_X1 U8340 ( .A1(n9065), .A2(P1_U3973), .ZN(n6595) );
  OAI21_X1 U8341 ( .B1(n6124), .B2(P1_U3973), .A(n6595), .ZN(P1_U3574) );
  XNOR2_X1 U8342 ( .A(n9300), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6613) );
  INV_X1 U8343 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6596) );
  MUX2_X1 U8344 ( .A(n6596), .B(P1_REG1_REG_1__SCAN_IN), .S(n6617), .Z(n9195)
         );
  AND2_X1 U8345 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9194) );
  NAND2_X1 U8346 ( .A1(n9195), .A2(n9194), .ZN(n9193) );
  NAND2_X1 U8347 ( .A1(n9199), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8348 ( .A1(n9193), .A2(n6597), .ZN(n6782) );
  INV_X1 U8349 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6598) );
  XNOR2_X1 U8350 ( .A(n6784), .B(n6598), .ZN(n6783) );
  NAND2_X1 U8351 ( .A1(n6782), .A2(n6783), .ZN(n6781) );
  NAND2_X1 U8352 ( .A1(n6784), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8353 ( .A1(n6781), .A2(n6599), .ZN(n9212) );
  INV_X1 U8354 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6600) );
  XNOR2_X1 U8355 ( .A(n9207), .B(n6600), .ZN(n9213) );
  NAND2_X1 U8356 ( .A1(n9212), .A2(n9213), .ZN(n9211) );
  NAND2_X1 U8357 ( .A1(n9207), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U8358 ( .A1(n9211), .A2(n6601), .ZN(n9222) );
  INV_X1 U8359 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U8360 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6602), .S(n6623), .Z(n9223)
         );
  NAND2_X1 U8361 ( .A1(n9222), .A2(n9223), .ZN(n9221) );
  NAND2_X1 U8362 ( .A1(n6623), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8363 ( .A1(n9221), .A2(n6603), .ZN(n9239) );
  INV_X1 U8364 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6604) );
  XNOR2_X1 U8365 ( .A(n9234), .B(n6604), .ZN(n9240) );
  NAND2_X1 U8366 ( .A1(n9239), .A2(n9240), .ZN(n9238) );
  NAND2_X1 U8367 ( .A1(n9234), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8368 ( .A1(n9238), .A2(n6605), .ZN(n9253) );
  XNOR2_X1 U8369 ( .A(n9244), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U8370 ( .A1(n9253), .A2(n9254), .ZN(n9252) );
  INV_X1 U8371 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6606) );
  OR2_X1 U8372 ( .A1(n9244), .A2(n6606), .ZN(n6607) );
  NAND2_X1 U8373 ( .A1(n9252), .A2(n6607), .ZN(n9266) );
  INV_X1 U8374 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9849) );
  MUX2_X1 U8375 ( .A(n9849), .B(P1_REG1_REG_7__SCAN_IN), .S(n6629), .Z(n9267)
         );
  NAND2_X1 U8376 ( .A1(n9266), .A2(n9267), .ZN(n9265) );
  NAND2_X1 U8377 ( .A1(n9261), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8378 ( .A1(n9265), .A2(n6608), .ZN(n9276) );
  INV_X1 U8379 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6609) );
  XNOR2_X1 U8380 ( .A(n9274), .B(n6609), .ZN(n9277) );
  NAND2_X1 U8381 ( .A1(n9276), .A2(n9277), .ZN(n9275) );
  NAND2_X1 U8382 ( .A1(n9274), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U8383 ( .A1(n9275), .A2(n6610), .ZN(n6612) );
  OR2_X1 U8384 ( .A1(n6612), .A2(n6613), .ZN(n9302) );
  INV_X1 U8385 ( .A(n9302), .ZN(n6611) );
  AOI21_X1 U8386 ( .B1(n6613), .B2(n6612), .A(n6611), .ZN(n6641) );
  NAND2_X1 U8387 ( .A1(n6615), .A2(n6614), .ZN(n9685) );
  OR2_X1 U8388 ( .A1(n9685), .A2(n6773), .ZN(n9795) );
  INV_X1 U8389 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8390 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7522) );
  OAI21_X1 U8391 ( .B1(n9799), .B2(n6616), .A(n7522), .ZN(n6639) );
  INV_X1 U8392 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7062) );
  MUX2_X1 U8393 ( .A(n7062), .B(P1_REG2_REG_1__SCAN_IN), .S(n6617), .Z(n9198)
         );
  AND2_X1 U8394 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9197) );
  NAND2_X1 U8395 ( .A1(n9198), .A2(n9197), .ZN(n9196) );
  NAND2_X1 U8396 ( .A1(n9199), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8397 ( .A1(n9196), .A2(n6618), .ZN(n6779) );
  INV_X1 U8398 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6619) );
  XNOR2_X1 U8399 ( .A(n6784), .B(n6619), .ZN(n6780) );
  NAND2_X1 U8400 ( .A1(n6779), .A2(n6780), .ZN(n6778) );
  NAND2_X1 U8401 ( .A1(n6784), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8402 ( .A1(n6778), .A2(n6620), .ZN(n9209) );
  INV_X1 U8403 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6621) );
  XNOR2_X1 U8404 ( .A(n9207), .B(n6621), .ZN(n9210) );
  NAND2_X1 U8405 ( .A1(n9209), .A2(n9210), .ZN(n9208) );
  NAND2_X1 U8406 ( .A1(n9207), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8407 ( .A1(n9208), .A2(n6622), .ZN(n9225) );
  INV_X1 U8408 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7053) );
  MUX2_X1 U8409 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7053), .S(n6623), .Z(n9226)
         );
  NAND2_X1 U8410 ( .A1(n9225), .A2(n9226), .ZN(n9224) );
  NAND2_X1 U8411 ( .A1(n6623), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U8412 ( .A1(n9224), .A2(n6624), .ZN(n9236) );
  INV_X1 U8413 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6625) );
  XNOR2_X1 U8414 ( .A(n9234), .B(n6625), .ZN(n9237) );
  NAND2_X1 U8415 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
  NAND2_X1 U8416 ( .A1(n9234), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8417 ( .A1(n9235), .A2(n6626), .ZN(n9250) );
  XNOR2_X1 U8418 ( .A(n9244), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U8419 ( .A1(n9250), .A2(n9251), .ZN(n9249) );
  INV_X1 U8420 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6627) );
  OR2_X1 U8421 ( .A1(n9244), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8422 ( .A1(n9249), .A2(n6628), .ZN(n9263) );
  INV_X1 U8423 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6630) );
  MUX2_X1 U8424 ( .A(n6630), .B(P1_REG2_REG_7__SCAN_IN), .S(n6629), .Z(n9264)
         );
  NAND2_X1 U8425 ( .A1(n9263), .A2(n9264), .ZN(n9262) );
  NAND2_X1 U8426 ( .A1(n9261), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8427 ( .A1(n9262), .A2(n6631), .ZN(n9279) );
  INV_X1 U8428 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6632) );
  XNOR2_X1 U8429 ( .A(n9274), .B(n6632), .ZN(n9280) );
  NAND2_X1 U8430 ( .A1(n9279), .A2(n9280), .ZN(n9278) );
  NAND2_X1 U8431 ( .A1(n9274), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8432 ( .A1(n9278), .A2(n6633), .ZN(n6635) );
  XNOR2_X1 U8433 ( .A(n9300), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6634) );
  OR2_X1 U8434 ( .A1(n6635), .A2(n6634), .ZN(n9287) );
  NAND2_X1 U8435 ( .A1(n6635), .A2(n6634), .ZN(n6637) );
  NAND2_X1 U8436 ( .A1(n6773), .A2(n6636), .ZN(n8049) );
  AOI21_X1 U8437 ( .B1(n9287), .B2(n6637), .A(n9758), .ZN(n6638) );
  AOI211_X1 U8438 ( .C1(n9777), .C2(n9300), .A(n6639), .B(n6638), .ZN(n6640)
         );
  OAI21_X1 U8439 ( .B1(n6641), .B2(n9764), .A(n6640), .ZN(P1_U3252) );
  INV_X1 U8440 ( .A(n6642), .ZN(n6676) );
  AOI22_X1 U8441 ( .A1(n9699), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9638), .ZN(n6643) );
  OAI21_X1 U8442 ( .B1(n6676), .B2(n9640), .A(n6643), .ZN(P1_U3343) );
  INV_X1 U8443 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8444 ( .A1(n8177), .A2(P2_U3893), .ZN(n6644) );
  OAI21_X1 U8445 ( .B1(P2_U3893), .B2(n6645), .A(n6644), .ZN(P2_U3511) );
  INV_X1 U8446 ( .A(n8540), .ZN(n6647) );
  INV_X1 U8447 ( .A(n8538), .ZN(n6646) );
  XNOR2_X1 U8448 ( .A(n8533), .B(n6888), .ZN(n8537) );
  AOI21_X1 U8449 ( .B1(n6955), .B2(n6648), .A(n6698), .ZN(n6675) );
  AOI22_X1 U8450 ( .A1(n6652), .A2(n6651), .B1(n6650), .B2(n6649), .ZN(n8531)
         );
  MUX2_X1 U8451 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8665), .Z(n6653) );
  NOR2_X1 U8452 ( .A1(n6653), .A2(n8533), .ZN(n6654) );
  AOI21_X1 U8453 ( .B1(n6653), .B2(n8533), .A(n6654), .ZN(n8530) );
  NAND2_X1 U8454 ( .A1(n8531), .A2(n8530), .ZN(n8529) );
  INV_X1 U8455 ( .A(n6654), .ZN(n6660) );
  MUX2_X1 U8456 ( .A(n6955), .B(n6655), .S(n8665), .Z(n6656) );
  NAND2_X1 U8457 ( .A1(n6656), .A2(n6697), .ZN(n6703) );
  INV_X1 U8458 ( .A(n6656), .ZN(n6657) );
  NAND2_X1 U8459 ( .A1(n6657), .A2(n4667), .ZN(n6658) );
  NAND2_X1 U8460 ( .A1(n6703), .A2(n6658), .ZN(n6659) );
  AOI21_X1 U8461 ( .B1(n8529), .B2(n6660), .A(n6659), .ZN(n6709) );
  AND3_X1 U8462 ( .A1(n8529), .A2(n6660), .A3(n6659), .ZN(n6661) );
  OAI21_X1 U8463 ( .B1(n6709), .B2(n6661), .A(n8683), .ZN(n6674) );
  NAND2_X1 U8464 ( .A1(n8533), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6666) );
  MUX2_X1 U8465 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6662), .S(n8533), .Z(n8547)
         );
  NAND2_X1 U8466 ( .A1(n8547), .A2(n8548), .ZN(n8546) );
  NAND2_X1 U8467 ( .A1(n6666), .A2(n8546), .ZN(n6712) );
  OAI21_X1 U8468 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n6667), .A(n6713), .ZN(
        n6672) );
  INV_X1 U8469 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U8470 ( .A1(n8587), .A2(n6697), .ZN(n6669) );
  AND2_X1 U8471 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6936) );
  INV_X1 U8472 ( .A(n6936), .ZN(n6668) );
  OAI211_X1 U8473 ( .C1(n6670), .C2(n8653), .A(n6669), .B(n6668), .ZN(n6671)
         );
  AOI21_X1 U8474 ( .B1(n6672), .B2(n8624), .A(n6671), .ZN(n6673) );
  OAI211_X1 U8475 ( .C1(n6675), .C2(n8685), .A(n6674), .B(n6673), .ZN(P2_U3189) );
  INV_X1 U8476 ( .A(n7546), .ZN(n7410) );
  OAI222_X1 U8477 ( .A1(P2_U3151), .A2(n7410), .B1(n9044), .B2(n6676), .C1(
        n10132), .C2(n9042), .ZN(P2_U3283) );
  INV_X1 U8478 ( .A(n6677), .ZN(n6695) );
  AOI22_X1 U8479 ( .A1(n9715), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9638), .ZN(n6678) );
  OAI21_X1 U8480 ( .B1(n6695), .B2(n9640), .A(n6678), .ZN(P1_U3342) );
  XNOR2_X1 U8481 ( .A(n8131), .B(n9882), .ZN(n6763) );
  XNOR2_X1 U8482 ( .A(n6763), .B(n9873), .ZN(n6687) );
  NAND2_X1 U8483 ( .A1(n6680), .A2(n8528), .ZN(n6681) );
  INV_X1 U8484 ( .A(n6686), .ZN(n6684) );
  INV_X1 U8485 ( .A(n6687), .ZN(n6683) );
  INV_X1 U8486 ( .A(n6767), .ZN(n6685) );
  AOI21_X1 U8487 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(n6693) );
  OAI22_X1 U8488 ( .A1(n5927), .A2(n8257), .B1(n8286), .B2(n9894), .ZN(n6688)
         );
  AOI211_X1 U8489 ( .C1(n6751), .C2(n8259), .A(n6689), .B(n6688), .ZN(n6692)
         );
  INV_X1 U8490 ( .A(n6690), .ZN(n6750) );
  NAND2_X1 U8491 ( .A1(n8267), .A2(n6750), .ZN(n6691) );
  OAI211_X1 U8492 ( .C1(n6693), .C2(n8280), .A(n6692), .B(n6691), .ZN(P2_U3170) );
  INV_X1 U8493 ( .A(n7630), .ZN(n7636) );
  INV_X1 U8494 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6694) );
  OAI222_X1 U8495 ( .A1(n7636), .A2(P2_U3151), .B1(n9044), .B2(n6695), .C1(
        n6694), .C2(n9042), .ZN(P2_U3282) );
  NOR2_X1 U8496 ( .A1(n6697), .A2(n6696), .ZN(n6699) );
  NOR2_X1 U8497 ( .A1(n6699), .A2(n6698), .ZN(n6702) );
  INV_X1 U8498 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6969) );
  MUX2_X1 U8499 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6969), .S(n6868), .Z(n6701)
         );
  INV_X1 U8500 ( .A(n6857), .ZN(n6700) );
  AOI21_X1 U8501 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(n6725) );
  INV_X1 U8502 ( .A(n6703), .ZN(n6708) );
  MUX2_X1 U8503 ( .A(n6969), .B(n6715), .S(n8665), .Z(n6704) );
  NAND2_X1 U8504 ( .A1(n6704), .A2(n6868), .ZN(n6864) );
  INV_X1 U8505 ( .A(n6704), .ZN(n6705) );
  NAND2_X1 U8506 ( .A1(n6705), .A2(n6720), .ZN(n6706) );
  AND2_X1 U8507 ( .A1(n6864), .A2(n6706), .ZN(n6707) );
  OAI21_X1 U8508 ( .B1(n6709), .B2(n6708), .A(n6707), .ZN(n6865) );
  INV_X1 U8509 ( .A(n6865), .ZN(n6711) );
  NOR3_X1 U8510 ( .A1(n6709), .A2(n6708), .A3(n6707), .ZN(n6710) );
  OAI21_X1 U8511 ( .B1(n6711), .B2(n6710), .A(n8683), .ZN(n6724) );
  NAND2_X1 U8512 ( .A1(n4667), .A2(n6712), .ZN(n6714) );
  MUX2_X1 U8513 ( .A(n6715), .B(P2_REG1_REG_8__SCAN_IN), .S(n6868), .Z(n6716)
         );
  OAI21_X1 U8514 ( .B1(n6717), .B2(n6716), .A(n6867), .ZN(n6722) );
  INV_X1 U8515 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U8516 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6718), .ZN(n7115) );
  AOI21_X1 U8517 ( .B1(n8669), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7115), .ZN(
        n6719) );
  OAI21_X1 U8518 ( .B1(n6720), .B2(n8673), .A(n6719), .ZN(n6721) );
  AOI21_X1 U8519 ( .B1(n6722), .B2(n8624), .A(n6721), .ZN(n6723) );
  OAI211_X1 U8520 ( .C1(n6725), .C2(n8685), .A(n6724), .B(n6723), .ZN(P2_U3190) );
  MUX2_X1 U8521 ( .A(n6728), .B(n6727), .S(n6726), .Z(n6730) );
  NAND2_X1 U8522 ( .A1(n6730), .A2(n6729), .ZN(n6735) );
  NAND2_X1 U8523 ( .A1(n8859), .A2(n9872), .ZN(n8727) );
  NAND3_X1 U8524 ( .A1(n6732), .A2(n6731), .A3(n9886), .ZN(n6733) );
  MUX2_X1 U8525 ( .A(n6734), .B(n6733), .S(n8859), .Z(n6738) );
  INV_X1 U8526 ( .A(n6735), .ZN(n6748) );
  INV_X1 U8527 ( .A(n8752), .ZN(n8871) );
  NAND2_X1 U8528 ( .A1(n6748), .A2(n8871), .ZN(n8885) );
  AOI22_X1 U8529 ( .A1(n8861), .A2(n6736), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8848), .ZN(n6737) );
  OAI211_X1 U8530 ( .C1(n6739), .C2(n8727), .A(n6738), .B(n6737), .ZN(P2_U3233) );
  INV_X1 U8531 ( .A(n6740), .ZN(n6762) );
  AOI22_X1 U8532 ( .A1(n9731), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9638), .ZN(n6741) );
  OAI21_X1 U8533 ( .B1(n6762), .B2(n9640), .A(n6741), .ZN(P1_U3341) );
  INV_X1 U8534 ( .A(n6803), .ZN(n6743) );
  OR2_X1 U8535 ( .A1(n6743), .A2(n8341), .ZN(n8477) );
  XNOR2_X1 U8536 ( .A(n6742), .B(n8477), .ZN(n6744) );
  AOI222_X1 U8537 ( .A1(n9902), .A2(n6744), .B1(n8527), .B2(n9872), .C1(n8528), 
        .C2(n9874), .ZN(n9881) );
  INV_X1 U8538 ( .A(n8477), .ZN(n8338) );
  XNOR2_X1 U8539 ( .A(n6745), .B(n8338), .ZN(n9885) );
  NOR2_X1 U8540 ( .A1(n4274), .A2(n6746), .ZN(n6747) );
  NAND2_X1 U8541 ( .A1(n6748), .A2(n6747), .ZN(n8700) );
  NAND2_X1 U8542 ( .A1(n8700), .A2(n9866), .ZN(n6749) );
  NAND2_X1 U8543 ( .A1(n6749), .A2(n8859), .ZN(n8864) );
  INV_X1 U8544 ( .A(n8864), .ZN(n8872) );
  AOI22_X1 U8545 ( .A1(n8861), .A2(n6751), .B1(n8848), .B2(n6750), .ZN(n6752)
         );
  OAI21_X1 U8546 ( .B1(n6753), .B2(n8859), .A(n6752), .ZN(n6754) );
  AOI21_X1 U8547 ( .B1(n9885), .B2(n8872), .A(n6754), .ZN(n6755) );
  OAI21_X1 U8548 ( .B1(n9881), .B2(n8890), .A(n6755), .ZN(P2_U3229) );
  XOR2_X1 U8549 ( .A(n6756), .B(n6757), .Z(n6777) );
  AOI22_X1 U8550 ( .A1(n6777), .A2(n9151), .B1(n9152), .B2(n5683), .ZN(n6760)
         );
  OR2_X1 U8551 ( .A1(n6758), .A2(n8051), .ZN(n8074) );
  AOI22_X1 U8552 ( .A1(n9675), .A2(n7008), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8074), .ZN(n6759) );
  NAND2_X1 U8553 ( .A1(n6760), .A2(n6759), .ZN(P1_U3232) );
  OAI222_X1 U8554 ( .A1(n8554), .A2(P2_U3151), .B1(n9044), .B2(n6762), .C1(
        n6761), .C2(n9042), .ZN(P2_U3281) );
  INV_X1 U8555 ( .A(n6763), .ZN(n6765) );
  NAND2_X1 U8556 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  XNOR2_X1 U8557 ( .A(n8131), .B(n9887), .ZN(n6913) );
  XNOR2_X1 U8558 ( .A(n6913), .B(n9894), .ZN(n6911) );
  XNOR2_X1 U8559 ( .A(n6911), .B(n6912), .ZN(n6768) );
  NAND2_X1 U8560 ( .A1(n6768), .A2(n8272), .ZN(n6772) );
  OAI22_X1 U8561 ( .A1(n8293), .A2(n9887), .B1(n8286), .B2(n9904), .ZN(n6769)
         );
  AOI211_X1 U8562 ( .C1(n8290), .C2(n9873), .A(n6770), .B(n6769), .ZN(n6771)
         );
  OAI211_X1 U8563 ( .C1(n6814), .C2(n8287), .A(n6772), .B(n6771), .ZN(P2_U3167) );
  NAND2_X1 U8564 ( .A1(n6773), .A2(n9681), .ZN(n6776) );
  INV_X1 U8565 ( .A(n8049), .ZN(n6774) );
  OAI21_X1 U8566 ( .B1(n9681), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6773), .ZN(
        n9679) );
  AOI22_X1 U8567 ( .A1(n6774), .A2(n9197), .B1(n9679), .B2(n4464), .ZN(n6775)
         );
  OAI211_X1 U8568 ( .C1(n6777), .C2(n6776), .A(P1_U3973), .B(n6775), .ZN(n9230) );
  INV_X1 U8569 ( .A(n9230), .ZN(n6790) );
  OAI211_X1 U8570 ( .C1(n6780), .C2(n6779), .A(n9784), .B(n6778), .ZN(n6788)
         );
  OAI211_X1 U8571 ( .C1(n6783), .C2(n6782), .A(n9788), .B(n6781), .ZN(n6787)
         );
  AOI22_X1 U8572 ( .A1(n9683), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6786) );
  NAND2_X1 U8573 ( .A1(n9777), .A2(n6784), .ZN(n6785) );
  NAND4_X1 U8574 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6789)
         );
  OR2_X1 U8575 ( .A1(n6790), .A2(n6789), .ZN(P1_U3245) );
  INV_X1 U8576 ( .A(n9866), .ZN(n9928) );
  INV_X1 U8577 ( .A(n8700), .ZN(n6817) );
  AOI21_X1 U8578 ( .B1(n9928), .B2(n8859), .A(n6817), .ZN(n8876) );
  XNOR2_X1 U8579 ( .A(n6791), .B(n6793), .ZN(n9867) );
  XNOR2_X1 U8580 ( .A(n6793), .B(n6792), .ZN(n6794) );
  NAND2_X1 U8581 ( .A1(n6794), .A2(n9902), .ZN(n9865) );
  OAI22_X1 U8582 ( .A1(n6796), .A2(n8752), .B1(n8882), .B2(n6795), .ZN(n6797)
         );
  INV_X1 U8583 ( .A(n6797), .ZN(n6798) );
  NAND2_X1 U8584 ( .A1(n9865), .A2(n6798), .ZN(n6799) );
  MUX2_X1 U8585 ( .A(n6799), .B(P2_REG2_REG_2__SCAN_IN), .S(n8890), .Z(n6800)
         );
  INV_X1 U8586 ( .A(n6800), .ZN(n6802) );
  NAND2_X1 U8587 ( .A1(n8859), .A2(n9874), .ZN(n8830) );
  INV_X1 U8588 ( .A(n8830), .ZN(n8880) );
  INV_X1 U8589 ( .A(n8727), .ZN(n8887) );
  AOI22_X1 U8590 ( .A1(n8880), .A2(n9863), .B1(n8887), .B2(n8528), .ZN(n6801)
         );
  OAI211_X1 U8591 ( .C1(n8876), .C2(n9867), .A(n6802), .B(n6801), .ZN(P2_U3231) );
  NAND2_X1 U8592 ( .A1(n6804), .A2(n6803), .ZN(n6805) );
  XNOR2_X1 U8593 ( .A(n6805), .B(n8476), .ZN(n9890) );
  NAND2_X1 U8594 ( .A1(n9890), .A2(n9928), .ZN(n6813) );
  OAI21_X1 U8595 ( .B1(n6807), .B2(n8476), .A(n6806), .ZN(n6811) );
  NAND2_X1 U8596 ( .A1(n8526), .A2(n9872), .ZN(n6809) );
  NAND2_X1 U8597 ( .A1(n9873), .A2(n9874), .ZN(n6808) );
  NAND2_X1 U8598 ( .A1(n6809), .A2(n6808), .ZN(n6810) );
  AOI21_X1 U8599 ( .B1(n6811), .B2(n9902), .A(n6810), .ZN(n6812) );
  AND2_X1 U8600 ( .A1(n6813), .A2(n6812), .ZN(n9892) );
  NOR2_X1 U8601 ( .A1(n8885), .A2(n9887), .ZN(n6816) );
  OAI22_X1 U8602 ( .A1(n8859), .A2(n5942), .B1(n6814), .B2(n8882), .ZN(n6815)
         );
  AOI211_X1 U8603 ( .C1(n9890), .C2(n6817), .A(n6816), .B(n6815), .ZN(n6818)
         );
  OAI21_X1 U8604 ( .B1(n9892), .B2(n8890), .A(n6818), .ZN(P2_U3228) );
  INV_X1 U8605 ( .A(n6819), .ZN(n6827) );
  INV_X1 U8606 ( .A(n9754), .ZN(n9307) );
  OAI222_X1 U8607 ( .A1(n9640), .A2(n6827), .B1(n9307), .B2(P1_U3086), .C1(
        n6820), .C2(n8084), .ZN(P1_U3340) );
  XOR2_X1 U8608 ( .A(n6822), .B(n6821), .Z(n6826) );
  NOR2_X1 U8609 ( .A1(n9157), .A2(n7910), .ZN(n6824) );
  OAI22_X1 U8610 ( .A1(n6832), .A2(n9662), .B1(n9661), .B2(n6833), .ZN(n6823)
         );
  AOI211_X1 U8611 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n8074), .A(n6824), .B(
        n6823), .ZN(n6825) );
  OAI21_X1 U8612 ( .B1(n9671), .B2(n6826), .A(n6825), .ZN(P1_U3237) );
  INV_X1 U8613 ( .A(n8577), .ZN(n8582) );
  OAI222_X1 U8614 ( .A1(P2_U3151), .A2(n8582), .B1(n9044), .B2(n6827), .C1(
        n10006), .C2(n9042), .ZN(P2_U3280) );
  OR2_X1 U8615 ( .A1(n6839), .A2(n7910), .ZN(n6829) );
  AND3_X1 U8616 ( .A1(n6879), .A2(n9551), .A3(n6829), .ZN(n7105) );
  INV_X1 U8617 ( .A(n9504), .ZN(n9453) );
  XNOR2_X1 U8618 ( .A(n6830), .B(n7991), .ZN(n6831) );
  OAI222_X1 U8619 ( .A1(n9458), .A2(n6833), .B1(n9456), .B2(n6832), .C1(n9453), 
        .C2(n6831), .ZN(n7104) );
  AOI211_X1 U8620 ( .C1(n9835), .C2(n7109), .A(n7105), .B(n7104), .ZN(n7347)
         );
  AOI22_X1 U8621 ( .A1(n7450), .A2(n6834), .B1(n5802), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6835) );
  OAI21_X1 U8622 ( .B1(n7347), .B2(n5802), .A(n6835), .ZN(P1_U3524) );
  OAI21_X1 U8623 ( .B1(n6836), .B2(n6838), .A(n6837), .ZN(n7066) );
  AOI211_X1 U8624 ( .C1(n7008), .C2(n6843), .A(n9509), .B(n6839), .ZN(n7065)
         );
  XNOR2_X1 U8625 ( .A(n7010), .B(n6836), .ZN(n6842) );
  INV_X1 U8626 ( .A(n7009), .ZN(n6840) );
  OAI22_X1 U8627 ( .A1(n6881), .A2(n9458), .B1(n6840), .B2(n9456), .ZN(n8075)
         );
  INV_X1 U8628 ( .A(n8075), .ZN(n6841) );
  OAI21_X1 U8629 ( .B1(n6842), .B2(n9453), .A(n6841), .ZN(n7060) );
  AOI211_X1 U8630 ( .C1(n9835), .C2(n7066), .A(n7065), .B(n7060), .ZN(n7340)
         );
  AOI22_X1 U8631 ( .A1(n7450), .A2(n6843), .B1(n5802), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6844) );
  OAI21_X1 U8632 ( .B1(n7340), .B2(n5802), .A(n6844), .ZN(P1_U3523) );
  NAND2_X1 U8633 ( .A1(n9170), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6845) );
  OAI21_X1 U8634 ( .B1(n6846), .B2(n9170), .A(n6845), .ZN(P1_U3583) );
  XNOR2_X1 U8635 ( .A(n6847), .B(n8473), .ZN(n9879) );
  INV_X1 U8636 ( .A(n9879), .ZN(n6855) );
  XNOR2_X1 U8637 ( .A(n6849), .B(n6848), .ZN(n9871) );
  AOI22_X1 U8638 ( .A1(n8880), .A2(n5910), .B1(n8887), .B2(n9873), .ZN(n6851)
         );
  AOI22_X1 U8639 ( .A1(n8861), .A2(n5926), .B1(n5827), .B2(n8848), .ZN(n6850)
         );
  OAI211_X1 U8640 ( .C1(n6852), .C2(n8859), .A(n6851), .B(n6850), .ZN(n6853)
         );
  AOI21_X1 U8641 ( .B1(n8826), .B2(n9871), .A(n6853), .ZN(n6854) );
  OAI21_X1 U8642 ( .B1(n6855), .B2(n8864), .A(n6854), .ZN(P2_U3230) );
  OR2_X1 U8643 ( .A1(n6868), .A2(n6969), .ZN(n6856) );
  AOI21_X1 U8644 ( .B1(n7036), .B2(n6858), .A(n6975), .ZN(n6875) );
  MUX2_X1 U8645 ( .A(n7036), .B(n6859), .S(n8665), .Z(n6860) );
  NAND2_X1 U8646 ( .A1(n6860), .A2(n6974), .ZN(n6980) );
  INV_X1 U8647 ( .A(n6860), .ZN(n6861) );
  NAND2_X1 U8648 ( .A1(n6861), .A2(n6990), .ZN(n6862) );
  NAND2_X1 U8649 ( .A1(n6980), .A2(n6862), .ZN(n6863) );
  AOI21_X1 U8650 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6986) );
  AND3_X1 U8651 ( .A1(n6865), .A2(n6864), .A3(n6863), .ZN(n6866) );
  OAI21_X1 U8652 ( .B1(n6986), .B2(n6866), .A(n8683), .ZN(n6874) );
  NAND2_X1 U8653 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n6869), .ZN(n6991) );
  OAI21_X1 U8654 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n6869), .A(n6991), .ZN(
        n6872) );
  AND2_X1 U8655 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7213) );
  AOI21_X1 U8656 ( .B1(n8669), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7213), .ZN(
        n6870) );
  OAI21_X1 U8657 ( .B1(n6990), .B2(n8673), .A(n6870), .ZN(n6871) );
  AOI21_X1 U8658 ( .B1(n6872), .B2(n8624), .A(n6871), .ZN(n6873) );
  OAI211_X1 U8659 ( .C1(n6875), .C2(n8685), .A(n6874), .B(n6873), .ZN(P2_U3191) );
  OAI21_X1 U8660 ( .B1(n6877), .B2(n7990), .A(n6876), .ZN(n7272) );
  INV_X1 U8661 ( .A(n6905), .ZN(n6878) );
  AOI211_X1 U8662 ( .C1(n6899), .C2(n6879), .A(n9509), .B(n6878), .ZN(n7267)
         );
  XNOR2_X1 U8663 ( .A(n7990), .B(n6880), .ZN(n6883) );
  OAI22_X1 U8664 ( .A1(n6881), .A2(n9456), .B1(n7132), .B2(n9458), .ZN(n6898)
         );
  INV_X1 U8665 ( .A(n6898), .ZN(n6882) );
  OAI21_X1 U8666 ( .B1(n6883), .B2(n9453), .A(n6882), .ZN(n7266) );
  AOI211_X1 U8667 ( .C1(n9835), .C2(n7272), .A(n7267), .B(n7266), .ZN(n7343)
         );
  OAI22_X1 U8668 ( .A1(n9590), .A2(n5686), .B1(n9854), .B2(n6600), .ZN(n6884)
         );
  INV_X1 U8669 ( .A(n6884), .ZN(n6885) );
  OAI21_X1 U8670 ( .B1(n7343), .B2(n5802), .A(n6885), .ZN(P1_U3525) );
  NAND2_X1 U8671 ( .A1(n9112), .A2(P1_U3973), .ZN(n6886) );
  OAI21_X1 U8672 ( .B1(n6166), .B2(P1_U3973), .A(n6886), .ZN(P1_U3579) );
  XNOR2_X1 U8673 ( .A(n6887), .B(n8478), .ZN(n9901) );
  OAI22_X1 U8674 ( .A1(n8859), .A2(n6888), .B1(n6922), .B2(n8882), .ZN(n6889)
         );
  AOI21_X1 U8675 ( .B1(n8887), .B2(n8525), .A(n6889), .ZN(n6891) );
  NAND2_X1 U8676 ( .A1(n8861), .A2(n9897), .ZN(n6890) );
  OAI211_X1 U8677 ( .C1(n9894), .C2(n8830), .A(n6891), .B(n6890), .ZN(n6894)
         );
  XNOR2_X1 U8678 ( .A(n6892), .B(n8478), .ZN(n9899) );
  NOR2_X1 U8679 ( .A1(n9899), .A2(n8864), .ZN(n6893) );
  AOI211_X1 U8680 ( .C1(n8826), .C2(n9901), .A(n6894), .B(n6893), .ZN(n6895)
         );
  INV_X1 U8681 ( .A(n6895), .ZN(P2_U3227) );
  XOR2_X1 U8682 ( .A(n6897), .B(n6896), .Z(n6902) );
  AOI22_X1 U8683 ( .A1(n9675), .A2(n6899), .B1(n9066), .B2(n6898), .ZN(n6901)
         );
  MUX2_X1 U8684 ( .A(n9678), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6900) );
  OAI211_X1 U8685 ( .C1(n6902), .C2(n9671), .A(n6901), .B(n6900), .ZN(P1_U3218) );
  OAI21_X1 U8686 ( .B1(n6904), .B2(n7997), .A(n6903), .ZN(n7050) );
  AOI211_X1 U8687 ( .C1(n6909), .C2(n6905), .A(n9509), .B(n7199), .ZN(n7056)
         );
  XNOR2_X1 U8688 ( .A(n6906), .B(n7997), .ZN(n6908) );
  AND2_X1 U8689 ( .A1(n9191), .A2(n9425), .ZN(n6907) );
  AOI21_X1 U8690 ( .B1(n9189), .B2(n9427), .A(n6907), .ZN(n7090) );
  OAI21_X1 U8691 ( .B1(n6908), .B2(n9453), .A(n7090), .ZN(n7051) );
  AOI211_X1 U8692 ( .C1(n9835), .C2(n7050), .A(n7056), .B(n7051), .ZN(n7332)
         );
  AOI22_X1 U8693 ( .A1(n7450), .A2(n6909), .B1(n5802), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6910) );
  OAI21_X1 U8694 ( .B1(n7332), .B2(n5802), .A(n6910), .ZN(P1_U3526) );
  XNOR2_X1 U8695 ( .A(n8131), .B(n9897), .ZN(n6930) );
  XNOR2_X1 U8696 ( .A(n6930), .B(n9904), .ZN(n6920) );
  INV_X1 U8697 ( .A(n6913), .ZN(n6914) );
  NAND2_X1 U8698 ( .A1(n6914), .A2(n9894), .ZN(n6915) );
  INV_X1 U8699 ( .A(n6919), .ZN(n6917) );
  INV_X1 U8700 ( .A(n6933), .ZN(n6918) );
  AOI211_X1 U8701 ( .C1(n6920), .C2(n6919), .A(n8280), .B(n6918), .ZN(n6929)
         );
  INV_X1 U8702 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8703 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6921), .ZN(n8534) );
  AOI21_X1 U8704 ( .B1(n8290), .B2(n8527), .A(n8534), .ZN(n6927) );
  NAND2_X1 U8705 ( .A1(n8259), .A2(n9897), .ZN(n6926) );
  INV_X1 U8706 ( .A(n6922), .ZN(n6923) );
  NAND2_X1 U8707 ( .A1(n8267), .A2(n6923), .ZN(n6925) );
  NAND2_X1 U8708 ( .A1(n8277), .A2(n8525), .ZN(n6924) );
  NAND4_X1 U8709 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n6928)
         );
  OR2_X1 U8710 ( .A1(n6929), .A2(n6928), .ZN(P2_U3179) );
  INV_X1 U8711 ( .A(n6930), .ZN(n6931) );
  NAND2_X1 U8712 ( .A1(n6931), .A2(n8526), .ZN(n6932) );
  XNOR2_X1 U8713 ( .A(n6937), .B(n8131), .ZN(n7112) );
  XNOR2_X1 U8714 ( .A(n7112), .B(n9895), .ZN(n6934) );
  OAI21_X1 U8715 ( .B1(n6935), .B2(n6934), .A(n7114), .ZN(n6944) );
  AOI21_X1 U8716 ( .B1(n8290), .B2(n8526), .A(n6936), .ZN(n6942) );
  INV_X1 U8717 ( .A(n6937), .ZN(n9906) );
  NAND2_X1 U8718 ( .A1(n8259), .A2(n9906), .ZN(n6941) );
  INV_X1 U8719 ( .A(n6938), .ZN(n6956) );
  NAND2_X1 U8720 ( .A1(n8267), .A2(n6956), .ZN(n6940) );
  NAND2_X1 U8721 ( .A1(n8277), .A2(n8524), .ZN(n6939) );
  NAND4_X1 U8722 ( .A1(n6942), .A2(n6941), .A3(n6940), .A4(n6939), .ZN(n6943)
         );
  AOI21_X1 U8723 ( .B1(n6944), .B2(n8272), .A(n6943), .ZN(n6945) );
  INV_X1 U8724 ( .A(n6945), .ZN(P2_U3153) );
  INV_X1 U8725 ( .A(n8612), .ZN(n8593) );
  INV_X1 U8726 ( .A(n6946), .ZN(n6948) );
  OAI222_X1 U8727 ( .A1(P2_U3151), .A2(n8593), .B1(n9044), .B2(n6948), .C1(
        n6947), .C2(n9042), .ZN(P2_U3279) );
  INV_X1 U8728 ( .A(n9309), .ZN(n9763) );
  OAI222_X1 U8729 ( .A1(n8084), .A2(n10114), .B1(n9763), .B2(P1_U3086), .C1(
        n9640), .C2(n6948), .ZN(P1_U3339) );
  INV_X1 U8730 ( .A(n6962), .ZN(n6949) );
  AOI21_X1 U8731 ( .B1(n6950), .B2(n6952), .A(n6949), .ZN(n9911) );
  INV_X1 U8732 ( .A(n9911), .ZN(n9908) );
  INV_X1 U8733 ( .A(n6952), .ZN(n8482) );
  XNOR2_X1 U8734 ( .A(n6951), .B(n8482), .ZN(n6953) );
  NOR2_X1 U8735 ( .A1(n6953), .A2(n8917), .ZN(n9910) );
  INV_X1 U8736 ( .A(n9910), .ZN(n6954) );
  MUX2_X1 U8737 ( .A(n6955), .B(n6954), .S(n8859), .Z(n6960) );
  AOI22_X1 U8738 ( .A1(n8887), .A2(n8524), .B1(n8848), .B2(n6956), .ZN(n6957)
         );
  OAI21_X1 U8739 ( .B1(n9904), .B2(n8830), .A(n6957), .ZN(n6958) );
  AOI21_X1 U8740 ( .B1(n8861), .B2(n9906), .A(n6958), .ZN(n6959) );
  OAI211_X1 U8741 ( .C1(n9908), .C2(n8876), .A(n6960), .B(n6959), .ZN(P2_U3226) );
  NAND2_X1 U8742 ( .A1(n6962), .A2(n6961), .ZN(n6963) );
  XNOR2_X1 U8743 ( .A(n6963), .B(n8481), .ZN(n9913) );
  NAND2_X1 U8744 ( .A1(n6964), .A2(n8481), .ZN(n6965) );
  NAND3_X1 U8745 ( .A1(n6966), .A2(n9902), .A3(n6965), .ZN(n6968) );
  AOI22_X1 U8746 ( .A1(n9874), .A2(n8525), .B1(n8523), .B2(n9872), .ZN(n6967)
         );
  NAND2_X1 U8747 ( .A1(n6968), .A2(n6967), .ZN(n9915) );
  NAND2_X1 U8748 ( .A1(n9915), .A2(n8859), .ZN(n6972) );
  OAI22_X1 U8749 ( .A1(n8859), .A2(n6969), .B1(n7116), .B2(n8882), .ZN(n6970)
         );
  AOI21_X1 U8750 ( .B1(n8861), .B2(n9916), .A(n6970), .ZN(n6971) );
  OAI211_X1 U8751 ( .C1(n9913), .C2(n8864), .A(n6972), .B(n6971), .ZN(P2_U3225) );
  NOR2_X1 U8752 ( .A1(n6974), .A2(n6973), .ZN(n6976) );
  NOR2_X1 U8753 ( .A1(n6976), .A2(n6975), .ZN(n6979) );
  INV_X1 U8754 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7145) );
  MUX2_X1 U8755 ( .A(n7145), .B(P2_REG2_REG_10__SCAN_IN), .S(n7149), .Z(n6978)
         );
  INV_X1 U8756 ( .A(n7151), .ZN(n6977) );
  AOI21_X1 U8757 ( .B1(n6979), .B2(n6978), .A(n6977), .ZN(n7002) );
  INV_X1 U8758 ( .A(n6980), .ZN(n6985) );
  MUX2_X1 U8759 ( .A(n7145), .B(n6993), .S(n8665), .Z(n6981) );
  NAND2_X1 U8760 ( .A1(n6981), .A2(n7154), .ZN(n7165) );
  INV_X1 U8761 ( .A(n6981), .ZN(n6982) );
  NAND2_X1 U8762 ( .A1(n6982), .A2(n7149), .ZN(n6983) );
  AND2_X1 U8763 ( .A1(n7165), .A2(n6983), .ZN(n6984) );
  OAI21_X1 U8764 ( .B1(n6986), .B2(n6985), .A(n6984), .ZN(n7166) );
  INV_X1 U8765 ( .A(n7166), .ZN(n6988) );
  NOR3_X1 U8766 ( .A1(n6986), .A2(n6985), .A3(n6984), .ZN(n6987) );
  OAI21_X1 U8767 ( .B1(n6988), .B2(n6987), .A(n8683), .ZN(n7001) );
  NAND2_X1 U8768 ( .A1(n6990), .A2(n6989), .ZN(n6992) );
  MUX2_X1 U8769 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6993), .S(n7149), .Z(n6994)
         );
  OAI21_X1 U8770 ( .B1(n6995), .B2(n6994), .A(n7153), .ZN(n6999) );
  INV_X1 U8771 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6996) );
  NOR2_X1 U8772 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6996), .ZN(n7362) );
  AOI21_X1 U8773 ( .B1(n8669), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7362), .ZN(
        n6997) );
  OAI21_X1 U8774 ( .B1(n7149), .B2(n8673), .A(n6997), .ZN(n6998) );
  AOI21_X1 U8775 ( .B1(n6999), .B2(n8624), .A(n6998), .ZN(n7000) );
  OAI211_X1 U8776 ( .C1(n7002), .C2(n8685), .A(n7001), .B(n7000), .ZN(P2_U3192) );
  INV_X1 U8777 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7016) );
  NAND3_X1 U8778 ( .A1(n7005), .A2(n7004), .A3(n7003), .ZN(n7006) );
  NOR2_X1 U8779 ( .A1(n9806), .A2(n9509), .ZN(n9432) );
  OR2_X2 U8780 ( .A1(n9813), .A2(n7007), .ZN(n9516) );
  INV_X1 U8781 ( .A(n9516), .ZN(n9803) );
  OAI21_X1 U8782 ( .B1(n9432), .B2(n9803), .A(n7008), .ZN(n7015) );
  INV_X1 U8783 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7012) );
  AND2_X1 U8784 ( .A1(n7009), .A2(n7029), .ZN(n7911) );
  NOR2_X1 U8785 ( .A1(n7010), .A2(n7911), .ZN(n7994) );
  INV_X1 U8786 ( .A(n7994), .ZN(n7026) );
  NAND3_X1 U8787 ( .A1(n7026), .A2(n8050), .A3(n7030), .ZN(n7011) );
  NAND2_X1 U8788 ( .A1(n5683), .A2(n9427), .ZN(n7027) );
  OAI211_X1 U8789 ( .C1(n7103), .C2(n7012), .A(n7011), .B(n7027), .ZN(n7013)
         );
  INV_X1 U8790 ( .A(n9813), .ZN(n9518) );
  NAND2_X1 U8791 ( .A1(n7013), .A2(n9518), .ZN(n7014) );
  OAI211_X1 U8792 ( .C1(n7016), .C2(n9518), .A(n7015), .B(n7014), .ZN(P1_U3293) );
  OAI21_X1 U8793 ( .B1(n7018), .B2(n7999), .A(n7017), .ZN(n9810) );
  INV_X1 U8794 ( .A(n9810), .ZN(n7023) );
  XNOR2_X1 U8795 ( .A(n7019), .B(n7999), .ZN(n7022) );
  NAND2_X1 U8796 ( .A1(n9187), .A2(n9427), .ZN(n7020) );
  OAI21_X1 U8797 ( .B1(n7021), .B2(n9456), .A(n7020), .ZN(n7248) );
  AOI21_X1 U8798 ( .B1(n7022), .B2(n9504), .A(n7248), .ZN(n9812) );
  OAI211_X1 U8799 ( .C1(n7200), .C2(n7373), .A(n9551), .B(n7185), .ZN(n9807)
         );
  OAI211_X1 U8800 ( .C1(n7023), .C2(n9583), .A(n9812), .B(n9807), .ZN(n7375)
         );
  OAI22_X1 U8801 ( .A1(n9590), .A2(n7373), .B1(n9854), .B2(n6606), .ZN(n7024)
         );
  AOI21_X1 U8802 ( .B1(n7375), .B2(n9854), .A(n7024), .ZN(n7025) );
  INV_X1 U8803 ( .A(n7025), .ZN(P1_U3528) );
  INV_X1 U8804 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7032) );
  OAI21_X1 U8805 ( .B1(n9835), .B2(n9504), .A(n7026), .ZN(n7028) );
  OAI211_X1 U8806 ( .C1(n7030), .C2(n7029), .A(n7028), .B(n7027), .ZN(n9591)
         );
  NAND2_X1 U8807 ( .A1(n9591), .A2(n9627), .ZN(n7031) );
  OAI21_X1 U8808 ( .B1(n9627), .B2(n7032), .A(n7031), .ZN(P1_U3453) );
  INV_X1 U8809 ( .A(n7033), .ZN(n7035) );
  INV_X1 U8810 ( .A(n7138), .ZN(n7034) );
  AOI21_X1 U8811 ( .B1(n4402), .B2(n7035), .A(n7034), .ZN(n9927) );
  INV_X1 U8812 ( .A(n9927), .ZN(n9924) );
  OAI22_X1 U8813 ( .A1(n8859), .A2(n7036), .B1(n7214), .B2(n8882), .ZN(n7037)
         );
  AOI21_X1 U8814 ( .B1(n8887), .B2(n8522), .A(n7037), .ZN(n7038) );
  OAI21_X1 U8815 ( .B1(n9918), .B2(n8830), .A(n7038), .ZN(n7039) );
  AOI21_X1 U8816 ( .B1(n8861), .B2(n9922), .A(n7039), .ZN(n7043) );
  XNOR2_X1 U8817 ( .A(n7040), .B(n4402), .ZN(n7041) );
  NOR2_X1 U8818 ( .A1(n7041), .A2(n8917), .ZN(n9925) );
  NAND2_X1 U8819 ( .A1(n9925), .A2(n8859), .ZN(n7042) );
  OAI211_X1 U8820 ( .C1(n9924), .C2(n8876), .A(n7043), .B(n7042), .ZN(P2_U3224) );
  INV_X1 U8821 ( .A(n7044), .ZN(n7046) );
  OAI222_X1 U8822 ( .A1(n8643), .A2(P2_U3151), .B1(n9044), .B2(n7046), .C1(
        n7045), .C2(n9042), .ZN(P2_U3278) );
  INV_X1 U8823 ( .A(n9778), .ZN(n9311) );
  OAI222_X1 U8824 ( .A1(n8084), .A2(n7047), .B1(n9640), .B2(n7046), .C1(
        P1_U3086), .C2(n9311), .ZN(P1_U3338) );
  OR2_X1 U8825 ( .A1(n7048), .A2(n5385), .ZN(n7049) );
  INV_X1 U8826 ( .A(n7050), .ZN(n7059) );
  NAND2_X1 U8827 ( .A1(n7051), .A2(n9518), .ZN(n7058) );
  NOR2_X1 U8828 ( .A1(n9516), .A2(n7329), .ZN(n7055) );
  INV_X1 U8829 ( .A(n7099), .ZN(n7052) );
  OAI22_X1 U8830 ( .A1(n9518), .A2(n7053), .B1(n7052), .B2(n7103), .ZN(n7054)
         );
  AOI211_X1 U8831 ( .C1(n7056), .C2(n9512), .A(n7055), .B(n7054), .ZN(n7057)
         );
  OAI211_X1 U8832 ( .C1(n9520), .C2(n7059), .A(n7058), .B(n7057), .ZN(P1_U3289) );
  INV_X1 U8833 ( .A(n7060), .ZN(n7069) );
  NOR2_X1 U8834 ( .A1(n9516), .A2(n4369), .ZN(n7064) );
  INV_X1 U8835 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7061) );
  OAI22_X1 U8836 ( .A1(n9518), .A2(n7062), .B1(n7061), .B2(n7103), .ZN(n7063)
         );
  AOI211_X1 U8837 ( .C1(n7065), .C2(n9512), .A(n7064), .B(n7063), .ZN(n7068)
         );
  NAND2_X1 U8838 ( .A1(n9809), .A2(n7066), .ZN(n7067) );
  OAI211_X1 U8839 ( .C1(n9813), .C2(n7069), .A(n7068), .B(n7067), .ZN(P1_U3292) );
  INV_X1 U8840 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U8841 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7070) );
  AOI21_X1 U8842 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7070), .ZN(n9968) );
  INV_X1 U8843 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9771) );
  INV_X1 U8844 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8590) );
  AOI22_X1 U8845 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n9771), .B2(n8590), .ZN(n9971) );
  NOR2_X1 U8846 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7071) );
  AOI21_X1 U8847 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7071), .ZN(n9974) );
  INV_X1 U8848 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10069) );
  INV_X1 U8849 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7072) );
  AOI22_X1 U8850 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .B1(n10069), .B2(n7072), .ZN(n9977) );
  NOR2_X1 U8851 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7073) );
  AOI21_X1 U8852 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7073), .ZN(n9980) );
  NOR2_X1 U8853 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7074) );
  AOI21_X1 U8854 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7074), .ZN(n9983) );
  NOR2_X1 U8855 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7075) );
  AOI21_X1 U8856 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7075), .ZN(n9986) );
  NOR2_X1 U8857 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7076) );
  AOI21_X1 U8858 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7076), .ZN(n9989) );
  NOR2_X1 U8859 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7077) );
  AOI21_X1 U8860 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7077), .ZN(n10158) );
  NOR2_X1 U8861 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7078) );
  AOI21_X1 U8862 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7078), .ZN(n10164) );
  NOR2_X1 U8863 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7079) );
  AOI21_X1 U8864 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7079), .ZN(n10161) );
  NOR2_X1 U8865 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7080) );
  AOI21_X1 U8866 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7080), .ZN(n10152) );
  NOR2_X1 U8867 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7081) );
  AOI21_X1 U8868 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7081), .ZN(n10155) );
  AND2_X1 U8869 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7082) );
  NOR2_X1 U8870 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7082), .ZN(n9958) );
  INV_X1 U8871 ( .A(n9958), .ZN(n9959) );
  NAND3_X1 U8872 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U8873 ( .A1(n9961), .A2(n9960), .ZN(n9957) );
  NAND2_X1 U8874 ( .A1(n9959), .A2(n9957), .ZN(n10167) );
  NAND2_X1 U8875 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7083) );
  OAI21_X1 U8876 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n7083), .ZN(n10166) );
  NOR2_X1 U8877 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10165), .ZN(n10170) );
  NAND2_X1 U8879 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7084) );
  OAI21_X1 U8880 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7084), .ZN(n10169) );
  NOR2_X1 U8881 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  AOI21_X1 U8882 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10168), .ZN(n10173) );
  NOR2_X1 U8883 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7085) );
  AOI21_X1 U8884 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7085), .ZN(n10172) );
  NAND2_X1 U8885 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  OAI21_X1 U8886 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10171), .ZN(n10154) );
  NAND2_X1 U8887 ( .A1(n10155), .A2(n10154), .ZN(n10153) );
  OAI21_X1 U8888 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10153), .ZN(n10151) );
  NAND2_X1 U8889 ( .A1(n10152), .A2(n10151), .ZN(n10150) );
  OAI21_X1 U8890 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10150), .ZN(n10160) );
  NAND2_X1 U8891 ( .A1(n10161), .A2(n10160), .ZN(n10159) );
  OAI21_X1 U8892 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10159), .ZN(n10163) );
  NAND2_X1 U8893 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  OAI21_X1 U8894 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10162), .ZN(n10157) );
  NAND2_X1 U8895 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  OAI21_X1 U8896 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10156), .ZN(n9988) );
  NAND2_X1 U8897 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  OAI21_X1 U8898 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9987), .ZN(n9985) );
  NAND2_X1 U8899 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  OAI21_X1 U8900 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9984), .ZN(n9982) );
  NAND2_X1 U8901 ( .A1(n9983), .A2(n9982), .ZN(n9981) );
  OAI21_X1 U8902 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9981), .ZN(n9979) );
  NAND2_X1 U8903 ( .A1(n9980), .A2(n9979), .ZN(n9978) );
  OAI21_X1 U8904 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9978), .ZN(n9976) );
  NAND2_X1 U8905 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  OAI21_X1 U8906 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9975), .ZN(n9973) );
  NAND2_X1 U8907 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  OAI21_X1 U8908 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9972), .ZN(n9970) );
  NAND2_X1 U8909 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  OAI21_X1 U8910 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9969), .ZN(n9967) );
  NAND2_X1 U8911 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  OAI21_X1 U8912 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9966), .ZN(n9963) );
  NAND2_X1 U8913 ( .A1(n9964), .A2(n9963), .ZN(n7086) );
  NOR2_X1 U8914 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  AOI21_X1 U8915 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7086), .A(n9962), .ZN(
        n7089) );
  XNOR2_X1 U8916 ( .A(n7087), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7088) );
  XNOR2_X1 U8917 ( .A(n7089), .B(n7088), .ZN(ADD_1068_U4) );
  INV_X1 U8918 ( .A(n7090), .ZN(n7091) );
  NAND2_X1 U8919 ( .A1(n9066), .A2(n7091), .ZN(n7092) );
  NAND2_X1 U8920 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9218) );
  OAI211_X1 U8921 ( .C1(n9157), .C2(n7329), .A(n7092), .B(n9218), .ZN(n7098)
         );
  INV_X1 U8922 ( .A(n7094), .ZN(n7095) );
  AOI211_X1 U8923 ( .C1(n7096), .C2(n7093), .A(n9671), .B(n7095), .ZN(n7097)
         );
  AOI211_X1 U8924 ( .C1(n7099), .C2(n9161), .A(n7098), .B(n7097), .ZN(n7100)
         );
  INV_X1 U8925 ( .A(n7100), .ZN(P1_U3230) );
  INV_X1 U8926 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7102) );
  INV_X1 U8927 ( .A(n7101), .ZN(n7125) );
  INV_X1 U8928 ( .A(n8663), .ZN(n8675) );
  OAI222_X1 U8929 ( .A1(n9042), .A2(n7102), .B1(n9044), .B2(n7125), .C1(
        P2_U3151), .C2(n8675), .ZN(P2_U3277) );
  INV_X2 U8930 ( .A(n7103), .ZN(n9800) );
  AOI21_X1 U8931 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9800), .A(n7104), .ZN(
        n7111) );
  NOR2_X1 U8932 ( .A1(n9516), .A2(n7910), .ZN(n7108) );
  INV_X1 U8933 ( .A(n7105), .ZN(n7106) );
  OAI22_X1 U8934 ( .A1(n9806), .A2(n7106), .B1(n9518), .B2(n6619), .ZN(n7107)
         );
  AOI211_X1 U8935 ( .C1(n9809), .C2(n7109), .A(n7108), .B(n7107), .ZN(n7110)
         );
  OAI21_X1 U8936 ( .B1(n7111), .B2(n9494), .A(n7110), .ZN(P1_U3291) );
  INV_X1 U8937 ( .A(n7112), .ZN(n7113) );
  XNOR2_X1 U8938 ( .A(n9916), .B(n8131), .ZN(n7352) );
  XOR2_X1 U8939 ( .A(n7209), .B(n7352), .Z(n7210) );
  XNOR2_X1 U8940 ( .A(n7210), .B(n9918), .ZN(n7123) );
  AOI21_X1 U8941 ( .B1(n8290), .B2(n8525), .A(n7115), .ZN(n7121) );
  NAND2_X1 U8942 ( .A1(n8259), .A2(n9916), .ZN(n7120) );
  INV_X1 U8943 ( .A(n7116), .ZN(n7117) );
  NAND2_X1 U8944 ( .A1(n8267), .A2(n7117), .ZN(n7119) );
  NAND2_X1 U8945 ( .A1(n8277), .A2(n8523), .ZN(n7118) );
  NAND4_X1 U8946 ( .A1(n7121), .A2(n7120), .A3(n7119), .A4(n7118), .ZN(n7122)
         );
  AOI21_X1 U8947 ( .B1(n7123), .B2(n8272), .A(n7122), .ZN(n7124) );
  INV_X1 U8948 ( .A(n7124), .ZN(P2_U3161) );
  INV_X1 U8949 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7126) );
  INV_X1 U8950 ( .A(n9313), .ZN(n9794) );
  OAI222_X1 U8951 ( .A1(n8084), .A2(n7126), .B1(n9794), .B2(P1_U3086), .C1(
        n9640), .C2(n7125), .ZN(P1_U3337) );
  NAND2_X1 U8952 ( .A1(n7127), .A2(n7128), .ZN(n7129) );
  XOR2_X1 U8953 ( .A(n7130), .B(n7129), .Z(n7136) );
  NAND2_X1 U8954 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9231) );
  OAI21_X1 U8955 ( .B1(n9157), .B2(n9817), .A(n9231), .ZN(n7134) );
  OAI22_X1 U8956 ( .A1(n7132), .A2(n9662), .B1(n9661), .B2(n7131), .ZN(n7133)
         );
  AOI211_X1 U8957 ( .C1(n7202), .C2(n9161), .A(n7134), .B(n7133), .ZN(n7135)
         );
  OAI21_X1 U8958 ( .B1(n7136), .B2(n9671), .A(n7135), .ZN(P1_U3227) );
  NAND2_X1 U8959 ( .A1(n7138), .A2(n7137), .ZN(n7139) );
  XNOR2_X1 U8960 ( .A(n9934), .B(n9920), .ZN(n8484) );
  XNOR2_X1 U8961 ( .A(n7139), .B(n8484), .ZN(n7141) );
  INV_X1 U8962 ( .A(n7141), .ZN(n9931) );
  XNOR2_X1 U8963 ( .A(n7140), .B(n8484), .ZN(n7144) );
  AOI22_X1 U8964 ( .A1(n8521), .A2(n9872), .B1(n9874), .B2(n8523), .ZN(n7143)
         );
  NAND2_X1 U8965 ( .A1(n7141), .A2(n9928), .ZN(n7142) );
  OAI211_X1 U8966 ( .C1(n7144), .C2(n8917), .A(n7143), .B(n7142), .ZN(n9932)
         );
  NAND2_X1 U8967 ( .A1(n9932), .A2(n8859), .ZN(n7148) );
  OAI22_X1 U8968 ( .A1(n8859), .A2(n7145), .B1(n7363), .B2(n8882), .ZN(n7146)
         );
  AOI21_X1 U8969 ( .B1(n9934), .B2(n8861), .A(n7146), .ZN(n7147) );
  OAI211_X1 U8970 ( .C1(n9931), .C2(n8700), .A(n7148), .B(n7147), .ZN(P2_U3223) );
  NAND2_X1 U8971 ( .A1(n7149), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7150) );
  AOI21_X1 U8972 ( .B1(n7160), .B2(n7152), .A(n7388), .ZN(n7173) );
  NAND2_X1 U8973 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7155), .ZN(n7396) );
  OAI21_X1 U8974 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7155), .A(n7396), .ZN(
        n7171) );
  INV_X1 U8975 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8976 ( .A1(n8587), .A2(n7387), .ZN(n7157) );
  AND2_X1 U8977 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7498) );
  INV_X1 U8978 ( .A(n7498), .ZN(n7156) );
  OAI211_X1 U8979 ( .C1(n7158), .C2(n8653), .A(n7157), .B(n7156), .ZN(n7170)
         );
  MUX2_X1 U8980 ( .A(n7160), .B(n7159), .S(n8665), .Z(n7161) );
  NAND2_X1 U8981 ( .A1(n7161), .A2(n7387), .ZN(n7406) );
  INV_X1 U8982 ( .A(n7161), .ZN(n7162) );
  NAND2_X1 U8983 ( .A1(n7162), .A2(n7395), .ZN(n7163) );
  NAND2_X1 U8984 ( .A1(n7406), .A2(n7163), .ZN(n7164) );
  AOI21_X1 U8985 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7414) );
  INV_X1 U8986 ( .A(n7414), .ZN(n7168) );
  NAND3_X1 U8987 ( .A1(n7166), .A2(n7165), .A3(n7164), .ZN(n7167) );
  AOI21_X1 U8988 ( .B1(n7168), .B2(n7167), .A(n8617), .ZN(n7169) );
  AOI211_X1 U8989 ( .C1(n8624), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7172)
         );
  OAI21_X1 U8990 ( .B1(n7173), .B2(n8685), .A(n7172), .ZN(P2_U3193) );
  OR2_X1 U8991 ( .A1(n7174), .A2(n7178), .ZN(n7175) );
  NAND2_X1 U8992 ( .A1(n7176), .A2(n7175), .ZN(n9822) );
  INV_X1 U8993 ( .A(n7622), .ZN(n7301) );
  NAND2_X1 U8994 ( .A1(n9822), .A2(n7301), .ZN(n7184) );
  INV_X1 U8995 ( .A(n7779), .ZN(n7784) );
  OR2_X1 U8996 ( .A1(n7019), .A2(n7784), .ZN(n7179) );
  NAND2_X1 U8997 ( .A1(n7179), .A2(n7919), .ZN(n7177) );
  INV_X1 U8998 ( .A(n7178), .ZN(n7785) );
  NAND2_X1 U8999 ( .A1(n7177), .A2(n7785), .ZN(n7230) );
  NAND3_X1 U9000 ( .A1(n7179), .A2(n7178), .A3(n7919), .ZN(n7180) );
  NAND2_X1 U9001 ( .A1(n7230), .A2(n7180), .ZN(n7181) );
  NAND2_X1 U9002 ( .A1(n7181), .A2(n9504), .ZN(n7183) );
  AOI22_X1 U9003 ( .A1(n9188), .A2(n9425), .B1(n9427), .B2(n9186), .ZN(n7182)
         );
  NAND3_X1 U9004 ( .A1(n7184), .A2(n7183), .A3(n7182), .ZN(n9827) );
  INV_X1 U9005 ( .A(n9827), .ZN(n7193) );
  INV_X1 U9006 ( .A(n7629), .ZN(n7307) );
  AOI21_X1 U9007 ( .B1(n7185), .B2(n7188), .A(n9509), .ZN(n7186) );
  NAND2_X1 U9008 ( .A1(n7186), .A2(n7225), .ZN(n9823) );
  AOI22_X1 U9009 ( .A1(n9494), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7187), .B2(
        n9800), .ZN(n7190) );
  NAND2_X1 U9010 ( .A1(n9803), .A2(n7188), .ZN(n7189) );
  OAI211_X1 U9011 ( .C1(n9823), .C2(n9806), .A(n7190), .B(n7189), .ZN(n7191)
         );
  AOI21_X1 U9012 ( .B1(n9822), .B2(n7307), .A(n7191), .ZN(n7192) );
  OAI21_X1 U9013 ( .B1(n7193), .B2(n9494), .A(n7192), .ZN(P1_U3286) );
  XNOR2_X1 U9014 ( .A(n7776), .B(n7996), .ZN(n7194) );
  NAND2_X1 U9015 ( .A1(n7194), .A2(n9504), .ZN(n7196) );
  AOI22_X1 U9016 ( .A1(n9188), .A2(n9427), .B1(n9425), .B2(n9190), .ZN(n7195)
         );
  NAND2_X1 U9017 ( .A1(n7196), .A2(n7195), .ZN(n9818) );
  INV_X1 U9018 ( .A(n9818), .ZN(n7208) );
  OAI21_X1 U9019 ( .B1(n7198), .B2(n7996), .A(n7197), .ZN(n9820) );
  OAI21_X1 U9020 ( .B1(n7199), .B2(n9817), .A(n9551), .ZN(n7201) );
  OR2_X1 U9021 ( .A1(n7201), .A2(n7200), .ZN(n9816) );
  AOI22_X1 U9022 ( .A1(n9494), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7202), .B2(
        n9800), .ZN(n7205) );
  NAND2_X1 U9023 ( .A1(n9803), .A2(n7203), .ZN(n7204) );
  OAI211_X1 U9024 ( .C1(n9816), .C2(n9806), .A(n7205), .B(n7204), .ZN(n7206)
         );
  AOI21_X1 U9025 ( .B1(n9820), .B2(n9809), .A(n7206), .ZN(n7207) );
  OAI21_X1 U9026 ( .B1(n7208), .B2(n9494), .A(n7207), .ZN(P1_U3288) );
  AOI22_X1 U9027 ( .A1(n7210), .A2(n9918), .B1(n7209), .B2(n7352), .ZN(n7212)
         );
  XOR2_X1 U9028 ( .A(n8131), .B(n9922), .Z(n7355) );
  XNOR2_X1 U9029 ( .A(n7355), .B(n8523), .ZN(n7211) );
  XNOR2_X1 U9030 ( .A(n7212), .B(n7211), .ZN(n7221) );
  AOI21_X1 U9031 ( .B1(n8290), .B2(n8524), .A(n7213), .ZN(n7219) );
  NAND2_X1 U9032 ( .A1(n8259), .A2(n9922), .ZN(n7218) );
  INV_X1 U9033 ( .A(n7214), .ZN(n7215) );
  NAND2_X1 U9034 ( .A1(n8267), .A2(n7215), .ZN(n7217) );
  NAND2_X1 U9035 ( .A1(n8277), .A2(n8522), .ZN(n7216) );
  NAND4_X1 U9036 ( .A1(n7219), .A2(n7218), .A3(n7217), .A4(n7216), .ZN(n7220)
         );
  AOI21_X1 U9037 ( .B1(n7221), .B2(n8272), .A(n7220), .ZN(n7222) );
  INV_X1 U9038 ( .A(n7222), .ZN(P2_U3171) );
  OAI21_X1 U9039 ( .B1(n7224), .B2(n7227), .A(n7223), .ZN(n7255) );
  AOI211_X1 U9040 ( .C1(n7226), .C2(n7225), .A(n9509), .B(n7283), .ZN(n7256)
         );
  INV_X1 U9041 ( .A(n7227), .ZN(n7228) );
  NAND3_X1 U9042 ( .A1(n7230), .A2(n7228), .A3(n7229), .ZN(n7275) );
  NAND2_X1 U9043 ( .A1(n7275), .A2(n9504), .ZN(n7233) );
  AOI21_X1 U9044 ( .B1(n7230), .B2(n7229), .A(n7228), .ZN(n7232) );
  AOI22_X1 U9045 ( .A1(n9185), .A2(n9427), .B1(n9425), .B2(n9187), .ZN(n7231)
         );
  OAI21_X1 U9046 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7260) );
  AOI211_X1 U9047 ( .C1(n9835), .C2(n7255), .A(n7256), .B(n7260), .ZN(n7336)
         );
  OAI22_X1 U9048 ( .A1(n9590), .A2(n7476), .B1(n9854), .B2(n6609), .ZN(n7234)
         );
  INV_X1 U9049 ( .A(n7234), .ZN(n7235) );
  OAI21_X1 U9050 ( .B1(n7336), .B2(n5802), .A(n7235), .ZN(P1_U3530) );
  NAND2_X1 U9051 ( .A1(n7236), .A2(n8362), .ZN(n7237) );
  XOR2_X1 U9052 ( .A(n8483), .B(n7237), .Z(n9936) );
  OAI211_X1 U9053 ( .C1(n4348), .C2(n6034), .A(n9902), .B(n7238), .ZN(n7240)
         );
  AOI22_X1 U9054 ( .A1(n9874), .A2(n8522), .B1(n8520), .B2(n9872), .ZN(n7239)
         );
  NAND2_X1 U9055 ( .A1(n7240), .A2(n7239), .ZN(n9937) );
  NAND2_X1 U9056 ( .A1(n9937), .A2(n8859), .ZN(n7243) );
  OAI22_X1 U9057 ( .A1(n8859), .A2(n7160), .B1(n7500), .B2(n8882), .ZN(n7241)
         );
  AOI21_X1 U9058 ( .B1(n9939), .B2(n8861), .A(n7241), .ZN(n7242) );
  OAI211_X1 U9059 ( .C1(n9936), .C2(n8864), .A(n7243), .B(n7242), .ZN(P2_U3222) );
  XNOR2_X1 U9060 ( .A(n7246), .B(n7245), .ZN(n7247) );
  XNOR2_X1 U9061 ( .A(n7244), .B(n7247), .ZN(n7253) );
  INV_X1 U9062 ( .A(n9801), .ZN(n7251) );
  NAND2_X1 U9063 ( .A1(n9675), .A2(n9802), .ZN(n7250) );
  AOI22_X1 U9064 ( .A1(n9066), .A2(n7248), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7249) );
  OAI211_X1 U9065 ( .C1(n9678), .C2(n7251), .A(n7250), .B(n7249), .ZN(n7252)
         );
  AOI21_X1 U9066 ( .B1(n7253), .B2(n9151), .A(n7252), .ZN(n7254) );
  INV_X1 U9067 ( .A(n7254), .ZN(P1_U3239) );
  INV_X1 U9068 ( .A(n7255), .ZN(n7262) );
  NAND2_X1 U9069 ( .A1(n7256), .A2(n9512), .ZN(n7258) );
  AOI22_X1 U9070 ( .A1(n9494), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7481), .B2(
        n9800), .ZN(n7257) );
  OAI211_X1 U9071 ( .C1(n7476), .C2(n9516), .A(n7258), .B(n7257), .ZN(n7259)
         );
  AOI21_X1 U9072 ( .B1(n7260), .B2(n9518), .A(n7259), .ZN(n7261) );
  OAI21_X1 U9073 ( .B1(n9520), .B2(n7262), .A(n7261), .ZN(P1_U3285) );
  INV_X1 U9074 ( .A(n7263), .ZN(n7265) );
  OAI222_X1 U9075 ( .A1(n8084), .A2(n10018), .B1(n9640), .B2(n7265), .C1(
        P1_U3086), .C2(n5385), .ZN(P1_U3336) );
  OAI222_X1 U9076 ( .A1(P2_U3151), .A2(n4274), .B1(n9044), .B2(n7265), .C1(
        n7264), .C2(n9042), .ZN(P2_U3276) );
  INV_X1 U9077 ( .A(n7266), .ZN(n7274) );
  NAND2_X1 U9078 ( .A1(n7267), .A2(n9512), .ZN(n7270) );
  AOI22_X1 U9079 ( .A1(n9813), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9800), .B2(
        n7268), .ZN(n7269) );
  OAI211_X1 U9080 ( .C1(n5686), .C2(n9516), .A(n7270), .B(n7269), .ZN(n7271)
         );
  AOI21_X1 U9081 ( .B1(n9809), .B2(n7272), .A(n7271), .ZN(n7273) );
  OAI21_X1 U9082 ( .B1(n9813), .B2(n7274), .A(n7273), .ZN(P1_U3290) );
  NAND2_X1 U9083 ( .A1(n7275), .A2(n7786), .ZN(n7276) );
  XNOR2_X1 U9084 ( .A(n7276), .B(n7281), .ZN(n7277) );
  AOI22_X1 U9085 ( .A1(n7277), .A2(n9504), .B1(n9425), .B2(n9186), .ZN(n9830)
         );
  INV_X1 U9086 ( .A(n9830), .ZN(n7278) );
  AOI21_X1 U9087 ( .B1(n7279), .B2(n9800), .A(n7278), .ZN(n7290) );
  OAI21_X1 U9088 ( .B1(n7282), .B2(n7281), .A(n7280), .ZN(n9834) );
  OAI21_X1 U9089 ( .B1(n7283), .B2(n9832), .A(n9551), .ZN(n7284) );
  OR2_X1 U9090 ( .A1(n7284), .A2(n7315), .ZN(n7286) );
  NAND2_X1 U9091 ( .A1(n9184), .A2(n9427), .ZN(n7285) );
  AND2_X1 U9092 ( .A1(n7286), .A2(n7285), .ZN(n9829) );
  AOI22_X1 U9093 ( .A1(n9803), .A2(n7527), .B1(n9813), .B2(
        P1_REG2_REG_9__SCAN_IN), .ZN(n7287) );
  OAI21_X1 U9094 ( .B1(n9829), .B2(n9806), .A(n7287), .ZN(n7288) );
  AOI21_X1 U9095 ( .B1(n9834), .B2(n9809), .A(n7288), .ZN(n7289) );
  OAI21_X1 U9096 ( .B1(n7290), .B2(n9494), .A(n7289), .ZN(P1_U3284) );
  OR2_X1 U9097 ( .A1(n7291), .A2(n8005), .ZN(n7292) );
  NAND2_X1 U9098 ( .A1(n7293), .A2(n7292), .ZN(n9843) );
  NAND2_X1 U9099 ( .A1(n7313), .A2(n7799), .ZN(n7294) );
  NAND2_X1 U9100 ( .A1(n7294), .A2(n8005), .ZN(n7296) );
  NAND3_X1 U9101 ( .A1(n7296), .A2(n7295), .A3(n9504), .ZN(n7299) );
  OAI22_X1 U9102 ( .A1(n9663), .A2(n9456), .B1(n9660), .B2(n9458), .ZN(n7297)
         );
  INV_X1 U9103 ( .A(n7297), .ZN(n7298) );
  NAND2_X1 U9104 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  AOI21_X1 U9105 ( .B1(n9843), .B2(n7301), .A(n7300), .ZN(n9845) );
  AOI21_X1 U9106 ( .B1(n7316), .B2(n9838), .A(n9509), .ZN(n7302) );
  NAND2_X1 U9107 ( .A1(n7302), .A2(n4349), .ZN(n9840) );
  AOI22_X1 U9108 ( .A1(n9494), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7303), .B2(
        n9800), .ZN(n7305) );
  NAND2_X1 U9109 ( .A1(n9838), .A2(n9803), .ZN(n7304) );
  OAI211_X1 U9110 ( .C1(n9840), .C2(n9806), .A(n7305), .B(n7304), .ZN(n7306)
         );
  AOI21_X1 U9111 ( .B1(n9843), .B2(n7307), .A(n7306), .ZN(n7308) );
  OAI21_X1 U9112 ( .B1(n9845), .B2(n9494), .A(n7308), .ZN(P1_U3282) );
  INV_X1 U9113 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7321) );
  OAI21_X1 U9114 ( .B1(n7310), .B2(n7312), .A(n7309), .ZN(n7311) );
  INV_X1 U9115 ( .A(n7311), .ZN(n7384) );
  OAI21_X1 U9116 ( .B1(n4352), .B2(n4612), .A(n7313), .ZN(n7314) );
  AOI222_X1 U9117 ( .A1(n9504), .A2(n7314), .B1(n9183), .B2(n9427), .C1(n9185), 
        .C2(n9425), .ZN(n7379) );
  INV_X1 U9118 ( .A(n7315), .ZN(n7317) );
  AOI21_X1 U9119 ( .B1(n7318), .B2(n7317), .A(n4527), .ZN(n7382) );
  AOI22_X1 U9120 ( .A1(n7382), .A2(n9551), .B1(n9837), .B2(n7318), .ZN(n7319)
         );
  OAI211_X1 U9121 ( .C1(n7384), .C2(n9583), .A(n7379), .B(n7319), .ZN(n7322)
         );
  NAND2_X1 U9122 ( .A1(n7322), .A2(n9854), .ZN(n7320) );
  OAI21_X1 U9123 ( .B1(n9854), .B2(n7321), .A(n7320), .ZN(P1_U3532) );
  INV_X1 U9124 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U9125 ( .A1(n7322), .A2(n9627), .ZN(n7323) );
  OAI21_X1 U9126 ( .B1(n9627), .B2(n7324), .A(n7323), .ZN(P1_U3483) );
  INV_X1 U9127 ( .A(n7325), .ZN(n7377) );
  NAND2_X1 U9128 ( .A1(n9638), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7326) );
  OAI211_X1 U9129 ( .C1(n7377), .C2(n9640), .A(n7327), .B(n7326), .ZN(P1_U3335) );
  INV_X1 U9130 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7328) );
  OAI22_X1 U9131 ( .A1(n9631), .A2(n7329), .B1(n9627), .B2(n7328), .ZN(n7330)
         );
  INV_X1 U9132 ( .A(n7330), .ZN(n7331) );
  OAI21_X1 U9133 ( .B1(n7332), .B2(n9846), .A(n7331), .ZN(P1_U3465) );
  INV_X1 U9134 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7333) );
  OAI22_X1 U9135 ( .A1(n9631), .A2(n7476), .B1(n9627), .B2(n7333), .ZN(n7334)
         );
  INV_X1 U9136 ( .A(n7334), .ZN(n7335) );
  OAI21_X1 U9137 ( .B1(n7336), .B2(n9846), .A(n7335), .ZN(P1_U3477) );
  INV_X1 U9138 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7337) );
  OAI22_X1 U9139 ( .A1(n9631), .A2(n4369), .B1(n9627), .B2(n7337), .ZN(n7338)
         );
  INV_X1 U9140 ( .A(n7338), .ZN(n7339) );
  OAI21_X1 U9141 ( .B1(n7340), .B2(n9846), .A(n7339), .ZN(P1_U3456) );
  OAI22_X1 U9142 ( .A1(n9631), .A2(n5686), .B1(n9627), .B2(n4978), .ZN(n7341)
         );
  INV_X1 U9143 ( .A(n7341), .ZN(n7342) );
  OAI21_X1 U9144 ( .B1(n7343), .B2(n9846), .A(n7342), .ZN(P1_U3462) );
  INV_X1 U9145 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7344) );
  OAI22_X1 U9146 ( .A1(n9631), .A2(n7910), .B1(n9627), .B2(n7344), .ZN(n7345)
         );
  INV_X1 U9147 ( .A(n7345), .ZN(n7346) );
  OAI21_X1 U9148 ( .B1(n7347), .B2(n9846), .A(n7346), .ZN(P1_U3459) );
  INV_X1 U9149 ( .A(n7348), .ZN(n7358) );
  NOR2_X1 U9150 ( .A1(n7355), .A2(n8523), .ZN(n7350) );
  OAI21_X1 U9151 ( .B1(n7352), .B2(n9918), .A(n8360), .ZN(n7354) );
  NOR3_X1 U9152 ( .A1(n7352), .A2(n8360), .A3(n9918), .ZN(n7353) );
  NOR2_X1 U9153 ( .A1(n7359), .A2(n9920), .ZN(n7486) );
  INV_X1 U9154 ( .A(n7486), .ZN(n7360) );
  NAND2_X1 U9155 ( .A1(n7359), .A2(n9920), .ZN(n7484) );
  NAND2_X1 U9156 ( .A1(n7360), .A2(n7484), .ZN(n7361) );
  XOR2_X1 U9157 ( .A(n8131), .B(n9934), .Z(n7485) );
  XNOR2_X1 U9158 ( .A(n7361), .B(n7485), .ZN(n7370) );
  AOI21_X1 U9159 ( .B1(n8290), .B2(n8523), .A(n7362), .ZN(n7368) );
  NAND2_X1 U9160 ( .A1(n9934), .A2(n8259), .ZN(n7367) );
  INV_X1 U9161 ( .A(n7363), .ZN(n7364) );
  NAND2_X1 U9162 ( .A1(n8267), .A2(n7364), .ZN(n7366) );
  NAND2_X1 U9163 ( .A1(n8277), .A2(n8521), .ZN(n7365) );
  NAND4_X1 U9164 ( .A1(n7368), .A2(n7367), .A3(n7366), .A4(n7365), .ZN(n7369)
         );
  AOI21_X1 U9165 ( .B1(n7370), .B2(n8272), .A(n7369), .ZN(n7371) );
  INV_X1 U9166 ( .A(n7371), .ZN(P2_U3157) );
  INV_X1 U9167 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7372) );
  OAI22_X1 U9168 ( .A1(n9631), .A2(n7373), .B1(n9627), .B2(n7372), .ZN(n7374)
         );
  AOI21_X1 U9169 ( .B1(n7375), .B2(n9627), .A(n7374), .ZN(n7376) );
  INV_X1 U9170 ( .A(n7376), .ZN(P1_U3471) );
  OAI222_X1 U9171 ( .A1(P2_U3151), .A2(n8462), .B1(n9042), .B2(n6124), .C1(
        n7377), .C2(n9048), .ZN(P2_U3275) );
  AOI22_X1 U9172 ( .A1(n9813), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7583), .B2(
        n9800), .ZN(n7378) );
  OAI21_X1 U9173 ( .B1(n7586), .B2(n9516), .A(n7378), .ZN(n7381) );
  NOR2_X1 U9174 ( .A1(n7379), .A2(n9494), .ZN(n7380) );
  AOI211_X1 U9175 ( .C1(n7382), .C2(n9432), .A(n7381), .B(n7380), .ZN(n7383)
         );
  OAI21_X1 U9176 ( .B1(n9520), .B2(n7384), .A(n7383), .ZN(P1_U3283) );
  INV_X1 U9177 ( .A(n7390), .ZN(n7393) );
  INV_X1 U9178 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7541) );
  MUX2_X1 U9179 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7541), .S(n7546), .Z(n7392)
         );
  INV_X1 U9180 ( .A(n7543), .ZN(n7391) );
  AOI21_X1 U9181 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7419) );
  NAND2_X1 U9182 ( .A1(n7395), .A2(n7394), .ZN(n7397) );
  MUX2_X1 U9183 ( .A(n7407), .B(P2_REG1_REG_12__SCAN_IN), .S(n7546), .Z(n7398)
         );
  OAI21_X1 U9184 ( .B1(n7399), .B2(n7398), .A(n7545), .ZN(n7405) );
  INV_X1 U9185 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9186 ( .A1(n8587), .A2(n7546), .ZN(n7402) );
  NOR2_X1 U9187 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7400), .ZN(n7490) );
  INV_X1 U9188 ( .A(n7490), .ZN(n7401) );
  OAI211_X1 U9189 ( .C1(n7403), .C2(n8653), .A(n7402), .B(n7401), .ZN(n7404)
         );
  AOI21_X1 U9190 ( .B1(n7405), .B2(n8624), .A(n7404), .ZN(n7418) );
  INV_X1 U9191 ( .A(n7406), .ZN(n7413) );
  MUX2_X1 U9192 ( .A(n7541), .B(n7407), .S(n8665), .Z(n7408) );
  NAND2_X1 U9193 ( .A1(n7408), .A2(n7546), .ZN(n7554) );
  INV_X1 U9194 ( .A(n7408), .ZN(n7409) );
  NAND2_X1 U9195 ( .A1(n7410), .A2(n7409), .ZN(n7411) );
  AND2_X1 U9196 ( .A1(n7554), .A2(n7411), .ZN(n7412) );
  OAI21_X1 U9197 ( .B1(n7414), .B2(n7413), .A(n7412), .ZN(n7555) );
  INV_X1 U9198 ( .A(n7555), .ZN(n7416) );
  NOR3_X1 U9199 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(n7415) );
  OAI21_X1 U9200 ( .B1(n7416), .B2(n7415), .A(n8683), .ZN(n7417) );
  OAI211_X1 U9201 ( .C1(n7419), .C2(n8685), .A(n7418), .B(n7417), .ZN(P2_U3194) );
  INV_X1 U9202 ( .A(n7420), .ZN(n7431) );
  OAI222_X1 U9203 ( .A1(n9640), .A2(n7431), .B1(n7993), .B2(P1_U3086), .C1(
        n7421), .C2(n8084), .ZN(P1_U3334) );
  XNOR2_X1 U9204 ( .A(n7422), .B(n8382), .ZN(n7423) );
  AOI222_X1 U9205 ( .A1(n9902), .A2(n7423), .B1(n8519), .B2(n9872), .C1(n8521), 
        .C2(n9874), .ZN(n7433) );
  MUX2_X1 U9206 ( .A(n7407), .B(n7433), .S(n9956), .Z(n7426) );
  INV_X1 U9207 ( .A(n8382), .ZN(n8486) );
  XNOR2_X1 U9208 ( .A(n7424), .B(n8486), .ZN(n7432) );
  NAND2_X1 U9209 ( .A1(n9956), .A2(n9884), .ZN(n8958) );
  INV_X1 U9210 ( .A(n8958), .ZN(n8954) );
  AOI22_X1 U9211 ( .A1(n7432), .A2(n8954), .B1(n8953), .B2(n7494), .ZN(n7425)
         );
  NAND2_X1 U9212 ( .A1(n7426), .A2(n7425), .ZN(P2_U3471) );
  MUX2_X1 U9213 ( .A(n7427), .B(n7433), .S(n9941), .Z(n7429) );
  INV_X1 U9214 ( .A(n9032), .ZN(n9025) );
  AOI22_X1 U9215 ( .A1(n7432), .A2(n9025), .B1(n9024), .B2(n7494), .ZN(n7428)
         );
  NAND2_X1 U9216 ( .A1(n7429), .A2(n7428), .ZN(P2_U3426) );
  OAI222_X1 U9217 ( .A1(n8323), .A2(P2_U3151), .B1(n9044), .B2(n7431), .C1(
        n7430), .C2(n9042), .ZN(P2_U3274) );
  INV_X1 U9218 ( .A(n7432), .ZN(n7437) );
  MUX2_X1 U9219 ( .A(n7541), .B(n7433), .S(n8859), .Z(n7436) );
  INV_X1 U9220 ( .A(n7492), .ZN(n7434) );
  AOI22_X1 U9221 ( .A1(n7494), .A2(n8861), .B1(n8848), .B2(n7434), .ZN(n7435)
         );
  OAI211_X1 U9222 ( .C1(n7437), .C2(n8864), .A(n7436), .B(n7435), .ZN(P2_U3221) );
  OAI21_X1 U9223 ( .B1(n7439), .B2(n7440), .A(n7438), .ZN(n7453) );
  AOI211_X1 U9224 ( .C1(n7454), .C2(n4349), .A(n9509), .B(n4290), .ZN(n7455)
         );
  XNOR2_X1 U9225 ( .A(n7441), .B(n7440), .ZN(n7442) );
  NAND2_X1 U9226 ( .A1(n7442), .A2(n9504), .ZN(n7445) );
  OAI22_X1 U9227 ( .A1(n7810), .A2(n9458), .B1(n7610), .B2(n9456), .ZN(n7443)
         );
  INV_X1 U9228 ( .A(n7443), .ZN(n7444) );
  NAND2_X1 U9229 ( .A1(n7445), .A2(n7444), .ZN(n7459) );
  AOI211_X1 U9230 ( .C1(n7453), .C2(n9835), .A(n7455), .B(n7459), .ZN(n7452)
         );
  INV_X1 U9231 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7446) );
  NOR2_X1 U9232 ( .A1(n9627), .A2(n7446), .ZN(n7447) );
  AOI21_X1 U9233 ( .B1(n7454), .B2(n7448), .A(n7447), .ZN(n7449) );
  OAI21_X1 U9234 ( .B1(n7452), .B2(n9846), .A(n7449), .ZN(P1_U3489) );
  INV_X1 U9235 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9304) );
  AOI22_X1 U9236 ( .A1(n7454), .A2(n7450), .B1(n5802), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7451) );
  OAI21_X1 U9237 ( .B1(n7452), .B2(n5802), .A(n7451), .ZN(P1_U3534) );
  INV_X1 U9238 ( .A(n7453), .ZN(n7461) );
  NAND2_X1 U9239 ( .A1(n7455), .A2(n9512), .ZN(n7457) );
  AOI22_X1 U9240 ( .A1(n9494), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7612), .B2(
        n9800), .ZN(n7456) );
  OAI211_X1 U9241 ( .C1(n5695), .C2(n9516), .A(n7457), .B(n7456), .ZN(n7458)
         );
  AOI21_X1 U9242 ( .B1(n9518), .B2(n7459), .A(n7458), .ZN(n7460) );
  OAI21_X1 U9243 ( .B1(n7461), .B2(n9520), .A(n7460), .ZN(P1_U3281) );
  INV_X1 U9244 ( .A(n8393), .ZN(n7462) );
  XNOR2_X1 U9245 ( .A(n7463), .B(n8487), .ZN(n7464) );
  AOI222_X1 U9246 ( .A1(n9902), .A2(n7464), .B1(n8855), .B2(n9872), .C1(n8520), 
        .C2(n9874), .ZN(n8867) );
  MUX2_X1 U9247 ( .A(n7550), .B(n8867), .S(n9956), .Z(n7467) );
  XOR2_X1 U9248 ( .A(n7465), .B(n8487), .Z(n8873) );
  AOI22_X1 U9249 ( .A1(n8873), .A2(n8954), .B1(n8953), .B2(n8870), .ZN(n7466)
         );
  NAND2_X1 U9250 ( .A1(n7467), .A2(n7466), .ZN(P2_U3472) );
  INV_X1 U9251 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7468) );
  MUX2_X1 U9252 ( .A(n7468), .B(n8867), .S(n9941), .Z(n7470) );
  AOI22_X1 U9253 ( .A1(n8873), .A2(n9025), .B1(n9024), .B2(n8870), .ZN(n7469)
         );
  NAND2_X1 U9254 ( .A1(n7470), .A2(n7469), .ZN(P2_U3429) );
  XNOR2_X1 U9255 ( .A(n7471), .B(n7472), .ZN(n7473) );
  NAND2_X1 U9256 ( .A1(n7473), .A2(n7474), .ZN(n7515) );
  OAI21_X1 U9257 ( .B1(n7474), .B2(n7473), .A(n7515), .ZN(n7475) );
  NAND2_X1 U9258 ( .A1(n7475), .A2(n9151), .ZN(n7483) );
  NOR2_X1 U9259 ( .A1(n9157), .A2(n7476), .ZN(n7480) );
  OR2_X1 U9260 ( .A1(n9662), .A2(n7477), .ZN(n7478) );
  NAND2_X1 U9261 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9271) );
  OAI211_X1 U9262 ( .C1(n9661), .C2(n7585), .A(n7478), .B(n9271), .ZN(n7479)
         );
  AOI211_X1 U9263 ( .C1(n7481), .C2(n9161), .A(n7480), .B(n7479), .ZN(n7482)
         );
  NAND2_X1 U9264 ( .A1(n7483), .A2(n7482), .ZN(P1_U3221) );
  XOR2_X1 U9265 ( .A(n8131), .B(n8483), .Z(n7503) );
  NOR2_X1 U9266 ( .A1(n7502), .A2(n7503), .ZN(n7501) );
  XOR2_X1 U9267 ( .A(n8131), .B(n7494), .Z(n8087) );
  XNOR2_X1 U9268 ( .A(n8087), .B(n8520), .ZN(n7487) );
  XNOR2_X1 U9269 ( .A(n8089), .B(n7487), .ZN(n7496) );
  NOR2_X1 U9270 ( .A1(n8257), .A2(n7488), .ZN(n7489) );
  AOI211_X1 U9271 ( .C1(n8277), .C2(n8519), .A(n7490), .B(n7489), .ZN(n7491)
         );
  OAI21_X1 U9272 ( .B1(n7492), .B2(n8287), .A(n7491), .ZN(n7493) );
  AOI21_X1 U9273 ( .B1(n7494), .B2(n8259), .A(n7493), .ZN(n7495) );
  OAI21_X1 U9274 ( .B1(n7496), .B2(n8280), .A(n7495), .ZN(P2_U3164) );
  NOR2_X1 U9275 ( .A1(n8257), .A2(n9920), .ZN(n7497) );
  AOI211_X1 U9276 ( .C1(n8277), .C2(n8520), .A(n7498), .B(n7497), .ZN(n7499)
         );
  OAI21_X1 U9277 ( .B1(n7500), .B2(n8287), .A(n7499), .ZN(n7505) );
  AOI211_X1 U9278 ( .C1(n7503), .C2(n7502), .A(n8280), .B(n7501), .ZN(n7504)
         );
  AOI211_X1 U9279 ( .C1(n9939), .C2(n8259), .A(n7505), .B(n7504), .ZN(n7506)
         );
  INV_X1 U9280 ( .A(n7506), .ZN(P2_U3176) );
  XNOR2_X1 U9281 ( .A(n7507), .B(n8395), .ZN(n9033) );
  OAI211_X1 U9282 ( .C1(n7509), .C2(n8395), .A(n7508), .B(n9902), .ZN(n7511)
         );
  AOI22_X1 U9283 ( .A1(n8518), .A2(n9872), .B1(n9874), .B2(n8519), .ZN(n7510)
         );
  NAND2_X1 U9284 ( .A1(n7511), .A2(n7510), .ZN(n9029) );
  INV_X1 U9285 ( .A(n8092), .ZN(n9031) );
  OAI22_X1 U9286 ( .A1(n9031), .A2(n8752), .B1(n8158), .B2(n8882), .ZN(n7512)
         );
  OAI21_X1 U9287 ( .B1(n9029), .B2(n7512), .A(n8859), .ZN(n7514) );
  NAND2_X1 U9288 ( .A1(n8890), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7513) );
  OAI211_X1 U9289 ( .C1(n9033), .C2(n8864), .A(n7514), .B(n7513), .ZN(P2_U3219) );
  OAI21_X1 U9290 ( .B1(n7516), .B2(n7471), .A(n7515), .ZN(n7520) );
  XNOR2_X1 U9291 ( .A(n7518), .B(n7517), .ZN(n7519) );
  XNOR2_X1 U9292 ( .A(n7520), .B(n7519), .ZN(n7529) );
  NOR2_X1 U9293 ( .A1(n9678), .A2(n7521), .ZN(n7526) );
  NAND2_X1 U9294 ( .A1(n9152), .A2(n9184), .ZN(n7523) );
  OAI211_X1 U9295 ( .C1(n7524), .C2(n9662), .A(n7523), .B(n7522), .ZN(n7525)
         );
  AOI211_X1 U9296 ( .C1(n7527), .C2(n9675), .A(n7526), .B(n7525), .ZN(n7528)
         );
  OAI21_X1 U9297 ( .B1(n7529), .B2(n9671), .A(n7528), .ZN(P1_U3231) );
  OAI21_X1 U9298 ( .B1(n7531), .B2(n8010), .A(n7530), .ZN(n7570) );
  INV_X1 U9299 ( .A(n7570), .ZN(n7540) );
  INV_X1 U9300 ( .A(n7532), .ZN(n7617) );
  AOI21_X1 U9301 ( .B1(n7533), .B2(n8010), .A(n7617), .ZN(n7534) );
  OAI222_X1 U9302 ( .A1(n9456), .A2(n9660), .B1(n9458), .B2(n7535), .C1(n9453), 
        .C2(n7534), .ZN(n7568) );
  INV_X1 U9303 ( .A(n7811), .ZN(n7812) );
  OAI211_X1 U9304 ( .C1(n7812), .C2(n4290), .A(n4350), .B(n9551), .ZN(n7567)
         );
  NOR2_X1 U9305 ( .A1(n7567), .A2(n9806), .ZN(n7538) );
  AOI22_X1 U9306 ( .A1(n9813), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n4861), .B2(
        n9800), .ZN(n7536) );
  OAI21_X1 U9307 ( .B1(n7812), .B2(n9516), .A(n7536), .ZN(n7537) );
  AOI211_X1 U9308 ( .C1(n7568), .C2(n9518), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9309 ( .B1(n9520), .B2(n7540), .A(n7539), .ZN(P1_U3280) );
  OR2_X1 U9310 ( .A1(n7546), .A2(n7541), .ZN(n7542) );
  AOI21_X1 U9311 ( .B1(n7551), .B2(n7544), .A(n7631), .ZN(n7562) );
  NAND2_X1 U9312 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7547), .ZN(n7637) );
  OAI21_X1 U9313 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7547), .A(n7637), .ZN(
        n7560) );
  INV_X1 U9314 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9315 ( .A1(n8587), .A2(n7630), .ZN(n7548) );
  NAND2_X1 U9316 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8243) );
  OAI211_X1 U9317 ( .C1(n7549), .C2(n8653), .A(n7548), .B(n8243), .ZN(n7559)
         );
  MUX2_X1 U9318 ( .A(n7551), .B(n7550), .S(n8665), .Z(n7552) );
  NAND2_X1 U9319 ( .A1(n7630), .A2(n7552), .ZN(n7641) );
  OAI21_X1 U9320 ( .B1(n7630), .B2(n7552), .A(n7641), .ZN(n7553) );
  AOI21_X1 U9321 ( .B1(n7555), .B2(n7554), .A(n7553), .ZN(n7647) );
  INV_X1 U9322 ( .A(n7647), .ZN(n7557) );
  NAND3_X1 U9323 ( .A1(n7555), .A2(n7554), .A3(n7553), .ZN(n7556) );
  AOI21_X1 U9324 ( .B1(n7557), .B2(n7556), .A(n8617), .ZN(n7558) );
  AOI211_X1 U9325 ( .C1(n7560), .C2(n8624), .A(n7559), .B(n7558), .ZN(n7561)
         );
  OAI21_X1 U9326 ( .B1(n7562), .B2(n8685), .A(n7561), .ZN(P2_U3195) );
  INV_X1 U9327 ( .A(n7563), .ZN(n7566) );
  OAI222_X1 U9328 ( .A1(n8084), .A2(n7565), .B1(n9640), .B2(n7566), .C1(
        P1_U3086), .C2(n7564), .ZN(P1_U3333) );
  OAI222_X1 U9329 ( .A1(P2_U3151), .A2(n8322), .B1(n9044), .B2(n7566), .C1(
        n10005), .C2(n9042), .ZN(P2_U3273) );
  OAI21_X1 U9330 ( .B1(n7812), .B2(n9831), .A(n7567), .ZN(n7569) );
  AOI211_X1 U9331 ( .C1(n9835), .C2(n7570), .A(n7569), .B(n7568), .ZN(n7573)
         );
  NAND2_X1 U9332 ( .A1(n5802), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7571) );
  OAI21_X1 U9333 ( .B1(n7573), .B2(n5802), .A(n7571), .ZN(P1_U3535) );
  NAND2_X1 U9334 ( .A1(n9846), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7572) );
  OAI21_X1 U9335 ( .B1(n7573), .B2(n9846), .A(n7572), .ZN(P1_U3492) );
  INV_X1 U9336 ( .A(n7577), .ZN(n7575) );
  NAND2_X1 U9337 ( .A1(n9638), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7574) );
  OAI211_X1 U9338 ( .C1(n7575), .C2(n9640), .A(n8054), .B(n7574), .ZN(P1_U3332) );
  NAND2_X1 U9339 ( .A1(n7577), .A2(n7576), .ZN(n7579) );
  NAND2_X1 U9340 ( .A1(n7578), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8511) );
  OAI211_X1 U9341 ( .C1(n10120), .C2(n9042), .A(n7579), .B(n8511), .ZN(
        P2_U3272) );
  XNOR2_X1 U9342 ( .A(n7580), .B(n9668), .ZN(n7582) );
  NOR2_X1 U9343 ( .A1(n7582), .A2(n7581), .ZN(n9667) );
  AOI21_X1 U9344 ( .B1(n7582), .B2(n7581), .A(n9667), .ZN(n7592) );
  INV_X1 U9345 ( .A(n7583), .ZN(n7584) );
  NOR2_X1 U9346 ( .A1(n9678), .A2(n7584), .ZN(n7590) );
  INV_X1 U9347 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9999) );
  OAI22_X1 U9348 ( .A1(n9661), .A2(n7610), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9999), .ZN(n7589) );
  NOR2_X1 U9349 ( .A1(n9662), .A2(n7585), .ZN(n7588) );
  NOR2_X1 U9350 ( .A1(n7586), .A2(n9157), .ZN(n7587) );
  NOR4_X1 U9351 ( .A1(n7590), .A2(n7589), .A3(n7588), .A4(n7587), .ZN(n7591)
         );
  OAI21_X1 U9352 ( .B1(n7592), .B2(n9671), .A(n7591), .ZN(P1_U3217) );
  INV_X1 U9353 ( .A(n7594), .ZN(n8013) );
  XNOR2_X1 U9354 ( .A(n7593), .B(n8013), .ZN(n7685) );
  INV_X1 U9355 ( .A(n7685), .ZN(n7605) );
  NAND2_X1 U9356 ( .A1(n7618), .A2(n7930), .ZN(n7595) );
  XNOR2_X1 U9357 ( .A(n7595), .B(n7594), .ZN(n7596) );
  NAND2_X1 U9358 ( .A1(n7596), .A2(n9504), .ZN(n7598) );
  AND2_X1 U9359 ( .A1(n9180), .A2(n9425), .ZN(n7597) );
  AOI21_X1 U9360 ( .B1(n9178), .B2(n9427), .A(n7597), .ZN(n9165) );
  NAND2_X1 U9361 ( .A1(n7598), .A2(n9165), .ZN(n7683) );
  INV_X1 U9362 ( .A(n7623), .ZN(n7600) );
  AOI211_X1 U9363 ( .C1(n9167), .C2(n7600), .A(n9509), .B(n7599), .ZN(n7684)
         );
  NAND2_X1 U9364 ( .A1(n7684), .A2(n9512), .ZN(n7602) );
  AOI22_X1 U9365 ( .A1(n9494), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9160), .B2(
        n9800), .ZN(n7601) );
  OAI211_X1 U9366 ( .C1(n7690), .C2(n9516), .A(n7602), .B(n7601), .ZN(n7603)
         );
  AOI21_X1 U9367 ( .B1(n9518), .B2(n7683), .A(n7603), .ZN(n7604) );
  OAI21_X1 U9368 ( .B1(n7605), .B2(n9520), .A(n7604), .ZN(P1_U3278) );
  OAI21_X1 U9369 ( .B1(n7607), .B2(n4351), .A(n7606), .ZN(n7608) );
  NAND2_X1 U9370 ( .A1(n7608), .A2(n9151), .ZN(n7614) );
  NAND2_X1 U9371 ( .A1(n9152), .A2(n9181), .ZN(n7609) );
  NAND2_X1 U9372 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9712) );
  OAI211_X1 U9373 ( .C1(n7610), .C2(n9662), .A(n7609), .B(n9712), .ZN(n7611)
         );
  AOI21_X1 U9374 ( .B1(n7612), .B2(n9161), .A(n7611), .ZN(n7613) );
  OAI211_X1 U9375 ( .C1(n5695), .C2(n9157), .A(n7614), .B(n7613), .ZN(P1_U3224) );
  INV_X1 U9376 ( .A(n7819), .ZN(n8012) );
  XNOR2_X1 U9377 ( .A(n7615), .B(n8012), .ZN(n7720) );
  AOI22_X1 U9378 ( .A1(n9181), .A2(n9425), .B1(n9427), .B2(n9179), .ZN(n7621)
         );
  OAI21_X1 U9379 ( .B1(n7617), .B2(n7616), .A(n7819), .ZN(n7619) );
  NAND3_X1 U9380 ( .A1(n7619), .A2(n7618), .A3(n9504), .ZN(n7620) );
  OAI211_X1 U9381 ( .C1(n7720), .C2(n7622), .A(n7621), .B(n7620), .ZN(n7721)
         );
  NAND2_X1 U9382 ( .A1(n7721), .A2(n9518), .ZN(n7628) );
  AOI211_X1 U9383 ( .C1(n7624), .C2(n4350), .A(n9509), .B(n7623), .ZN(n7722)
         );
  AOI22_X1 U9384 ( .A1(n9494), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7745), .B2(
        n9800), .ZN(n7625) );
  OAI21_X1 U9385 ( .B1(n7742), .B2(n9516), .A(n7625), .ZN(n7626) );
  AOI21_X1 U9386 ( .B1(n7722), .B2(n9512), .A(n7626), .ZN(n7627) );
  OAI211_X1 U9387 ( .C1(n7720), .C2(n7629), .A(n7628), .B(n7627), .ZN(P1_U3279) );
  NOR2_X1 U9388 ( .A1(n7630), .A2(n4316), .ZN(n7632) );
  AOI22_X1 U9389 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8558), .B1(n8554), .B2(
        n7642), .ZN(n7633) );
  NOR2_X1 U9390 ( .A1(n7634), .A2(n7633), .ZN(n8553) );
  AOI21_X1 U9391 ( .B1(n7634), .B2(n7633), .A(n8553), .ZN(n7656) );
  AOI22_X1 U9392 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8554), .B1(n8558), .B2(
        n8557), .ZN(n7640) );
  NAND2_X1 U9393 ( .A1(n7636), .A2(n7635), .ZN(n7638) );
  NAND2_X1 U9394 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  OAI21_X1 U9395 ( .B1(n7640), .B2(n7639), .A(n8556), .ZN(n7654) );
  INV_X1 U9396 ( .A(n7641), .ZN(n7646) );
  MUX2_X1 U9397 ( .A(n7642), .B(n8557), .S(n8665), .Z(n7643) );
  OR2_X1 U9398 ( .A1(n8558), .A2(n7643), .ZN(n7644) );
  NAND2_X1 U9399 ( .A1(n8558), .A2(n7643), .ZN(n8567) );
  AND2_X1 U9400 ( .A1(n7644), .A2(n8567), .ZN(n7645) );
  OAI21_X1 U9401 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n8568) );
  INV_X1 U9402 ( .A(n8568), .ZN(n7649) );
  NOR3_X1 U9403 ( .A1(n7647), .A2(n7646), .A3(n7645), .ZN(n7648) );
  OAI21_X1 U9404 ( .B1(n7649), .B2(n7648), .A(n8683), .ZN(n7652) );
  INV_X1 U9405 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7650) );
  NOR2_X1 U9406 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7650), .ZN(n8159) );
  AOI21_X1 U9407 ( .B1(n8669), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n8159), .ZN(
        n7651) );
  OAI211_X1 U9408 ( .C1(n8673), .C2(n8554), .A(n7652), .B(n7651), .ZN(n7653)
         );
  AOI21_X1 U9409 ( .B1(n8624), .B2(n7654), .A(n7653), .ZN(n7655) );
  OAI21_X1 U9410 ( .B1(n7656), .B2(n8685), .A(n7655), .ZN(P2_U3196) );
  INV_X1 U9411 ( .A(n7657), .ZN(n8069) );
  OAI222_X1 U9412 ( .A1(n7659), .A2(P2_U3151), .B1(n9048), .B2(n8069), .C1(
        n7658), .C2(n9042), .ZN(P2_U3271) );
  XNOR2_X1 U9413 ( .A(n7660), .B(n7661), .ZN(n9587) );
  INV_X1 U9414 ( .A(n9587), .ZN(n7674) );
  XNOR2_X1 U9415 ( .A(n7662), .B(n7661), .ZN(n7663) );
  NAND2_X1 U9416 ( .A1(n7663), .A2(n9504), .ZN(n7666) );
  NAND2_X1 U9417 ( .A1(n9179), .A2(n9425), .ZN(n7665) );
  NAND2_X1 U9418 ( .A1(n9177), .A2(n9427), .ZN(n7664) );
  AND2_X1 U9419 ( .A1(n7665), .A2(n7664), .ZN(n9089) );
  NAND2_X1 U9420 ( .A1(n7666), .A2(n9089), .ZN(n9585) );
  INV_X1 U9421 ( .A(n7599), .ZN(n7668) );
  INV_X1 U9422 ( .A(n7715), .ZN(n7667) );
  AOI211_X1 U9423 ( .C1(n7669), .C2(n7668), .A(n9509), .B(n7667), .ZN(n9586)
         );
  NAND2_X1 U9424 ( .A1(n9586), .A2(n9512), .ZN(n7671) );
  AOI22_X1 U9425 ( .A1(n9494), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9091), .B2(
        n9800), .ZN(n7670) );
  OAI211_X1 U9426 ( .C1(n9632), .C2(n9516), .A(n7671), .B(n7670), .ZN(n7672)
         );
  AOI21_X1 U9427 ( .B1(n9518), .B2(n9585), .A(n7672), .ZN(n7673) );
  OAI21_X1 U9428 ( .B1(n7674), .B2(n9520), .A(n7673), .ZN(P1_U3277) );
  OAI21_X1 U9429 ( .B1(n7677), .B2(n7676), .A(n7675), .ZN(n7678) );
  NAND2_X1 U9430 ( .A1(n7678), .A2(n9151), .ZN(n7682) );
  NAND2_X1 U9431 ( .A1(n9152), .A2(n9180), .ZN(n7679) );
  NAND2_X1 U9432 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9728) );
  OAI211_X1 U9433 ( .C1(n9660), .C2(n9662), .A(n7679), .B(n9728), .ZN(n7680)
         );
  AOI21_X1 U9434 ( .B1(n4861), .B2(n9161), .A(n7680), .ZN(n7681) );
  OAI211_X1 U9435 ( .C1(n7812), .C2(n9157), .A(n7682), .B(n7681), .ZN(P1_U3234) );
  INV_X1 U9436 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9747) );
  AOI211_X1 U9437 ( .C1(n7685), .C2(n9835), .A(n7684), .B(n7683), .ZN(n7687)
         );
  MUX2_X1 U9438 ( .A(n9747), .B(n7687), .S(n9854), .Z(n7686) );
  OAI21_X1 U9439 ( .B1(n7690), .B2(n9590), .A(n7686), .ZN(P1_U3537) );
  INV_X1 U9440 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7688) );
  MUX2_X1 U9441 ( .A(n7688), .B(n7687), .S(n9627), .Z(n7689) );
  OAI21_X1 U9442 ( .B1(n7690), .B2(n9631), .A(n7689), .ZN(P1_U3498) );
  INV_X1 U9443 ( .A(n7691), .ZN(n7732) );
  OAI222_X1 U9444 ( .A1(n8084), .A2(n7693), .B1(n9640), .B2(n7732), .C1(
        P1_U3086), .C2(n7692), .ZN(P1_U3330) );
  OAI211_X1 U9445 ( .C1(n7695), .C2(n8491), .A(n7694), .B(n9902), .ZN(n7698)
         );
  OAI22_X1 U9446 ( .A1(n8095), .A2(n9917), .B1(n8831), .B2(n9919), .ZN(n7696)
         );
  INV_X1 U9447 ( .A(n7696), .ZN(n7697) );
  NAND2_X1 U9448 ( .A1(n7698), .A2(n7697), .ZN(n7705) );
  MUX2_X1 U9449 ( .A(n7705), .B(P2_REG0_REG_16__SCAN_IN), .S(n9943), .Z(n7702)
         );
  INV_X1 U9450 ( .A(n8491), .ZN(n7700) );
  XNOR2_X1 U9451 ( .A(n7699), .B(n7700), .ZN(n7707) );
  INV_X1 U9452 ( .A(n8098), .ZN(n8210) );
  OAI22_X1 U9453 ( .A1(n7707), .A2(n9032), .B1(n8210), .B2(n9030), .ZN(n7701)
         );
  OR2_X1 U9454 ( .A1(n7702), .A2(n7701), .ZN(P2_U3438) );
  MUX2_X1 U9455 ( .A(n7705), .B(P2_REG1_REG_16__SCAN_IN), .S(n4414), .Z(n7704)
         );
  OAI22_X1 U9456 ( .A1(n7707), .A2(n8958), .B1(n8210), .B2(n8957), .ZN(n7703)
         );
  OR2_X1 U9457 ( .A1(n7704), .A2(n7703), .ZN(P2_U3475) );
  MUX2_X1 U9458 ( .A(n7705), .B(P2_REG2_REG_16__SCAN_IN), .S(n8890), .Z(n7709)
         );
  AOI22_X1 U9459 ( .A1(n8098), .A2(n8861), .B1(n8848), .B2(n8213), .ZN(n7706)
         );
  OAI21_X1 U9460 ( .B1(n7707), .B2(n8864), .A(n7706), .ZN(n7708) );
  OR2_X1 U9461 ( .A1(n7709), .A2(n7708), .ZN(P2_U3217) );
  XNOR2_X1 U9462 ( .A(n7710), .B(n4294), .ZN(n9584) );
  OAI211_X1 U9463 ( .C1(n4859), .C2(n4294), .A(n9504), .B(n7711), .ZN(n7713)
         );
  AOI22_X1 U9464 ( .A1(n9178), .A2(n9425), .B1(n9427), .B2(n9176), .ZN(n7712)
         );
  NAND2_X1 U9465 ( .A1(n7713), .A2(n7712), .ZN(n9579) );
  INV_X1 U9466 ( .A(n9510), .ZN(n7714) );
  AOI211_X1 U9467 ( .C1(n9581), .C2(n7715), .A(n9509), .B(n7714), .ZN(n9580)
         );
  NAND2_X1 U9468 ( .A1(n9580), .A2(n9512), .ZN(n7717) );
  AOI22_X1 U9469 ( .A1(n9494), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9103), .B2(
        n9800), .ZN(n7716) );
  OAI211_X1 U9470 ( .C1(n9100), .C2(n9516), .A(n7717), .B(n7716), .ZN(n7718)
         );
  AOI21_X1 U9471 ( .B1(n9518), .B2(n9579), .A(n7718), .ZN(n7719) );
  OAI21_X1 U9472 ( .B1(n9584), .B2(n9520), .A(n7719), .ZN(P1_U3276) );
  INV_X1 U9473 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7724) );
  INV_X1 U9474 ( .A(n7720), .ZN(n7723) );
  AOI211_X1 U9475 ( .C1(n9842), .C2(n7723), .A(n7722), .B(n7721), .ZN(n7726)
         );
  MUX2_X1 U9476 ( .A(n7724), .B(n7726), .S(n9854), .Z(n7725) );
  OAI21_X1 U9477 ( .B1(n7742), .B2(n9590), .A(n7725), .ZN(P1_U3536) );
  INV_X1 U9478 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7727) );
  MUX2_X1 U9479 ( .A(n7727), .B(n7726), .S(n9627), .Z(n7728) );
  OAI21_X1 U9480 ( .B1(n7742), .B2(n9631), .A(n7728), .ZN(P1_U3495) );
  INV_X1 U9481 ( .A(n7729), .ZN(n7737) );
  OAI222_X1 U9482 ( .A1(n9640), .A2(n7737), .B1(n7731), .B2(P1_U3086), .C1(
        n7730), .C2(n8084), .ZN(P1_U3329) );
  OAI222_X1 U9483 ( .A1(P2_U3151), .A2(n7733), .B1(n9048), .B2(n7732), .C1(
        n9042), .C2(n6166), .ZN(P2_U3270) );
  INV_X1 U9484 ( .A(n7734), .ZN(n8066) );
  AOI21_X1 U9485 ( .B1(n9046), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7735), .ZN(
        n7736) );
  OAI21_X1 U9486 ( .B1(n8066), .B2(n9048), .A(n7736), .ZN(P2_U3268) );
  OAI222_X1 U9487 ( .A1(n7738), .A2(P2_U3151), .B1(n9048), .B2(n7737), .C1(
        n10076), .C2(n9042), .ZN(P2_U3269) );
  AOI21_X1 U9488 ( .B1(n7740), .B2(n7739), .A(n4342), .ZN(n7747) );
  NAND2_X1 U9489 ( .A1(n9152), .A2(n9179), .ZN(n7741) );
  NAND2_X1 U9490 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9744) );
  OAI211_X1 U9491 ( .C1(n7810), .C2(n9662), .A(n7741), .B(n9744), .ZN(n7744)
         );
  NOR2_X1 U9492 ( .A1(n7742), .A2(n9157), .ZN(n7743) );
  AOI211_X1 U9493 ( .C1(n7745), .C2(n9161), .A(n7744), .B(n7743), .ZN(n7746)
         );
  OAI21_X1 U9494 ( .B1(n7747), .B2(n9671), .A(n7746), .ZN(P1_U3215) );
  INV_X1 U9495 ( .A(n7748), .ZN(n7749) );
  NAND2_X1 U9496 ( .A1(n7749), .A2(SI_29_), .ZN(n7753) );
  NAND2_X1 U9497 ( .A1(n7753), .A2(n7752), .ZN(n7886) );
  INV_X1 U9498 ( .A(n7886), .ZN(n7760) );
  INV_X1 U9499 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7754) );
  INV_X1 U9500 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9043) );
  MUX2_X1 U9501 ( .A(n7754), .B(n9043), .S(n8295), .Z(n7756) );
  INV_X1 U9502 ( .A(SI_30_), .ZN(n7755) );
  NAND2_X1 U9503 ( .A1(n7756), .A2(n7755), .ZN(n7761) );
  INV_X1 U9504 ( .A(n7756), .ZN(n7757) );
  NAND2_X1 U9505 ( .A1(n7757), .A2(SI_30_), .ZN(n7758) );
  NAND2_X1 U9506 ( .A1(n7761), .A2(n7758), .ZN(n7885) );
  INV_X1 U9507 ( .A(n7885), .ZN(n7759) );
  INV_X1 U9508 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7762) );
  MUX2_X1 U9509 ( .A(n7762), .B(n6592), .S(n8295), .Z(n7763) );
  XNOR2_X1 U9510 ( .A(n7763), .B(SI_31_), .ZN(n7764) );
  NAND2_X1 U9511 ( .A1(n9036), .A2(n7889), .ZN(n7767) );
  NAND2_X1 U9512 ( .A1(n7890), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7766) );
  AOI211_X1 U9513 ( .C1(n8042), .C2(n9321), .A(n5651), .B(n7768), .ZN(n7906)
         );
  NAND3_X1 U9514 ( .A1(n7839), .A2(n9622), .A3(n7836), .ZN(n7769) );
  OAI21_X1 U9515 ( .B1(n7770), .B2(n7905), .A(n7769), .ZN(n7772) );
  NAND2_X1 U9516 ( .A1(n7772), .A2(n7771), .ZN(n7774) );
  NAND3_X1 U9517 ( .A1(n7839), .A2(n7905), .A3(n7836), .ZN(n7773) );
  NAND2_X1 U9518 ( .A1(n7774), .A2(n7773), .ZN(n7847) );
  INV_X1 U9519 ( .A(n7775), .ZN(n7777) );
  MUX2_X1 U9520 ( .A(n7777), .B(n7776), .S(n7905), .Z(n7783) );
  INV_X1 U9521 ( .A(n7917), .ZN(n7778) );
  NAND2_X1 U9522 ( .A1(n7781), .A2(n7780), .ZN(n7782) );
  INV_X1 U9523 ( .A(n7905), .ZN(n7897) );
  AND2_X1 U9524 ( .A1(n7786), .A2(n8000), .ZN(n7788) );
  MUX2_X1 U9525 ( .A(n7788), .B(n7787), .S(n7897), .Z(n7793) );
  NAND2_X1 U9526 ( .A1(n7795), .A2(n7789), .ZN(n7790) );
  MUX2_X1 U9527 ( .A(n7791), .B(n7790), .S(n7905), .Z(n7792) );
  AOI21_X1 U9528 ( .B1(n7794), .B2(n7793), .A(n7792), .ZN(n7801) );
  INV_X1 U9529 ( .A(n7795), .ZN(n7796) );
  OAI21_X1 U9530 ( .B1(n7801), .B2(n7796), .A(n7922), .ZN(n7797) );
  AND2_X1 U9531 ( .A1(n7804), .A2(n7799), .ZN(n7926) );
  NAND2_X1 U9532 ( .A1(n7806), .A2(n7802), .ZN(n7925) );
  AOI21_X1 U9533 ( .B1(n7797), .B2(n7926), .A(n7925), .ZN(n7824) );
  NAND4_X1 U9534 ( .A1(n7815), .A2(n7928), .A3(n7929), .A4(n7897), .ZN(n7823)
         );
  INV_X1 U9535 ( .A(n7798), .ZN(n7800) );
  OAI21_X1 U9536 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7803) );
  NAND3_X1 U9537 ( .A1(n7803), .A2(n7802), .A3(n7922), .ZN(n7805) );
  NAND3_X1 U9538 ( .A1(n7805), .A2(n7804), .A3(n7928), .ZN(n7809) );
  NAND3_X1 U9539 ( .A1(n7931), .A2(n7905), .A3(n7806), .ZN(n7807) );
  NOR2_X1 U9540 ( .A1(n7819), .A2(n7807), .ZN(n7808) );
  NAND2_X1 U9541 ( .A1(n7809), .A2(n7808), .ZN(n7822) );
  NAND3_X1 U9542 ( .A1(n7811), .A2(n7810), .A3(n7905), .ZN(n7818) );
  NAND4_X1 U9543 ( .A1(n7815), .A2(n7812), .A3(n9181), .A4(n7897), .ZN(n7813)
         );
  OAI211_X1 U9544 ( .C1(n7905), .C2(n7930), .A(n7825), .B(n7813), .ZN(n7814)
         );
  INV_X1 U9545 ( .A(n7814), .ZN(n7817) );
  NAND2_X1 U9546 ( .A1(n7827), .A2(n7815), .ZN(n7934) );
  NAND2_X1 U9547 ( .A1(n7934), .A2(n7905), .ZN(n7816) );
  OAI211_X1 U9548 ( .C1(n7819), .C2(n7818), .A(n7817), .B(n7816), .ZN(n7820)
         );
  NOR2_X1 U9549 ( .A1(n8015), .A2(n7820), .ZN(n7821) );
  OAI211_X1 U9550 ( .C1(n7824), .C2(n7823), .A(n7822), .B(n7821), .ZN(n7833)
         );
  INV_X1 U9551 ( .A(n7825), .ZN(n7935) );
  NAND2_X1 U9552 ( .A1(n7938), .A2(n7935), .ZN(n7826) );
  AND2_X1 U9553 ( .A1(n7826), .A2(n7939), .ZN(n7831) );
  INV_X1 U9554 ( .A(n7827), .ZN(n7828) );
  NAND2_X1 U9555 ( .A1(n7939), .A2(n7828), .ZN(n7829) );
  AND2_X1 U9556 ( .A1(n7829), .A2(n7938), .ZN(n7830) );
  MUX2_X1 U9557 ( .A(n7831), .B(n7830), .S(n7897), .Z(n7832) );
  NAND2_X1 U9558 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  NAND2_X1 U9559 ( .A1(n7834), .A2(n4294), .ZN(n7843) );
  AND2_X1 U9560 ( .A1(n7844), .A2(n7835), .ZN(n7946) );
  NAND2_X1 U9561 ( .A1(n7843), .A2(n7946), .ZN(n7837) );
  AND2_X1 U9562 ( .A1(n7836), .A2(n7842), .ZN(n7943) );
  NAND2_X1 U9563 ( .A1(n7837), .A2(n7943), .ZN(n7838) );
  NAND2_X1 U9564 ( .A1(n7847), .A2(n7838), .ZN(n7840) );
  AND2_X1 U9565 ( .A1(n7851), .A2(n7839), .ZN(n7954) );
  NAND3_X1 U9566 ( .A1(n7843), .A2(n7940), .A3(n7842), .ZN(n7845) );
  NAND3_X1 U9567 ( .A1(n7845), .A2(n7909), .A3(n7844), .ZN(n7846) );
  NAND2_X1 U9568 ( .A1(n7847), .A2(n7846), .ZN(n7850) );
  INV_X1 U9569 ( .A(n7848), .ZN(n7849) );
  OR2_X1 U9570 ( .A1(n9613), .A2(n9426), .ZN(n7852) );
  AND2_X1 U9571 ( .A1(n9400), .A2(n7852), .ZN(n7963) );
  INV_X1 U9572 ( .A(n7854), .ZN(n7853) );
  AOI21_X1 U9573 ( .B1(n7857), .B2(n7963), .A(n7853), .ZN(n7859) );
  INV_X1 U9574 ( .A(n9421), .ZN(n7855) );
  AND2_X1 U9575 ( .A1(n7855), .A2(n7854), .ZN(n7947) );
  AOI21_X1 U9576 ( .B1(n7857), .B2(n7947), .A(n7856), .ZN(n7858) );
  MUX2_X1 U9577 ( .A(n7964), .B(n7950), .S(n7905), .Z(n7861) );
  INV_X1 U9578 ( .A(n7952), .ZN(n7863) );
  NAND2_X1 U9579 ( .A1(n9355), .A2(n7965), .ZN(n7873) );
  INV_X1 U9580 ( .A(n7873), .ZN(n7862) );
  OR2_X1 U9581 ( .A1(n9374), .A2(n9387), .ZN(n7959) );
  NAND2_X1 U9582 ( .A1(n7864), .A2(n7959), .ZN(n7865) );
  NAND2_X1 U9583 ( .A1(n7865), .A2(n7876), .ZN(n7866) );
  NAND2_X1 U9584 ( .A1(n7866), .A2(n4860), .ZN(n7867) );
  NAND2_X1 U9585 ( .A1(n7867), .A2(n7877), .ZN(n7868) );
  NAND2_X1 U9586 ( .A1(n7868), .A2(n8024), .ZN(n7872) );
  INV_X1 U9587 ( .A(n7869), .ZN(n7870) );
  AOI21_X1 U9588 ( .B1(n7952), .B2(n7874), .A(n7873), .ZN(n7875) );
  NAND2_X1 U9589 ( .A1(n7973), .A2(n7959), .ZN(n8032) );
  NOR2_X1 U9590 ( .A1(n7875), .A2(n8032), .ZN(n7878) );
  NAND2_X1 U9591 ( .A1(n7877), .A2(n7876), .ZN(n7969) );
  OAI21_X1 U9592 ( .B1(n7878), .B2(n7969), .A(n7974), .ZN(n7879) );
  NAND2_X1 U9593 ( .A1(n8024), .A2(n7879), .ZN(n7882) );
  INV_X1 U9594 ( .A(n7975), .ZN(n7880) );
  NAND2_X1 U9595 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  NAND2_X1 U9596 ( .A1(n9041), .A2(n7889), .ZN(n7892) );
  NAND2_X1 U9597 ( .A1(n7890), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7891) );
  INV_X1 U9598 ( .A(n7901), .ZN(n7895) );
  OAI211_X1 U9599 ( .C1(n9326), .C2(n7897), .A(n9330), .B(n9171), .ZN(n7893)
         );
  INV_X1 U9600 ( .A(n7893), .ZN(n7894) );
  INV_X1 U9601 ( .A(n7896), .ZN(n7900) );
  AOI22_X1 U9602 ( .A1(n9326), .A2(n7897), .B1(n9329), .B2(n9171), .ZN(n7899)
         );
  OAI211_X1 U9603 ( .C1(n7901), .C2(n7900), .A(n7899), .B(n7898), .ZN(n7902)
         );
  NAND2_X1 U9604 ( .A1(n7903), .A2(n7902), .ZN(n7988) );
  INV_X1 U9605 ( .A(n7988), .ZN(n7904) );
  NOR2_X1 U9606 ( .A1(n5385), .A2(n7907), .ZN(n7983) );
  INV_X1 U9607 ( .A(n9171), .ZN(n7976) );
  NOR2_X1 U9608 ( .A1(n9326), .A2(n7976), .ZN(n8037) );
  INV_X1 U9609 ( .A(n8037), .ZN(n7908) );
  NAND2_X1 U9610 ( .A1(n8040), .A2(n7908), .ZN(n8026) );
  INV_X1 U9611 ( .A(n8026), .ZN(n7981) );
  INV_X1 U9612 ( .A(n7909), .ZN(n7958) );
  AOI21_X1 U9613 ( .B1(n9192), .B2(n7910), .A(n7993), .ZN(n7915) );
  INV_X1 U9614 ( .A(n7911), .ZN(n7913) );
  NAND2_X1 U9615 ( .A1(n5683), .A2(n4369), .ZN(n7912) );
  AND4_X1 U9616 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n7918)
         );
  NAND3_X1 U9617 ( .A1(n7918), .A2(n7917), .A3(n7916), .ZN(n7920) );
  NAND2_X1 U9618 ( .A1(n7920), .A2(n7919), .ZN(n7923) );
  OAI211_X1 U9619 ( .C1(n7924), .C2(n7923), .A(n7922), .B(n7921), .ZN(n7927)
         );
  AOI21_X1 U9620 ( .B1(n7927), .B2(n7926), .A(n7925), .ZN(n7933) );
  NAND2_X1 U9621 ( .A1(n7929), .A2(n7928), .ZN(n7932) );
  OAI211_X1 U9622 ( .C1(n7933), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7937)
         );
  INV_X1 U9623 ( .A(n7934), .ZN(n7936) );
  AOI21_X1 U9624 ( .B1(n7937), .B2(n7936), .A(n7935), .ZN(n7942) );
  INV_X1 U9625 ( .A(n7938), .ZN(n7941) );
  OAI211_X1 U9626 ( .C1(n7942), .C2(n7941), .A(n7940), .B(n7939), .ZN(n7945)
         );
  INV_X1 U9627 ( .A(n7943), .ZN(n7944) );
  AOI21_X1 U9628 ( .B1(n7946), .B2(n7945), .A(n7944), .ZN(n7957) );
  INV_X1 U9629 ( .A(n7947), .ZN(n7948) );
  NAND2_X1 U9630 ( .A1(n7948), .A2(n9400), .ZN(n7949) );
  NAND2_X1 U9631 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  NAND2_X1 U9632 ( .A1(n7951), .A2(n7964), .ZN(n7953) );
  AND2_X1 U9633 ( .A1(n7953), .A2(n7952), .ZN(n7968) );
  INV_X1 U9634 ( .A(n7968), .ZN(n7956) );
  INV_X1 U9635 ( .A(n7954), .ZN(n7955) );
  NOR2_X1 U9636 ( .A1(n7956), .A2(n7955), .ZN(n8031) );
  OAI21_X1 U9637 ( .B1(n7958), .B2(n7957), .A(n8031), .ZN(n7961) );
  INV_X1 U9638 ( .A(n7959), .ZN(n7960) );
  OAI21_X1 U9639 ( .B1(n7961), .B2(n7960), .A(n9355), .ZN(n7972) );
  NAND3_X1 U9640 ( .A1(n7964), .A2(n7963), .A3(n7962), .ZN(n7967) );
  INV_X1 U9641 ( .A(n7965), .ZN(n7966) );
  AOI21_X1 U9642 ( .B1(n7968), .B2(n7967), .A(n7966), .ZN(n7971) );
  INV_X1 U9643 ( .A(n7969), .ZN(n7970) );
  OAI21_X1 U9644 ( .B1(n7971), .B2(n8032), .A(n7970), .ZN(n8035) );
  AOI21_X1 U9645 ( .B1(n7973), .B2(n7972), .A(n8035), .ZN(n7979) );
  AND2_X1 U9646 ( .A1(n7975), .A2(n7974), .ZN(n8034) );
  INV_X1 U9647 ( .A(n8034), .ZN(n7978) );
  NAND2_X1 U9648 ( .A1(n9326), .A2(n7976), .ZN(n8021) );
  NAND2_X1 U9649 ( .A1(n8021), .A2(n7869), .ZN(n8029) );
  INV_X1 U9650 ( .A(n8029), .ZN(n7977) );
  OAI21_X1 U9651 ( .B1(n7979), .B2(n7978), .A(n7977), .ZN(n7980) );
  AOI21_X1 U9652 ( .B1(n7981), .B2(n7980), .A(n8042), .ZN(n7982) );
  MUX2_X1 U9653 ( .A(n7984), .B(n7983), .S(n7982), .Z(n7985) );
  INV_X1 U9654 ( .A(n7985), .ZN(n8048) );
  INV_X1 U9655 ( .A(n7986), .ZN(n7987) );
  OR2_X1 U9656 ( .A1(n5385), .A2(n7989), .ZN(n8027) );
  INV_X1 U9657 ( .A(n9420), .ZN(n9412) );
  NOR2_X1 U9658 ( .A1(n7991), .A2(n7990), .ZN(n7995) );
  NAND4_X1 U9659 ( .A1(n7995), .A2(n7994), .A3(n7993), .A4(n7992), .ZN(n7998)
         );
  NOR3_X1 U9660 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n8003) );
  INV_X1 U9661 ( .A(n7999), .ZN(n8001) );
  NAND4_X1 U9662 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(n8004)
         );
  NOR2_X1 U9663 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  NAND4_X1 U9664 ( .A1(n8008), .A2(n8007), .A3(n4612), .A4(n8006), .ZN(n8009)
         );
  NOR2_X1 U9665 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  NAND3_X1 U9666 ( .A1(n8013), .A2(n8012), .A3(n8011), .ZN(n8014) );
  NOR2_X1 U9667 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND4_X1 U9668 ( .A1(n9486), .A2(n4294), .A3(n4390), .A4(n8016), .ZN(n8017)
         );
  NOR2_X1 U9669 ( .A1(n9469), .A2(n8017), .ZN(n8018) );
  INV_X1 U9670 ( .A(n9449), .ZN(n9451) );
  NAND4_X1 U9671 ( .A1(n9412), .A2(n8018), .A3(n9436), .A4(n9451), .ZN(n8019)
         );
  NOR2_X1 U9672 ( .A1(n9385), .A2(n8019), .ZN(n8020) );
  AND4_X1 U9673 ( .A1(n9354), .A2(n9399), .A3(n8020), .A4(n9371), .ZN(n8022)
         );
  NAND4_X1 U9674 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n8025)
         );
  AOI21_X1 U9675 ( .B1(n8030), .B2(n9326), .A(n8029), .ZN(n8039) );
  NAND2_X1 U9676 ( .A1(n8031), .A2(n9471), .ZN(n8033) );
  AOI21_X1 U9677 ( .B1(n9355), .B2(n8033), .A(n8032), .ZN(n8036) );
  OAI21_X1 U9678 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8038) );
  AOI22_X1 U9679 ( .A1(n8039), .A2(n8038), .B1(n8037), .B2(n9329), .ZN(n8043)
         );
  OAI211_X1 U9680 ( .C1(n8043), .C2(n8042), .A(n8041), .B(n8040), .ZN(n8045)
         );
  AOI21_X1 U9681 ( .B1(n8045), .B2(n8044), .A(n9321), .ZN(n8047) );
  NOR3_X1 U9682 ( .A1(n8051), .A2(n8050), .A3(n8049), .ZN(n8053) );
  OAI21_X1 U9683 ( .B1(n8054), .B2(n5651), .A(P1_B_REG_SCAN_IN), .ZN(n8052) );
  INV_X1 U9684 ( .A(n8055), .ZN(n8062) );
  AOI22_X1 U9685 ( .A1(n9494), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8056), .B2(
        n9800), .ZN(n8057) );
  OAI21_X1 U9686 ( .B1(n8058), .B2(n9516), .A(n8057), .ZN(n8061) );
  NOR2_X1 U9687 ( .A1(n8059), .A2(n9494), .ZN(n8060) );
  AOI211_X1 U9688 ( .C1(n9512), .C2(n8062), .A(n8061), .B(n8060), .ZN(n8063)
         );
  OAI21_X1 U9689 ( .B1(n8064), .B2(n9520), .A(n8063), .ZN(P1_U3265) );
  OAI222_X1 U9690 ( .A1(n9640), .A2(n8066), .B1(n9681), .B2(P1_U3086), .C1(
        n8065), .C2(n8084), .ZN(P1_U3328) );
  OAI222_X1 U9691 ( .A1(n9640), .A2(n8069), .B1(n8068), .B2(P1_U3086), .C1(
        n8067), .C2(n8084), .ZN(P1_U3331) );
  OAI21_X1 U9692 ( .B1(n8070), .B2(n8072), .A(n8071), .ZN(n8073) );
  NAND2_X1 U9693 ( .A1(n8073), .A2(n9151), .ZN(n8077) );
  AOI22_X1 U9694 ( .A1(n9066), .A2(n8075), .B1(n8074), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8076) );
  OAI211_X1 U9695 ( .C1(n4369), .C2(n9157), .A(n8077), .B(n8076), .ZN(P1_U3222) );
  INV_X1 U9696 ( .A(n8078), .ZN(n9049) );
  OAI222_X1 U9697 ( .A1(n9640), .A2(n9049), .B1(n8080), .B2(P1_U3086), .C1(
        n8079), .C2(n8084), .ZN(P1_U3327) );
  INV_X1 U9698 ( .A(n8081), .ZN(n8086) );
  OAI222_X1 U9699 ( .A1(P2_U3151), .A2(n8083), .B1(n9048), .B2(n8086), .C1(
        n8082), .C2(n9042), .ZN(P2_U3266) );
  OAI222_X1 U9700 ( .A1(n9640), .A2(n8086), .B1(n8085), .B2(P1_U3086), .C1(
        n9991), .C2(n8084), .ZN(P1_U3326) );
  INV_X1 U9701 ( .A(n8087), .ZN(n8088) );
  XNOR2_X1 U9702 ( .A(n8870), .B(n8131), .ZN(n8090) );
  NAND2_X1 U9703 ( .A1(n8090), .A2(n8161), .ZN(n8091) );
  OAI21_X1 U9704 ( .B1(n8090), .B2(n8161), .A(n8091), .ZN(n8242) );
  INV_X1 U9705 ( .A(n8091), .ZN(n8155) );
  XNOR2_X1 U9706 ( .A(n8092), .B(n8131), .ZN(n8093) );
  XNOR2_X1 U9707 ( .A(n8093), .B(n8855), .ZN(n8154) );
  OAI21_X1 U9708 ( .B1(n8153), .B2(n8155), .A(n8154), .ZN(n8152) );
  XNOR2_X1 U9709 ( .A(n9023), .B(n8131), .ZN(n8096) );
  XNOR2_X1 U9710 ( .A(n8096), .B(n8095), .ZN(n8281) );
  XNOR2_X1 U9711 ( .A(n8098), .B(n8131), .ZN(n8099) );
  NAND2_X1 U9712 ( .A1(n8099), .A2(n8841), .ZN(n8205) );
  NAND2_X1 U9713 ( .A1(n8207), .A2(n8205), .ZN(n8101) );
  INV_X1 U9714 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U9715 ( .A1(n8100), .A2(n8856), .ZN(n8206) );
  XNOR2_X1 U9716 ( .A(n9018), .B(n8131), .ZN(n8102) );
  XNOR2_X1 U9717 ( .A(n8102), .B(n8831), .ZN(n8217) );
  NAND2_X1 U9718 ( .A1(n8102), .A2(n8831), .ZN(n8103) );
  XNOR2_X1 U9719 ( .A(n8833), .B(n8131), .ZN(n8104) );
  XNOR2_X1 U9720 ( .A(n8104), .B(n8517), .ZN(n8263) );
  INV_X1 U9721 ( .A(n8263), .ZN(n8106) );
  INV_X1 U9722 ( .A(n8104), .ZN(n8105) );
  XNOR2_X1 U9723 ( .A(n9007), .B(n8131), .ZN(n8109) );
  XNOR2_X1 U9724 ( .A(n8109), .B(n8933), .ZN(n8175) );
  NAND2_X1 U9725 ( .A1(n8174), .A2(n8108), .ZN(n8183) );
  NAND2_X1 U9726 ( .A1(n8109), .A2(n8933), .ZN(n8231) );
  XNOR2_X1 U9727 ( .A(n8931), .B(n8131), .ZN(n8113) );
  NAND2_X1 U9728 ( .A1(n8113), .A2(n8924), .ZN(n8112) );
  AND2_X1 U9729 ( .A1(n8231), .A2(n8112), .ZN(n8184) );
  XNOR2_X1 U9730 ( .A(n8792), .B(n8131), .ZN(n8111) );
  NAND2_X1 U9731 ( .A1(n8111), .A2(n8934), .ZN(n8110) );
  AND2_X1 U9732 ( .A1(n8184), .A2(n8110), .ZN(n8117) );
  INV_X1 U9733 ( .A(n8110), .ZN(n8116) );
  XOR2_X1 U9734 ( .A(n8934), .B(n8111), .Z(n8188) );
  INV_X1 U9735 ( .A(n8112), .ZN(n8114) );
  XNOR2_X1 U9736 ( .A(n8113), .B(n8177), .ZN(n8234) );
  OR2_X1 U9737 ( .A1(n8114), .A2(n8234), .ZN(n8185) );
  AND2_X1 U9738 ( .A1(n8188), .A2(n8185), .ZN(n8115) );
  XNOR2_X1 U9739 ( .A(n8921), .B(n8126), .ZN(n8118) );
  NAND2_X1 U9740 ( .A1(n8118), .A2(n8787), .ZN(n8251) );
  INV_X1 U9741 ( .A(n8118), .ZN(n8119) );
  NAND2_X1 U9742 ( .A1(n8119), .A2(n8925), .ZN(n8252) );
  NAND2_X1 U9743 ( .A1(n8166), .A2(n8916), .ZN(n8122) );
  NAND2_X1 U9744 ( .A1(n8122), .A2(n8167), .ZN(n8224) );
  XNOR2_X1 U9745 ( .A(n8123), .B(n8126), .ZN(n8124) );
  NOR2_X1 U9746 ( .A1(n8124), .A2(n8759), .ZN(n8195) );
  AOI21_X1 U9747 ( .B1(n8124), .B2(n8759), .A(n8195), .ZN(n8225) );
  XNOR2_X1 U9748 ( .A(n8978), .B(n8131), .ZN(n8125) );
  XNOR2_X1 U9749 ( .A(n8125), .B(n8516), .ZN(n8194) );
  XNOR2_X1 U9750 ( .A(n8732), .B(n8126), .ZN(n8127) );
  NAND2_X1 U9751 ( .A1(n8271), .A2(n8715), .ZN(n8270) );
  INV_X1 U9752 ( .A(n8127), .ZN(n8128) );
  NAND2_X1 U9753 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  XNOR2_X1 U9754 ( .A(n8968), .B(n8131), .ZN(n8133) );
  XNOR2_X1 U9755 ( .A(n8133), .B(n8902), .ZN(n8143) );
  INV_X1 U9756 ( .A(n8143), .ZN(n8132) );
  INV_X1 U9757 ( .A(n8133), .ZN(n8134) );
  INV_X1 U9758 ( .A(n8902), .ZN(n8515) );
  NAND2_X1 U9759 ( .A1(n8134), .A2(n8515), .ZN(n8135) );
  XOR2_X1 U9760 ( .A(n6679), .B(n8469), .Z(n8136) );
  XNOR2_X1 U9761 ( .A(n8137), .B(n8136), .ZN(n8142) );
  NOR2_X1 U9762 ( .A1(n9990), .A2(n8286), .ZN(n8140) );
  AOI22_X1 U9763 ( .A1(n8703), .A2(n8267), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8138) );
  OAI21_X1 U9764 ( .B1(n8902), .B2(n8257), .A(n8138), .ZN(n8139) );
  AOI211_X1 U9765 ( .C1(n6336), .C2(n8259), .A(n8140), .B(n8139), .ZN(n8141)
         );
  OAI21_X1 U9766 ( .B1(n8142), .B2(n8280), .A(n8141), .ZN(P2_U3160) );
  AOI21_X1 U9767 ( .B1(n8144), .B2(n8143), .A(n8280), .ZN(n8146) );
  NAND2_X1 U9768 ( .A1(n8146), .A2(n8145), .ZN(n8150) );
  AOI22_X1 U9769 ( .A1(n8721), .A2(n8267), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8147) );
  OAI21_X1 U9770 ( .B1(n8715), .B2(n8257), .A(n8147), .ZN(n8148) );
  AOI21_X1 U9771 ( .B1(n8514), .B2(n8277), .A(n8148), .ZN(n8149) );
  OAI211_X1 U9772 ( .C1(n8151), .C2(n8293), .A(n8150), .B(n8149), .ZN(P2_U3154) );
  INV_X1 U9773 ( .A(n8152), .ZN(n8157) );
  NOR3_X1 U9774 ( .A1(n8240), .A2(n8155), .A3(n8154), .ZN(n8156) );
  OAI21_X1 U9775 ( .B1(n8157), .B2(n8156), .A(n8272), .ZN(n8165) );
  INV_X1 U9776 ( .A(n8158), .ZN(n8163) );
  AOI21_X1 U9777 ( .B1(n8277), .B2(n8518), .A(n8159), .ZN(n8160) );
  OAI21_X1 U9778 ( .B1(n8161), .B2(n8257), .A(n8160), .ZN(n8162) );
  AOI21_X1 U9779 ( .B1(n8163), .B2(n8267), .A(n8162), .ZN(n8164) );
  OAI211_X1 U9780 ( .C1(n9031), .C2(n8293), .A(n8165), .B(n8164), .ZN(P2_U3155) );
  NAND2_X1 U9781 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  XNOR2_X1 U9782 ( .A(n8168), .B(n8916), .ZN(n8173) );
  AOI22_X1 U9783 ( .A1(n8759), .A2(n8277), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8170) );
  NAND2_X1 U9784 ( .A1(n8762), .A2(n8267), .ZN(n8169) );
  OAI211_X1 U9785 ( .C1(n8925), .C2(n8257), .A(n8170), .B(n8169), .ZN(n8171)
         );
  AOI21_X1 U9786 ( .B1(n8989), .B2(n8259), .A(n8171), .ZN(n8172) );
  OAI21_X1 U9787 ( .B1(n8173), .B2(n8280), .A(n8172), .ZN(P2_U3156) );
  XOR2_X1 U9788 ( .A(n8176), .B(n8175), .Z(n8182) );
  NAND2_X1 U9789 ( .A1(n8277), .A2(n8177), .ZN(n8178) );
  NAND2_X1 U9790 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8670) );
  OAI211_X1 U9791 ( .C1(n8842), .C2(n8257), .A(n8178), .B(n8670), .ZN(n8179)
         );
  AOI21_X1 U9792 ( .B1(n8816), .B2(n8267), .A(n8179), .ZN(n8181) );
  NAND2_X1 U9793 ( .A1(n9007), .A2(n8259), .ZN(n8180) );
  OAI211_X1 U9794 ( .C1(n8182), .C2(n8280), .A(n8181), .B(n8180), .ZN(P2_U3159) );
  NAND2_X1 U9795 ( .A1(n8232), .A2(n8184), .ZN(n8186) );
  AND2_X1 U9796 ( .A1(n8186), .A2(n8185), .ZN(n8187) );
  XOR2_X1 U9797 ( .A(n8188), .B(n8187), .Z(n8193) );
  AOI22_X1 U9798 ( .A1(n8787), .A2(n8277), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8190) );
  NAND2_X1 U9799 ( .A1(n8267), .A2(n8788), .ZN(n8189) );
  OAI211_X1 U9800 ( .C1(n8924), .C2(n8257), .A(n8190), .B(n8189), .ZN(n8191)
         );
  AOI21_X1 U9801 ( .B1(n8792), .B2(n8259), .A(n8191), .ZN(n8192) );
  OAI21_X1 U9802 ( .B1(n8193), .B2(n8280), .A(n8192), .ZN(P2_U3163) );
  INV_X1 U9803 ( .A(n8978), .ZN(n8741) );
  INV_X1 U9804 ( .A(n8223), .ZN(n8196) );
  NOR3_X1 U9805 ( .A1(n8196), .A2(n8195), .A3(n8194), .ZN(n8199) );
  INV_X1 U9806 ( .A(n8197), .ZN(n8198) );
  OAI21_X1 U9807 ( .B1(n8199), .B2(n8198), .A(n8272), .ZN(n8204) );
  INV_X1 U9808 ( .A(n8200), .ZN(n8740) );
  AOI22_X1 U9809 ( .A1(n8759), .A2(n8290), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8201) );
  OAI21_X1 U9810 ( .B1(n8740), .B2(n8287), .A(n8201), .ZN(n8202) );
  AOI21_X1 U9811 ( .B1(n8277), .B2(n8738), .A(n8202), .ZN(n8203) );
  OAI211_X1 U9812 ( .C1(n8741), .C2(n8293), .A(n8204), .B(n8203), .ZN(P2_U3165) );
  NAND2_X1 U9813 ( .A1(n8206), .A2(n8205), .ZN(n8208) );
  XOR2_X1 U9814 ( .A(n8208), .B(n8207), .Z(n8215) );
  NAND2_X1 U9815 ( .A1(n8290), .A2(n8518), .ZN(n8209) );
  NAND2_X1 U9816 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8588) );
  OAI211_X1 U9817 ( .C1(n8831), .C2(n8286), .A(n8209), .B(n8588), .ZN(n8212)
         );
  NOR2_X1 U9818 ( .A1(n8210), .A2(n8293), .ZN(n8211) );
  AOI211_X1 U9819 ( .C1(n8213), .C2(n8267), .A(n8212), .B(n8211), .ZN(n8214)
         );
  OAI21_X1 U9820 ( .B1(n8215), .B2(n8280), .A(n8214), .ZN(P2_U3166) );
  XOR2_X1 U9821 ( .A(n8216), .B(n8217), .Z(n8222) );
  NAND2_X1 U9822 ( .A1(n8290), .A2(n8856), .ZN(n8218) );
  NAND2_X1 U9823 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U9824 ( .C1(n8842), .C2(n8286), .A(n8218), .B(n8620), .ZN(n8220)
         );
  INV_X1 U9825 ( .A(n9018), .ZN(n8950) );
  NOR2_X1 U9826 ( .A1(n8950), .A2(n8293), .ZN(n8219) );
  AOI211_X1 U9827 ( .C1(n8847), .C2(n8267), .A(n8220), .B(n8219), .ZN(n8221)
         );
  OAI21_X1 U9828 ( .B1(n8222), .B2(n8280), .A(n8221), .ZN(P2_U3168) );
  OAI21_X1 U9829 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8226) );
  NAND2_X1 U9830 ( .A1(n8226), .A2(n8272), .ZN(n8230) );
  AOI22_X1 U9831 ( .A1(n8775), .A2(n8290), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8227) );
  OAI21_X1 U9832 ( .B1(n8901), .B2(n8286), .A(n8227), .ZN(n8228) );
  AOI21_X1 U9833 ( .B1(n8750), .B2(n8267), .A(n8228), .ZN(n8229) );
  OAI211_X1 U9834 ( .C1(n8983), .C2(n8293), .A(n8230), .B(n8229), .ZN(P2_U3169) );
  NAND2_X1 U9835 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  XOR2_X1 U9836 ( .A(n8234), .B(n8233), .Z(n8239) );
  INV_X1 U9837 ( .A(n8934), .ZN(n8798) );
  AOI22_X1 U9838 ( .A1(n8798), .A2(n8277), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8236) );
  NAND2_X1 U9839 ( .A1(n8267), .A2(n8799), .ZN(n8235) );
  OAI211_X1 U9840 ( .C1(n8933), .C2(n8257), .A(n8236), .B(n8235), .ZN(n8237)
         );
  AOI21_X1 U9841 ( .B1(n8931), .B2(n8259), .A(n8237), .ZN(n8238) );
  OAI21_X1 U9842 ( .B1(n8239), .B2(n8280), .A(n8238), .ZN(P2_U3173) );
  AOI21_X1 U9843 ( .B1(n8242), .B2(n8241), .A(n8240), .ZN(n8249) );
  OAI21_X1 U9844 ( .B1(n8257), .B2(n8244), .A(n8243), .ZN(n8245) );
  AOI21_X1 U9845 ( .B1(n8277), .B2(n8855), .A(n8245), .ZN(n8246) );
  OAI21_X1 U9846 ( .B1(n8866), .B2(n8287), .A(n8246), .ZN(n8247) );
  AOI21_X1 U9847 ( .B1(n8870), .B2(n8259), .A(n8247), .ZN(n8248) );
  OAI21_X1 U9848 ( .B1(n8249), .B2(n8280), .A(n8248), .ZN(P2_U3174) );
  NAND2_X1 U9849 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  XNOR2_X1 U9850 ( .A(n8254), .B(n8253), .ZN(n8261) );
  AOI22_X1 U9851 ( .A1(n8775), .A2(n8277), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8256) );
  NAND2_X1 U9852 ( .A1(n8267), .A2(n8771), .ZN(n8255) );
  OAI211_X1 U9853 ( .C1(n8934), .C2(n8257), .A(n8256), .B(n8255), .ZN(n8258)
         );
  AOI21_X1 U9854 ( .B1(n8921), .B2(n8259), .A(n8258), .ZN(n8260) );
  OAI21_X1 U9855 ( .B1(n8261), .B2(n8280), .A(n8260), .ZN(P2_U3175) );
  XOR2_X1 U9856 ( .A(n8262), .B(n8263), .Z(n8269) );
  NAND2_X1 U9857 ( .A1(n8290), .A2(n8943), .ZN(n8264) );
  NAND2_X1 U9858 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8650) );
  OAI211_X1 U9859 ( .C1(n8933), .C2(n8286), .A(n8264), .B(n8650), .ZN(n8266)
         );
  INV_X1 U9860 ( .A(n8833), .ZN(n8946) );
  NOR2_X1 U9861 ( .A1(n8946), .A2(n8293), .ZN(n8265) );
  AOI211_X1 U9862 ( .C1(n8827), .C2(n8267), .A(n8266), .B(n8265), .ZN(n8268)
         );
  OAI21_X1 U9863 ( .B1(n8269), .B2(n8280), .A(n8268), .ZN(P2_U3178) );
  OAI21_X1 U9864 ( .B1(n8715), .B2(n8271), .A(n8270), .ZN(n8273) );
  NAND2_X1 U9865 ( .A1(n8273), .A2(n8272), .ZN(n8279) );
  INV_X1 U9866 ( .A(n8728), .ZN(n8275) );
  AOI22_X1 U9867 ( .A1(n8516), .A2(n8290), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8274) );
  OAI21_X1 U9868 ( .B1(n8275), .B2(n8287), .A(n8274), .ZN(n8276) );
  AOI21_X1 U9869 ( .B1(n8515), .B2(n8277), .A(n8276), .ZN(n8278) );
  OAI211_X1 U9870 ( .C1(n8975), .C2(n8293), .A(n8279), .B(n8278), .ZN(P2_U3180) );
  INV_X1 U9871 ( .A(n9023), .ZN(n8294) );
  AOI21_X1 U9872 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8284) );
  NAND2_X1 U9873 ( .A1(n8284), .A2(n8283), .ZN(n8292) );
  NAND2_X1 U9874 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8560) );
  OAI21_X1 U9875 ( .B1(n8286), .B2(n8841), .A(n8560), .ZN(n8289) );
  NOR2_X1 U9876 ( .A1(n8287), .A2(n8858), .ZN(n8288) );
  AOI211_X1 U9877 ( .C1(n8290), .C2(n8855), .A(n8289), .B(n8288), .ZN(n8291)
         );
  OAI211_X1 U9878 ( .C1(n8294), .C2(n8293), .A(n8292), .B(n8291), .ZN(P2_U3181) );
  MUX2_X1 U9879 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9036), .S(n8295), .Z(n8297) );
  NAND2_X1 U9880 ( .A1(n8297), .A2(n8296), .ZN(n8691) );
  NAND2_X1 U9881 ( .A1(n9041), .A2(n8298), .ZN(n8301) );
  OR2_X1 U9882 ( .A1(n8299), .A2(n9043), .ZN(n8300) );
  NOR2_X1 U9883 ( .A1(n8961), .A2(n4696), .ZN(n8313) );
  INV_X1 U9884 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U9885 ( .A1(n5913), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8304) );
  INV_X1 U9886 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8302) );
  OR2_X1 U9887 ( .A1(n5897), .A2(n8302), .ZN(n8303) );
  OAI211_X1 U9888 ( .C1(n8306), .C2(n4275), .A(n8304), .B(n8303), .ZN(n8307)
         );
  INV_X1 U9889 ( .A(n8307), .ZN(n8308) );
  NAND2_X1 U9890 ( .A1(n8309), .A2(n8308), .ZN(n8688) );
  NAND2_X1 U9891 ( .A1(n8691), .A2(n8688), .ZN(n8467) );
  INV_X1 U9892 ( .A(n8513), .ZN(n8315) );
  INV_X1 U9893 ( .A(n8318), .ZN(n8457) );
  MUX2_X1 U9894 ( .A(n8320), .B(n8319), .S(n4495), .Z(n8452) );
  INV_X1 U9895 ( .A(n8710), .ZN(n8713) );
  INV_X1 U9896 ( .A(n8321), .ZN(n8472) );
  AND2_X1 U9897 ( .A1(n8327), .A2(n8322), .ZN(n8324) );
  MUX2_X1 U9898 ( .A(n8459), .B(n8326), .S(n6232), .Z(n8337) );
  NAND2_X1 U9899 ( .A1(n8879), .A2(n8327), .ZN(n8328) );
  OAI21_X1 U9900 ( .B1(n8329), .B2(n8328), .A(n8474), .ZN(n8336) );
  NAND2_X1 U9901 ( .A1(n6234), .A2(n8330), .ZN(n8333) );
  NAND2_X1 U9902 ( .A1(n8340), .A2(n8331), .ZN(n8332) );
  MUX2_X1 U9903 ( .A(n8333), .B(n8332), .S(n8459), .Z(n8334) );
  INV_X1 U9904 ( .A(n8334), .ZN(n8335) );
  OAI21_X1 U9905 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n8339) );
  INV_X1 U9906 ( .A(n8340), .ZN(n8342) );
  OAI211_X1 U9907 ( .C1(n8347), .C2(n8342), .A(n8348), .B(n6236), .ZN(n8344)
         );
  AND3_X1 U9908 ( .A1(n8344), .A2(n8343), .A3(n8350), .ZN(n8353) );
  INV_X1 U9909 ( .A(n6234), .ZN(n8346) );
  OAI21_X1 U9910 ( .B1(n8347), .B2(n8346), .A(n8345), .ZN(n8349) );
  NAND2_X1 U9911 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  MUX2_X1 U9912 ( .A(n8354), .B(n8359), .S(n4495), .Z(n8355) );
  OAI211_X1 U9913 ( .C1(n8459), .C2(n8357), .A(n4487), .B(n8482), .ZN(n8368)
         );
  AND2_X1 U9914 ( .A1(n8359), .A2(n8358), .ZN(n8363) );
  NAND2_X1 U9915 ( .A1(n9922), .A2(n8360), .ZN(n8361) );
  INV_X1 U9916 ( .A(n8375), .ZN(n8370) );
  NOR2_X1 U9917 ( .A1(n8371), .A2(n8370), .ZN(n8378) );
  INV_X1 U9918 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U9919 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  NAND2_X1 U9920 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  MUX2_X1 U9921 ( .A(n8378), .B(n8377), .S(n8459), .Z(n8379) );
  INV_X1 U9922 ( .A(n8379), .ZN(n8380) );
  NAND2_X1 U9923 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  NAND2_X1 U9924 ( .A1(n8383), .A2(n8382), .ZN(n8387) );
  MUX2_X1 U9925 ( .A(n8385), .B(n8384), .S(n4495), .Z(n8386) );
  NAND2_X1 U9926 ( .A1(n8387), .A2(n8386), .ZN(n8391) );
  INV_X1 U9927 ( .A(n8391), .ZN(n8394) );
  INV_X1 U9928 ( .A(n8388), .ZN(n8390) );
  MUX2_X1 U9929 ( .A(n8519), .B(n8870), .S(n4495), .Z(n8389) );
  OAI21_X1 U9930 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8392) );
  INV_X1 U9931 ( .A(n8395), .ZN(n8489) );
  MUX2_X1 U9932 ( .A(n8397), .B(n8396), .S(n8459), .Z(n8398) );
  AND2_X1 U9933 ( .A1(n8405), .A2(n8400), .ZN(n8401) );
  MUX2_X1 U9934 ( .A(n8402), .B(n8401), .S(n8459), .Z(n8403) );
  INV_X1 U9935 ( .A(n8839), .ZN(n8836) );
  NOR2_X1 U9936 ( .A1(n8408), .A2(n4744), .ZN(n8410) );
  INV_X1 U9937 ( .A(n8405), .ZN(n8407) );
  OAI211_X1 U9938 ( .C1(n8408), .C2(n8407), .A(n8414), .B(n8406), .ZN(n8409)
         );
  NAND3_X1 U9939 ( .A1(n8417), .A2(n8418), .A3(n8413), .ZN(n8411) );
  NAND3_X1 U9940 ( .A1(n8411), .A2(n8415), .A3(n8420), .ZN(n8419) );
  NAND2_X1 U9941 ( .A1(n8413), .A2(n8412), .ZN(n8416) );
  INV_X1 U9942 ( .A(n8782), .ZN(n8424) );
  AND2_X1 U9943 ( .A1(n8427), .A2(n8420), .ZN(n8421) );
  MUX2_X1 U9944 ( .A(n8422), .B(n8421), .S(n8459), .Z(n8423) );
  OAI21_X1 U9945 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8429) );
  MUX2_X1 U9946 ( .A(n8427), .B(n8426), .S(n8459), .Z(n8428) );
  AND2_X1 U9947 ( .A1(n8471), .A2(n8430), .ZN(n8431) );
  MUX2_X1 U9948 ( .A(n8432), .B(n8431), .S(n4495), .Z(n8433) );
  OAI21_X1 U9949 ( .B1(n8434), .B2(n4428), .A(n8435), .ZN(n8438) );
  NAND2_X1 U9950 ( .A1(n8435), .A2(n8472), .ZN(n8436) );
  NAND2_X1 U9951 ( .A1(n6250), .A2(n8436), .ZN(n8437) );
  MUX2_X1 U9952 ( .A(n8438), .B(n8437), .S(n4495), .Z(n8442) );
  INV_X1 U9953 ( .A(n8439), .ZN(n8441) );
  MUX2_X1 U9954 ( .A(n8443), .B(n4334), .S(n8459), .Z(n8445) );
  INV_X1 U9955 ( .A(n8448), .ZN(n8444) );
  INV_X1 U9956 ( .A(n8446), .ZN(n8447) );
  MUX2_X1 U9957 ( .A(n8448), .B(n8447), .S(n4495), .Z(n8449) );
  NAND3_X1 U9958 ( .A1(n8713), .A2(n8450), .A3(n8449), .ZN(n8451) );
  MUX2_X1 U9959 ( .A(n8716), .B(n8455), .S(n4495), .Z(n8454) );
  MUX2_X1 U9960 ( .A(n8716), .B(n8455), .S(n8459), .Z(n8456) );
  AOI21_X1 U9961 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8460) );
  OR2_X1 U9962 ( .A1(n8691), .A2(n8688), .ZN(n8461) );
  INV_X1 U9963 ( .A(n8461), .ZN(n8463) );
  NAND2_X1 U9964 ( .A1(n8466), .A2(n8465), .ZN(n8503) );
  INV_X1 U9965 ( .A(n8467), .ZN(n8501) );
  INV_X1 U9966 ( .A(n8468), .ZN(n8498) );
  INV_X1 U9967 ( .A(n8725), .ZN(n8497) );
  INV_X1 U9968 ( .A(n8767), .ZN(n8765) );
  NAND2_X1 U9969 ( .A1(n8472), .A2(n8471), .ZN(n8757) );
  INV_X1 U9970 ( .A(n8785), .ZN(n8494) );
  INV_X1 U9971 ( .A(n8797), .ZN(n8493) );
  NAND4_X1 U9972 ( .A1(n8475), .A2(n8879), .A3(n8474), .A4(n8473), .ZN(n8479)
         );
  NOR4_X1 U9973 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n8480)
         );
  NAND4_X1 U9974 ( .A1(n8483), .A2(n8482), .A3(n8481), .A4(n8480), .ZN(n8485)
         );
  NOR4_X1 U9975 ( .A1(n8486), .A2(n8485), .A3(n4402), .A4(n8484), .ZN(n8488)
         );
  NAND4_X1 U9976 ( .A1(n8853), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8490)
         );
  NOR4_X1 U9977 ( .A1(n8824), .A2(n8839), .A3(n8491), .A4(n8490), .ZN(n8492)
         );
  NAND4_X1 U9978 ( .A1(n8494), .A2(n8493), .A3(n8808), .A4(n8492), .ZN(n8495)
         );
  NOR4_X1 U9979 ( .A1(n8737), .A2(n8765), .A3(n8757), .A4(n8495), .ZN(n8496)
         );
  NAND4_X1 U9980 ( .A1(n8498), .A2(n6317), .A3(n8311), .A4(n4850), .ZN(n8500)
         );
  OAI21_X1 U9981 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8502) );
  NOR3_X1 U9982 ( .A1(n8507), .A2(n8506), .A3(n6257), .ZN(n8510) );
  OAI21_X1 U9983 ( .B1(n8511), .B2(n8508), .A(P2_B_REG_SCAN_IN), .ZN(n8509) );
  OAI22_X1 U9984 ( .A1(n8512), .A2(n8511), .B1(n8510), .B2(n8509), .ZN(
        P2_U3296) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8688), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8513), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8514), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8515), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9989 ( .A(n8738), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8641), .Z(
        P2_U3517) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8516), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8759), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9992 ( .A(n8775), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8641), .Z(
        P2_U3514) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8787), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9994 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8798), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8944), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8517), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8943), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8856), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8518), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8855), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10001 ( .A(n8519), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8641), .Z(
        P2_U3504) );
  MUX2_X1 U10002 ( .A(n8520), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8641), .Z(
        P2_U3503) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8521), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10004 ( .A(n8522), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8641), .Z(
        P2_U3501) );
  MUX2_X1 U10005 ( .A(n8523), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8641), .Z(
        P2_U3500) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8524), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10007 ( .A(n8525), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8641), .Z(
        P2_U3498) );
  MUX2_X1 U10008 ( .A(n8526), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8641), .Z(
        P2_U3497) );
  MUX2_X1 U10009 ( .A(n8527), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8641), .Z(
        P2_U3496) );
  MUX2_X1 U10010 ( .A(n9873), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8641), .Z(
        P2_U3495) );
  MUX2_X1 U10011 ( .A(n8528), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8641), .Z(
        P2_U3494) );
  MUX2_X1 U10012 ( .A(n5910), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8641), .Z(
        P2_U3493) );
  MUX2_X1 U10013 ( .A(n9863), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8641), .Z(
        P2_U3492) );
  MUX2_X1 U10014 ( .A(n6415), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8641), .Z(
        P2_U3491) );
  OAI21_X1 U10015 ( .B1(n8531), .B2(n8530), .A(n8529), .ZN(n8532) );
  NAND2_X1 U10016 ( .A1(n8532), .A2(n8683), .ZN(n8552) );
  INV_X1 U10017 ( .A(n8533), .ZN(n8545) );
  INV_X1 U10018 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8536) );
  INV_X1 U10019 ( .A(n8534), .ZN(n8535) );
  OAI21_X1 U10020 ( .B1(n8653), .B2(n8536), .A(n8535), .ZN(n8544) );
  INV_X1 U10021 ( .A(n8537), .ZN(n8539) );
  NAND3_X1 U10022 ( .A1(n8540), .A2(n8539), .A3(n8538), .ZN(n8541) );
  AOI21_X1 U10023 ( .B1(n8542), .B2(n8541), .A(n8685), .ZN(n8543) );
  AOI211_X1 U10024 ( .C1(n8587), .C2(n8545), .A(n8544), .B(n8543), .ZN(n8551)
         );
  OAI21_X1 U10025 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8549) );
  NAND2_X1 U10026 ( .A1(n8549), .A2(n8624), .ZN(n8550) );
  NAND3_X1 U10027 ( .A1(n8552), .A2(n8551), .A3(n8550), .ZN(P2_U3188) );
  XOR2_X1 U10028 ( .A(n8576), .B(n8582), .Z(n8555) );
  AOI21_X1 U10029 ( .B1(n8563), .B2(n8555), .A(n8578), .ZN(n8575) );
  OAI21_X1 U10030 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8559), .A(n8583), .ZN(
        n8573) );
  INV_X1 U10031 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10032 ( .A1(n8587), .A2(n8577), .ZN(n8561) );
  OAI211_X1 U10033 ( .C1(n8562), .C2(n8653), .A(n8561), .B(n8560), .ZN(n8572)
         );
  MUX2_X1 U10034 ( .A(n8563), .B(n10113), .S(n8665), .Z(n8564) );
  NAND2_X1 U10035 ( .A1(n8577), .A2(n8564), .ZN(n8591) );
  OR2_X1 U10036 ( .A1(n8577), .A2(n8564), .ZN(n8565) );
  NAND2_X1 U10037 ( .A1(n8591), .A2(n8565), .ZN(n8566) );
  AOI21_X1 U10038 ( .B1(n8568), .B2(n8567), .A(n8566), .ZN(n8598) );
  INV_X1 U10039 ( .A(n8598), .ZN(n8570) );
  NAND3_X1 U10040 ( .A1(n8568), .A2(n8567), .A3(n8566), .ZN(n8569) );
  AOI21_X1 U10041 ( .B1(n8570), .B2(n8569), .A(n8617), .ZN(n8571) );
  AOI211_X1 U10042 ( .C1(n8573), .C2(n8624), .A(n8572), .B(n8571), .ZN(n8574)
         );
  OAI21_X1 U10043 ( .B1(n8575), .B2(n8685), .A(n8574), .ZN(P2_U3197) );
  NOR2_X1 U10044 ( .A1(n8577), .A2(n8576), .ZN(n8579) );
  AOI22_X1 U10045 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8612), .B1(n8593), .B2(
        n8605), .ZN(n8580) );
  AOI21_X1 U10046 ( .B1(n4310), .B2(n8580), .A(n8606), .ZN(n8604) );
  AOI22_X1 U10047 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8593), .B1(n8612), .B2(
        n8611), .ZN(n8586) );
  NAND2_X1 U10048 ( .A1(n8582), .A2(n8581), .ZN(n8584) );
  NAND2_X1 U10049 ( .A1(n8584), .A2(n8583), .ZN(n8585) );
  NAND2_X1 U10050 ( .A1(n8586), .A2(n8585), .ZN(n8610) );
  OAI21_X1 U10051 ( .B1(n8586), .B2(n8585), .A(n8610), .ZN(n8602) );
  NAND2_X1 U10052 ( .A1(n8587), .A2(n8612), .ZN(n8589) );
  OAI211_X1 U10053 ( .C1(n8590), .C2(n8653), .A(n8589), .B(n8588), .ZN(n8601)
         );
  INV_X1 U10054 ( .A(n8591), .ZN(n8597) );
  MUX2_X1 U10055 ( .A(n8605), .B(n8611), .S(n8665), .Z(n8592) );
  NAND2_X1 U10056 ( .A1(n8592), .A2(n8612), .ZN(n8614) );
  INV_X1 U10057 ( .A(n8592), .ZN(n8594) );
  NAND2_X1 U10058 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  AND2_X1 U10059 ( .A1(n8614), .A2(n8595), .ZN(n8596) );
  OAI21_X1 U10060 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8616) );
  OR3_X1 U10061 ( .A1(n8598), .A2(n8597), .A3(n8596), .ZN(n8599) );
  AOI21_X1 U10062 ( .B1(n8616), .B2(n8599), .A(n8617), .ZN(n8600) );
  AOI211_X1 U10063 ( .C1(n8602), .C2(n8624), .A(n8601), .B(n8600), .ZN(n8603)
         );
  OAI21_X1 U10064 ( .B1(n8604), .B2(n8685), .A(n8603), .ZN(P2_U3198) );
  OAI21_X1 U10065 ( .B1(n8607), .B2(n8643), .A(n8631), .ZN(n8609) );
  INV_X1 U10066 ( .A(n8632), .ZN(n8608) );
  AOI21_X1 U10067 ( .B1(n10130), .B2(n8609), .A(n8608), .ZN(n8627) );
  OAI21_X1 U10068 ( .B1(n8612), .B2(n8611), .A(n8610), .ZN(n8642) );
  XNOR2_X1 U10069 ( .A(n8642), .B(n8637), .ZN(n8613) );
  OAI21_X1 U10070 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8613), .A(n8646), .ZN(
        n8625) );
  MUX2_X1 U10071 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8665), .Z(n8634) );
  XNOR2_X1 U10072 ( .A(n8634), .B(n8643), .ZN(n8615) );
  AOI21_X1 U10073 ( .B1(n8616), .B2(n8614), .A(n8615), .ZN(n8635) );
  INV_X1 U10074 ( .A(n8635), .ZN(n8619) );
  NAND3_X1 U10075 ( .A1(n8616), .A2(n8615), .A3(n8614), .ZN(n8618) );
  AOI21_X1 U10076 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(n8623) );
  NAND2_X1 U10077 ( .A1(n8669), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8621) );
  OAI211_X1 U10078 ( .C1(n8673), .C2(n8643), .A(n8621), .B(n8620), .ZN(n8622)
         );
  AOI211_X1 U10079 ( .C1(n8625), .C2(n8624), .A(n8623), .B(n8622), .ZN(n8626)
         );
  OAI21_X1 U10080 ( .B1(n8627), .B2(n8685), .A(n8626), .ZN(P2_U3199) );
  INV_X1 U10081 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8628) );
  OR2_X1 U10082 ( .A1(n8663), .A2(n8628), .ZN(n8659) );
  NAND2_X1 U10083 ( .A1(n8663), .A2(n8628), .ZN(n8629) );
  NAND2_X1 U10084 ( .A1(n8659), .A2(n8629), .ZN(n8630) );
  AND3_X1 U10085 ( .A1(n8632), .A2(n8631), .A3(n8630), .ZN(n8633) );
  NOR2_X1 U10086 ( .A1(n8633), .A2(n8661), .ZN(n8658) );
  INV_X1 U10087 ( .A(n8634), .ZN(n8636) );
  AOI21_X1 U10088 ( .B1(n8637), .B2(n8636), .A(n8635), .ZN(n8639) );
  MUX2_X1 U10089 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8665), .Z(n8638) );
  NOR2_X1 U10090 ( .A1(n8639), .A2(n8638), .ZN(n8664) );
  INV_X1 U10091 ( .A(n8664), .ZN(n8640) );
  NAND2_X1 U10092 ( .A1(n8639), .A2(n8638), .ZN(n8662) );
  NAND2_X1 U10093 ( .A1(n8640), .A2(n8662), .ZN(n8649) );
  OAI21_X1 U10094 ( .B1(n8649), .B2(n8641), .A(n8673), .ZN(n8656) );
  NAND2_X1 U10095 ( .A1(n8643), .A2(n8642), .ZN(n8645) );
  XNOR2_X1 U10096 ( .A(n8663), .B(n9997), .ZN(n8644) );
  AOI21_X1 U10097 ( .B1(n8646), .B2(n8645), .A(n8644), .ZN(n8674) );
  INV_X1 U10098 ( .A(n8674), .ZN(n8648) );
  NAND3_X1 U10099 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n8647) );
  AOI21_X1 U10100 ( .B1(n8648), .B2(n8647), .A(n8678), .ZN(n8655) );
  INV_X1 U10101 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8652) );
  NAND3_X1 U10102 ( .A1(n8649), .A2(n8683), .A3(n8675), .ZN(n8651) );
  OAI211_X1 U10103 ( .C1(n8653), .C2(n8652), .A(n8651), .B(n8650), .ZN(n8654)
         );
  AOI211_X1 U10104 ( .C1(n8663), .C2(n8656), .A(n8655), .B(n8654), .ZN(n8657)
         );
  OAI21_X1 U10105 ( .B1(n8658), .B2(n8685), .A(n8657), .ZN(P2_U3200) );
  INV_X1 U10106 ( .A(n8659), .ZN(n8660) );
  XNOR2_X1 U10107 ( .A(n4274), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8666) );
  OAI21_X1 U10108 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8668) );
  XNOR2_X1 U10109 ( .A(n4274), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8677) );
  MUX2_X1 U10110 ( .A(n8666), .B(n8677), .S(n8665), .Z(n8667) );
  XNOR2_X1 U10111 ( .A(n8668), .B(n8667), .ZN(n8682) );
  NAND2_X1 U10112 ( .A1(n8669), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8671) );
  OAI211_X1 U10113 ( .C1(n8673), .C2(n4274), .A(n8671), .B(n8670), .ZN(n8681)
         );
  AOI21_X1 U10114 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8675), .A(n8674), .ZN(
        n8676) );
  XOR2_X1 U10115 ( .A(n8677), .B(n8676), .Z(n8679) );
  NOR2_X1 U10116 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  OAI21_X1 U10117 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(P2_U3201) );
  NOR2_X1 U10118 ( .A1(n8689), .A2(n8882), .ZN(n8697) );
  AOI21_X1 U10119 ( .B1(n8962), .B2(n8859), .A(n8697), .ZN(n8693) );
  NAND2_X1 U10120 ( .A1(n8890), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U10121 ( .C1(n8691), .C2(n8885), .A(n8693), .B(n8690), .ZN(
        P2_U3202) );
  NAND2_X1 U10122 ( .A1(n8890), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8692) );
  OAI211_X1 U10123 ( .C1(n4696), .C2(n8885), .A(n8693), .B(n8692), .ZN(
        P2_U3203) );
  NAND2_X1 U10124 ( .A1(n8694), .A2(n8859), .ZN(n8699) );
  NOR2_X1 U10125 ( .A1(n8695), .A2(n8885), .ZN(n8696) );
  AOI211_X1 U10126 ( .C1(n8890), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8697), .B(
        n8696), .ZN(n8698) );
  OAI211_X1 U10127 ( .C1(n8701), .C2(n8700), .A(n8699), .B(n8698), .ZN(
        P2_U3204) );
  NAND2_X1 U10128 ( .A1(n8702), .A2(n8826), .ZN(n8708) );
  NOR2_X1 U10129 ( .A1(n9990), .A2(n8727), .ZN(n8706) );
  AOI22_X1 U10130 ( .A1(n8703), .A2(n8848), .B1(n8890), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8704) );
  OAI21_X1 U10131 ( .B1(n8902), .B2(n8830), .A(n8704), .ZN(n8705) );
  AOI211_X1 U10132 ( .C1(n6336), .C2(n8861), .A(n8706), .B(n8705), .ZN(n8707)
         );
  OAI211_X1 U10133 ( .C1(n8709), .C2(n8864), .A(n8708), .B(n8707), .ZN(
        P2_U3205) );
  XOR2_X1 U10134 ( .A(n8711), .B(n8710), .Z(n8971) );
  INV_X1 U10135 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8720) );
  INV_X1 U10136 ( .A(n8712), .ZN(n8714) );
  AOI21_X1 U10137 ( .B1(n8714), .B2(n8713), .A(n8917), .ZN(n8719) );
  OAI22_X1 U10138 ( .A1(n8716), .A2(n9919), .B1(n8715), .B2(n9917), .ZN(n8717)
         );
  AOI21_X1 U10139 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8966) );
  MUX2_X1 U10140 ( .A(n8720), .B(n8966), .S(n8859), .Z(n8723) );
  AOI22_X1 U10141 ( .A1(n8968), .A2(n8861), .B1(n8848), .B2(n8721), .ZN(n8722)
         );
  OAI211_X1 U10142 ( .C1(n8971), .C2(n8864), .A(n8723), .B(n8722), .ZN(
        P2_U3206) );
  XNOR2_X1 U10143 ( .A(n8724), .B(n8725), .ZN(n8900) );
  XNOR2_X1 U10144 ( .A(n8726), .B(n8725), .ZN(n8905) );
  NAND2_X1 U10145 ( .A1(n8905), .A2(n8826), .ZN(n8734) );
  NOR2_X1 U10146 ( .A1(n8902), .A2(n8727), .ZN(n8731) );
  AOI22_X1 U10147 ( .A1(n8728), .A2(n8848), .B1(n8890), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8729) );
  OAI21_X1 U10148 ( .B1(n8901), .B2(n8830), .A(n8729), .ZN(n8730) );
  AOI211_X1 U10149 ( .C1(n8732), .C2(n8861), .A(n8731), .B(n8730), .ZN(n8733)
         );
  OAI211_X1 U10150 ( .C1(n8864), .C2(n8900), .A(n8734), .B(n8733), .ZN(
        P2_U3207) );
  XOR2_X1 U10151 ( .A(n8737), .B(n8735), .Z(n8981) );
  XOR2_X1 U10152 ( .A(n8737), .B(n8736), .Z(n8739) );
  AOI222_X1 U10153 ( .A1(n9902), .A2(n8739), .B1(n8738), .B2(n9872), .C1(n8759), .C2(n9874), .ZN(n8976) );
  INV_X1 U10154 ( .A(n8976), .ZN(n8743) );
  OAI22_X1 U10155 ( .A1(n8741), .A2(n8752), .B1(n8740), .B2(n8882), .ZN(n8742)
         );
  OAI21_X1 U10156 ( .B1(n8743), .B2(n8742), .A(n8859), .ZN(n8745) );
  NAND2_X1 U10157 ( .A1(n8890), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8744) );
  OAI211_X1 U10158 ( .C1(n8981), .C2(n8864), .A(n8745), .B(n8744), .ZN(
        P2_U3208) );
  XOR2_X1 U10159 ( .A(n8746), .B(n8747), .Z(n8984) );
  XOR2_X1 U10160 ( .A(n8748), .B(n8747), .Z(n8749) );
  OAI222_X1 U10161 ( .A1(n9919), .A2(n8901), .B1(n9917), .B2(n8916), .C1(n8749), .C2(n8917), .ZN(n8982) );
  INV_X1 U10162 ( .A(n8750), .ZN(n8751) );
  OAI22_X1 U10163 ( .A1(n8983), .A2(n8752), .B1(n8751), .B2(n8882), .ZN(n8753)
         );
  OAI21_X1 U10164 ( .B1(n8982), .B2(n8753), .A(n8859), .ZN(n8755) );
  NAND2_X1 U10165 ( .A1(n8890), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8754) );
  OAI211_X1 U10166 ( .C1(n8984), .C2(n8864), .A(n8755), .B(n8754), .ZN(
        P2_U3209) );
  XOR2_X1 U10167 ( .A(n8757), .B(n8756), .Z(n8992) );
  XNOR2_X1 U10168 ( .A(n8758), .B(n8757), .ZN(n8760) );
  AOI222_X1 U10169 ( .A1(n9902), .A2(n8760), .B1(n8759), .B2(n9872), .C1(n8787), .C2(n9874), .ZN(n8987) );
  MUX2_X1 U10170 ( .A(n8761), .B(n8987), .S(n8859), .Z(n8764) );
  AOI22_X1 U10171 ( .A1(n8989), .A2(n8861), .B1(n8848), .B2(n8762), .ZN(n8763)
         );
  OAI211_X1 U10172 ( .C1(n8992), .C2(n8864), .A(n8764), .B(n8763), .ZN(
        P2_U3210) );
  XNOR2_X1 U10173 ( .A(n8766), .B(n8765), .ZN(n8918) );
  INV_X1 U10174 ( .A(n8826), .ZN(n8781) );
  OR2_X1 U10175 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  NAND2_X1 U10176 ( .A1(n8770), .A2(n8769), .ZN(n8996) );
  INV_X1 U10177 ( .A(n8996), .ZN(n8779) );
  NAND2_X1 U10178 ( .A1(n8921), .A2(n8861), .ZN(n8777) );
  NAND2_X1 U10179 ( .A1(n8848), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U10180 ( .A1(n8890), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10181 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  AOI21_X1 U10182 ( .B1(n8775), .B2(n8887), .A(n8774), .ZN(n8776) );
  OAI211_X1 U10183 ( .C1(n8934), .C2(n8830), .A(n8777), .B(n8776), .ZN(n8778)
         );
  AOI21_X1 U10184 ( .B1(n8779), .B2(n8872), .A(n8778), .ZN(n8780) );
  OAI21_X1 U10185 ( .B1(n8918), .B2(n8781), .A(n8780), .ZN(P2_U3211) );
  NAND2_X1 U10186 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  XNOR2_X1 U10187 ( .A(n8784), .B(n8785), .ZN(n8923) );
  XNOR2_X1 U10188 ( .A(n8786), .B(n8785), .ZN(n8928) );
  NAND2_X1 U10189 ( .A1(n8928), .A2(n8826), .ZN(n8794) );
  NAND2_X1 U10190 ( .A1(n8787), .A2(n8887), .ZN(n8790) );
  AOI22_X1 U10191 ( .A1(n8890), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8848), .B2(
        n8788), .ZN(n8789) );
  OAI211_X1 U10192 ( .C1(n8924), .C2(n8830), .A(n8790), .B(n8789), .ZN(n8791)
         );
  AOI21_X1 U10193 ( .B1(n8792), .B2(n8861), .A(n8791), .ZN(n8793) );
  OAI211_X1 U10194 ( .C1(n8923), .C2(n8864), .A(n8794), .B(n8793), .ZN(
        P2_U3212) );
  XNOR2_X1 U10195 ( .A(n8795), .B(n8797), .ZN(n8932) );
  OAI21_X1 U10196 ( .B1(n4340), .B2(n8797), .A(n8796), .ZN(n8937) );
  NAND2_X1 U10197 ( .A1(n8937), .A2(n8826), .ZN(n8804) );
  NAND2_X1 U10198 ( .A1(n8798), .A2(n8887), .ZN(n8801) );
  AOI22_X1 U10199 ( .A1(n8890), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8848), .B2(
        n8799), .ZN(n8800) );
  OAI211_X1 U10200 ( .C1(n8933), .C2(n8830), .A(n8801), .B(n8800), .ZN(n8802)
         );
  AOI21_X1 U10201 ( .B1(n8931), .B2(n8861), .A(n8802), .ZN(n8803) );
  OAI211_X1 U10202 ( .C1(n8932), .C2(n8864), .A(n8804), .B(n8803), .ZN(
        P2_U3213) );
  INV_X1 U10203 ( .A(n8808), .ZN(n8805) );
  XNOR2_X1 U10204 ( .A(n8806), .B(n8805), .ZN(n9008) );
  INV_X1 U10205 ( .A(n9008), .ZN(n8819) );
  NAND2_X1 U10206 ( .A1(n8807), .A2(n8808), .ZN(n8809) );
  NAND2_X1 U10207 ( .A1(n8809), .A2(n9902), .ZN(n8810) );
  OR2_X1 U10208 ( .A1(n8811), .A2(n8810), .ZN(n8814) );
  OAI22_X1 U10209 ( .A1(n8924), .A2(n9919), .B1(n8842), .B2(n9917), .ZN(n8812)
         );
  INV_X1 U10210 ( .A(n8812), .ZN(n8813) );
  NAND2_X1 U10211 ( .A1(n8814), .A2(n8813), .ZN(n9005) );
  MUX2_X1 U10212 ( .A(n9005), .B(P2_REG2_REG_19__SCAN_IN), .S(n8890), .Z(n8815) );
  INV_X1 U10213 ( .A(n8815), .ZN(n8818) );
  AOI22_X1 U10214 ( .A1(n9007), .A2(n8861), .B1(n8848), .B2(n8816), .ZN(n8817)
         );
  OAI211_X1 U10215 ( .C1(n8819), .C2(n8864), .A(n8818), .B(n8817), .ZN(
        P2_U3214) );
  NAND2_X1 U10216 ( .A1(n8820), .A2(n8824), .ZN(n8821) );
  NAND2_X1 U10217 ( .A1(n8822), .A2(n8821), .ZN(n9014) );
  OAI21_X1 U10218 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8948) );
  NAND2_X1 U10219 ( .A1(n8948), .A2(n8826), .ZN(n8835) );
  AOI22_X1 U10220 ( .A1(n8890), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8848), .B2(
        n8827), .ZN(n8829) );
  NAND2_X1 U10221 ( .A1(n8887), .A2(n8944), .ZN(n8828) );
  OAI211_X1 U10222 ( .C1(n8831), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8832)
         );
  AOI21_X1 U10223 ( .B1(n8833), .B2(n8861), .A(n8832), .ZN(n8834) );
  OAI211_X1 U10224 ( .C1(n9014), .C2(n8864), .A(n8835), .B(n8834), .ZN(
        P2_U3215) );
  XNOR2_X1 U10225 ( .A(n8837), .B(n8836), .ZN(n9021) );
  OAI211_X1 U10226 ( .C1(n8840), .C2(n8839), .A(n8838), .B(n9902), .ZN(n8845)
         );
  OAI22_X1 U10227 ( .A1(n8842), .A2(n9919), .B1(n8841), .B2(n9917), .ZN(n8843)
         );
  INV_X1 U10228 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U10229 ( .A1(n8845), .A2(n8844), .ZN(n9015) );
  MUX2_X1 U10230 ( .A(n9015), .B(P2_REG2_REG_17__SCAN_IN), .S(n8890), .Z(n8846) );
  INV_X1 U10231 ( .A(n8846), .ZN(n8850) );
  AOI22_X1 U10232 ( .A1(n9018), .A2(n8861), .B1(n8848), .B2(n8847), .ZN(n8849)
         );
  OAI211_X1 U10233 ( .C1(n9021), .C2(n8864), .A(n8850), .B(n8849), .ZN(
        P2_U3216) );
  XOR2_X1 U10234 ( .A(n8853), .B(n8851), .Z(n9026) );
  INV_X1 U10235 ( .A(n9026), .ZN(n8865) );
  OAI21_X1 U10236 ( .B1(n8852), .B2(n6085), .A(n8854), .ZN(n8857) );
  AOI222_X1 U10237 ( .A1(n9902), .A2(n8857), .B1(n8856), .B2(n9872), .C1(n8855), .C2(n9874), .ZN(n9022) );
  OAI21_X1 U10238 ( .B1(n8858), .B2(n8882), .A(n9022), .ZN(n8860) );
  NAND2_X1 U10239 ( .A1(n8860), .A2(n8859), .ZN(n8863) );
  AOI22_X1 U10240 ( .A1(n9023), .A2(n8861), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n8890), .ZN(n8862) );
  OAI211_X1 U10241 ( .C1(n8865), .C2(n8864), .A(n8863), .B(n8862), .ZN(
        P2_U3218) );
  NOR2_X1 U10242 ( .A1(n8882), .A2(n8866), .ZN(n8869) );
  INV_X1 U10243 ( .A(n8867), .ZN(n8868) );
  AOI211_X1 U10244 ( .C1(n8871), .C2(n8870), .A(n8869), .B(n8868), .ZN(n8875)
         );
  AOI22_X1 U10245 ( .A1(n8873), .A2(n8872), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8890), .ZN(n8874) );
  OAI21_X1 U10246 ( .B1(n8875), .B2(n8890), .A(n8874), .ZN(P2_U3220) );
  INV_X1 U10247 ( .A(n8876), .ZN(n8881) );
  OAI21_X1 U10248 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n9861) );
  AOI22_X1 U10249 ( .A1(n8881), .A2(n9861), .B1(n8880), .B2(n6415), .ZN(n8893)
         );
  OAI22_X1 U10250 ( .A1(n8885), .A2(n8884), .B1(n8883), .B2(n8882), .ZN(n8886)
         );
  AOI21_X1 U10251 ( .B1(n8887), .B2(n5910), .A(n8886), .ZN(n8892) );
  XNOR2_X1 U10252 ( .A(n8888), .B(n6231), .ZN(n8889) );
  NAND2_X1 U10253 ( .A1(n8889), .A2(n9902), .ZN(n9855) );
  MUX2_X1 U10254 ( .A(n9855), .B(n10102), .S(n8890), .Z(n8891) );
  NAND3_X1 U10255 ( .A1(n8893), .A2(n8892), .A3(n8891), .ZN(P2_U3232) );
  NAND2_X1 U10256 ( .A1(n8961), .A2(n8953), .ZN(n8894) );
  NAND2_X1 U10257 ( .A1(n8962), .A2(n9956), .ZN(n8896) );
  OAI211_X1 U10258 ( .C1(n9956), .C2(n8306), .A(n8894), .B(n8896), .ZN(
        P2_U3490) );
  NAND2_X1 U10259 ( .A1(n8895), .A2(n8953), .ZN(n8897) );
  OAI211_X1 U10260 ( .C1(n9956), .C2(n6262), .A(n8897), .B(n8896), .ZN(
        P2_U3489) );
  MUX2_X1 U10261 ( .A(n10058), .B(n8966), .S(n9956), .Z(n8899) );
  NAND2_X1 U10262 ( .A1(n8968), .A2(n8953), .ZN(n8898) );
  OAI211_X1 U10263 ( .C1(n8971), .C2(n8958), .A(n8899), .B(n8898), .ZN(
        P2_U3486) );
  NOR2_X1 U10264 ( .A1(n8900), .A2(n9935), .ZN(n8904) );
  OAI22_X1 U10265 ( .A1(n8902), .A2(n9919), .B1(n8901), .B2(n9917), .ZN(n8903)
         );
  AOI211_X1 U10266 ( .C1(n8905), .C2(n9902), .A(n8904), .B(n8903), .ZN(n8972)
         );
  MUX2_X1 U10267 ( .A(n8906), .B(n8972), .S(n9956), .Z(n8907) );
  OAI21_X1 U10268 ( .B1(n8975), .B2(n8957), .A(n8907), .ZN(P2_U3485) );
  MUX2_X1 U10269 ( .A(n8908), .B(n8976), .S(n9956), .Z(n8910) );
  NAND2_X1 U10270 ( .A1(n8978), .A2(n8953), .ZN(n8909) );
  OAI211_X1 U10271 ( .C1(n8958), .C2(n8981), .A(n8910), .B(n8909), .ZN(
        P2_U3484) );
  MUX2_X1 U10272 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8982), .S(n9956), .Z(n8912) );
  OAI22_X1 U10273 ( .A1(n8984), .A2(n8958), .B1(n8983), .B2(n8957), .ZN(n8911)
         );
  OR2_X1 U10274 ( .A1(n8912), .A2(n8911), .ZN(P2_U3483) );
  INV_X1 U10275 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8913) );
  MUX2_X1 U10276 ( .A(n8913), .B(n8987), .S(n9956), .Z(n8915) );
  NAND2_X1 U10277 ( .A1(n8989), .A2(n8953), .ZN(n8914) );
  OAI211_X1 U10278 ( .C1(n8992), .C2(n8958), .A(n8915), .B(n8914), .ZN(
        P2_U3482) );
  OAI22_X1 U10279 ( .A1(n8916), .A2(n9919), .B1(n8934), .B2(n9917), .ZN(n8920)
         );
  NOR2_X1 U10280 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  AOI211_X1 U10281 ( .C1(n9940), .C2(n8921), .A(n8920), .B(n8919), .ZN(n8993)
         );
  MUX2_X1 U10282 ( .A(n10104), .B(n8993), .S(n9956), .Z(n8922) );
  OAI21_X1 U10283 ( .B1(n8958), .B2(n8996), .A(n8922), .ZN(P2_U3481) );
  NOR2_X1 U10284 ( .A1(n8923), .A2(n9935), .ZN(n8927) );
  OAI22_X1 U10285 ( .A1(n8925), .A2(n9919), .B1(n8924), .B2(n9917), .ZN(n8926)
         );
  AOI211_X1 U10286 ( .C1(n8928), .C2(n9902), .A(n8927), .B(n8926), .ZN(n8997)
         );
  MUX2_X1 U10287 ( .A(n8929), .B(n8997), .S(n9956), .Z(n8930) );
  OAI21_X1 U10288 ( .B1(n9000), .B2(n8957), .A(n8930), .ZN(P2_U3480) );
  INV_X1 U10289 ( .A(n8931), .ZN(n9004) );
  INV_X1 U10290 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8938) );
  NOR2_X1 U10291 ( .A1(n8932), .A2(n9935), .ZN(n8936) );
  OAI22_X1 U10292 ( .A1(n8934), .A2(n9919), .B1(n8933), .B2(n9917), .ZN(n8935)
         );
  AOI211_X1 U10293 ( .C1(n8937), .C2(n9902), .A(n8936), .B(n8935), .ZN(n9001)
         );
  MUX2_X1 U10294 ( .A(n8938), .B(n9001), .S(n9956), .Z(n8939) );
  OAI21_X1 U10295 ( .B1(n9004), .B2(n8957), .A(n8939), .ZN(P2_U3479) );
  MUX2_X1 U10296 ( .A(n9005), .B(P2_REG1_REG_19__SCAN_IN), .S(n4414), .Z(n8940) );
  INV_X1 U10297 ( .A(n8940), .ZN(n8942) );
  AOI22_X1 U10298 ( .A1(n9008), .A2(n8954), .B1(n8953), .B2(n9007), .ZN(n8941)
         );
  NAND2_X1 U10299 ( .A1(n8942), .A2(n8941), .ZN(P2_U3478) );
  AOI22_X1 U10300 ( .A1(n8944), .A2(n9872), .B1(n9874), .B2(n8943), .ZN(n8945)
         );
  OAI21_X1 U10301 ( .B1(n8946), .B2(n9886), .A(n8945), .ZN(n8947) );
  AOI21_X1 U10302 ( .B1(n8948), .B2(n9902), .A(n8947), .ZN(n9011) );
  MUX2_X1 U10303 ( .A(n9997), .B(n9011), .S(n9956), .Z(n8949) );
  OAI21_X1 U10304 ( .B1(n8958), .B2(n9014), .A(n8949), .ZN(P2_U3477) );
  MUX2_X1 U10305 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9015), .S(n9956), .Z(n8952) );
  OAI22_X1 U10306 ( .A1(n9021), .A2(n8958), .B1(n8950), .B2(n8957), .ZN(n8951)
         );
  OR2_X1 U10307 ( .A1(n8952), .A2(n8951), .ZN(P2_U3476) );
  MUX2_X1 U10308 ( .A(n10113), .B(n9022), .S(n9956), .Z(n8956) );
  AOI22_X1 U10309 ( .A1(n9026), .A2(n8954), .B1(n8953), .B2(n9023), .ZN(n8955)
         );
  NAND2_X1 U10310 ( .A1(n8956), .A2(n8955), .ZN(P2_U3474) );
  MUX2_X1 U10311 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9029), .S(n9956), .Z(n8960) );
  OAI22_X1 U10312 ( .A1(n9033), .A2(n8958), .B1(n9031), .B2(n8957), .ZN(n8959)
         );
  OR2_X1 U10313 ( .A1(n8960), .A2(n8959), .ZN(P2_U3473) );
  NAND2_X1 U10314 ( .A1(n8961), .A2(n9024), .ZN(n8963) );
  NAND2_X1 U10315 ( .A1(n8962), .A2(n9941), .ZN(n8964) );
  OAI211_X1 U10316 ( .C1(n8302), .C2(n9941), .A(n8963), .B(n8964), .ZN(
        P2_U3458) );
  NAND2_X1 U10317 ( .A1(n9943), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8965) );
  OAI211_X1 U10318 ( .C1(n4696), .C2(n9030), .A(n8965), .B(n8964), .ZN(
        P2_U3457) );
  INV_X1 U10319 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8967) );
  MUX2_X1 U10320 ( .A(n8967), .B(n8966), .S(n9941), .Z(n8970) );
  NAND2_X1 U10321 ( .A1(n8968), .A2(n9024), .ZN(n8969) );
  OAI211_X1 U10322 ( .C1(n8971), .C2(n9032), .A(n8970), .B(n8969), .ZN(
        P2_U3454) );
  INV_X1 U10323 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U10324 ( .A(n8973), .B(n8972), .S(n9941), .Z(n8974) );
  OAI21_X1 U10325 ( .B1(n8975), .B2(n9030), .A(n8974), .ZN(P2_U3453) );
  INV_X1 U10326 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8977) );
  MUX2_X1 U10327 ( .A(n8977), .B(n8976), .S(n9941), .Z(n8980) );
  NAND2_X1 U10328 ( .A1(n8978), .A2(n9024), .ZN(n8979) );
  OAI211_X1 U10329 ( .C1(n8981), .C2(n9032), .A(n8980), .B(n8979), .ZN(
        P2_U3452) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8982), .S(n9941), .Z(n8986) );
  OAI22_X1 U10331 ( .A1(n8984), .A2(n9032), .B1(n8983), .B2(n9030), .ZN(n8985)
         );
  OR2_X1 U10332 ( .A1(n8986), .A2(n8985), .ZN(P2_U3451) );
  INV_X1 U10333 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U10334 ( .A(n8988), .B(n8987), .S(n9941), .Z(n8991) );
  NAND2_X1 U10335 ( .A1(n8989), .A2(n9024), .ZN(n8990) );
  OAI211_X1 U10336 ( .C1(n8992), .C2(n9032), .A(n8991), .B(n8990), .ZN(
        P2_U3450) );
  INV_X1 U10337 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8994) );
  MUX2_X1 U10338 ( .A(n8994), .B(n8993), .S(n9941), .Z(n8995) );
  OAI21_X1 U10339 ( .B1(n8996), .B2(n9032), .A(n8995), .ZN(P2_U3449) );
  INV_X1 U10340 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8998) );
  MUX2_X1 U10341 ( .A(n8998), .B(n8997), .S(n9941), .Z(n8999) );
  OAI21_X1 U10342 ( .B1(n9000), .B2(n9030), .A(n8999), .ZN(P2_U3448) );
  INV_X1 U10343 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9002) );
  MUX2_X1 U10344 ( .A(n9002), .B(n9001), .S(n9941), .Z(n9003) );
  OAI21_X1 U10345 ( .B1(n9004), .B2(n9030), .A(n9003), .ZN(P2_U3447) );
  MUX2_X1 U10346 ( .A(n9005), .B(P2_REG0_REG_19__SCAN_IN), .S(n9943), .Z(n9006) );
  INV_X1 U10347 ( .A(n9006), .ZN(n9010) );
  AOI22_X1 U10348 ( .A1(n9008), .A2(n9025), .B1(n9024), .B2(n9007), .ZN(n9009)
         );
  NAND2_X1 U10349 ( .A1(n9010), .A2(n9009), .ZN(P2_U3446) );
  INV_X1 U10350 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9012) );
  MUX2_X1 U10351 ( .A(n9012), .B(n9011), .S(n9941), .Z(n9013) );
  OAI21_X1 U10352 ( .B1(n9014), .B2(n9032), .A(n9013), .ZN(P2_U3444) );
  INV_X1 U10353 ( .A(n9015), .ZN(n9017) );
  MUX2_X1 U10354 ( .A(n9017), .B(n9016), .S(n9943), .Z(n9020) );
  NAND2_X1 U10355 ( .A1(n9018), .A2(n9024), .ZN(n9019) );
  OAI211_X1 U10356 ( .C1(n9021), .C2(n9032), .A(n9020), .B(n9019), .ZN(
        P2_U3441) );
  MUX2_X1 U10357 ( .A(n10119), .B(n9022), .S(n9941), .Z(n9028) );
  AOI22_X1 U10358 ( .A1(n9026), .A2(n9025), .B1(n9024), .B2(n9023), .ZN(n9027)
         );
  NAND2_X1 U10359 ( .A1(n9028), .A2(n9027), .ZN(P2_U3435) );
  MUX2_X1 U10360 ( .A(n9029), .B(P2_REG0_REG_14__SCAN_IN), .S(n9943), .Z(n9035) );
  OAI22_X1 U10361 ( .A1(n9033), .A2(n9032), .B1(n9031), .B2(n9030), .ZN(n9034)
         );
  OR2_X1 U10362 ( .A1(n9035), .A2(n9034), .ZN(P2_U3432) );
  INV_X1 U10363 ( .A(n9036), .ZN(n9637) );
  NOR4_X1 U10364 ( .A1(n9037), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5849), .ZN(n9038) );
  AOI21_X1 U10365 ( .B1(n9046), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9038), .ZN(
        n9039) );
  OAI21_X1 U10366 ( .B1(n9637), .B2(n9048), .A(n9039), .ZN(P2_U3264) );
  INV_X1 U10367 ( .A(n9041), .ZN(n9641) );
  OAI222_X1 U10368 ( .A1(n9040), .A2(P2_U3151), .B1(n9044), .B2(n9641), .C1(
        n9043), .C2(n9042), .ZN(P2_U3265) );
  AOI21_X1 U10369 ( .B1(n9046), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9045), .ZN(
        n9047) );
  OAI21_X1 U10370 ( .B1(n9049), .B2(n9048), .A(n9047), .ZN(P2_U3267) );
  MUX2_X1 U10371 ( .A(n9050), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10372 ( .A(n9108), .ZN(n9053) );
  NOR3_X1 U10373 ( .A1(n9127), .A2(n9131), .A3(n9051), .ZN(n9052) );
  OAI21_X1 U10374 ( .B1(n9053), .B2(n9052), .A(n9151), .ZN(n9057) );
  AOI22_X1 U10375 ( .A1(n9152), .A2(n9428), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9054) );
  OAI21_X1 U10376 ( .B1(n9457), .B2(n9662), .A(n9054), .ZN(n9055) );
  AOI21_X1 U10377 ( .B1(n9417), .B2(n9161), .A(n9055), .ZN(n9056) );
  OAI211_X1 U10378 ( .C1(n9419), .C2(n9157), .A(n9057), .B(n9056), .ZN(
        P1_U3216) );
  XNOR2_X1 U10379 ( .A(n9058), .B(n9059), .ZN(n9140) );
  NOR2_X1 U10380 ( .A1(n9140), .A2(n9139), .ZN(n9138) );
  AOI21_X1 U10381 ( .B1(n9059), .B2(n9058), .A(n9138), .ZN(n9063) );
  XNOR2_X1 U10382 ( .A(n9061), .B(n9060), .ZN(n9062) );
  XNOR2_X1 U10383 ( .A(n9063), .B(n9062), .ZN(n9070) );
  AND2_X1 U10384 ( .A1(n9176), .A2(n9425), .ZN(n9064) );
  AOI21_X1 U10385 ( .B1(n9065), .B2(n9427), .A(n9064), .ZN(n9489) );
  INV_X1 U10386 ( .A(n9066), .ZN(n9164) );
  NAND2_X1 U10387 ( .A1(n9161), .A2(n9493), .ZN(n9067) );
  NAND2_X1 U10388 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9324) );
  OAI211_X1 U10389 ( .C1(n9489), .C2(n9164), .A(n9067), .B(n9324), .ZN(n9068)
         );
  AOI21_X1 U10390 ( .B1(n9492), .B2(n9675), .A(n9068), .ZN(n9069) );
  OAI21_X1 U10391 ( .B1(n9070), .B2(n9671), .A(n9069), .ZN(P1_U3219) );
  XOR2_X1 U10392 ( .A(n9072), .B(n9071), .Z(n9077) );
  NOR2_X1 U10393 ( .A1(n9678), .A2(n9461), .ZN(n9075) );
  AOI22_X1 U10394 ( .A1(n9152), .A2(n9426), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9073) );
  OAI21_X1 U10395 ( .B1(n9455), .B2(n9662), .A(n9073), .ZN(n9074) );
  AOI211_X1 U10396 ( .C1(n9562), .C2(n9675), .A(n9075), .B(n9074), .ZN(n9076)
         );
  OAI21_X1 U10397 ( .B1(n9077), .B2(n9671), .A(n9076), .ZN(P1_U3223) );
  AOI21_X1 U10398 ( .B1(n9079), .B2(n9078), .A(n9149), .ZN(n9084) );
  AOI22_X1 U10399 ( .A1(n9152), .A2(n9358), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9081) );
  NAND2_X1 U10400 ( .A1(n9161), .A2(n9391), .ZN(n9080) );
  OAI211_X1 U10401 ( .C1(n9388), .C2(n9662), .A(n9081), .B(n9080), .ZN(n9082)
         );
  AOI21_X1 U10402 ( .B1(n9542), .B2(n9675), .A(n9082), .ZN(n9083) );
  OAI21_X1 U10403 ( .B1(n9084), .B2(n9671), .A(n9083), .ZN(P1_U3225) );
  OAI21_X1 U10404 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(n9088) );
  NAND2_X1 U10405 ( .A1(n9088), .A2(n9151), .ZN(n9093) );
  NAND2_X1 U10406 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9769) );
  OAI21_X1 U10407 ( .B1(n9164), .B2(n9089), .A(n9769), .ZN(n9090) );
  AOI21_X1 U10408 ( .B1(n9091), .B2(n9161), .A(n9090), .ZN(n9092) );
  OAI211_X1 U10409 ( .C1(n9632), .C2(n9157), .A(n9093), .B(n9092), .ZN(
        P1_U3226) );
  NAND2_X1 U10410 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  XNOR2_X1 U10411 ( .A(n9097), .B(n9096), .ZN(n9105) );
  NAND2_X1 U10412 ( .A1(n9152), .A2(n9176), .ZN(n9098) );
  NAND2_X1 U10413 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9781) );
  OAI211_X1 U10414 ( .C1(n9099), .C2(n9662), .A(n9098), .B(n9781), .ZN(n9102)
         );
  NOR2_X1 U10415 ( .A1(n9100), .A2(n9157), .ZN(n9101) );
  AOI211_X1 U10416 ( .C1(n9103), .C2(n9161), .A(n9102), .B(n9101), .ZN(n9104)
         );
  OAI21_X1 U10417 ( .B1(n9105), .B2(n9671), .A(n9104), .ZN(P1_U3228) );
  AND3_X1 U10418 ( .A1(n9108), .A2(n9107), .A3(n9106), .ZN(n9109) );
  OAI21_X1 U10419 ( .B1(n9110), .B2(n9109), .A(n9151), .ZN(n9116) );
  AND2_X1 U10420 ( .A1(n9173), .A2(n9425), .ZN(n9111) );
  AOI21_X1 U10421 ( .B1(n9112), .B2(n9427), .A(n9111), .ZN(n9401) );
  OAI22_X1 U10422 ( .A1(n9164), .A2(n9401), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9113), .ZN(n9114) );
  AOI21_X1 U10423 ( .B1(n9406), .B2(n9161), .A(n9114), .ZN(n9115) );
  OAI211_X1 U10424 ( .C1(n9608), .C2(n9157), .A(n9116), .B(n9115), .ZN(
        P1_U3229) );
  XNOR2_X1 U10425 ( .A(n9118), .B(n9117), .ZN(n9119) );
  XNOR2_X1 U10426 ( .A(n9120), .B(n9119), .ZN(n9126) );
  NOR2_X1 U10427 ( .A1(n9678), .A2(n9478), .ZN(n9124) );
  AND2_X1 U10428 ( .A1(n9175), .A2(n9425), .ZN(n9121) );
  AOI21_X1 U10429 ( .B1(n9174), .B2(n9427), .A(n9121), .ZN(n9473) );
  OAI22_X1 U10430 ( .A1(n9164), .A2(n9473), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9122), .ZN(n9123) );
  OAI21_X1 U10431 ( .B1(n9126), .B2(n9671), .A(n9125), .ZN(P1_U3233) );
  INV_X1 U10432 ( .A(n9127), .ZN(n9132) );
  OAI21_X1 U10433 ( .B1(n9129), .B2(n9131), .A(n9128), .ZN(n9130) );
  OAI21_X1 U10434 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(n9133) );
  NAND2_X1 U10435 ( .A1(n9133), .A2(n9151), .ZN(n9137) );
  AND2_X1 U10436 ( .A1(n9173), .A2(n9427), .ZN(n9134) );
  AOI21_X1 U10437 ( .B1(n9174), .B2(n9425), .A(n9134), .ZN(n9438) );
  OAI22_X1 U10438 ( .A1(n9164), .A2(n9438), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10115), .ZN(n9135) );
  AOI21_X1 U10439 ( .B1(n9442), .B2(n9161), .A(n9135), .ZN(n9136) );
  OAI211_X1 U10440 ( .C1(n9613), .C2(n9157), .A(n9137), .B(n9136), .ZN(
        P1_U3235) );
  AOI21_X1 U10441 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9146) );
  NAND2_X1 U10442 ( .A1(n9175), .A2(n9427), .ZN(n9142) );
  NAND2_X1 U10443 ( .A1(n9177), .A2(n9425), .ZN(n9141) );
  AND2_X1 U10444 ( .A1(n9142), .A2(n9141), .ZN(n9506) );
  NAND2_X1 U10445 ( .A1(n9161), .A2(n9513), .ZN(n9143) );
  NAND2_X1 U10446 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9797) );
  OAI211_X1 U10447 ( .C1(n9506), .C2(n9164), .A(n9143), .B(n9797), .ZN(n9144)
         );
  AOI21_X1 U10448 ( .B1(n9511), .B2(n9675), .A(n9144), .ZN(n9145) );
  OAI21_X1 U10449 ( .B1(n9146), .B2(n9671), .A(n9145), .ZN(P1_U3238) );
  OAI21_X1 U10450 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9150) );
  NAND3_X1 U10451 ( .A1(n4526), .A2(n9151), .A3(n9150), .ZN(n9156) );
  AOI22_X1 U10452 ( .A1(n9152), .A2(n9172), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9153) );
  OAI21_X1 U10453 ( .B1(n9366), .B2(n9662), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10454 ( .B1(n9375), .B2(n9161), .A(n9154), .ZN(n9155) );
  OAI211_X1 U10455 ( .C1(n9603), .C2(n9157), .A(n9156), .B(n9155), .ZN(
        P1_U3240) );
  AOI21_X1 U10456 ( .B1(n9158), .B2(n9159), .A(n4289), .ZN(n9169) );
  NAND2_X1 U10457 ( .A1(n9161), .A2(n9160), .ZN(n9163) );
  NAND2_X1 U10458 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9755) );
  OAI211_X1 U10459 ( .C1(n9165), .C2(n9164), .A(n9163), .B(n9755), .ZN(n9166)
         );
  AOI21_X1 U10460 ( .B1(n9167), .B2(n9675), .A(n9166), .ZN(n9168) );
  OAI21_X1 U10461 ( .B1(n9169), .B2(n9671), .A(n9168), .ZN(P1_U3241) );
  MUX2_X1 U10462 ( .A(n9171), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9170), .Z(
        P1_U3584) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9359), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9172), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9358), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9428), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9173), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9426), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9174), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9176), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9177), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9180), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9181), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9182), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9183), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9184), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9186), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9187), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9188), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9189), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9190), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9192), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5683), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10489 ( .C1(n9195), .C2(n9194), .A(n9788), .B(n9193), .ZN(n9203)
         );
  OAI211_X1 U10490 ( .C1(n9198), .C2(n9197), .A(n9784), .B(n9196), .ZN(n9202)
         );
  AOI22_X1 U10491 ( .A1(n9683), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9201) );
  NAND2_X1 U10492 ( .A1(n9777), .A2(n9199), .ZN(n9200) );
  NAND4_X1 U10493 ( .A1(n9203), .A2(n9202), .A3(n9201), .A4(n9200), .ZN(
        P1_U3244) );
  INV_X1 U10494 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U10495 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9204) );
  OAI21_X1 U10496 ( .B1(n9799), .B2(n9205), .A(n9204), .ZN(n9206) );
  AOI21_X1 U10497 ( .B1(n9207), .B2(n9777), .A(n9206), .ZN(n9216) );
  OAI211_X1 U10498 ( .C1(n9210), .C2(n9209), .A(n9784), .B(n9208), .ZN(n9215)
         );
  OAI211_X1 U10499 ( .C1(n9213), .C2(n9212), .A(n9788), .B(n9211), .ZN(n9214)
         );
  NAND3_X1 U10500 ( .A1(n9216), .A2(n9215), .A3(n9214), .ZN(P1_U3246) );
  NAND2_X1 U10501 ( .A1(n9683), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9217) );
  OAI211_X1 U10502 ( .C1(n9795), .C2(n9219), .A(n9218), .B(n9217), .ZN(n9220)
         );
  INV_X1 U10503 ( .A(n9220), .ZN(n9229) );
  OAI211_X1 U10504 ( .C1(n9223), .C2(n9222), .A(n9788), .B(n9221), .ZN(n9228)
         );
  OAI211_X1 U10505 ( .C1(n9226), .C2(n9225), .A(n9784), .B(n9224), .ZN(n9227)
         );
  NAND4_X1 U10506 ( .A1(n9230), .A2(n9229), .A3(n9228), .A4(n9227), .ZN(
        P1_U3247) );
  INV_X1 U10507 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9232) );
  OAI21_X1 U10508 ( .B1(n9799), .B2(n9232), .A(n9231), .ZN(n9233) );
  AOI21_X1 U10509 ( .B1(n9234), .B2(n9777), .A(n9233), .ZN(n9243) );
  OAI211_X1 U10510 ( .C1(n9237), .C2(n9236), .A(n9784), .B(n9235), .ZN(n9242)
         );
  OAI211_X1 U10511 ( .C1(n9240), .C2(n9239), .A(n9788), .B(n9238), .ZN(n9241)
         );
  NAND3_X1 U10512 ( .A1(n9243), .A2(n9242), .A3(n9241), .ZN(P1_U3248) );
  INV_X1 U10513 ( .A(n9244), .ZN(n9248) );
  INV_X1 U10514 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U10515 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9245) );
  OAI21_X1 U10516 ( .B1(n9799), .B2(n9246), .A(n9245), .ZN(n9247) );
  AOI21_X1 U10517 ( .B1(n9248), .B2(n9777), .A(n9247), .ZN(n9257) );
  OAI211_X1 U10518 ( .C1(n9251), .C2(n9250), .A(n9784), .B(n9249), .ZN(n9256)
         );
  OAI211_X1 U10519 ( .C1(n9254), .C2(n9253), .A(n9788), .B(n9252), .ZN(n9255)
         );
  NAND3_X1 U10520 ( .A1(n9257), .A2(n9256), .A3(n9255), .ZN(P1_U3249) );
  INV_X1 U10521 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U10522 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9258) );
  OAI21_X1 U10523 ( .B1(n9799), .B2(n9259), .A(n9258), .ZN(n9260) );
  AOI21_X1 U10524 ( .B1(n9261), .B2(n9777), .A(n9260), .ZN(n9270) );
  OAI211_X1 U10525 ( .C1(n9264), .C2(n9263), .A(n9784), .B(n9262), .ZN(n9269)
         );
  OAI211_X1 U10526 ( .C1(n9267), .C2(n9266), .A(n9788), .B(n9265), .ZN(n9268)
         );
  NAND3_X1 U10527 ( .A1(n9270), .A2(n9269), .A3(n9268), .ZN(P1_U3250) );
  INV_X1 U10528 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9272) );
  OAI21_X1 U10529 ( .B1(n9799), .B2(n9272), .A(n9271), .ZN(n9273) );
  AOI21_X1 U10530 ( .B1(n9274), .B2(n9777), .A(n9273), .ZN(n9283) );
  OAI211_X1 U10531 ( .C1(n9277), .C2(n9276), .A(n9788), .B(n9275), .ZN(n9282)
         );
  OAI211_X1 U10532 ( .C1(n9280), .C2(n9279), .A(n9784), .B(n9278), .ZN(n9281)
         );
  NAND3_X1 U10533 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(P1_U3251) );
  NAND2_X1 U10534 ( .A1(n9715), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9284) );
  OAI21_X1 U10535 ( .B1(n9715), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9284), .ZN(
        n9718) );
  NOR2_X1 U10536 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9699), .ZN(n9285) );
  AOI21_X1 U10537 ( .B1(n9699), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9285), .ZN(
        n9706) );
  OR2_X1 U10538 ( .A1(n9300), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U10539 ( .A1(n9287), .A2(n9286), .ZN(n9644) );
  OR2_X1 U10540 ( .A1(n9651), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U10541 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9651), .ZN(n9288) );
  NAND2_X1 U10542 ( .A1(n9289), .A2(n9288), .ZN(n9643) );
  NOR2_X1 U10543 ( .A1(n9644), .A2(n9643), .ZN(n9655) );
  AOI21_X1 U10544 ( .B1(n9651), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9655), .ZN(
        n9689) );
  NAND2_X1 U10545 ( .A1(n9695), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9290) );
  OAI21_X1 U10546 ( .B1(n9695), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9290), .ZN(
        n9688) );
  NOR2_X1 U10547 ( .A1(n9689), .A2(n9688), .ZN(n9687) );
  AOI21_X1 U10548 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9695), .A(n9687), .ZN(
        n9705) );
  NAND2_X1 U10549 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  OAI21_X1 U10550 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9699), .A(n9704), .ZN(
        n9717) );
  NOR2_X1 U10551 ( .A1(n9718), .A2(n9717), .ZN(n9716) );
  AOI21_X1 U10552 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9715), .A(n9716), .ZN(
        n9733) );
  NAND2_X1 U10553 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9731), .ZN(n9291) );
  OAI21_X1 U10554 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9731), .A(n9291), .ZN(
        n9734) );
  NOR2_X1 U10555 ( .A1(n9733), .A2(n9734), .ZN(n9732) );
  AOI21_X1 U10556 ( .B1(n9731), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9732), .ZN(
        n9292) );
  NOR2_X1 U10557 ( .A1(n9292), .A2(n9307), .ZN(n9293) );
  INV_X1 U10558 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9750) );
  XOR2_X1 U10559 ( .A(n9754), .B(n9292), .Z(n9751) );
  NOR2_X1 U10560 ( .A1(n9750), .A2(n9751), .ZN(n9749) );
  NOR2_X1 U10561 ( .A1(n9293), .A2(n9749), .ZN(n9760) );
  XNOR2_X1 U10562 ( .A(n9309), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9759) );
  OR2_X1 U10563 ( .A1(n9760), .A2(n9759), .ZN(n9767) );
  NAND2_X1 U10564 ( .A1(n9309), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9294) );
  AND2_X1 U10565 ( .A1(n9767), .A2(n9294), .ZN(n9773) );
  INV_X1 U10566 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9295) );
  XNOR2_X1 U10567 ( .A(n9778), .B(n9295), .ZN(n9774) );
  NAND2_X1 U10568 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  OR2_X1 U10569 ( .A1(n9778), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U10570 ( .A1(n9313), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9298) );
  OR2_X1 U10571 ( .A1(n9313), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9297) );
  AND2_X1 U10572 ( .A1(n9298), .A2(n9297), .ZN(n9786) );
  NAND2_X1 U10573 ( .A1(n9787), .A2(n9786), .ZN(n9785) );
  NAND2_X1 U10574 ( .A1(n9785), .A2(n9298), .ZN(n9299) );
  XNOR2_X1 U10575 ( .A(n9299), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9320) );
  INV_X1 U10576 ( .A(n9320), .ZN(n9317) );
  XNOR2_X1 U10577 ( .A(n9715), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9722) );
  OR2_X1 U10578 ( .A1(n9699), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9305) );
  OR2_X1 U10579 ( .A1(n9300), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U10580 ( .A1(n9302), .A2(n9301), .ZN(n9648) );
  MUX2_X1 U10581 ( .A(n7321), .B(P1_REG1_REG_10__SCAN_IN), .S(n9651), .Z(n9647) );
  NOR2_X1 U10582 ( .A1(n9648), .A2(n9647), .ZN(n9646) );
  AOI21_X1 U10583 ( .B1(n9651), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9646), .ZN(
        n9692) );
  INV_X1 U10584 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9303) );
  MUX2_X1 U10585 ( .A(n9303), .B(P1_REG1_REG_11__SCAN_IN), .S(n9695), .Z(n9691) );
  NOR2_X1 U10586 ( .A1(n9692), .A2(n9691), .ZN(n9690) );
  AOI21_X1 U10587 ( .B1(n9695), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9690), .ZN(
        n9701) );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9304), .S(n9699), .Z(n9702) );
  NAND2_X1 U10589 ( .A1(n9701), .A2(n9702), .ZN(n9700) );
  NAND2_X1 U10590 ( .A1(n9305), .A2(n9700), .ZN(n9721) );
  NOR2_X1 U10591 ( .A1(n9722), .A2(n9721), .ZN(n9720) );
  AOI21_X1 U10592 ( .B1(n9715), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9720), .ZN(
        n9738) );
  XNOR2_X1 U10593 ( .A(n9731), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9737) );
  NOR2_X1 U10594 ( .A1(n9738), .A2(n9737), .ZN(n9736) );
  AOI21_X1 U10595 ( .B1(n9731), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9736), .ZN(
        n9306) );
  NOR2_X1 U10596 ( .A1(n9306), .A2(n9307), .ZN(n9308) );
  XNOR2_X1 U10597 ( .A(n9307), .B(n9306), .ZN(n9748) );
  NOR2_X1 U10598 ( .A1(n9747), .A2(n9748), .ZN(n9746) );
  NOR2_X1 U10599 ( .A1(n9308), .A2(n9746), .ZN(n9762) );
  INV_X1 U10600 ( .A(n9762), .ZN(n9310) );
  XNOR2_X1 U10601 ( .A(n9309), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9761) );
  OAI22_X1 U10602 ( .A1(n9310), .A2(n9761), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n9309), .ZN(n9776) );
  INV_X1 U10603 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9312) );
  XNOR2_X1 U10604 ( .A(n9778), .B(n9312), .ZN(n9775) );
  AOI22_X1 U10605 ( .A1(n9776), .A2(n9775), .B1(n9312), .B2(n9311), .ZN(n9791)
         );
  INV_X1 U10606 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9577) );
  AND2_X1 U10607 ( .A1(n9313), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9314) );
  AOI21_X1 U10608 ( .B1(n9577), .B2(n9794), .A(n9314), .ZN(n9790) );
  NAND2_X1 U10609 ( .A1(n9791), .A2(n9790), .ZN(n9789) );
  INV_X1 U10610 ( .A(n9314), .ZN(n9315) );
  NAND2_X1 U10611 ( .A1(n9789), .A2(n9315), .ZN(n9316) );
  INV_X1 U10612 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10028) );
  XNOR2_X1 U10613 ( .A(n9316), .B(n10028), .ZN(n9318) );
  AOI22_X1 U10614 ( .A1(n9317), .A2(n9784), .B1(n9788), .B2(n9318), .ZN(n9323)
         );
  OAI21_X1 U10615 ( .B1(n9318), .B2(n9764), .A(n9795), .ZN(n9319) );
  AOI21_X1 U10616 ( .B1(n9320), .B2(n9784), .A(n9319), .ZN(n9322) );
  MUX2_X1 U10617 ( .A(n9323), .B(n9322), .S(n9321), .Z(n9325) );
  OAI211_X1 U10618 ( .C1(n4907), .C2(n9799), .A(n9325), .B(n9324), .ZN(
        P1_U3262) );
  NAND2_X1 U10619 ( .A1(n9329), .A2(n9328), .ZN(n9525) );
  NOR2_X1 U10620 ( .A1(n9494), .A2(n9525), .ZN(n9336) );
  NOR2_X1 U10621 ( .A1(n9595), .A2(n9516), .ZN(n9331) );
  AOI211_X1 U10622 ( .C1(n9813), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9336), .B(
        n9331), .ZN(n9332) );
  OAI21_X1 U10623 ( .B1(n9522), .B2(n9806), .A(n9332), .ZN(P1_U3263) );
  XNOR2_X1 U10624 ( .A(n9333), .B(n9598), .ZN(n9334) );
  NAND2_X1 U10625 ( .A1(n9527), .A2(n9512), .ZN(n9338) );
  AND2_X1 U10626 ( .A1(n9813), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9335) );
  NOR2_X1 U10627 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  OAI211_X1 U10628 ( .C1(n9598), .C2(n9516), .A(n9338), .B(n9337), .ZN(
        P1_U3264) );
  NAND2_X1 U10629 ( .A1(n9339), .A2(n9809), .ZN(n9346) );
  INV_X1 U10630 ( .A(n5776), .ZN(n9342) );
  AOI22_X1 U10631 ( .A1(n9813), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9340), .B2(
        n9800), .ZN(n9341) );
  OAI21_X1 U10632 ( .B1(n9342), .B2(n9516), .A(n9341), .ZN(n9343) );
  AOI21_X1 U10633 ( .B1(n9344), .B2(n9512), .A(n9343), .ZN(n9345) );
  OAI211_X1 U10634 ( .C1(n4864), .C2(n9494), .A(n9346), .B(n9345), .ZN(
        P1_U3356) );
  XOR2_X1 U10635 ( .A(n9354), .B(n9347), .Z(n9534) );
  INV_X1 U10636 ( .A(n9373), .ZN(n9349) );
  AOI211_X1 U10637 ( .C1(n9531), .C2(n9349), .A(n9509), .B(n9348), .ZN(n9530)
         );
  AOI22_X1 U10638 ( .A1(n9813), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9350), .B2(
        n9800), .ZN(n9351) );
  OAI21_X1 U10639 ( .B1(n9352), .B2(n9516), .A(n9351), .ZN(n9362) );
  NAND3_X1 U10640 ( .A1(n9353), .A2(n9355), .A3(n4623), .ZN(n9356) );
  NAND2_X1 U10641 ( .A1(n9357), .A2(n9356), .ZN(n9360) );
  AOI222_X1 U10642 ( .A1(n9504), .A2(n9360), .B1(n9359), .B2(n9427), .C1(n9358), .C2(n9425), .ZN(n9533) );
  NOR2_X1 U10643 ( .A1(n9533), .A2(n9494), .ZN(n9361) );
  AOI211_X1 U10644 ( .C1(n9512), .C2(n9530), .A(n9362), .B(n9361), .ZN(n9363)
         );
  OAI21_X1 U10645 ( .B1(n9534), .B2(n9520), .A(n9363), .ZN(P1_U3266) );
  OAI21_X1 U10646 ( .B1(n9364), .B2(n9371), .A(n9353), .ZN(n9365) );
  NAND2_X1 U10647 ( .A1(n9365), .A2(n9504), .ZN(n9370) );
  OAI22_X1 U10648 ( .A1(n9367), .A2(n9458), .B1(n9366), .B2(n9456), .ZN(n9368)
         );
  INV_X1 U10649 ( .A(n9368), .ZN(n9369) );
  NAND2_X1 U10650 ( .A1(n9370), .A2(n9369), .ZN(n9535) );
  INV_X1 U10651 ( .A(n9535), .ZN(n9380) );
  XOR2_X1 U10652 ( .A(n9372), .B(n9371), .Z(n9537) );
  NAND2_X1 U10653 ( .A1(n9537), .A2(n9809), .ZN(n9379) );
  AOI211_X1 U10654 ( .C1(n9374), .C2(n9389), .A(n9509), .B(n9373), .ZN(n9536)
         );
  AOI22_X1 U10655 ( .A1(n9813), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9375), .B2(
        n9800), .ZN(n9376) );
  OAI21_X1 U10656 ( .B1(n9603), .B2(n9516), .A(n9376), .ZN(n9377) );
  AOI21_X1 U10657 ( .B1(n9536), .B2(n9512), .A(n9377), .ZN(n9378) );
  OAI211_X1 U10658 ( .C1(n9813), .C2(n9380), .A(n9379), .B(n9378), .ZN(
        P1_U3267) );
  XNOR2_X1 U10659 ( .A(n9381), .B(n9385), .ZN(n9544) );
  INV_X1 U10660 ( .A(n9382), .ZN(n9383) );
  AOI21_X1 U10661 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9386) );
  OAI222_X1 U10662 ( .A1(n9456), .A2(n9388), .B1(n9458), .B2(n9387), .C1(n9453), .C2(n9386), .ZN(n9540) );
  INV_X1 U10663 ( .A(n9389), .ZN(n9390) );
  AOI211_X1 U10664 ( .C1(n9542), .C2(n9404), .A(n9509), .B(n9390), .ZN(n9541)
         );
  NAND2_X1 U10665 ( .A1(n9541), .A2(n9512), .ZN(n9393) );
  AOI22_X1 U10666 ( .A1(n9813), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9391), .B2(
        n9800), .ZN(n9392) );
  OAI211_X1 U10667 ( .C1(n9394), .C2(n9516), .A(n9393), .B(n9392), .ZN(n9395)
         );
  AOI21_X1 U10668 ( .B1(n9540), .B2(n9518), .A(n9395), .ZN(n9396) );
  OAI21_X1 U10669 ( .B1(n9544), .B2(n9520), .A(n9396), .ZN(P1_U3268) );
  XNOR2_X1 U10670 ( .A(n9397), .B(n9399), .ZN(n9547) );
  INV_X1 U10671 ( .A(n9547), .ZN(n9411) );
  NAND2_X1 U10672 ( .A1(n9398), .A2(n9504), .ZN(n9403) );
  AOI21_X1 U10673 ( .B1(n9423), .B2(n9400), .A(n9399), .ZN(n9402) );
  OAI21_X1 U10674 ( .B1(n9403), .B2(n9402), .A(n9401), .ZN(n9545) );
  AOI211_X1 U10675 ( .C1(n9405), .C2(n9414), .A(n9509), .B(n4541), .ZN(n9546)
         );
  NAND2_X1 U10676 ( .A1(n9546), .A2(n9512), .ZN(n9408) );
  AOI22_X1 U10677 ( .A1(n9813), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9406), .B2(
        n9800), .ZN(n9407) );
  OAI211_X1 U10678 ( .C1(n9608), .C2(n9516), .A(n9408), .B(n9407), .ZN(n9409)
         );
  AOI21_X1 U10679 ( .B1(n9518), .B2(n9545), .A(n9409), .ZN(n9410) );
  OAI21_X1 U10680 ( .B1(n9411), .B2(n9520), .A(n9410), .ZN(P1_U3269) );
  XNOR2_X1 U10681 ( .A(n9413), .B(n9412), .ZN(n9555) );
  INV_X1 U10682 ( .A(n9440), .ZN(n9416) );
  INV_X1 U10683 ( .A(n9414), .ZN(n9415) );
  AOI21_X1 U10684 ( .B1(n9550), .B2(n9416), .A(n9415), .ZN(n9552) );
  AOI22_X1 U10685 ( .A1(n9813), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9417), .B2(
        n9800), .ZN(n9418) );
  OAI21_X1 U10686 ( .B1(n9419), .B2(n9516), .A(n9418), .ZN(n9431) );
  INV_X1 U10687 ( .A(n9435), .ZN(n9422) );
  OAI21_X1 U10688 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9424) );
  NAND2_X1 U10689 ( .A1(n9424), .A2(n9423), .ZN(n9429) );
  AOI222_X1 U10690 ( .A1(n9504), .A2(n9429), .B1(n9428), .B2(n9427), .C1(n9426), .C2(n9425), .ZN(n9554) );
  NOR2_X1 U10691 ( .A1(n9554), .A2(n9494), .ZN(n9430) );
  AOI211_X1 U10692 ( .C1(n9552), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9433)
         );
  OAI21_X1 U10693 ( .B1(n9555), .B2(n9520), .A(n9433), .ZN(P1_U3270) );
  XNOR2_X1 U10694 ( .A(n9434), .B(n9436), .ZN(n9558) );
  INV_X1 U10695 ( .A(n9558), .ZN(n9447) );
  OAI211_X1 U10696 ( .C1(n9437), .C2(n9436), .A(n9435), .B(n9504), .ZN(n9439)
         );
  NAND2_X1 U10697 ( .A1(n9439), .A2(n9438), .ZN(n9556) );
  AOI211_X1 U10698 ( .C1(n9441), .C2(n9459), .A(n9509), .B(n9440), .ZN(n9557)
         );
  NAND2_X1 U10699 ( .A1(n9557), .A2(n9512), .ZN(n9444) );
  AOI22_X1 U10700 ( .A1(n9813), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9442), .B2(
        n9800), .ZN(n9443) );
  OAI211_X1 U10701 ( .C1(n9613), .C2(n9516), .A(n9444), .B(n9443), .ZN(n9445)
         );
  AOI21_X1 U10702 ( .B1(n9556), .B2(n9518), .A(n9445), .ZN(n9446) );
  OAI21_X1 U10703 ( .B1(n9447), .B2(n9520), .A(n9446), .ZN(P1_U3271) );
  XNOR2_X1 U10704 ( .A(n9450), .B(n9449), .ZN(n9564) );
  XNOR2_X1 U10705 ( .A(n9452), .B(n9451), .ZN(n9454) );
  OAI222_X1 U10706 ( .A1(n9458), .A2(n9457), .B1(n9456), .B2(n9455), .C1(n9454), .C2(n9453), .ZN(n9560) );
  INV_X1 U10707 ( .A(n9459), .ZN(n9460) );
  AOI211_X1 U10708 ( .C1(n9562), .C2(n9475), .A(n9509), .B(n9460), .ZN(n9561)
         );
  NAND2_X1 U10709 ( .A1(n9561), .A2(n9512), .ZN(n9464) );
  INV_X1 U10710 ( .A(n9461), .ZN(n9462) );
  AOI22_X1 U10711 ( .A1(n9494), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9462), .B2(
        n9800), .ZN(n9463) );
  OAI211_X1 U10712 ( .C1(n9465), .C2(n9516), .A(n9464), .B(n9463), .ZN(n9466)
         );
  AOI21_X1 U10713 ( .B1(n9560), .B2(n9518), .A(n9466), .ZN(n9467) );
  OAI21_X1 U10714 ( .B1(n9564), .B2(n9520), .A(n9467), .ZN(P1_U3272) );
  XOR2_X1 U10715 ( .A(n9468), .B(n9469), .Z(n9567) );
  INV_X1 U10716 ( .A(n9567), .ZN(n9484) );
  INV_X1 U10717 ( .A(n9469), .ZN(n9470) );
  XNOR2_X1 U10718 ( .A(n9471), .B(n9470), .ZN(n9472) );
  NAND2_X1 U10719 ( .A1(n9472), .A2(n9504), .ZN(n9474) );
  NAND2_X1 U10720 ( .A1(n9474), .A2(n9473), .ZN(n9565) );
  INV_X1 U10721 ( .A(n9491), .ZN(n9477) );
  INV_X1 U10722 ( .A(n9475), .ZN(n9476) );
  NAND2_X1 U10723 ( .A1(n9566), .A2(n9512), .ZN(n9481) );
  INV_X1 U10724 ( .A(n9478), .ZN(n9479) );
  AOI22_X1 U10725 ( .A1(n9494), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9479), .B2(
        n9800), .ZN(n9480) );
  OAI211_X1 U10726 ( .C1(n9618), .C2(n9516), .A(n9481), .B(n9480), .ZN(n9482)
         );
  AOI21_X1 U10727 ( .B1(n9565), .B2(n9518), .A(n9482), .ZN(n9483) );
  OAI21_X1 U10728 ( .B1(n9484), .B2(n9520), .A(n9483), .ZN(P1_U3273) );
  XNOR2_X1 U10729 ( .A(n9485), .B(n9486), .ZN(n9572) );
  INV_X1 U10730 ( .A(n9572), .ZN(n9499) );
  XNOR2_X1 U10731 ( .A(n9487), .B(n9486), .ZN(n9488) );
  NAND2_X1 U10732 ( .A1(n9488), .A2(n9504), .ZN(n9490) );
  NAND2_X1 U10733 ( .A1(n9490), .A2(n9489), .ZN(n9570) );
  AOI211_X1 U10734 ( .C1(n9492), .C2(n4547), .A(n9509), .B(n9491), .ZN(n9571)
         );
  NAND2_X1 U10735 ( .A1(n9571), .A2(n9512), .ZN(n9496) );
  AOI22_X1 U10736 ( .A1(n9494), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9493), .B2(
        n9800), .ZN(n9495) );
  OAI211_X1 U10737 ( .C1(n9622), .C2(n9516), .A(n9496), .B(n9495), .ZN(n9497)
         );
  AOI21_X1 U10738 ( .B1(n9570), .B2(n9518), .A(n9497), .ZN(n9498) );
  OAI21_X1 U10739 ( .B1(n9499), .B2(n9520), .A(n9498), .ZN(P1_U3274) );
  XNOR2_X1 U10740 ( .A(n9501), .B(n4390), .ZN(n9576) );
  INV_X1 U10741 ( .A(n9576), .ZN(n9521) );
  XNOR2_X1 U10742 ( .A(n9503), .B(n9502), .ZN(n9505) );
  NAND2_X1 U10743 ( .A1(n9505), .A2(n9504), .ZN(n9507) );
  NAND2_X1 U10744 ( .A1(n9507), .A2(n9506), .ZN(n9574) );
  AOI211_X1 U10745 ( .C1(n9511), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9575)
         );
  NAND2_X1 U10746 ( .A1(n9575), .A2(n9512), .ZN(n9515) );
  AOI22_X1 U10747 ( .A1(n9813), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9513), .B2(
        n9800), .ZN(n9514) );
  OAI211_X1 U10748 ( .C1(n4545), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9517)
         );
  AOI21_X1 U10749 ( .B1(n9574), .B2(n9518), .A(n9517), .ZN(n9519) );
  OAI21_X1 U10750 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(P1_U3275) );
  INV_X1 U10751 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9523) );
  MUX2_X1 U10752 ( .A(n9523), .B(n9592), .S(n9854), .Z(n9524) );
  OAI21_X1 U10753 ( .B1(n9595), .B2(n9590), .A(n9524), .ZN(P1_U3553) );
  INV_X1 U10754 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9528) );
  INV_X1 U10755 ( .A(n9525), .ZN(n9526) );
  NOR2_X1 U10756 ( .A1(n9527), .A2(n9526), .ZN(n9596) );
  MUX2_X1 U10757 ( .A(n9528), .B(n9596), .S(n9854), .Z(n9529) );
  OAI21_X1 U10758 ( .B1(n9598), .B2(n9590), .A(n9529), .ZN(P1_U3552) );
  AOI21_X1 U10759 ( .B1(n9837), .B2(n9531), .A(n9530), .ZN(n9532) );
  OAI211_X1 U10760 ( .C1(n9534), .C2(n9583), .A(n9533), .B(n9532), .ZN(n9599)
         );
  MUX2_X1 U10761 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9599), .S(n9854), .Z(
        P1_U3549) );
  INV_X1 U10762 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9538) );
  AOI211_X1 U10763 ( .C1(n9537), .C2(n9835), .A(n9536), .B(n9535), .ZN(n9600)
         );
  MUX2_X1 U10764 ( .A(n9538), .B(n9600), .S(n9854), .Z(n9539) );
  OAI21_X1 U10765 ( .B1(n9603), .B2(n9590), .A(n9539), .ZN(P1_U3548) );
  AOI211_X1 U10766 ( .C1(n9837), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9543)
         );
  OAI21_X1 U10767 ( .B1(n9544), .B2(n9583), .A(n9543), .ZN(n9604) );
  MUX2_X1 U10768 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9604), .S(n9854), .Z(
        P1_U3547) );
  INV_X1 U10769 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9548) );
  AOI211_X1 U10770 ( .C1(n9547), .C2(n9835), .A(n9546), .B(n9545), .ZN(n9605)
         );
  MUX2_X1 U10771 ( .A(n9548), .B(n9605), .S(n9854), .Z(n9549) );
  OAI21_X1 U10772 ( .B1(n9608), .B2(n9590), .A(n9549), .ZN(P1_U3546) );
  AOI22_X1 U10773 ( .A1(n9552), .A2(n9551), .B1(n9837), .B2(n9550), .ZN(n9553)
         );
  OAI211_X1 U10774 ( .C1(n9555), .C2(n9583), .A(n9554), .B(n9553), .ZN(n9609)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9609), .S(n9854), .Z(
        P1_U3545) );
  INV_X1 U10776 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10046) );
  AOI211_X1 U10777 ( .C1(n9558), .C2(n9835), .A(n9557), .B(n9556), .ZN(n9610)
         );
  MUX2_X1 U10778 ( .A(n10046), .B(n9610), .S(n9854), .Z(n9559) );
  OAI21_X1 U10779 ( .B1(n9613), .B2(n9590), .A(n9559), .ZN(P1_U3544) );
  AOI211_X1 U10780 ( .C1(n9837), .C2(n9562), .A(n9561), .B(n9560), .ZN(n9563)
         );
  OAI21_X1 U10781 ( .B1(n9564), .B2(n9583), .A(n9563), .ZN(n9614) );
  MUX2_X1 U10782 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9614), .S(n9854), .Z(
        P1_U3543) );
  INV_X1 U10783 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9568) );
  AOI211_X1 U10784 ( .C1(n9567), .C2(n9835), .A(n9566), .B(n9565), .ZN(n9615)
         );
  MUX2_X1 U10785 ( .A(n9568), .B(n9615), .S(n9854), .Z(n9569) );
  OAI21_X1 U10786 ( .B1(n9618), .B2(n9590), .A(n9569), .ZN(P1_U3542) );
  AOI211_X1 U10787 ( .C1(n9572), .C2(n9835), .A(n9571), .B(n9570), .ZN(n9619)
         );
  MUX2_X1 U10788 ( .A(n10028), .B(n9619), .S(n9854), .Z(n9573) );
  OAI21_X1 U10789 ( .B1(n9622), .B2(n9590), .A(n9573), .ZN(P1_U3541) );
  AOI211_X1 U10790 ( .C1(n9576), .C2(n9835), .A(n9575), .B(n9574), .ZN(n9623)
         );
  MUX2_X1 U10791 ( .A(n9577), .B(n9623), .S(n9854), .Z(n9578) );
  OAI21_X1 U10792 ( .B1(n4545), .B2(n9590), .A(n9578), .ZN(P1_U3540) );
  AOI211_X1 U10793 ( .C1(n9837), .C2(n9581), .A(n9580), .B(n9579), .ZN(n9582)
         );
  OAI21_X1 U10794 ( .B1(n9584), .B2(n9583), .A(n9582), .ZN(n9626) );
  MUX2_X1 U10795 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9626), .S(n9854), .Z(
        P1_U3539) );
  INV_X1 U10796 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9588) );
  AOI211_X1 U10797 ( .C1(n9587), .C2(n9835), .A(n9586), .B(n9585), .ZN(n9628)
         );
  MUX2_X1 U10798 ( .A(n9588), .B(n9628), .S(n9854), .Z(n9589) );
  OAI21_X1 U10799 ( .B1(n9632), .B2(n9590), .A(n9589), .ZN(P1_U3538) );
  MUX2_X1 U10800 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9591), .S(n9854), .Z(
        P1_U3522) );
  INV_X1 U10801 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9593) );
  MUX2_X1 U10802 ( .A(n9593), .B(n9592), .S(n9627), .Z(n9594) );
  OAI21_X1 U10803 ( .B1(n9595), .B2(n9631), .A(n9594), .ZN(P1_U3521) );
  INV_X1 U10804 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10129) );
  MUX2_X1 U10805 ( .A(n10129), .B(n9596), .S(n9627), .Z(n9597) );
  OAI21_X1 U10806 ( .B1(n9598), .B2(n9631), .A(n9597), .ZN(P1_U3520) );
  MUX2_X1 U10807 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9599), .S(n9627), .Z(
        P1_U3517) );
  INV_X1 U10808 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9601) );
  MUX2_X1 U10809 ( .A(n9601), .B(n9600), .S(n9627), .Z(n9602) );
  OAI21_X1 U10810 ( .B1(n9603), .B2(n9631), .A(n9602), .ZN(P1_U3516) );
  MUX2_X1 U10811 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9604), .S(n9627), .Z(
        P1_U3515) );
  INV_X1 U10812 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9606) );
  MUX2_X1 U10813 ( .A(n9606), .B(n9605), .S(n9627), .Z(n9607) );
  OAI21_X1 U10814 ( .B1(n9608), .B2(n9631), .A(n9607), .ZN(P1_U3514) );
  MUX2_X1 U10815 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9609), .S(n9627), .Z(
        P1_U3513) );
  INV_X1 U10816 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U10817 ( .A(n9611), .B(n9610), .S(n9627), .Z(n9612) );
  OAI21_X1 U10818 ( .B1(n9613), .B2(n9631), .A(n9612), .ZN(P1_U3512) );
  MUX2_X1 U10819 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9614), .S(n9627), .Z(
        P1_U3511) );
  INV_X1 U10820 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9616) );
  MUX2_X1 U10821 ( .A(n9616), .B(n9615), .S(n9627), .Z(n9617) );
  OAI21_X1 U10822 ( .B1(n9618), .B2(n9631), .A(n9617), .ZN(P1_U3510) );
  INV_X1 U10823 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9620) );
  MUX2_X1 U10824 ( .A(n9620), .B(n9619), .S(n9627), .Z(n9621) );
  OAI21_X1 U10825 ( .B1(n9622), .B2(n9631), .A(n9621), .ZN(P1_U3509) );
  INV_X1 U10826 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U10827 ( .A(n9624), .B(n9623), .S(n9627), .Z(n9625) );
  OAI21_X1 U10828 ( .B1(n4545), .B2(n9631), .A(n9625), .ZN(P1_U3507) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9626), .S(n9627), .Z(
        P1_U3504) );
  INV_X1 U10830 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9629) );
  MUX2_X1 U10831 ( .A(n9629), .B(n9628), .S(n9627), .Z(n9630) );
  OAI21_X1 U10832 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(P1_U3501) );
  MUX2_X1 U10833 ( .A(n9633), .B(P1_D_REG_1__SCAN_IN), .S(n9815), .Z(P1_U3440)
         );
  MUX2_X1 U10834 ( .A(n9634), .B(P1_D_REG_0__SCAN_IN), .S(n9815), .Z(P1_U3439)
         );
  NOR4_X1 U10835 ( .A1(n4924), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n4875), .ZN(n9635) );
  AOI21_X1 U10836 ( .B1(n9638), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9635), .ZN(
        n9636) );
  OAI21_X1 U10837 ( .B1(n9637), .B2(n9640), .A(n9636), .ZN(P1_U3324) );
  AOI22_X1 U10838 ( .A1(n4928), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9638), .ZN(n9639) );
  OAI21_X1 U10839 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(P1_U3325) );
  MUX2_X1 U10840 ( .A(n9642), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10841 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U10842 ( .A1(n9644), .A2(n9643), .ZN(n9645) );
  NAND2_X1 U10843 ( .A1(n9784), .A2(n9645), .ZN(n9654) );
  INV_X1 U10844 ( .A(n9646), .ZN(n9650) );
  NAND2_X1 U10845 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  NAND3_X1 U10846 ( .A1(n9650), .A2(n9788), .A3(n9649), .ZN(n9653) );
  NAND2_X1 U10847 ( .A1(n9777), .A2(n9651), .ZN(n9652) );
  OAI211_X1 U10848 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9656)
         );
  INV_X1 U10849 ( .A(n9656), .ZN(n9658) );
  NAND2_X1 U10850 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9657) );
  OAI211_X1 U10851 ( .C1(n9799), .C2(n9659), .A(n9658), .B(n9657), .ZN(
        P1_U3253) );
  OAI22_X1 U10852 ( .A1(n9663), .A2(n9662), .B1(n9661), .B2(n9660), .ZN(n9674)
         );
  OAI21_X1 U10853 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9670) );
  AOI21_X1 U10854 ( .B1(n9668), .B2(n7580), .A(n9667), .ZN(n9669) );
  XOR2_X1 U10855 ( .A(n9670), .B(n9669), .Z(n9672) );
  NOR2_X1 U10856 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  AOI211_X1 U10857 ( .C1(n9838), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  NAND2_X1 U10858 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9696) );
  OAI211_X1 U10859 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9696), .ZN(
        P1_U3236) );
  XNOR2_X1 U10860 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10861 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10862 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9680) );
  AOI21_X1 U10863 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9682) );
  XNOR2_X1 U10864 ( .A(n9682), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9686) );
  AOI22_X1 U10865 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9683), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9684) );
  OAI21_X1 U10866 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(P1_U3243) );
  INV_X1 U10867 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9698) );
  AOI211_X1 U10868 ( .C1(n9689), .C2(n9688), .A(n9687), .B(n9758), .ZN(n9694)
         );
  AOI211_X1 U10869 ( .C1(n9692), .C2(n9691), .A(n9690), .B(n9764), .ZN(n9693)
         );
  AOI211_X1 U10870 ( .C1(n9777), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9697)
         );
  OAI211_X1 U10871 ( .C1(n9799), .C2(n9698), .A(n9697), .B(n9696), .ZN(
        P1_U3254) );
  INV_X1 U10872 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9714) );
  INV_X1 U10873 ( .A(n9699), .ZN(n9710) );
  OAI21_X1 U10874 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9703) );
  NAND2_X1 U10875 ( .A1(n9788), .A2(n9703), .ZN(n9709) );
  OAI21_X1 U10876 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  NAND2_X1 U10877 ( .A1(n9784), .A2(n9707), .ZN(n9708) );
  OAI211_X1 U10878 ( .C1(n9795), .C2(n9710), .A(n9709), .B(n9708), .ZN(n9711)
         );
  INV_X1 U10879 ( .A(n9711), .ZN(n9713) );
  OAI211_X1 U10880 ( .C1(n9799), .C2(n9714), .A(n9713), .B(n9712), .ZN(
        P1_U3255) );
  INV_X1 U10881 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9730) );
  INV_X1 U10882 ( .A(n9715), .ZN(n9726) );
  AOI21_X1 U10883 ( .B1(n9718), .B2(n9717), .A(n9716), .ZN(n9719) );
  NAND2_X1 U10884 ( .A1(n9784), .A2(n9719), .ZN(n9725) );
  AOI21_X1 U10885 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  NAND2_X1 U10886 ( .A1(n9788), .A2(n9723), .ZN(n9724) );
  OAI211_X1 U10887 ( .C1(n9795), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9727)
         );
  INV_X1 U10888 ( .A(n9727), .ZN(n9729) );
  OAI211_X1 U10889 ( .C1(n9799), .C2(n9730), .A(n9729), .B(n9728), .ZN(
        P1_U3256) );
  INV_X1 U10890 ( .A(n9731), .ZN(n9742) );
  AOI21_X1 U10891 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  NAND2_X1 U10892 ( .A1(n9784), .A2(n9735), .ZN(n9741) );
  AOI21_X1 U10893 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(n9739) );
  NAND2_X1 U10894 ( .A1(n9788), .A2(n9739), .ZN(n9740) );
  OAI211_X1 U10895 ( .C1(n9795), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9743)
         );
  INV_X1 U10896 ( .A(n9743), .ZN(n9745) );
  OAI211_X1 U10897 ( .C1(n9799), .C2(n10069), .A(n9745), .B(n9744), .ZN(
        P1_U3257) );
  INV_X1 U10898 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9757) );
  AOI211_X1 U10899 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n9764), .ZN(n9753)
         );
  AOI211_X1 U10900 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9758), .ZN(n9752)
         );
  AOI211_X1 U10901 ( .C1(n9777), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9756)
         );
  OAI211_X1 U10902 ( .C1(n9799), .C2(n9757), .A(n9756), .B(n9755), .ZN(
        P1_U3258) );
  AOI21_X1 U10903 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9768) );
  XNOR2_X1 U10904 ( .A(n9762), .B(n9761), .ZN(n9765) );
  OAI22_X1 U10905 ( .A1(n9765), .A2(n9764), .B1(n9763), .B2(n9795), .ZN(n9766)
         );
  AOI21_X1 U10906 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(n9770) );
  OAI211_X1 U10907 ( .C1(n9799), .C2(n9771), .A(n9770), .B(n9769), .ZN(
        P1_U3259) );
  INV_X1 U10908 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9783) );
  OAI21_X1 U10909 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9780) );
  XNOR2_X1 U10910 ( .A(n9776), .B(n9775), .ZN(n9779) );
  AOI222_X1 U10911 ( .A1(n9780), .A2(n9784), .B1(n9788), .B2(n9779), .C1(n9778), .C2(n9777), .ZN(n9782) );
  OAI211_X1 U10912 ( .C1(n9799), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P1_U3260) );
  OAI211_X1 U10913 ( .C1(n9787), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9793)
         );
  OAI211_X1 U10914 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9792)
         );
  OAI211_X1 U10915 ( .C1(n9795), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9796)
         );
  INV_X1 U10916 ( .A(n9796), .ZN(n9798) );
  OAI211_X1 U10917 ( .C1(n9799), .C2(n9964), .A(n9798), .B(n9797), .ZN(
        P1_U3261) );
  AOI22_X1 U10918 ( .A1(n9813), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9801), .B2(
        n9800), .ZN(n9805) );
  NAND2_X1 U10919 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  OAI211_X1 U10920 ( .C1(n9807), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9808)
         );
  AOI21_X1 U10921 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9811) );
  OAI21_X1 U10922 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(P1_U3287) );
  AND2_X1 U10923 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9815), .ZN(P1_U3294) );
  INV_X1 U10924 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U10925 ( .A1(n9814), .A2(n10044), .ZN(P1_U3295) );
  AND2_X1 U10926 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9815), .ZN(P1_U3296) );
  AND2_X1 U10927 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9815), .ZN(P1_U3297) );
  AND2_X1 U10928 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9815), .ZN(P1_U3298) );
  AND2_X1 U10929 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9815), .ZN(P1_U3299) );
  AND2_X1 U10930 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9815), .ZN(P1_U3300) );
  AND2_X1 U10931 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9815), .ZN(P1_U3301) );
  INV_X1 U10932 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U10933 ( .A1(n9814), .A2(n10047), .ZN(P1_U3302) );
  AND2_X1 U10934 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9815), .ZN(P1_U3303) );
  AND2_X1 U10935 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9815), .ZN(P1_U3304) );
  AND2_X1 U10936 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9815), .ZN(P1_U3305) );
  AND2_X1 U10937 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9815), .ZN(P1_U3306) );
  AND2_X1 U10938 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9815), .ZN(P1_U3307) );
  AND2_X1 U10939 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9815), .ZN(P1_U3308) );
  AND2_X1 U10940 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9815), .ZN(P1_U3309) );
  INV_X1 U10941 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U10942 ( .A1(n9814), .A2(n10052), .ZN(P1_U3310) );
  AND2_X1 U10943 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9815), .ZN(P1_U3311) );
  AND2_X1 U10944 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9815), .ZN(P1_U3312) );
  AND2_X1 U10945 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9815), .ZN(P1_U3313) );
  INV_X1 U10946 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10111) );
  NOR2_X1 U10947 ( .A1(n9814), .A2(n10111), .ZN(P1_U3314) );
  AND2_X1 U10948 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9815), .ZN(P1_U3315) );
  AND2_X1 U10949 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9815), .ZN(P1_U3316) );
  AND2_X1 U10950 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9815), .ZN(P1_U3317) );
  AND2_X1 U10951 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9815), .ZN(P1_U3318) );
  AND2_X1 U10952 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9815), .ZN(P1_U3319) );
  AND2_X1 U10953 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9815), .ZN(P1_U3320) );
  INV_X1 U10954 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U10955 ( .A1(n9814), .A2(n10017), .ZN(P1_U3321) );
  AND2_X1 U10956 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9815), .ZN(P1_U3322) );
  AND2_X1 U10957 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9815), .ZN(P1_U3323) );
  OAI21_X1 U10958 ( .B1(n9817), .B2(n9831), .A(n9816), .ZN(n9819) );
  AOI211_X1 U10959 ( .C1(n9835), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9848)
         );
  INV_X1 U10960 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U10961 ( .A1(n9627), .A2(n9848), .B1(n9821), .B2(n9846), .ZN(
        P1_U3468) );
  NAND2_X1 U10962 ( .A1(n9822), .A2(n9842), .ZN(n9824) );
  OAI211_X1 U10963 ( .C1(n9825), .C2(n9831), .A(n9824), .B(n9823), .ZN(n9826)
         );
  NOR2_X1 U10964 ( .A1(n9827), .A2(n9826), .ZN(n9850) );
  INV_X1 U10965 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10966 ( .A1(n9627), .A2(n9850), .B1(n9828), .B2(n9846), .ZN(
        P1_U3474) );
  OAI211_X1 U10967 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  AOI21_X1 U10968 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9852) );
  INV_X1 U10969 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10970 ( .A1(n9627), .A2(n9852), .B1(n9836), .B2(n9846), .ZN(
        P1_U3480) );
  NAND2_X1 U10971 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  NAND2_X1 U10972 ( .A1(n9840), .A2(n9839), .ZN(n9841) );
  AOI21_X1 U10973 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  AND2_X1 U10974 ( .A1(n9845), .A2(n9844), .ZN(n9853) );
  INV_X1 U10975 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10976 ( .A1(n9627), .A2(n9853), .B1(n9847), .B2(n9846), .ZN(
        P1_U3486) );
  AOI22_X1 U10977 ( .A1(n9854), .A2(n9848), .B1(n6604), .B2(n5802), .ZN(
        P1_U3527) );
  AOI22_X1 U10978 ( .A1(n9854), .A2(n9850), .B1(n9849), .B2(n5802), .ZN(
        P1_U3529) );
  INV_X1 U10979 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10980 ( .A1(n9854), .A2(n9852), .B1(n9851), .B2(n5802), .ZN(
        P1_U3531) );
  AOI22_X1 U10981 ( .A1(n9854), .A2(n9853), .B1(n9303), .B2(n5802), .ZN(
        P1_U3533) );
  INV_X1 U10982 ( .A(n9855), .ZN(n9860) );
  INV_X1 U10983 ( .A(n6415), .ZN(n9858) );
  INV_X1 U10984 ( .A(n9930), .ZN(n9889) );
  NAND2_X1 U10985 ( .A1(n9861), .A2(n9889), .ZN(n9857) );
  AOI22_X1 U10986 ( .A1(n5910), .A2(n9872), .B1(n9940), .B2(n5883), .ZN(n9856)
         );
  OAI211_X1 U10987 ( .C1(n9858), .C2(n9917), .A(n9857), .B(n9856), .ZN(n9859)
         );
  AOI211_X1 U10988 ( .C1(n9928), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9944)
         );
  AOI22_X1 U10989 ( .A1(n9943), .A2(n5872), .B1(n9944), .B2(n9941), .ZN(
        P2_U3393) );
  INV_X1 U10990 ( .A(n9867), .ZN(n9870) );
  AOI22_X1 U10991 ( .A1(n9863), .A2(n9874), .B1(n9862), .B2(n9940), .ZN(n9864)
         );
  OAI211_X1 U10992 ( .C1(n5927), .C2(n9919), .A(n9865), .B(n9864), .ZN(n9869)
         );
  NOR2_X1 U10993 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  AOI211_X1 U10994 ( .C1(n9870), .C2(n9889), .A(n9869), .B(n9868), .ZN(n9946)
         );
  AOI22_X1 U10995 ( .A1(n9943), .A2(n5896), .B1(n9946), .B2(n9941), .ZN(
        P2_U3396) );
  INV_X1 U10996 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U10997 ( .A1(n9871), .A2(n9902), .ZN(n9876) );
  AOI22_X1 U10998 ( .A1(n9874), .A2(n5910), .B1(n9873), .B2(n9872), .ZN(n9875)
         );
  OAI211_X1 U10999 ( .C1(n9877), .C2(n9886), .A(n9876), .B(n9875), .ZN(n9878)
         );
  AOI21_X1 U11000 ( .B1(n9879), .B2(n9884), .A(n9878), .ZN(n9947) );
  AOI22_X1 U11001 ( .A1(n9943), .A2(n9880), .B1(n9947), .B2(n9941), .ZN(
        P2_U3399) );
  OAI21_X1 U11002 ( .B1(n9882), .B2(n9886), .A(n9881), .ZN(n9883) );
  AOI21_X1 U11003 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9948) );
  AOI22_X1 U11004 ( .A1(n9943), .A2(n5931), .B1(n9948), .B2(n9941), .ZN(
        P2_U3402) );
  INV_X1 U11005 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9893) );
  NOR2_X1 U11006 ( .A1(n9887), .A2(n9886), .ZN(n9888) );
  AOI21_X1 U11007 ( .B1(n9890), .B2(n9889), .A(n9888), .ZN(n9891) );
  AND2_X1 U11008 ( .A1(n9892), .A2(n9891), .ZN(n9949) );
  AOI22_X1 U11009 ( .A1(n9943), .A2(n9893), .B1(n9949), .B2(n9941), .ZN(
        P2_U3405) );
  INV_X1 U11010 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9903) );
  OAI22_X1 U11011 ( .A1(n9895), .A2(n9919), .B1(n9894), .B2(n9917), .ZN(n9896)
         );
  AOI21_X1 U11012 ( .B1(n9940), .B2(n9897), .A(n9896), .ZN(n9898) );
  OAI21_X1 U11013 ( .B1(n9899), .B2(n9935), .A(n9898), .ZN(n9900) );
  AOI21_X1 U11014 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(n9950) );
  AOI22_X1 U11015 ( .A1(n9943), .A2(n9903), .B1(n9950), .B2(n9941), .ZN(
        P2_U3408) );
  INV_X1 U11016 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9912) );
  OAI22_X1 U11017 ( .A1(n9904), .A2(n9917), .B1(n9918), .B2(n9919), .ZN(n9905)
         );
  AOI21_X1 U11018 ( .B1(n9940), .B2(n9906), .A(n9905), .ZN(n9907) );
  OAI21_X1 U11019 ( .B1(n9908), .B2(n9930), .A(n9907), .ZN(n9909) );
  AOI211_X1 U11020 ( .C1(n9928), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9951)
         );
  AOI22_X1 U11021 ( .A1(n9943), .A2(n9912), .B1(n9951), .B2(n9941), .ZN(
        P2_U3411) );
  NOR2_X1 U11022 ( .A1(n9913), .A2(n9935), .ZN(n9914) );
  AOI211_X1 U11023 ( .C1(n9940), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9952)
         );
  AOI22_X1 U11024 ( .A1(n9943), .A2(n5987), .B1(n9952), .B2(n9941), .ZN(
        P2_U3414) );
  INV_X1 U11025 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9929) );
  OAI22_X1 U11026 ( .A1(n9920), .A2(n9919), .B1(n9918), .B2(n9917), .ZN(n9921)
         );
  AOI21_X1 U11027 ( .B1(n9940), .B2(n9922), .A(n9921), .ZN(n9923) );
  OAI21_X1 U11028 ( .B1(n9924), .B2(n9930), .A(n9923), .ZN(n9926) );
  AOI211_X1 U11029 ( .C1(n9928), .C2(n9927), .A(n9926), .B(n9925), .ZN(n9953)
         );
  AOI22_X1 U11030 ( .A1(n9943), .A2(n9929), .B1(n9953), .B2(n9941), .ZN(
        P2_U3417) );
  NOR2_X1 U11031 ( .A1(n9931), .A2(n9930), .ZN(n9933) );
  AOI211_X1 U11032 ( .C1(n9940), .C2(n9934), .A(n9933), .B(n9932), .ZN(n9954)
         );
  AOI22_X1 U11033 ( .A1(n9943), .A2(n6014), .B1(n9954), .B2(n9941), .ZN(
        P2_U3420) );
  INV_X1 U11034 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U11035 ( .A1(n9936), .A2(n9935), .ZN(n9938) );
  AOI211_X1 U11036 ( .C1(n9940), .C2(n9939), .A(n9938), .B(n9937), .ZN(n9955)
         );
  AOI22_X1 U11037 ( .A1(n9943), .A2(n9942), .B1(n9955), .B2(n9941), .ZN(
        P2_U3423) );
  AOI22_X1 U11038 ( .A1(n9956), .A2(n9944), .B1(n6429), .B2(n4414), .ZN(
        P2_U3460) );
  INV_X1 U11039 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9945) );
  AOI22_X1 U11040 ( .A1(n9956), .A2(n9946), .B1(n9945), .B2(n4414), .ZN(
        P2_U3461) );
  AOI22_X1 U11041 ( .A1(n9956), .A2(n9947), .B1(n5914), .B2(n4414), .ZN(
        P2_U3462) );
  AOI22_X1 U11042 ( .A1(n9956), .A2(n9948), .B1(n5933), .B2(n4414), .ZN(
        P2_U3463) );
  AOI22_X1 U11043 ( .A1(n9956), .A2(n9949), .B1(n6663), .B2(n4414), .ZN(
        P2_U3464) );
  AOI22_X1 U11044 ( .A1(n9956), .A2(n9950), .B1(n6662), .B2(n4414), .ZN(
        P2_U3465) );
  AOI22_X1 U11045 ( .A1(n9956), .A2(n9951), .B1(n6655), .B2(n4414), .ZN(
        P2_U3466) );
  AOI22_X1 U11046 ( .A1(n9956), .A2(n9952), .B1(n6715), .B2(n4414), .ZN(
        P2_U3467) );
  AOI22_X1 U11047 ( .A1(n9956), .A2(n9953), .B1(n6859), .B2(n4414), .ZN(
        P2_U3468) );
  AOI22_X1 U11048 ( .A1(n9956), .A2(n9954), .B1(n6993), .B2(n4414), .ZN(
        P2_U3469) );
  AOI22_X1 U11049 ( .A1(n9956), .A2(n9955), .B1(n7159), .B2(n4414), .ZN(
        P2_U3470) );
  OAI222_X1 U11050 ( .A1(n9961), .A2(n9960), .B1(n9961), .B2(n9959), .C1(n9958), .C2(n9957), .ZN(ADD_1068_U5) );
  XOR2_X1 U11051 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11052 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  XOR2_X1 U11053 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n9965), .Z(ADD_1068_U55) );
  OAI21_X1 U11054 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(ADD_1068_U56) );
  OAI21_X1 U11055 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(ADD_1068_U57) );
  OAI21_X1 U11056 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(ADD_1068_U58) );
  OAI21_X1 U11057 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(ADD_1068_U59) );
  OAI21_X1 U11058 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(ADD_1068_U60) );
  OAI21_X1 U11059 ( .B1(n9983), .B2(n9982), .A(n9981), .ZN(ADD_1068_U61) );
  OAI21_X1 U11060 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(ADD_1068_U62) );
  OAI21_X1 U11061 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(ADD_1068_U63) );
  MUX2_X1 U11062 ( .A(n9991), .B(n9990), .S(P2_U3893), .Z(n10149) );
  INV_X1 U11063 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11064 ( .A1(n10121), .A2(keyinput50), .B1(n9993), .B2(keyinput28), 
        .ZN(n9992) );
  OAI221_X1 U11065 ( .B1(n10121), .B2(keyinput50), .C1(n9993), .C2(keyinput28), 
        .A(n9992), .ZN(n10003) );
  AOI22_X1 U11066 ( .A1(n10129), .A2(keyinput29), .B1(n10131), .B2(keyinput48), 
        .ZN(n9994) );
  OAI221_X1 U11067 ( .B1(n10129), .B2(keyinput29), .C1(n10131), .C2(keyinput48), .A(n9994), .ZN(n10002) );
  AOI22_X1 U11068 ( .A1(n9997), .A2(keyinput51), .B1(n9996), .B2(keyinput19), 
        .ZN(n9995) );
  OAI221_X1 U11069 ( .B1(n9997), .B2(keyinput51), .C1(n9996), .C2(keyinput19), 
        .A(n9995), .ZN(n10001) );
  AOI22_X1 U11070 ( .A1(n9999), .A2(keyinput3), .B1(keyinput61), .B2(n10130), 
        .ZN(n9998) );
  OAI221_X1 U11071 ( .B1(n9999), .B2(keyinput3), .C1(n10130), .C2(keyinput61), 
        .A(n9998), .ZN(n10000) );
  NOR4_X1 U11072 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10042) );
  AOI22_X1 U11073 ( .A1(n10006), .A2(keyinput24), .B1(n10005), .B2(keyinput47), 
        .ZN(n10004) );
  OAI221_X1 U11074 ( .B1(n10006), .B2(keyinput24), .C1(n10005), .C2(keyinput47), .A(n10004), .ZN(n10014) );
  AOI22_X1 U11075 ( .A1(n10119), .A2(keyinput54), .B1(n10120), .B2(keyinput0), 
        .ZN(n10007) );
  OAI221_X1 U11076 ( .B1(n10119), .B2(keyinput54), .C1(n10120), .C2(keyinput0), 
        .A(n10007), .ZN(n10013) );
  INV_X1 U11077 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U11078 ( .A1(n10126), .A2(keyinput5), .B1(n10128), .B2(keyinput18), 
        .ZN(n10008) );
  OAI221_X1 U11079 ( .B1(n10126), .B2(keyinput5), .C1(n10128), .C2(keyinput18), 
        .A(n10008), .ZN(n10012) );
  INV_X1 U11080 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10127) );
  INV_X1 U11081 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11082 ( .A1(n10127), .A2(keyinput13), .B1(n10010), .B2(keyinput49), 
        .ZN(n10009) );
  OAI221_X1 U11083 ( .B1(n10127), .B2(keyinput13), .C1(n10010), .C2(keyinput49), .A(n10009), .ZN(n10011) );
  NOR4_X1 U11084 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10041) );
  AOI22_X1 U11085 ( .A1(n10104), .A2(keyinput62), .B1(keyinput25), .B2(n7551), 
        .ZN(n10015) );
  OAI221_X1 U11086 ( .B1(n10104), .B2(keyinput62), .C1(n7551), .C2(keyinput25), 
        .A(n10015), .ZN(n10026) );
  AOI22_X1 U11087 ( .A1(n10018), .A2(keyinput12), .B1(n10017), .B2(keyinput36), 
        .ZN(n10016) );
  OAI221_X1 U11088 ( .B1(n10018), .B2(keyinput12), .C1(n10017), .C2(keyinput36), .A(n10016), .ZN(n10025) );
  AOI22_X1 U11089 ( .A1(n10114), .A2(keyinput10), .B1(keyinput42), .B2(n10020), 
        .ZN(n10019) );
  OAI221_X1 U11090 ( .B1(n10114), .B2(keyinput10), .C1(n10020), .C2(keyinput42), .A(n10019), .ZN(n10024) );
  XNOR2_X1 U11091 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput11), .ZN(n10022) );
  XNOR2_X1 U11092 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput27), .ZN(n10021)
         );
  NAND2_X1 U11093 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  NOR4_X1 U11094 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10040) );
  INV_X1 U11095 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11096 ( .A1(n10028), .A2(keyinput4), .B1(n10103), .B2(keyinput43), 
        .ZN(n10027) );
  OAI221_X1 U11097 ( .B1(n10028), .B2(keyinput4), .C1(n10103), .C2(keyinput43), 
        .A(n10027), .ZN(n10032) );
  XOR2_X1 U11098 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput58), .Z(n10031) );
  INV_X1 U11099 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10029) );
  XNOR2_X1 U11100 ( .A(keyinput41), .B(n10029), .ZN(n10030) );
  NOR3_X1 U11101 ( .A1(n10032), .A2(n10031), .A3(n10030), .ZN(n10036) );
  XOR2_X1 U11102 ( .A(n5896), .B(keyinput21), .Z(n10035) );
  XNOR2_X1 U11103 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput2), .ZN(n10034) );
  XNOR2_X1 U11104 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput45), .ZN(n10033)
         );
  NAND4_X1 U11105 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10038) );
  XNOR2_X1 U11106 ( .A(n10109), .B(keyinput14), .ZN(n10037) );
  NOR2_X1 U11107 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NAND4_X1 U11108 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10100) );
  INV_X1 U11109 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11110 ( .A1(n10044), .A2(keyinput1), .B1(keyinput44), .B2(n10101), 
        .ZN(n10043) );
  OAI221_X1 U11111 ( .B1(n10044), .B2(keyinput1), .C1(n10101), .C2(keyinput44), 
        .A(n10043), .ZN(n10051) );
  AOI22_X1 U11112 ( .A1(n10047), .A2(keyinput52), .B1(keyinput33), .B2(n10046), 
        .ZN(n10045) );
  OAI221_X1 U11113 ( .B1(n10047), .B2(keyinput52), .C1(n10046), .C2(keyinput33), .A(n10045), .ZN(n10050) );
  XOR2_X1 U11114 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput15), .Z(n10049) );
  XNOR2_X1 U11115 ( .A(n10102), .B(keyinput53), .ZN(n10048) );
  OR4_X1 U11116 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10055) );
  XNOR2_X1 U11117 ( .A(n10111), .B(keyinput60), .ZN(n10054) );
  XNOR2_X1 U11118 ( .A(n10052), .B(keyinput22), .ZN(n10053) );
  NOR3_X1 U11119 ( .A1(n10055), .A2(n10054), .A3(n10053), .ZN(n10098) );
  INV_X1 U11120 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U11121 ( .A1(n10058), .A2(keyinput37), .B1(n10057), .B2(keyinput7), 
        .ZN(n10056) );
  OAI221_X1 U11122 ( .B1(n10058), .B2(keyinput37), .C1(n10057), .C2(keyinput7), 
        .A(n10056), .ZN(n10067) );
  INV_X1 U11123 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11124 ( .A1(n10133), .A2(keyinput20), .B1(keyinput38), .B2(n6663), 
        .ZN(n10059) );
  OAI221_X1 U11125 ( .B1(n10133), .B2(keyinput20), .C1(n6663), .C2(keyinput38), 
        .A(n10059), .ZN(n10066) );
  INV_X1 U11126 ( .A(SI_18_), .ZN(n10061) );
  AOI22_X1 U11127 ( .A1(n10132), .A2(keyinput23), .B1(n10061), .B2(keyinput26), 
        .ZN(n10060) );
  OAI221_X1 U11128 ( .B1(n10132), .B2(keyinput23), .C1(n10061), .C2(keyinput26), .A(n10060), .ZN(n10065) );
  XNOR2_X1 U11129 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput31), .ZN(n10063) );
  XNOR2_X1 U11130 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput8), .ZN(n10062) );
  NAND2_X1 U11131 ( .A1(n10063), .A2(n10062), .ZN(n10064) );
  NOR4_X1 U11132 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n10097) );
  AOI22_X1 U11133 ( .A1(n10069), .A2(keyinput46), .B1(n10115), .B2(keyinput56), 
        .ZN(n10068) );
  OAI221_X1 U11134 ( .B1(n10069), .B2(keyinput46), .C1(n10115), .C2(keyinput56), .A(n10068), .ZN(n10080) );
  AOI22_X1 U11135 ( .A1(n8761), .A2(keyinput57), .B1(n10071), .B2(keyinput63), 
        .ZN(n10070) );
  OAI221_X1 U11136 ( .B1(n8761), .B2(keyinput57), .C1(n10071), .C2(keyinput63), 
        .A(n10070), .ZN(n10079) );
  AOI22_X1 U11137 ( .A1(n10074), .A2(keyinput59), .B1(n10073), .B2(keyinput17), 
        .ZN(n10072) );
  OAI221_X1 U11138 ( .B1(n10074), .B2(keyinput59), .C1(n10073), .C2(keyinput17), .A(n10072), .ZN(n10078) );
  AOI22_X1 U11139 ( .A1(n10076), .A2(keyinput40), .B1(keyinput16), .B2(n10124), 
        .ZN(n10075) );
  OAI221_X1 U11140 ( .B1(n10076), .B2(keyinput40), .C1(n10124), .C2(keyinput16), .A(n10075), .ZN(n10077) );
  NOR4_X1 U11141 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10096) );
  INV_X1 U11142 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11143 ( .A1(n10083), .A2(keyinput35), .B1(n10082), .B2(keyinput55), 
        .ZN(n10081) );
  OAI221_X1 U11144 ( .B1(n10083), .B2(keyinput35), .C1(n10082), .C2(keyinput55), .A(n10081), .ZN(n10094) );
  INV_X1 U11145 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10086) );
  INV_X1 U11146 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11147 ( .A1(n10086), .A2(keyinput39), .B1(keyinput9), .B2(n10085), 
        .ZN(n10084) );
  OAI221_X1 U11148 ( .B1(n10086), .B2(keyinput39), .C1(n10085), .C2(keyinput9), 
        .A(n10084), .ZN(n10093) );
  AOI22_X1 U11149 ( .A1(n10113), .A2(keyinput34), .B1(n10088), .B2(keyinput30), 
        .ZN(n10087) );
  OAI221_X1 U11150 ( .B1(n10113), .B2(keyinput34), .C1(n10088), .C2(keyinput30), .A(n10087), .ZN(n10092) );
  XOR2_X1 U11151 ( .A(n5906), .B(keyinput6), .Z(n10090) );
  XNOR2_X1 U11152 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput32), .ZN(n10089) );
  NAND2_X1 U11153 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  NOR4_X1 U11154 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n10091), .ZN(
        n10095) );
  NAND4_X1 U11155 ( .A1(n10098), .A2(n10097), .A3(n10096), .A4(n10095), .ZN(
        n10099) );
  NOR2_X1 U11156 ( .A1(n10100), .A2(n10099), .ZN(n10147) );
  AND4_X1 U11157 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(P2_DATAO_REG_4__SCAN_IN), 
        .A3(n10101), .A4(n5896), .ZN(n10112) );
  NAND4_X1 U11158 ( .A1(n10102), .A2(P1_REG1_REG_19__SCAN_IN), .A3(
        P1_REG2_REG_26__SCAN_IN), .A4(P1_REG1_REG_2__SCAN_IN), .ZN(n10108) );
  AND4_X1 U11159 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P2_REG2_REG_13__SCAN_IN), 
        .A3(n10104), .A4(n10103), .ZN(n10105) );
  NAND3_X1 U11160 ( .A1(n10106), .A2(P1_D_REG_23__SCAN_IN), .A3(n10105), .ZN(
        n10107) );
  NOR2_X1 U11161 ( .A1(n10108), .A2(n10107), .ZN(n10110) );
  AND4_X1 U11162 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10145) );
  NOR4_X1 U11163 ( .A1(SI_17_), .A2(P1_REG2_REG_29__SCAN_IN), .A3(
        P1_REG0_REG_13__SCAN_IN), .A4(n10113), .ZN(n10144) );
  NAND4_X1 U11164 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), 
        .A3(P1_DATAO_REG_8__SCAN_IN), .A4(n10114), .ZN(n10118) );
  NAND4_X1 U11165 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_DATAO_REG_27__SCAN_IN), 
        .A3(P2_DATAO_REG_9__SCAN_IN), .A4(P2_REG2_REG_23__SCAN_IN), .ZN(n10117) );
  NAND4_X1 U11166 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(P2_REG0_REG_16__SCAN_IN), .A3(P1_ADDR_REG_14__SCAN_IN), .A4(n10115), .ZN(n10116) );
  NOR3_X1 U11167 ( .A1(n10118), .A2(n10117), .A3(n10116), .ZN(n10143) );
  NAND4_X1 U11168 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .A3(P2_REG3_REG_22__SCAN_IN), .A4(P2_REG3_REG_19__SCAN_IN), .ZN(n10141) );
  NAND4_X1 U11169 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_15__SCAN_IN), .A3(n10120), .A4(n10119), .ZN(n10140) );
  NAND3_X1 U11170 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), 
        .A3(n10121), .ZN(n10122) );
  NOR3_X1 U11171 ( .A1(n10122), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n10123) );
  NAND3_X1 U11172 ( .A1(n10125), .A2(n10124), .A3(n10123), .ZN(n10139) );
  NOR4_X1 U11173 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(n10128), .A3(n10127), 
        .A4(n10126), .ZN(n10137) );
  NOR4_X1 U11174 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(n10131), .A3(n10130), 
        .A4(n10129), .ZN(n10136) );
  NOR4_X1 U11175 ( .A1(SI_18_), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_REG1_REG_18__SCAN_IN), .A4(n10132), .ZN(n10135) );
  NOR4_X1 U11176 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(P1_REG2_REG_9__SCAN_IN), 
        .A3(n10133), .A4(n6663), .ZN(n10134) );
  NAND4_X1 U11177 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NOR4_X1 U11178 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10142) );
  NAND4_X1 U11179 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10146) );
  XNOR2_X1 U11180 ( .A(n10147), .B(n10146), .ZN(n10148) );
  XNOR2_X1 U11181 ( .A(n10149), .B(n10148), .ZN(P2_U3520) );
  OAI21_X1 U11182 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(ADD_1068_U50) );
  OAI21_X1 U11183 ( .B1(n10155), .B2(n10154), .A(n10153), .ZN(ADD_1068_U51) );
  OAI21_X1 U11184 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(ADD_1068_U47) );
  OAI21_X1 U11185 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(ADD_1068_U49) );
  OAI21_X1 U11186 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(ADD_1068_U48) );
  AOI21_X1 U11187 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(ADD_1068_U54) );
  AOI21_X1 U11188 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(ADD_1068_U53) );
  OAI21_X1 U11189 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4795 ( .A(n8672), .Z(n4274) );
endmodule

