

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748;

  INV_X2 U3697 ( .A(n6697), .ZN(n3783) );
  AND2_X1 U3698 ( .A1(n4242), .A2(n3899), .ZN(n4234) );
  CLKBUF_X2 U3699 ( .A(n4610), .Z(n4587) );
  CLKBUF_X1 U3700 ( .A(n3925), .Z(n4778) );
  CLKBUF_X2 U3701 ( .A(n3987), .Z(n4711) );
  CLKBUF_X2 U3702 ( .A(n4022), .Z(n4785) );
  CLKBUF_X2 U3703 ( .A(n3677), .Z(n3992) );
  CLKBUF_X2 U3704 ( .A(n3703), .Z(n4710) );
  CLKBUF_X1 U3705 ( .A(n4784), .Z(n4751) );
  CLKBUF_X2 U3706 ( .A(n3673), .Z(n4757) );
  CLKBUF_X1 U3707 ( .A(n3710), .Z(n5050) );
  CLKBUF_X2 U3708 ( .A(n3939), .Z(n3698) );
  CLKBUF_X1 U3709 ( .A(n3700), .Z(n3673) );
  AND2_X2 U3710 ( .A1(n5123), .A2(n4912), .ZN(n4411) );
  NAND2_X1 U3711 ( .A1(n5093), .A2(n4299), .ZN(n3969) );
  AND4_X1 U3712 ( .A1(n3857), .A2(n3859), .A3(n3858), .A4(n3860), .ZN(n3715)
         );
  AND4_X1 U3713 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  INV_X1 U3714 ( .A(n6029), .ZN(n6058) );
  NOR2_X1 U3715 ( .A1(n5721), .A2(n5206), .ZN(n6103) );
  INV_X1 U3716 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7522) );
  INV_X1 U3717 ( .A(n7304), .ZN(n4065) );
  OR2_X1 U3718 ( .A1(n4064), .A2(n4063), .ZN(n4308) );
  INV_X1 U3719 ( .A(n7475), .ZN(n7420) );
  NAND2_X2 U3720 ( .A1(n3741), .A2(n3739), .ZN(n5642) );
  AOI21_X2 U3721 ( .B1(n5805), .B2(n5804), .A(n3717), .ZN(n5934) );
  OAI22_X2 U3722 ( .A1(n5630), .A2(n5629), .B1(n4177), .B2(n5337), .ZN(n5805)
         );
  INV_X1 U3723 ( .A(n4332), .ZN(n3663) );
  INV_X1 U3724 ( .A(n3663), .ZN(n3664) );
  NAND3_X1 U3725 ( .A1(n3754), .A2(n3755), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U3726 ( .A1(n3683), .A2(n4357), .ZN(n5521) );
  CLKBUF_X2 U3727 ( .A(n5157), .Z(n3706) );
  NAND2_X1 U3728 ( .A1(n5147), .A2(n4085), .ZN(n5129) );
  CLKBUF_X2 U3729 ( .A(n5042), .Z(n5065) );
  INV_X2 U3730 ( .A(n5721), .ZN(n3971) );
  NAND2_X2 U3731 ( .A1(n5225), .A2(n5165), .ZN(n4865) );
  INV_X1 U3732 ( .A(n3671), .ZN(n4295) );
  INV_X2 U3733 ( .A(n3710), .ZN(n3899) );
  AND4_X1 U3734 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  CLKBUF_X2 U3735 ( .A(n3939), .Z(n3697) );
  CLKBUF_X1 U3736 ( .A(n4114), .Z(n3695) );
  CLKBUF_X1 U3737 ( .A(n4114), .Z(n3696) );
  INV_X1 U3738 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3676) );
  NOR2_X4 U3739 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3839) );
  NOR2_X1 U3740 ( .A1(n4810), .A2(n4809), .ZN(n4811) );
  OAI21_X1 U3741 ( .B1(n6406), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n6407), 
        .ZN(n6609) );
  INV_X1 U3742 ( .A(n6412), .ZN(n6369) );
  AOI211_X1 U3743 ( .C1(n6513), .C2(n6429), .A(n6428), .B(n6427), .ZN(n6430)
         );
  AOI211_X1 U3744 ( .C1(n6513), .C2(n6422), .A(n6421), .B(n6420), .ZN(n6423)
         );
  AND2_X1 U3745 ( .A1(n6144), .A2(n4817), .ZN(n6412) );
  OR2_X1 U3746 ( .A1(n6142), .A2(n6156), .ZN(n6419) );
  OR2_X1 U3747 ( .A1(n6221), .A2(n6220), .ZN(n6482) );
  AOI21_X1 U3748 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3783), .A(n6471), 
        .ZN(n6464) );
  AND2_X1 U3749 ( .A1(n3687), .A2(n3790), .ZN(n6399) );
  NAND2_X1 U3750 ( .A1(n3810), .A2(n4563), .ZN(n6330) );
  NOR2_X2 U3751 ( .A1(n6329), .A2(n3808), .ZN(n6207) );
  NAND2_X1 U3752 ( .A1(n6457), .A2(n4224), .ZN(n6441) );
  AND2_X1 U3753 ( .A1(n3784), .A2(n3786), .ZN(n6493) );
  NAND2_X1 U3754 ( .A1(n3787), .A2(n3785), .ZN(n6457) );
  AND2_X1 U3755 ( .A1(n5915), .A2(n5958), .ZN(n5977) );
  NOR2_X1 U3756 ( .A1(n3813), .A2(n5521), .ZN(n5915) );
  NAND2_X1 U3757 ( .A1(n3776), .A2(n3716), .ZN(n3775) );
  OR2_X1 U3758 ( .A1(n3779), .A2(n3778), .ZN(n3776) );
  NOR2_X1 U3759 ( .A1(n4221), .A2(n3751), .ZN(n3750) );
  NOR2_X2 U3760 ( .A1(n5155), .A2(n5334), .ZN(n3683) );
  OR2_X1 U3761 ( .A1(n5557), .A2(n3727), .ZN(n3813) );
  INV_X1 U3762 ( .A(n4358), .ZN(n4365) );
  OAI21_X1 U3763 ( .B1(n4339), .B2(n4470), .A(n4338), .ZN(n5156) );
  AOI21_X1 U3764 ( .B1(n4347), .B2(n4480), .A(n4346), .ZN(n5334) );
  XNOR2_X1 U3765 ( .A(n4212), .B(n4205), .ZN(n4358) );
  AOI21_X1 U3766 ( .B1(n3833), .B2(n4480), .A(n4356), .ZN(n5522) );
  OAI21_X1 U3767 ( .B1(n4339), .B2(n4210), .A(n4160), .ZN(n4162) );
  NAND2_X1 U3768 ( .A1(n4194), .A2(n4190), .ZN(n4212) );
  OR2_X1 U3769 ( .A1(n4194), .A2(n4193), .ZN(n3833) );
  NAND2_X1 U3770 ( .A1(n4300), .A2(n4498), .ZN(n5077) );
  NAND2_X1 U3771 ( .A1(n4151), .A2(n4152), .ZN(n4179) );
  AND2_X1 U3772 ( .A1(n4138), .A2(n4137), .ZN(n4151) );
  XNOR2_X1 U3773 ( .A(n4137), .B(n4136), .ZN(n4332) );
  XNOR2_X1 U3774 ( .A(n4128), .B(n4127), .ZN(n5157) );
  NAND2_X1 U3775 ( .A1(n4100), .A2(n4099), .ZN(n4128) );
  NAND2_X2 U3776 ( .A1(n3796), .A2(n3801), .ZN(n5854) );
  AND2_X1 U3777 ( .A1(n4940), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4954)
         );
  INV_X1 U3778 ( .A(n5129), .ZN(n3665) );
  NAND2_X1 U3780 ( .A1(n4074), .A2(n4073), .ZN(n4076) );
  NAND2_X2 U3781 ( .A1(n6391), .A2(n5057), .ZN(n7570) );
  CLKBUF_X1 U3782 ( .A(n4309), .Z(n4310) );
  NAND2_X2 U3783 ( .A1(n6352), .A2(n5219), .ZN(n6355) );
  AOI21_X1 U3784 ( .B1(n4107), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4081), 
        .ZN(n4083) );
  CLKBUF_X1 U3785 ( .A(n4077), .Z(n4107) );
  NAND2_X1 U3786 ( .A1(n3984), .A2(n4874), .ZN(n4053) );
  AND2_X1 U3787 ( .A1(n3981), .A2(n3980), .ZN(n3984) );
  OAI211_X1 U3788 ( .C1(n4853), .C2(n4042), .A(n4882), .B(n4971), .ZN(n4043)
         );
  AND3_X1 U3789 ( .A1(n4866), .A2(n4033), .A3(n4032), .ZN(n4858) );
  NAND2_X1 U3790 ( .A1(n6054), .A2(n6049), .ZN(n6114) );
  OR2_X1 U3791 ( .A1(n3976), .A2(n5214), .ZN(n4294) );
  AND2_X1 U3792 ( .A1(n6018), .A2(n5523), .ZN(n6029) );
  AND2_X1 U3793 ( .A1(n5721), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4242) );
  INV_X1 U3794 ( .A(n5170), .ZN(n4868) );
  OR2_X1 U3795 ( .A1(n3998), .A2(n3997), .ZN(n4213) );
  OR2_X1 U3796 ( .A1(n4011), .A2(n4010), .ZN(n4066) );
  AND2_X2 U3797 ( .A1(n5721), .A2(n5206), .ZN(n6018) );
  OR2_X2 U3798 ( .A1(n3897), .A2(n3896), .ZN(n5214) );
  CLKBUF_X1 U3799 ( .A(n4031), .Z(n5049) );
  AND2_X1 U3800 ( .A1(n3956), .A2(n3959), .ZN(n3732) );
  AND4_X1 U3801 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3957)
         );
  AND4_X1 U3802 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3935)
         );
  AND4_X1 U3803 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3958)
         );
  AND4_X1 U3804 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3937)
         );
  AND4_X1 U3805 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3936)
         );
  NAND2_X2 U3806 ( .A1(n3856), .A2(n3855), .ZN(n4302) );
  AND4_X1 U3807 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3886)
         );
  BUF_X2 U3808 ( .A(n4411), .Z(n4569) );
  AND4_X1 U3809 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3885)
         );
  AND4_X1 U3810 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  AND4_X1 U3811 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3959)
         );
  AND4_X1 U3812 ( .A1(n3867), .A2(n3868), .A3(n3866), .A4(n3865), .ZN(n3874)
         );
  AND4_X1 U3813 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3855)
         );
  AND4_X1 U3814 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3856)
         );
  AND4_X1 U3815 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3846)
         );
  NAND2_X2 U3816 ( .A1(n7569), .A2(n7562), .ZN(n7242) );
  NAND2_X2 U3817 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7569), .ZN(n7252) );
  BUF_X2 U3818 ( .A(n3999), .Z(n4779) );
  BUF_X2 U3819 ( .A(n4564), .Z(n4730) );
  CLKBUF_X3 U3820 ( .A(n3939), .Z(n4752) );
  AND2_X2 U3821 ( .A1(n3840), .A2(n4906), .ZN(n3705) );
  AND2_X2 U3822 ( .A1(n4912), .A2(n3774), .ZN(n4610) );
  BUF_X2 U3823 ( .A(n4582), .Z(n4611) );
  AND2_X1 U3824 ( .A1(n4912), .A2(n3839), .ZN(n3700) );
  AND2_X2 U3825 ( .A1(n3834), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5123)
         );
  AND2_X2 U3826 ( .A1(n4311), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4912)
         );
  AND2_X1 U3827 ( .A1(n3676), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3670)
         );
  AND2_X2 U3828 ( .A1(n3729), .A2(n4914), .ZN(n4001) );
  AND3_X1 U3829 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .ZN(n3729) );
  INV_X2 U3830 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4914) );
  INV_X1 U3831 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4311) );
  AND2_X2 U3832 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4906) );
  AND2_X2 U3833 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3774) );
  AND2_X1 U3834 ( .A1(n4043), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3666) );
  INV_X1 U3835 ( .A(n4114), .ZN(n3667) );
  INV_X1 U3836 ( .A(n3667), .ZN(n3668) );
  INV_X1 U3837 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3669) );
  AND2_X1 U3838 ( .A1(n3676), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4910)
         );
  AND2_X2 U3839 ( .A1(n5170), .A2(n5206), .ZN(n5093) );
  OR2_X2 U3840 ( .A1(n3915), .A2(n3914), .ZN(n5170) );
  AND2_X2 U3841 ( .A1(n3905), .A2(n4302), .ZN(n3671) );
  INV_X1 U3842 ( .A(n4040), .ZN(n3672) );
  NAND2_X1 U3843 ( .A1(n4031), .A2(n4302), .ZN(n4039) );
  AND2_X1 U3844 ( .A1(n3963), .A2(n5050), .ZN(n4866) );
  AND2_X1 U3845 ( .A1(n3840), .A2(n4906), .ZN(n3674) );
  AND2_X1 U3846 ( .A1(n3840), .A2(n4906), .ZN(n3704) );
  NAND2_X1 U3847 ( .A1(n3671), .A2(n3899), .ZN(n3970) );
  AND2_X2 U3848 ( .A1(n3886), .A2(n3885), .ZN(n3710) );
  AND3_X1 U3849 ( .A1(n4866), .A2(n4033), .A3(n4032), .ZN(n3675) );
  INV_X1 U3850 ( .A(n4036), .ZN(n4033) );
  AND2_X1 U3851 ( .A1(n3670), .A2(n3840), .ZN(n3677) );
  AND2_X1 U3852 ( .A1(n3670), .A2(n3840), .ZN(n3678) );
  AND2_X1 U3853 ( .A1(n3670), .A2(n3840), .ZN(n4088) );
  OR2_X1 U3854 ( .A1(n4295), .A2(n3710), .ZN(n3679) );
  NOR2_X1 U3855 ( .A1(n5521), .A2(n3813), .ZN(n3680) );
  NAND2_X1 U3856 ( .A1(n3680), .A2(n3681), .ZN(n5975) );
  AND2_X1 U3857 ( .A1(n5976), .A2(n5958), .ZN(n3681) );
  CLKBUF_X1 U3858 ( .A(n6457), .Z(n3682) );
  INV_X1 U3859 ( .A(n3683), .ZN(n5332) );
  INV_X1 U3860 ( .A(n6432), .ZN(n3684) );
  INV_X1 U3861 ( .A(n6431), .ZN(n3733) );
  INV_X1 U3862 ( .A(n3688), .ZN(n3689) );
  NAND2_X1 U3863 ( .A1(n4102), .A2(n4057), .ZN(n4301) );
  NAND2_X1 U3865 ( .A1(n3685), .A2(n6405), .ZN(U2955) );
  AOI21_X1 U3866 ( .B1(n6404), .B2(n6534), .A(n6403), .ZN(n6405) );
  AND2_X2 U3867 ( .A1(n3670), .A2(n3839), .ZN(n3987) );
  AND2_X2 U3868 ( .A1(n6154), .A2(n6155), .ZN(n6142) );
  NAND2_X1 U3869 ( .A1(n3733), .A2(n4228), .ZN(n3686) );
  NAND2_X1 U3870 ( .A1(n3733), .A2(n4228), .ZN(n3687) );
  INV_X1 U3871 ( .A(n4301), .ZN(n3688) );
  AOI21_X1 U3872 ( .B1(n5950), .B2(n5951), .A(n4219), .ZN(n3690) );
  CLKBUF_X1 U3873 ( .A(n5080), .Z(n3691) );
  NAND2_X1 U3874 ( .A1(n3733), .A2(n4228), .ZN(n6414) );
  AOI21_X1 U3875 ( .B1(n5950), .B2(n5951), .A(n4219), .ZN(n5961) );
  XNOR2_X1 U3876 ( .A(n4106), .B(n5937), .ZN(n5080) );
  INV_X1 U3877 ( .A(n4895), .ZN(n3692) );
  OAI22_X1 U3879 ( .A1(n5630), .A2(n5629), .B1(n4177), .B2(n5337), .ZN(n3694)
         );
  NAND2_X1 U3880 ( .A1(n4843), .A2(n4955), .ZN(n4882) );
  NAND2_X1 U3881 ( .A1(n4051), .A2(n4075), .ZN(n4072) );
  AND2_X2 U3882 ( .A1(n4038), .A2(n4037), .ZN(n4843) );
  INV_X2 U3883 ( .A(n3900), .ZN(n5165) );
  AND2_X1 U3884 ( .A1(n3840), .A2(n4905), .ZN(n3920) );
  NAND2_X1 U3885 ( .A1(n4865), .A2(n5170), .ZN(n4036) );
  INV_X2 U3886 ( .A(n3905), .ZN(n4031) );
  BUF_X8 U3887 ( .A(n4001), .Z(n3891) );
  INV_X2 U3888 ( .A(n4903), .ZN(n4054) );
  AND2_X4 U3889 ( .A1(n5116), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3840)
         );
  INV_X2 U3890 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5116) );
  NOR2_X4 U3891 ( .A1(n4817), .A2(n4818), .ZN(n6118) );
  NOR2_X2 U3893 ( .A1(n5112), .A2(n5111), .ZN(n5113) );
  AND2_X1 U3894 ( .A1(n3670), .A2(n3839), .ZN(n3699) );
  AND2_X4 U3895 ( .A1(n4905), .A2(n3774), .ZN(n3925) );
  AND2_X1 U3896 ( .A1(n4912), .A2(n3774), .ZN(n3701) );
  AND2_X1 U3897 ( .A1(n3840), .A2(n4905), .ZN(n3702) );
  AND2_X1 U3898 ( .A1(n3840), .A2(n4905), .ZN(n3703) );
  AOI21_X2 U3899 ( .B1(n5643), .B2(n5642), .A(n4163), .ZN(n5630) );
  NOR2_X2 U3900 ( .A1(n6208), .A2(n3820), .ZN(n6154) );
  NAND2_X2 U3901 ( .A1(n6207), .A2(n6209), .ZN(n6208) );
  NOR3_X2 U3902 ( .A1(n6414), .A2(n6601), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n6397) );
  NAND2_X2 U3903 ( .A1(n6337), .A2(n6338), .ZN(n6329) );
  OAI211_X2 U3904 ( .C1(n4050), .C2(n4914), .A(n4049), .B(n4048), .ZN(n4075)
         );
  XNOR2_X2 U3905 ( .A(n6118), .B(n6117), .ZN(n6005) );
  OAI21_X1 U3906 ( .B1(n4274), .B2(n4150), .A(n4149), .ZN(n4152) );
  NAND2_X1 U3907 ( .A1(n3737), .A2(n4128), .ZN(n4136) );
  INV_X1 U3908 ( .A(n4234), .ZN(n4274) );
  OR2_X1 U3909 ( .A1(n5721), .A2(n3966), .ZN(n4086) );
  NAND2_X1 U3910 ( .A1(n3762), .A2(n6333), .ZN(n3761) );
  INV_X1 U3911 ( .A(n6344), .ZN(n3762) );
  INV_X1 U3912 ( .A(n3750), .ZN(n3749) );
  NAND2_X1 U3913 ( .A1(n3750), .A2(n3748), .ZN(n3747) );
  OR2_X1 U3914 ( .A1(n3899), .A2(n3966), .ZN(n4087) );
  NAND2_X1 U3915 ( .A1(n7522), .A2(n7303), .ZN(n5704) );
  INV_X1 U3916 ( .A(n6157), .ZN(n3768) );
  INV_X2 U3917 ( .A(n4348), .ZN(n4766) );
  NAND2_X1 U3918 ( .A1(n6167), .A2(n3821), .ZN(n3820) );
  INV_X1 U3919 ( .A(n3823), .ZN(n3821) );
  NAND2_X1 U3920 ( .A1(n3822), .A2(n3825), .ZN(n6178) );
  INV_X1 U3921 ( .A(n6208), .ZN(n3822) );
  NAND2_X1 U3922 ( .A1(n4227), .A2(n3738), .ZN(n6431) );
  OAI21_X1 U3923 ( .B1(n6441), .B2(n4226), .A(n3783), .ZN(n3738) );
  NOR2_X1 U3924 ( .A1(n4210), .A2(n4209), .ZN(n4211) );
  OR2_X1 U3925 ( .A1(n4189), .A2(n4188), .ZN(n4198) );
  AOI22_X1 U3926 ( .A1(n4234), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4290), 
        .B2(n4195), .ZN(n4178) );
  AND2_X1 U3927 ( .A1(n4290), .A2(n4198), .ZN(n4190) );
  NOR2_X2 U3928 ( .A1(n4179), .A2(n4178), .ZN(n4194) );
  OR2_X1 U3929 ( .A1(n4028), .A2(n4027), .ZN(n4058) );
  AND2_X1 U3930 ( .A1(n4914), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U3931 ( .A1(n3824), .A2(n3825), .ZN(n3823) );
  INV_X1 U3932 ( .A(n6179), .ZN(n3824) );
  AND2_X1 U3933 ( .A1(n4669), .A2(n3826), .ZN(n3825) );
  INV_X1 U3934 ( .A(n6309), .ZN(n3826) );
  INV_X1 U3935 ( .A(n6195), .ZN(n4669) );
  AND2_X1 U3936 ( .A1(n4454), .A2(n6274), .ZN(n3805) );
  NOR2_X1 U3937 ( .A1(n5557), .A2(n3818), .ZN(n3817) );
  NAND2_X1 U3938 ( .A1(n4155), .A2(n4179), .ZN(n4339) );
  INV_X1 U3939 ( .A(n5704), .ZN(n4798) );
  NAND2_X1 U3940 ( .A1(n6487), .A2(n6442), .ZN(n6445) );
  INV_X1 U3941 ( .A(n6520), .ZN(n3751) );
  AND2_X1 U3942 ( .A1(n3772), .A2(n3771), .ZN(n3770) );
  INV_X1 U3943 ( .A(n6750), .ZN(n3771) );
  AND2_X1 U3944 ( .A1(n5919), .A2(n3773), .ZN(n3772) );
  INV_X1 U3945 ( .A(n5983), .ZN(n3773) );
  AND2_X1 U3946 ( .A1(n5093), .A2(n6018), .ZN(n6052) );
  INV_X1 U3947 ( .A(n6052), .ZN(n6107) );
  NAND2_X1 U3948 ( .A1(n4309), .A2(n3966), .ZN(n3736) );
  NOR2_X1 U3949 ( .A1(n6170), .A2(n3767), .ZN(n3764) );
  NAND2_X1 U3950 ( .A1(n3769), .A2(n3768), .ZN(n3767) );
  NOR2_X1 U3951 ( .A1(n6146), .A2(EBX_REG_29__SCAN_IN), .ZN(n3769) );
  OR2_X1 U3952 ( .A1(n4896), .A2(n4956), .ZN(n6100) );
  INV_X1 U3953 ( .A(n4498), .ZN(n6119) );
  OR2_X1 U3954 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  OR2_X1 U3955 ( .A1(n4772), .A2(n6134), .ZN(n5709) );
  NOR2_X1 U3956 ( .A1(n4724), .A2(n6425), .ZN(n4725) );
  NAND2_X1 U3957 ( .A1(n4725), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4771)
         );
  OR2_X1 U3958 ( .A1(n4687), .A2(n6180), .ZN(n4724) );
  OR2_X1 U3959 ( .A1(n4599), .A2(n6475), .ZN(n4649) );
  NAND2_X1 U3960 ( .A1(n6320), .A2(n3809), .ZN(n3808) );
  INV_X1 U3961 ( .A(n3811), .ZN(n3809) );
  INV_X1 U3962 ( .A(n6329), .ZN(n3810) );
  OR2_X1 U3963 ( .A1(n7421), .A2(n5704), .ZN(n4524) );
  NAND2_X1 U3964 ( .A1(n3815), .A2(n4393), .ZN(n3814) );
  OR2_X1 U3965 ( .A1(n6099), .A2(n7546), .ZN(n4920) );
  OR2_X1 U3966 ( .A1(n6190), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U3967 ( .A1(n6203), .A2(n6188), .ZN(n6190) );
  AND2_X1 U3968 ( .A1(n3786), .A2(n3831), .ZN(n3785) );
  NOR2_X2 U3969 ( .A1(n6345), .A2(n3723), .ZN(n6322) );
  NOR2_X1 U3970 ( .A1(n6345), .A2(n6344), .ZN(n6346) );
  NOR3_X1 U3971 ( .A1(n6345), .A2(n3763), .A3(n6344), .ZN(n6341) );
  NAND2_X1 U3972 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4222) );
  NOR2_X1 U3973 ( .A1(n3679), .A2(n3972), .ZN(n4980) );
  NAND2_X1 U3974 ( .A1(n3693), .A2(n6529), .ZN(n3752) );
  NAND2_X1 U3975 ( .A1(n3752), .A2(n3750), .ZN(n6519) );
  AOI21_X1 U3976 ( .B1(n3707), .B2(n3780), .A(n3709), .ZN(n3779) );
  INV_X1 U3977 ( .A(n6543), .ZN(n3780) );
  NOR2_X1 U3978 ( .A1(n6543), .A2(n3782), .ZN(n3781) );
  INV_X1 U3979 ( .A(n5989), .ZN(n3782) );
  NOR2_X1 U3980 ( .A1(n4218), .A2(n4216), .ZN(n4219) );
  NAND2_X1 U3981 ( .A1(n3743), .A2(n3742), .ZN(n3741) );
  AND2_X1 U3982 ( .A1(n7348), .A2(n6732), .ZN(n6727) );
  NAND2_X1 U3983 ( .A1(n4966), .A2(n5175), .ZN(n4986) );
  NAND2_X1 U3984 ( .A1(n4102), .A2(n4101), .ZN(n4127) );
  INV_X1 U3985 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7506) );
  NAND2_X1 U3986 ( .A1(n5142), .A2(n3774), .ZN(n5143) );
  NAND2_X1 U3987 ( .A1(n7426), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6124) );
  AND2_X1 U3988 ( .A1(n7426), .A2(n5712), .ZN(n7477) );
  NAND2_X1 U3989 ( .A1(n5054), .A2(n5053), .ZN(n6391) );
  OR2_X2 U3990 ( .A1(n4920), .A2(n7509), .ZN(n7482) );
  NAND2_X1 U3991 ( .A1(n3803), .A2(n5146), .ZN(n3801) );
  NOR2_X1 U3992 ( .A1(n5219), .A2(n7522), .ZN(n4312) );
  INV_X1 U3993 ( .A(n6529), .ZN(n3748) );
  OAI211_X1 U3994 ( .C1(n4865), .C2(n3899), .A(n5170), .B(n3963), .ZN(n3976)
         );
  OR2_X1 U3995 ( .A1(n4173), .A2(n4172), .ZN(n4195) );
  OR2_X1 U3996 ( .A1(n4148), .A2(n4147), .ZN(n4158) );
  AND2_X1 U3997 ( .A1(n4955), .A2(n3758), .ZN(n4042) );
  INV_X1 U3998 ( .A(n4822), .ZN(n3758) );
  AOI22_X1 U3999 ( .A1(n4411), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4000 ( .A1(n3730), .A2(n3968), .ZN(n4052) );
  NAND2_X1 U4001 ( .A1(n4077), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4002 ( .A1(n4598), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4599)
         );
  NAND2_X1 U4003 ( .A1(n3812), .A2(n4563), .ZN(n3811) );
  INV_X1 U4004 ( .A(n6219), .ZN(n3812) );
  INV_X1 U4005 ( .A(n6332), .ZN(n4563) );
  NAND2_X1 U4006 ( .A1(n4487), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4518)
         );
  NOR2_X1 U4007 ( .A1(n4410), .A2(n4409), .ZN(n4424) );
  INV_X1 U4008 ( .A(n5916), .ZN(n3815) );
  INV_X1 U4009 ( .A(n5698), .ZN(n3818) );
  AND2_X1 U4010 ( .A1(n3788), .A2(n3719), .ZN(n3786) );
  INV_X1 U4011 ( .A(n6538), .ZN(n3778) );
  NAND2_X1 U4012 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  AOI21_X1 U4013 ( .B1(n4301), .B2(n5206), .A(n4060), .ZN(n4070) );
  NOR2_X1 U4014 ( .A1(n3711), .A2(n3735), .ZN(n3734) );
  INV_X1 U4015 ( .A(n4016), .ZN(n3735) );
  OR2_X1 U4016 ( .A1(n4098), .A2(n4097), .ZN(n4130) );
  OR2_X1 U4017 ( .A1(n4046), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4047)
         );
  OR2_X1 U4018 ( .A1(n4124), .A2(n4123), .ZN(n4133) );
  AOI21_X1 U4019 ( .B1(n4784), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n3955), 
        .ZN(n3956) );
  NAND2_X1 U4020 ( .A1(n3728), .A2(n3729), .ZN(n3952) );
  AOI21_X1 U4021 ( .B1(n7536), .B2(n7542), .A(n6087), .ZN(n5164) );
  NAND2_X1 U4022 ( .A1(n4087), .A2(n4086), .ZN(n4290) );
  INV_X1 U4023 ( .A(n4276), .ZN(n4287) );
  INV_X1 U4024 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7501) );
  INV_X1 U4025 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U4026 ( .A1(n3971), .A2(n5206), .ZN(n5752) );
  AND2_X1 U4027 ( .A1(n6028), .A2(n6027), .ZN(n6344) );
  AND2_X1 U4028 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  OR2_X1 U4029 ( .A1(n5097), .A2(n5096), .ZN(n5293) );
  INV_X1 U4030 ( .A(n7196), .ZN(n4921) );
  AND2_X1 U4031 ( .A1(n6074), .A2(n4798), .ZN(n4799) );
  AND2_X1 U4032 ( .A1(n6408), .A2(n4798), .ZN(n4746) );
  AND2_X1 U4033 ( .A1(n6429), .A2(n4798), .ZN(n4705) );
  NAND2_X1 U4034 ( .A1(n4686), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4687)
         );
  INV_X1 U4035 ( .A(n4685), .ZN(n4686) );
  NAND2_X1 U4036 ( .A1(n4690), .A2(n4689), .ZN(n6179) );
  OR2_X1 U4037 ( .A1(n6437), .A2(n5704), .ZN(n4689) );
  AND3_X1 U4038 ( .A1(n4668), .A2(n4667), .A3(n4666), .ZN(n6195) );
  AND2_X1 U4039 ( .A1(n6469), .A2(n4798), .ZN(n4620) );
  AND2_X1 U4040 ( .A1(n4556), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4557)
         );
  NOR2_X1 U4041 ( .A1(n4518), .A2(n6503), .ZN(n4519) );
  AND2_X1 U4042 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4519), .ZN(n4556)
         );
  NOR2_X1 U4043 ( .A1(n3795), .A2(n6348), .ZN(n3793) );
  NOR2_X1 U4044 ( .A1(n4471), .A2(n6261), .ZN(n4487) );
  AOI21_X1 U4045 ( .B1(n3807), .B2(n6274), .A(n4454), .ZN(n3806) );
  NAND2_X1 U4046 ( .A1(n5975), .A2(n3805), .ZN(n3804) );
  NAND2_X1 U4047 ( .A1(n4424), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4451)
         );
  NAND2_X1 U4048 ( .A1(n4394), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4410)
         );
  NOR2_X1 U4049 ( .A1(n4380), .A2(n5952), .ZN(n4394) );
  NAND2_X1 U4050 ( .A1(n4359), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4380)
         );
  INV_X1 U4051 ( .A(n4363), .ZN(n4364) );
  AND2_X1 U4052 ( .A1(n4349), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4359)
         );
  NAND2_X1 U4053 ( .A1(n4333), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4342)
         );
  AND3_X1 U4054 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4333) );
  NAND2_X1 U4055 ( .A1(n5157), .A2(n4480), .ZN(n4300) );
  NOR2_X1 U4056 ( .A1(n3791), .A2(n6622), .ZN(n3790) );
  INV_X1 U4057 ( .A(n3830), .ZN(n3791) );
  NOR3_X1 U4058 ( .A1(n6170), .A2(n6157), .A3(n6146), .ZN(n6145) );
  NOR2_X1 U4059 ( .A1(n6310), .A2(n6204), .ZN(n6203) );
  NAND2_X1 U4060 ( .A1(n3760), .A2(n3759), .ZN(n6310) );
  INV_X1 U4061 ( .A(n6313), .ZN(n3759) );
  NAND2_X1 U4062 ( .A1(n6445), .A2(n6444), .ZN(n6473) );
  NAND2_X1 U4063 ( .A1(n3783), .A2(n3829), .ZN(n4224) );
  NOR2_X1 U4064 ( .A1(n6441), .A2(n6488), .ZN(n6487) );
  NAND2_X1 U4065 ( .A1(n3712), .A2(n3789), .ZN(n3788) );
  INV_X1 U4066 ( .A(n6510), .ZN(n3789) );
  OR2_X1 U4067 ( .A1(n6259), .A2(n6024), .ZN(n6345) );
  AND2_X1 U4068 ( .A1(n5920), .A2(n3726), .ZN(n6277) );
  AND2_X1 U4069 ( .A1(n6015), .A2(n6014), .ZN(n6258) );
  NAND2_X1 U4070 ( .A1(n6277), .A2(n6258), .ZN(n6259) );
  AND2_X1 U4071 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  NAND2_X1 U4072 ( .A1(n5920), .A2(n3772), .ZN(n6749) );
  NAND2_X1 U4073 ( .A1(n5920), .A2(n5919), .ZN(n5984) );
  AND2_X1 U4074 ( .A1(n5832), .A2(n5831), .ZN(n5920) );
  NOR2_X1 U4075 ( .A1(n5700), .A2(n5701), .ZN(n5832) );
  AND2_X1 U4076 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U4077 ( .A1(n3757), .A2(n3756), .ZN(n5700) );
  INV_X1 U4078 ( .A(n5566), .ZN(n3756) );
  NAND2_X1 U4079 ( .A1(n5480), .A2(n5341), .ZN(n5525) );
  AND2_X1 U4080 ( .A1(n5336), .A2(n5335), .ZN(n5477) );
  AND2_X1 U4081 ( .A1(n5478), .A2(n5477), .ZN(n5480) );
  NOR2_X1 U4082 ( .A1(n5293), .A2(n5292), .ZN(n5478) );
  XNOR2_X1 U4083 ( .A(n4162), .B(n4161), .ZN(n5643) );
  NAND2_X1 U4084 ( .A1(n3746), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3745)
         );
  OR2_X1 U4085 ( .A1(n6100), .A2(n4986), .ZN(n6683) );
  NAND2_X1 U4086 ( .A1(n3736), .A2(n4016), .ZN(n4064) );
  NAND2_X1 U4087 ( .A1(n4082), .A2(n4075), .ZN(n3803) );
  INV_X1 U4088 ( .A(n4083), .ZN(n4082) );
  NOR2_X1 U4089 ( .A1(n4295), .A2(n4296), .ZN(n4960) );
  INV_X1 U4090 ( .A(n5206), .ZN(n4955) );
  NAND2_X1 U4091 ( .A1(n3800), .A2(n4076), .ZN(n5147) );
  INV_X1 U4092 ( .A(n3803), .ZN(n3800) );
  INV_X1 U4093 ( .A(n7546), .ZN(n5175) );
  INV_X1 U4094 ( .A(n5396), .ZN(n5227) );
  AND2_X1 U4095 ( .A1(n3706), .A2(n5158), .ZN(n5163) );
  INV_X1 U4096 ( .A(n5456), .ZN(n5575) );
  CLKBUF_X1 U4097 ( .A(n4302), .Z(n5219) );
  INV_X1 U4098 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7098) );
  OR2_X1 U4099 ( .A1(n4920), .A2(n4853), .ZN(n4861) );
  INV_X1 U4100 ( .A(n7472), .ZN(n7450) );
  AND2_X1 U4101 ( .A1(n7426), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7472) );
  OR3_X1 U4102 ( .A1(n6124), .A2(n5724), .A3(n5723), .ZN(n7446) );
  INV_X1 U4103 ( .A(n7467), .ZN(n7473) );
  INV_X1 U4104 ( .A(n7370), .ZN(n7354) );
  NOR2_X1 U4105 ( .A1(n6111), .A2(n3765), .ZN(n6061) );
  NOR3_X1 U4106 ( .A1(n6170), .A2(n6146), .A3(n3766), .ZN(n3765) );
  NAND2_X1 U4107 ( .A1(n3768), .A2(n6060), .ZN(n3766) );
  INV_X1 U4108 ( .A(n6359), .ZN(n7284) );
  NAND2_X1 U4109 ( .A1(n6352), .A2(n3901), .ZN(n6359) );
  INV_X1 U4110 ( .A(n6391), .ZN(n7583) );
  AND2_X1 U4111 ( .A1(n6391), .A2(n6006), .ZN(n7584) );
  NAND2_X1 U4112 ( .A1(n6391), .A2(n5056), .ZN(n6394) );
  XNOR2_X1 U4113 ( .A(n5710), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6402)
         );
  AND2_X1 U4114 ( .A1(n5709), .A2(n4773), .ZN(n6132) );
  AND2_X1 U4115 ( .A1(n4771), .A2(n4727), .ZN(n6422) );
  INV_X1 U4116 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6503) );
  INV_X1 U4117 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5952) );
  NOR2_X1 U4118 ( .A1(n5718), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6546) );
  AND2_X1 U4119 ( .A1(n7482), .A2(n4803), .ZN(n7289) );
  XNOR2_X1 U4120 ( .A(n3753), .B(n4816), .ZN(n6600) );
  AND2_X1 U4121 ( .A1(n6627), .A2(n6618), .ZN(n6603) );
  INV_X1 U4122 ( .A(n3687), .ZN(n6433) );
  NAND2_X1 U4123 ( .A1(n6519), .A2(n4222), .ZN(n6511) );
  OR2_X1 U4124 ( .A1(n4986), .A2(n4982), .ZN(n6732) );
  AND2_X1 U4125 ( .A1(n3752), .A2(n4220), .ZN(n6521) );
  NAND2_X1 U4126 ( .A1(n5990), .A2(n3781), .ZN(n3777) );
  AOI21_X1 U4127 ( .B1(n5990), .B2(n5989), .A(n3707), .ZN(n6544) );
  OR2_X1 U4128 ( .A1(n6727), .A2(n5087), .ZN(n6741) );
  AND2_X1 U4129 ( .A1(n7348), .A2(n7349), .ZN(n5087) );
  INV_X1 U4130 ( .A(n6546), .ZN(n6759) );
  OR2_X1 U4131 ( .A1(n4986), .A2(n5134), .ZN(n7348) );
  INV_X1 U4132 ( .A(n6765), .ZN(n7344) );
  INV_X1 U4133 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7557) );
  INV_X1 U4134 ( .A(n4308), .ZN(n7554) );
  CLKBUF_X1 U4135 ( .A(n4903), .Z(n4904) );
  NOR2_X1 U4136 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6081) );
  INV_X1 U4137 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7490) );
  INV_X1 U4138 ( .A(n5367), .ZN(n7722) );
  INV_X1 U4139 ( .A(n7646), .ZN(n7642) );
  OAI21_X1 U4140 ( .B1(n5585), .B2(n5584), .A(n5583), .ZN(n7710) );
  AND2_X1 U4141 ( .A1(n5163), .A2(n4308), .ZN(n5822) );
  INV_X1 U4142 ( .A(n5498), .ZN(n7608) );
  INV_X1 U4143 ( .A(n5790), .ZN(n7631) );
  INV_X1 U4144 ( .A(n5785), .ZN(n7652) );
  INV_X1 U4145 ( .A(n7144), .ZN(n7697) );
  INV_X1 U4146 ( .A(n5768), .ZN(n7747) );
  INV_X1 U4147 ( .A(n7147), .ZN(n5432) );
  OR2_X1 U4148 ( .A1(n6099), .A2(n7534), .ZN(n7543) );
  OR4_X1 U4149 ( .A1(n7515), .A2(n7514), .A3(n7513), .A4(n7512), .ZN(n7535) );
  NAND2_X1 U4150 ( .A1(n4808), .A2(n4807), .ZN(n4809) );
  AND2_X2 U4151 ( .A1(n5123), .A2(n4910), .ZN(n3999) );
  AND2_X1 U4152 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3707)
         );
  NAND2_X1 U4153 ( .A1(n6697), .A2(n6730), .ZN(n4220) );
  NAND2_X1 U4154 ( .A1(n3816), .A2(n3817), .ZN(n5697) );
  AND2_X1 U4155 ( .A1(n4486), .A2(n4485), .ZN(n3708) );
  INV_X1 U4156 ( .A(n4220), .ZN(n4221) );
  AND2_X1 U4157 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3709)
         );
  AOI21_X1 U4158 ( .B1(n3684), .B2(n3725), .A(n6697), .ZN(n4815) );
  AND2_X1 U4159 ( .A1(n4486), .A2(n3793), .ZN(n6337) );
  NOR2_X1 U4160 ( .A1(n6208), .A2(n6309), .ZN(n6193) );
  OR2_X1 U4161 ( .A1(n4030), .A2(n4029), .ZN(n3711) );
  AND2_X1 U4162 ( .A1(n3755), .A2(n3754), .ZN(n6406) );
  NAND2_X1 U4163 ( .A1(n4486), .A2(n3794), .ZN(n6234) );
  OR2_X1 U4164 ( .A1(n4223), .A2(n6697), .ZN(n3712) );
  NAND2_X1 U4165 ( .A1(n3784), .A2(n3788), .ZN(n6501) );
  NAND2_X1 U4166 ( .A1(n5165), .A2(n3710), .ZN(n4034) );
  AND2_X1 U4167 ( .A1(n3781), .A2(n6538), .ZN(n3713) );
  OR2_X1 U4168 ( .A1(n6170), .A2(n6157), .ZN(n3714) );
  NAND2_X1 U4169 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3716) );
  AND2_X1 U4170 ( .A1(n4204), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3717)
         );
  NOR2_X1 U4171 ( .A1(n6329), .A2(n3811), .ZN(n6220) );
  AND2_X1 U4172 ( .A1(n3712), .A2(n4222), .ZN(n3718) );
  NAND2_X1 U4173 ( .A1(n3736), .A2(n3734), .ZN(n4101) );
  NAND2_X1 U4174 ( .A1(n6697), .A2(n7335), .ZN(n3719) );
  OR2_X1 U4175 ( .A1(n4055), .A2(n4087), .ZN(n3720) );
  AND2_X1 U4176 ( .A1(n3718), .A2(n3747), .ZN(n3721) );
  OAI22_X1 U4177 ( .A1(n5961), .A2(n5962), .B1(n6551), .B2(n6697), .ZN(n5990)
         );
  NOR2_X1 U4178 ( .A1(n5521), .A2(n5557), .ZN(n5556) );
  AND2_X1 U4179 ( .A1(n5920), .A2(n3770), .ZN(n3722) );
  OR3_X1 U4180 ( .A1(n3761), .A2(n3763), .A3(n6222), .ZN(n3723) );
  XNOR2_X1 U4181 ( .A(n5975), .B(n4454), .ZN(n6273) );
  NAND2_X1 U4182 ( .A1(n3777), .A2(n3779), .ZN(n6537) );
  OR3_X1 U4183 ( .A1(n6345), .A2(n3761), .A3(n3763), .ZN(n3724) );
  AND2_X1 U4184 ( .A1(n4228), .A2(n4813), .ZN(n3725) );
  INV_X1 U4185 ( .A(n5521), .ZN(n3816) );
  INV_X1 U4186 ( .A(n3760), .ZN(n6312) );
  NOR2_X1 U4187 ( .A1(n6324), .A2(n6210), .ZN(n3760) );
  AOI21_X1 U4188 ( .B1(n5992), .B2(n4798), .A(n4408), .ZN(n5916) );
  AND2_X1 U4189 ( .A1(n3770), .A2(n6275), .ZN(n3726) );
  OR2_X1 U4190 ( .A1(n3814), .A2(n3818), .ZN(n3727) );
  INV_X1 U4191 ( .A(n4454), .ZN(n3807) );
  OR2_X1 U4192 ( .A1(n5525), .A2(n5526), .ZN(n5567) );
  INV_X1 U4193 ( .A(n5567), .ZN(n3757) );
  INV_X1 U4194 ( .A(n4233), .ZN(n4210) );
  AND2_X1 U4195 ( .A1(n5165), .A2(n5206), .ZN(n4233) );
  INV_X1 U4196 ( .A(n3795), .ZN(n3794) );
  NAND2_X1 U4197 ( .A1(n4485), .A2(n4503), .ZN(n3795) );
  NAND2_X1 U4198 ( .A1(n4113), .A2(n4112), .ZN(n5146) );
  INV_X1 U4199 ( .A(n5146), .ZN(n3802) );
  AND2_X2 U4200 ( .A1(n3731), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4077) );
  NAND3_X1 U4201 ( .A1(n3965), .A2(n3967), .A3(n3964), .ZN(n3731) );
  NAND3_X4 U4202 ( .A1(n3732), .A2(n3957), .A3(n3958), .ZN(n5206) );
  INV_X1 U4203 ( .A(n4136), .ZN(n4138) );
  INV_X1 U4204 ( .A(n4127), .ZN(n3737) );
  XNOR2_X1 U4205 ( .A(n3744), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5508)
         );
  NAND2_X1 U4206 ( .A1(n3740), .A2(n3744), .ZN(n3739) );
  OAI21_X1 U4207 ( .B1(n5509), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5515), 
        .ZN(n3740) );
  NOR2_X1 U4208 ( .A1(n5509), .A2(n5515), .ZN(n3742) );
  INV_X1 U4209 ( .A(n3744), .ZN(n3743) );
  OAI21_X2 U4210 ( .B1(n5080), .B2(n5081), .A(n3745), .ZN(n3744) );
  INV_X1 U4211 ( .A(n4106), .ZN(n3746) );
  OAI21_X1 U4212 ( .B1(n6530), .B2(n3749), .A(n3721), .ZN(n3787) );
  NAND2_X1 U4213 ( .A1(n6407), .A2(n3755), .ZN(n3753) );
  NAND2_X1 U4214 ( .A1(n4814), .A2(n6697), .ZN(n3754) );
  INV_X1 U4215 ( .A(n4815), .ZN(n3755) );
  AND2_X2 U4216 ( .A1(n4955), .A2(n5721), .ZN(n7304) );
  INV_X1 U4217 ( .A(n6339), .ZN(n3763) );
  NOR2_X1 U4218 ( .A1(n3764), .A2(n5523), .ZN(n6111) );
  AND2_X2 U4219 ( .A1(n4906), .A2(n3774), .ZN(n4582) );
  AOI21_X2 U4220 ( .B1(n5990), .B2(n3713), .A(n3775), .ZN(n6530) );
  CLKBUF_X1 U4221 ( .A(n3787), .Z(n3784) );
  NAND2_X1 U4222 ( .A1(n3686), .A2(n3830), .ZN(n3792) );
  XNOR2_X1 U4223 ( .A(n3792), .B(n6424), .ZN(n6626) );
  NAND2_X1 U4224 ( .A1(n3798), .A2(n3797), .ZN(n3796) );
  OAI21_X1 U4225 ( .B1(n5146), .B2(n3803), .A(n4076), .ZN(n3797) );
  NAND2_X1 U4226 ( .A1(n3799), .A2(n3802), .ZN(n3798) );
  INV_X1 U4227 ( .A(n4076), .ZN(n3799) );
  NAND2_X1 U4228 ( .A1(n4076), .A2(n4075), .ZN(n4084) );
  OAI21_X2 U4229 ( .B1(n5975), .B2(n3806), .A(n3804), .ZN(n6257) );
  NAND2_X1 U4230 ( .A1(n6257), .A2(n6256), .ZN(n6248) );
  NAND3_X1 U4231 ( .A1(n3816), .A2(n3817), .A3(n4393), .ZN(n3819) );
  INV_X1 U4232 ( .A(n3819), .ZN(n5826) );
  NOR2_X1 U4233 ( .A1(n6208), .A2(n3823), .ZN(n6165) );
  NAND2_X1 U4234 ( .A1(n4054), .A2(n3966), .ZN(n4056) );
  NAND3_X1 U4235 ( .A1(n4101), .A2(n4056), .A3(n3720), .ZN(n4102) );
  NAND2_X1 U4236 ( .A1(n4784), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3864) );
  AND2_X1 U4237 ( .A1(n5311), .A2(n3664), .ZN(n5319) );
  NAND2_X1 U4238 ( .A1(n4325), .A2(n4324), .ZN(n5112) );
  OR2_X1 U4239 ( .A1(n5077), .A2(n5076), .ZN(n4324) );
  CLKBUF_X1 U4240 ( .A(n5155), .Z(n5333) );
  OAI22_X2 U4241 ( .A1(n5934), .A2(n5935), .B1(n4208), .B2(n5560), .ZN(n5950)
         );
  INV_X1 U4242 ( .A(n6233), .ZN(n4503) );
  AND3_X1 U4243 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3827) );
  NAND2_X1 U4244 ( .A1(n4199), .A2(n4198), .ZN(n3828) );
  INV_X1 U4245 ( .A(n4312), .ZN(n4348) );
  OR3_X1 U4246 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3829) );
  OR2_X1 U4247 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3830)
         );
  OR2_X1 U4248 ( .A1(n3783), .A2(n6554), .ZN(n3831) );
  AND3_X1 U4249 ( .A1(n6565), .A2(n6572), .A3(n6570), .ZN(n3832) );
  INV_X1 U4250 ( .A(n6565), .ZN(n6443) );
  INV_X1 U4251 ( .A(n6352), .ZN(n6353) );
  INV_X1 U4252 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4223) );
  INV_X1 U4253 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3966) );
  INV_X1 U4254 ( .A(n6193), .ZN(n6308) );
  AND2_X1 U4255 ( .A1(n4261), .A2(n4256), .ZN(n4257) );
  OR2_X1 U4256 ( .A1(n4236), .A2(n4241), .ZN(n4255) );
  OAI21_X1 U4257 ( .B1(n3978), .B2(n4065), .A(n3977), .ZN(n3979) );
  INV_X1 U4258 ( .A(n4058), .ZN(n4055) );
  AND2_X1 U4259 ( .A1(n7490), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4281)
         );
  NAND2_X1 U4260 ( .A1(n4234), .A2(n4233), .ZN(n4276) );
  AND2_X1 U4261 ( .A1(n4045), .A2(n4044), .ZN(n4049) );
  INV_X1 U4262 ( .A(n4843), .ZN(n4887) );
  INV_X1 U4263 ( .A(n4649), .ZN(n4650) );
  AOI22_X1 U4264 ( .A1(n3920), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3987), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3849) );
  AND2_X1 U4265 ( .A1(n4480), .A2(n4450), .ZN(n4454) );
  INV_X1 U4266 ( .A(n4597), .ZN(n4598) );
  NAND2_X1 U4267 ( .A1(n4465), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4471)
         );
  INV_X1 U4268 ( .A(n5522), .ZN(n4357) );
  NAND2_X1 U4269 ( .A1(n3783), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6442) );
  NOR2_X1 U4270 ( .A1(n4200), .A2(n4065), .ZN(n4201) );
  NAND2_X1 U4271 ( .A1(n4650), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4651)
         );
  INV_X1 U4272 ( .A(n4342), .ZN(n4341) );
  AND2_X1 U4273 ( .A1(n6032), .A2(n6031), .ZN(n6339) );
  NOR2_X1 U4274 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  NAND2_X1 U4275 ( .A1(n4960), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4768) );
  NOR2_X1 U4276 ( .A1(n4451), .A2(n7413), .ZN(n4465) );
  INV_X1 U4277 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4409) );
  INV_X1 U4278 ( .A(n4355), .ZN(n4356) );
  NOR2_X2 U4279 ( .A1(n5049), .A2(n7522), .ZN(n4480) );
  NAND2_X1 U4280 ( .A1(n6697), .A2(n6443), .ZN(n6444) );
  OR2_X1 U4281 ( .A1(n3706), .A2(n3689), .ZN(n5395) );
  INV_X1 U4282 ( .A(n5226), .ZN(n5220) );
  OR2_X1 U4283 ( .A1(n4651), .A2(n6460), .ZN(n4685) );
  INV_X1 U4284 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n7413) );
  AND2_X1 U4285 ( .A1(n6402), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5713) );
  AND2_X1 U4286 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4341), .ZN(n4349)
         );
  NAND2_X1 U4287 ( .A1(n7306), .A2(n5707), .ZN(n7426) );
  OR2_X1 U4288 ( .A1(n4967), .A2(READY_N), .ZN(n4881) );
  NAND2_X1 U4289 ( .A1(n4557), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4597)
         );
  INV_X1 U4290 ( .A(n4480), .ZN(n4470) );
  INV_X1 U4291 ( .A(n7289), .ZN(n6516) );
  OR2_X1 U4292 ( .A1(n6659), .A2(n6571), .ZN(n6645) );
  AND2_X1 U4293 ( .A1(n4162), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4163)
         );
  OR2_X1 U4294 ( .A1(n5542), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5399) );
  NOR2_X1 U4295 ( .A1(n3664), .A2(n5395), .ZN(n5459) );
  OR2_X1 U4296 ( .A1(n5280), .A2(n7554), .ZN(n5367) );
  OR2_X1 U4297 ( .A1(n5442), .A2(n7554), .ZN(n5620) );
  INV_X1 U4299 ( .A(n5822), .ZN(n5691) );
  AOI21_X1 U4300 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7557), .A(n5227), .ZN(
        n5461) );
  NAND2_X1 U4301 ( .A1(n7534), .A2(n7522), .ZN(n5456) );
  NAND2_X1 U4302 ( .A1(n4292), .A2(n4291), .ZN(n6099) );
  OR2_X1 U4303 ( .A1(n5836), .A2(n7388), .ZN(n6281) );
  INV_X1 U4304 ( .A(n7443), .ZN(n7471) );
  AND2_X1 U4305 ( .A1(n7426), .A2(n5713), .ZN(n7475) );
  INV_X1 U4306 ( .A(n7446), .ZN(n7470) );
  OAI21_X1 U4307 ( .B1(n7304), .B2(n7516), .A(n4862), .ZN(n5042) );
  INV_X1 U4308 ( .A(n5014), .ZN(n5015) );
  INV_X1 U4309 ( .A(n7294), .ZN(n6513) );
  NAND2_X1 U4310 ( .A1(n6322), .A2(n6321), .ZN(n6324) );
  INV_X1 U4311 ( .A(n6759), .ZN(n7330) );
  INV_X1 U4312 ( .A(n7342), .ZN(n7332) );
  INV_X1 U4313 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5711) );
  INV_X1 U4314 ( .A(n7543), .ZN(n6087) );
  INV_X1 U4315 ( .A(n7740), .ZN(n7694) );
  AND2_X1 U4316 ( .A1(n5459), .A2(n7554), .ZN(n7742) );
  AND2_X1 U4317 ( .A1(n5354), .A2(n4308), .ZN(n7731) );
  AND2_X1 U4318 ( .A1(n5346), .A2(n5345), .ZN(n5354) );
  INV_X1 U4319 ( .A(n5627), .ZN(n7723) );
  OAI211_X1 U4320 ( .C1(n5592), .C2(n7534), .A(n5546), .B(n5545), .ZN(n5619)
         );
  INV_X1 U4321 ( .A(n5620), .ZN(n5745) );
  OAI211_X1 U4322 ( .C1(n5872), .C2(n7534), .A(n5871), .B(n5870), .ZN(n5907)
         );
  INV_X1 U4323 ( .A(n5914), .ZN(n7715) );
  AND2_X1 U4324 ( .A1(n5319), .A2(n7554), .ZN(n7716) );
  INV_X1 U4325 ( .A(n7708), .ZN(n7701) );
  AND2_X1 U4326 ( .A1(n5345), .A2(n3664), .ZN(n5302) );
  INV_X1 U4327 ( .A(n7699), .ZN(n7676) );
  NOR2_X1 U4328 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5164), .ZN(n5396) );
  INV_X1 U4329 ( .A(n5537), .ZN(n5231) );
  AND2_X1 U4330 ( .A1(n5711), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4293) );
  OR2_X1 U4331 ( .A1(n5456), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5718) );
  AND2_X1 U4332 ( .A1(n4861), .A2(n4855), .ZN(n7306) );
  INV_X1 U4333 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7303) );
  OR3_X1 U4334 ( .A1(n6124), .A2(n6113), .A3(n5717), .ZN(n7467) );
  INV_X1 U4335 ( .A(n7477), .ZN(n7437) );
  OR2_X1 U4336 ( .A1(n6124), .A2(n5716), .ZN(n7443) );
  NOR2_X1 U4337 ( .A1(n7182), .A2(n4921), .ZN(n7172) );
  OR2_X1 U4338 ( .A1(n4920), .A2(n4919), .ZN(n7196) );
  INV_X1 U4339 ( .A(n5015), .ZN(n5068) );
  NAND2_X1 U4340 ( .A1(n4860), .A2(n4859), .ZN(n5014) );
  OR2_X1 U4341 ( .A1(n7289), .A2(n4947), .ZN(n7294) );
  NAND2_X1 U4342 ( .A1(n4832), .A2(n5575), .ZN(n6509) );
  OR2_X1 U4343 ( .A1(n4986), .A2(n4973), .ZN(n7342) );
  INV_X1 U4344 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5348) );
  INV_X1 U4345 ( .A(n7731), .ZN(n5793) );
  NAND2_X1 U4346 ( .A1(n5354), .A2(n7554), .ZN(n7643) );
  OR2_X1 U4347 ( .A1(n5280), .A2(n4308), .ZN(n5627) );
  NAND2_X1 U4348 ( .A1(n5319), .A2(n4308), .ZN(n5914) );
  AND2_X1 U4349 ( .A1(n5318), .A2(n5317), .ZN(n7720) );
  AOI22_X1 U4350 ( .A1(n5580), .A2(n5584), .B1(n5874), .B2(n5579), .ZN(n7713)
         );
  INV_X1 U4351 ( .A(n5773), .ZN(n7673) );
  NAND2_X1 U4352 ( .A1(n5163), .A2(n7554), .ZN(n5537) );
  OR2_X1 U4353 ( .A1(n5238), .A2(n7554), .ZN(n5271) );
  INV_X1 U4354 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7534) );
  NOR2_X4 U4355 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U4356 ( .A1(n3703), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3987), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3838) );
  AND2_X4 U4357 ( .A1(n4905), .A2(n3839), .ZN(n4784) );
  AOI22_X1 U4358 ( .A1(n4784), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3837) );
  AND2_X4 U4359 ( .A1(n4912), .A2(n3840), .ZN(n4564) );
  AOI22_X1 U4360 ( .A1(n4564), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3836) );
  INV_X2 U4361 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3834) );
  AND2_X2 U4362 ( .A1(n5123), .A2(n4906), .ZN(n3939) );
  AND2_X2 U4363 ( .A1(n3839), .A2(n4906), .ZN(n4022) );
  AOI22_X1 U4364 ( .A1(n3939), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3835) );
  AND2_X2 U4365 ( .A1(n5123), .A2(n4905), .ZN(n4114) );
  AOI22_X1 U4366 ( .A1(n4114), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3844) );
  AND2_X4 U4367 ( .A1(n3840), .A2(n4906), .ZN(n3986) );
  AOI22_X1 U4368 ( .A1(n3678), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4369 ( .A1(n3999), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3841) );
  AND2_X2 U4370 ( .A1(n3846), .A2(n3845), .ZN(n3905) );
  AOI22_X1 U4371 ( .A1(n4784), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4372 ( .A1(n4564), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4373 ( .A1(n3939), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4374 ( .A1(n4114), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4375 ( .A1(n4411), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4376 ( .A1(n3677), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4377 ( .A1(n3999), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3851) );
  NAND2_X1 U4378 ( .A1(n3699), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4379 ( .A1(n4001), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U4380 ( .A1(n3702), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4381 ( .A1(n4564), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4382 ( .A1(n4582), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3863)
         );
  NAND2_X1 U4383 ( .A1(n4022), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4384 ( .A1(n3939), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3861)
         );
  NAND3_X1 U4385 ( .A1(n3715), .A2(n3864), .A3(n3827), .ZN(n3876) );
  NAND2_X1 U4386 ( .A1(n4114), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3868) );
  NAND2_X1 U4387 ( .A1(n3999), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3867) );
  NAND2_X1 U4388 ( .A1(n3701), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4389 ( .A1(n3925), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3865)
         );
  NAND2_X1 U4390 ( .A1(n4411), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3872)
         );
  NAND2_X1 U4391 ( .A1(n3700), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4392 ( .A1(n4088), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3870) );
  NAND2_X1 U4393 ( .A1(n3704), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4394 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  NOR2_X2 U4395 ( .A1(n3876), .A2(n3875), .ZN(n3900) );
  AOI22_X1 U4396 ( .A1(n3939), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4397 ( .A1(n3678), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4398 ( .A1(n4114), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4399 ( .A1(n3987), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4400 ( .A1(n4411), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4401 ( .A1(n4564), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4402 ( .A1(n3999), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4403 ( .A1(n3703), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3881) );
  OAI21_X1 U4404 ( .B1(n4039), .B2(n5165), .A(n3970), .ZN(n3898) );
  AOI22_X1 U4405 ( .A1(n3999), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4406 ( .A1(n3677), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4407 ( .A1(n4752), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4408 ( .A1(n4564), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4409 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3897)
         );
  AOI22_X1 U4410 ( .A1(n4411), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4411 ( .A1(n3920), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3987), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4412 ( .A1(n3668), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4413 ( .A1(n3891), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4414 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  INV_X2 U4415 ( .A(n5214), .ZN(n4957) );
  NAND2_X1 U4416 ( .A1(n3898), .A2(n4957), .ZN(n3904) );
  NOR2_X1 U4417 ( .A1(n3671), .A2(n3899), .ZN(n3902) );
  INV_X1 U4418 ( .A(n4302), .ZN(n3901) );
  AOI21_X2 U4419 ( .B1(n3900), .B2(n4031), .A(n3901), .ZN(n3963) );
  NAND3_X1 U4420 ( .A1(n3902), .A2(n5214), .A3(n3963), .ZN(n3903) );
  NAND2_X1 U4421 ( .A1(n3904), .A2(n3903), .ZN(n4038) );
  AOI22_X1 U4422 ( .A1(n3678), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4423 ( .A1(n3920), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3987), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4424 ( .A1(n3695), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4425 ( .A1(n3891), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4426 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3915)
         );
  AOI22_X1 U4427 ( .A1(n3698), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4428 ( .A1(n4411), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4429 ( .A1(n3999), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4430 ( .A1(n4564), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4431 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  NAND2_X1 U4432 ( .A1(n4038), .A2(n4036), .ZN(n3938) );
  NAND2_X1 U4433 ( .A1(n4411), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3919)
         );
  NAND2_X1 U4434 ( .A1(n3673), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U4435 ( .A1(n3678), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3917) );
  NAND2_X1 U4436 ( .A1(n3986), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4437 ( .A1(n4001), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3924)
         );
  NAND2_X1 U4438 ( .A1(n4564), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U4439 ( .A1(n3703), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4440 ( .A1(n3987), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3921) );
  NAND2_X1 U4441 ( .A1(n3668), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4442 ( .A1(n3999), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3928) );
  NAND2_X1 U4443 ( .A1(n4610), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3927)
         );
  NAND2_X1 U4444 ( .A1(n3925), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3926)
         );
  NAND2_X1 U4445 ( .A1(n3697), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3933)
         );
  NAND2_X1 U4446 ( .A1(n4784), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4447 ( .A1(n4022), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4448 ( .A1(n4582), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3930)
         );
  NAND4_X4 U4449 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n5721)
         );
  NAND2_X1 U4450 ( .A1(n3938), .A2(n3971), .ZN(n3960) );
  NAND2_X1 U4451 ( .A1(n4411), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3943)
         );
  NAND2_X1 U4452 ( .A1(n4610), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3942)
         );
  NAND2_X1 U4453 ( .A1(n3677), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4454 ( .A1(n3939), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3940)
         );
  NAND2_X1 U4455 ( .A1(n4564), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U4456 ( .A1(n3920), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4457 ( .A1(n3987), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4458 ( .A1(n4022), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U4459 ( .A1(n3999), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3951) );
  NAND2_X1 U4460 ( .A1(n3668), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4461 ( .A1(n3673), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3949) );
  NAND2_X1 U4462 ( .A1(n3925), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3948)
         );
  NAND2_X1 U4463 ( .A1(n4582), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3954)
         );
  NAND2_X1 U4464 ( .A1(n3705), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3953) );
  NAND3_X1 U4465 ( .A1(n3954), .A2(n3953), .A3(n3952), .ZN(n3955) );
  NAND2_X1 U4466 ( .A1(n3960), .A2(n5752), .ZN(n3983) );
  INV_X1 U4467 ( .A(n3983), .ZN(n3967) );
  INV_X1 U4468 ( .A(n4866), .ZN(n3962) );
  XNOR2_X1 U4469 ( .A(n7098), .B(STATE_REG_2__SCAN_IN), .ZN(n4822) );
  INV_X1 U4470 ( .A(n4034), .ZN(n4299) );
  NAND2_X1 U4471 ( .A1(n4865), .A2(n3899), .ZN(n3974) );
  OAI211_X1 U4472 ( .C1(n4042), .C2(n5165), .A(n3969), .B(n3974), .ZN(n3961)
         );
  AOI21_X1 U4473 ( .B1(n7304), .B2(n3962), .A(n3961), .ZN(n3965) );
  INV_X1 U4474 ( .A(n4294), .ZN(n3964) );
  NAND2_X1 U4475 ( .A1(n6081), .A2(n3966), .ZN(n4802) );
  MUX2_X1 U4476 ( .A(n4802), .B(n4293), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3968) );
  NAND2_X1 U4477 ( .A1(n6081), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7527) );
  AOI21_X1 U4478 ( .B1(n5214), .B2(n5721), .A(n7527), .ZN(n3973) );
  NAND3_X1 U4479 ( .A1(n4868), .A2(n4957), .A3(n3971), .ZN(n3972) );
  INV_X1 U4480 ( .A(n4980), .ZN(n5132) );
  AND3_X1 U4481 ( .A1(n3969), .A2(n3973), .A3(n5132), .ZN(n3981) );
  AND2_X1 U4482 ( .A1(n4866), .A2(n4033), .ZN(n3978) );
  INV_X1 U4483 ( .A(n3974), .ZN(n3975) );
  OAI21_X1 U4484 ( .B1(n3976), .B2(n3975), .A(n5206), .ZN(n3977) );
  INV_X1 U4485 ( .A(n3979), .ZN(n3980) );
  NAND2_X1 U4486 ( .A1(n4233), .A2(n5050), .ZN(n3982) );
  NAND2_X1 U4487 ( .A1(n3983), .A2(n3982), .ZN(n4874) );
  INV_X1 U4488 ( .A(n4053), .ZN(n3985) );
  XNOR2_X1 U4489 ( .A(n4052), .B(n3985), .ZN(n4309) );
  INV_X1 U4490 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4491 ( .A1(n4779), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4492 ( .A1(n4730), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4493 ( .A1(n4710), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4494 ( .A1(n3698), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4495 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3998)
         );
  AOI22_X1 U4496 ( .A1(n4569), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3996) );
  BUF_X1 U4497 ( .A(n3668), .Z(n4000) );
  AOI22_X1 U4498 ( .A1(n4000), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4610), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4499 ( .A1(n4757), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4500 ( .A1(n4784), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4501 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3997)
         );
  AOI21_X1 U4502 ( .B1(n5050), .B2(n4213), .A(n3966), .ZN(n4013) );
  AOI22_X1 U4503 ( .A1(n4779), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4504 ( .A1(n4730), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4505 ( .A1(n4710), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4506 ( .A1(n3992), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4507 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4011)
         );
  AOI22_X1 U4508 ( .A1(n4569), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4509 ( .A1(n4610), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4510 ( .A1(n4711), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4511 ( .A1(n3986), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4512 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  NAND2_X1 U4513 ( .A1(n3971), .A2(n4066), .ZN(n4012) );
  OAI211_X1 U4514 ( .C1(n4274), .C2(n4014), .A(n4013), .B(n4012), .ZN(n4062)
         );
  XNOR2_X1 U4515 ( .A(n4213), .B(n4066), .ZN(n4015) );
  NOR2_X1 U4516 ( .A1(n4015), .A2(n4087), .ZN(n4061) );
  NAND2_X1 U4517 ( .A1(n4062), .A2(n4061), .ZN(n4016) );
  INV_X1 U4518 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4017) );
  NOR2_X1 U4519 ( .A1(n4274), .A2(n4017), .ZN(n4030) );
  AOI22_X1 U4520 ( .A1(n3696), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4521 ( .A1(n4710), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4522 ( .A1(n4569), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4523 ( .A1(n3992), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4524 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4028)
         );
  AOI22_X1 U4525 ( .A1(n4779), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4526 ( .A1(n3891), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4527 ( .A1(n3705), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4528 ( .A1(n4730), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4529 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  OAI21_X1 U4530 ( .B1(n4055), .B2(n4086), .A(n4087), .ZN(n4029) );
  NOR2_X1 U4531 ( .A1(n5049), .A2(n5214), .ZN(n4032) );
  NAND2_X1 U4532 ( .A1(n4858), .A2(n5721), .ZN(n4853) );
  NOR2_X1 U4533 ( .A1(n4034), .A2(n5721), .ZN(n4035) );
  AND2_X1 U4534 ( .A1(n4036), .A2(n4035), .ZN(n4037) );
  NAND3_X1 U4535 ( .A1(n3900), .A2(n4868), .A3(n4957), .ZN(n5052) );
  INV_X1 U4536 ( .A(n5052), .ZN(n4041) );
  INV_X1 U4537 ( .A(n4039), .ZN(n4040) );
  NAND3_X1 U4538 ( .A1(n4041), .A2(n4040), .A3(n6103), .ZN(n4971) );
  NAND2_X1 U4539 ( .A1(n4043), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4048) );
  NAND2_X1 U4540 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4079) );
  OAI21_X1 U4541 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4079), .ZN(n5652) );
  OR2_X1 U4542 ( .A1(n4802), .A2(n5652), .ZN(n4045) );
  INV_X1 U4543 ( .A(n4293), .ZN(n4110) );
  NAND2_X1 U4544 ( .A1(n4110), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4044) );
  INV_X1 U4545 ( .A(n4049), .ZN(n4046) );
  NAND2_X1 U4546 ( .A1(n3666), .A2(n4047), .ZN(n4051) );
  INV_X1 U4547 ( .A(n4077), .ZN(n4050) );
  NAND2_X1 U4548 ( .A1(n4053), .A2(n4052), .ZN(n4073) );
  XNOR2_X1 U4549 ( .A(n4072), .B(n4073), .ZN(n4903) );
  OR2_X2 U4550 ( .A1(n4056), .A2(n4064), .ZN(n4057) );
  NAND2_X1 U4551 ( .A1(n4066), .A2(n4058), .ZN(n4132) );
  OAI211_X1 U4552 ( .C1(n4066), .C2(n4058), .A(n7304), .B(n4132), .ZN(n4059)
         );
  NAND3_X1 U4553 ( .A1(n4059), .A2(n4957), .A3(n5165), .ZN(n4060) );
  XNOR2_X1 U4554 ( .A(n4070), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4953)
         );
  NOR2_X1 U4555 ( .A1(n4062), .A2(n4061), .ZN(n4063) );
  OR2_X1 U4556 ( .A1(n4308), .A2(n4210), .ZN(n4069) );
  NAND2_X1 U4557 ( .A1(n3971), .A2(n5170), .ZN(n4103) );
  OAI21_X1 U4558 ( .B1(n4065), .B2(n4066), .A(n4103), .ZN(n4067) );
  INV_X1 U4559 ( .A(n4067), .ZN(n4068) );
  NAND2_X1 U4560 ( .A1(n4069), .A2(n4068), .ZN(n4940) );
  INV_X1 U4561 ( .A(n4070), .ZN(n4071) );
  AOI22_X2 U4562 ( .A1(n4953), .A2(n4954), .B1(n4071), .B2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4106) );
  INV_X1 U4563 ( .A(n4072), .ZN(n4074) );
  INV_X1 U4564 ( .A(n4079), .ZN(n4078) );
  NAND2_X1 U4565 ( .A1(n4078), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U4566 ( .A1(n4079), .A2(n7501), .ZN(n4080) );
  NAND2_X1 U4567 ( .A1(n5234), .A2(n4080), .ZN(n5193) );
  OAI22_X1 U4568 ( .A1(n5193), .A2(n4802), .B1(n4293), .B2(n7501), .ZN(n4081)
         );
  NAND2_X1 U4569 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  NAND2_X1 U4570 ( .A1(n3665), .A2(n3966), .ZN(n4100) );
  AOI22_X1 U4571 ( .A1(n4569), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4572 ( .A1(n3986), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4752), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4573 ( .A1(n3891), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U4574 ( .A1(n4730), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U4575 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4098)
         );
  AOI22_X1 U4576 ( .A1(n4000), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U4577 ( .A1(n4779), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4578 ( .A1(n4757), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4579 ( .A1(n4710), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U4580 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4097)
         );
  AOI22_X1 U4581 ( .A1(n4234), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4290), 
        .B2(n4130), .ZN(n4099) );
  XNOR2_X1 U4582 ( .A(n4132), .B(n4130), .ZN(n4104) );
  OAI21_X1 U4583 ( .B1(n4104), .B2(n4065), .A(n4103), .ZN(n4105) );
  AOI21_X1 U4584 ( .B1(n3706), .B2(n4233), .A(n4105), .ZN(n5081) );
  INV_X1 U4585 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U4586 ( .A1(n4107), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4113) );
  INV_X1 U4587 ( .A(n5234), .ZN(n4108) );
  NAND2_X1 U4588 ( .A1(n4108), .A2(n7506), .ZN(n5742) );
  NAND2_X1 U4589 ( .A1(n5234), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4109) );
  NAND2_X1 U4590 ( .A1(n5742), .A2(n4109), .ZN(n5653) );
  INV_X1 U4591 ( .A(n4802), .ZN(n4111) );
  AOI22_X1 U4592 ( .A1(n5653), .A2(n4111), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4110), .ZN(n4112) );
  NAND2_X1 U4593 ( .A1(n5854), .A2(n3966), .ZN(n4126) );
  AOI22_X1 U4594 ( .A1(n4000), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4595 ( .A1(n4569), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4596 ( .A1(n3992), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U4597 ( .A1(n4779), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U4598 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4124)
         );
  AOI22_X1 U4599 ( .A1(n4730), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U4600 ( .A1(n4710), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U4601 ( .A1(n4751), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U4602 ( .A1(n3698), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U4603 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  AOI22_X1 U4604 ( .A1(n4234), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4290), 
        .B2(n4133), .ZN(n4125) );
  NAND2_X1 U4605 ( .A1(n4126), .A2(n4125), .ZN(n4137) );
  NOR2_X1 U4606 ( .A1(n4130), .A2(n4133), .ZN(n4129) );
  AOI21_X1 U4607 ( .B1(n4129), .B2(n4132), .A(n4065), .ZN(n4135) );
  INV_X1 U4608 ( .A(n4130), .ZN(n4131) );
  NAND2_X1 U4609 ( .A1(n4132), .A2(n4131), .ZN(n4134) );
  NAND2_X1 U4610 ( .A1(n4134), .A2(n4133), .ZN(n4157) );
  AOI22_X1 U4611 ( .A1(n3664), .A2(n4233), .B1(n4135), .B2(n4157), .ZN(n5509)
         );
  INV_X1 U4612 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5515) );
  INV_X1 U4613 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U4614 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4000), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4615 ( .A1(n4569), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U4616 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3992), .B1(n3705), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4617 ( .A1(n4779), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U4618 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4148)
         );
  AOI22_X1 U4619 ( .A1(n4564), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4711), .B1(n4710), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U4621 ( .A1(n4784), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U4622 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4752), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U4623 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4147)
         );
  NAND2_X1 U4624 ( .A1(n4290), .A2(n4158), .ZN(n4149) );
  INV_X1 U4625 ( .A(n4151), .ZN(n4154) );
  INV_X1 U4626 ( .A(n4152), .ZN(n4153) );
  NAND2_X1 U4627 ( .A1(n4154), .A2(n4153), .ZN(n4155) );
  INV_X1 U4628 ( .A(n4157), .ZN(n4159) );
  INV_X1 U4629 ( .A(n4158), .ZN(n4156) );
  OR2_X1 U4630 ( .A1(n4157), .A2(n4156), .ZN(n4197) );
  OAI211_X1 U4631 ( .C1(n4159), .C2(n4158), .A(n7304), .B(n4197), .ZN(n4160)
         );
  INV_X1 U4632 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U4633 ( .A1(n4000), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U4634 ( .A1(n4569), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4635 ( .A1(n3992), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4636 ( .A1(n4779), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4164) );
  NAND4_X1 U4637 ( .A1(n4167), .A2(n4166), .A3(n4165), .A4(n4164), .ZN(n4173)
         );
  AOI22_X1 U4638 ( .A1(n4730), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U4639 ( .A1(n4710), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4640 ( .A1(n4784), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4641 ( .A1(n3698), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U4642 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4172)
         );
  XNOR2_X1 U4643 ( .A(n4179), .B(n4178), .ZN(n4340) );
  INV_X1 U4644 ( .A(n4197), .ZN(n4174) );
  XNOR2_X1 U4645 ( .A(n4174), .B(n4195), .ZN(n4175) );
  OAI22_X1 U4646 ( .A1(n4340), .A2(n4210), .B1(n4175), .B2(n4065), .ZN(n4176)
         );
  XNOR2_X1 U4647 ( .A(n4176), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5629)
         );
  INV_X1 U4648 ( .A(n4176), .ZN(n4177) );
  INV_X1 U4649 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5337) );
  AOI22_X1 U4650 ( .A1(n4000), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U4651 ( .A1(n4569), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U4652 ( .A1(n3992), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U4653 ( .A1(n4779), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4180) );
  NAND4_X1 U4654 ( .A1(n4183), .A2(n4182), .A3(n4181), .A4(n4180), .ZN(n4189)
         );
  AOI22_X1 U4655 ( .A1(n4730), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4656 ( .A1(n4710), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4657 ( .A1(n4784), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4658 ( .A1(n3698), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U4659 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4188)
         );
  INV_X1 U4660 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4192) );
  INV_X1 U4661 ( .A(n4190), .ZN(n4191) );
  OAI21_X1 U4662 ( .B1(n4274), .B2(n4192), .A(n4191), .ZN(n4193) );
  NAND3_X1 U4663 ( .A1(n4212), .A2(n3833), .A3(n4233), .ZN(n4203) );
  INV_X1 U4664 ( .A(n4195), .ZN(n4196) );
  NOR2_X1 U4665 ( .A1(n4197), .A2(n4196), .ZN(n4199) );
  NOR2_X1 U4666 ( .A1(n4199), .A2(n4198), .ZN(n4200) );
  NAND2_X1 U4667 ( .A1(n3828), .A2(n4201), .ZN(n4202) );
  XOR2_X1 U4668 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .B(n4204), .Z(n5804) );
  AOI22_X1 U4669 ( .A1(n4234), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4290), 
        .B2(n4213), .ZN(n4205) );
  XOR2_X1 U4670 ( .A(n4213), .B(n3828), .Z(n4206) );
  OAI22_X1 U4671 ( .A1(n4358), .A2(n4210), .B1(n4206), .B2(n4065), .ZN(n4207)
         );
  XNOR2_X1 U4672 ( .A(n4207), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5935)
         );
  INV_X1 U4673 ( .A(n4207), .ZN(n4208) );
  INV_X1 U4674 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5560) );
  INV_X1 U4675 ( .A(n4213), .ZN(n4209) );
  NAND2_X4 U4676 ( .A1(n4212), .A2(n4211), .ZN(n6697) );
  NAND2_X1 U4677 ( .A1(n7304), .A2(n4213), .ZN(n4214) );
  OR2_X1 U4678 ( .A1(n3828), .A2(n4214), .ZN(n4215) );
  NAND2_X1 U4679 ( .A1(n6697), .A2(n4215), .ZN(n4217) );
  INV_X1 U4680 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4216) );
  XNOR2_X1 U4681 ( .A(n4217), .B(n4216), .ZN(n5951) );
  INV_X1 U4682 ( .A(n4217), .ZN(n4218) );
  XOR2_X1 U4683 ( .A(n6697), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .Z(n5962) );
  INV_X1 U4684 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6551) );
  XNOR2_X1 U4685 ( .A(n6697), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5989)
         );
  XOR2_X1 U4686 ( .A(n6697), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n6543) );
  INV_X1 U4687 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6752) );
  XNOR2_X1 U4688 ( .A(n6697), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6538)
         );
  XNOR2_X1 U4689 ( .A(n6697), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6529)
         );
  INV_X1 U4690 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6730) );
  XNOR2_X1 U4691 ( .A(n6697), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6520)
         );
  INV_X1 U4692 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6712) );
  XNOR2_X1 U4693 ( .A(n6697), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6510)
         );
  INV_X1 U4694 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7335) );
  AND2_X1 U4695 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6554) );
  NOR4_X1 U4696 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4225) );
  NOR2_X1 U4697 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U4698 ( .A1(n4225), .A2(n6446), .ZN(n4226) );
  AND2_X1 U4699 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6565) );
  AND2_X1 U4700 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6572) );
  AND2_X1 U4701 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U4702 ( .A1(n6441), .A2(n3832), .ZN(n4227) );
  XOR2_X1 U4703 ( .A(n6697), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n6434) );
  INV_X1 U4704 ( .A(n6434), .ZN(n4228) );
  INV_X1 U4705 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U4706 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6602) );
  INV_X1 U4707 ( .A(n6602), .ZN(n6593) );
  NAND3_X1 U4708 ( .A1(n6399), .A2(n6593), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4231) );
  OR2_X1 U4709 ( .A1(n6697), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6395)
         );
  INV_X1 U4710 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6416) );
  INV_X1 U4711 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4229) );
  NAND2_X1 U4712 ( .A1(n6416), .A2(n4229), .ZN(n6601) );
  NOR2_X1 U4713 ( .A1(n6397), .A2(n6697), .ZN(n4230) );
  AOI21_X2 U4714 ( .B1(n4231), .B2(n6395), .A(n4230), .ZN(n4232) );
  XNOR2_X1 U4715 ( .A(n4232), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6583)
         );
  NAND2_X1 U4716 ( .A1(n5348), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U4717 ( .A1(n4914), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U4718 ( .A1(n4254), .A2(n4235), .ZN(n4236) );
  NAND2_X1 U4719 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7557), .ZN(n4241) );
  NAND2_X1 U4720 ( .A1(n4236), .A2(n4241), .ZN(n4237) );
  NAND2_X1 U4721 ( .A1(n4255), .A2(n4237), .ZN(n4845) );
  INV_X1 U4722 ( .A(n4845), .ZN(n4240) );
  NAND2_X1 U4723 ( .A1(n4240), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U4724 ( .A1(n4276), .A2(n4238), .ZN(n4251) );
  NAND2_X1 U4725 ( .A1(n4290), .A2(n5206), .ZN(n4239) );
  OAI211_X1 U4726 ( .C1(n4274), .C2(n4240), .A(n5165), .B(n4239), .ZN(n4250)
         );
  OAI21_X1 U4727 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7557), .A(n4241), 
        .ZN(n4246) );
  INV_X1 U4728 ( .A(n4246), .ZN(n4244) );
  INV_X1 U4729 ( .A(n4242), .ZN(n4243) );
  AOI21_X1 U4730 ( .B1(n4034), .B2(n4244), .A(n4243), .ZN(n4245) );
  AOI21_X1 U4731 ( .B1(n3900), .B2(n5721), .A(n5206), .ZN(n4265) );
  OR2_X1 U4732 ( .A1(n4245), .A2(n4265), .ZN(n4249) );
  INV_X1 U4733 ( .A(n4290), .ZN(n4247) );
  OAI21_X1 U4734 ( .B1(n4247), .B2(n4246), .A(n4276), .ZN(n4248) );
  OAI211_X1 U4735 ( .C1(n4251), .C2(n4250), .A(n4249), .B(n4248), .ZN(n4253)
         );
  NAND2_X1 U4736 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  NAND2_X1 U4737 ( .A1(n4253), .A2(n4252), .ZN(n4270) );
  NAND2_X1 U4738 ( .A1(n4255), .A2(n4254), .ZN(n4258) );
  NAND2_X1 U4739 ( .A1(n7501), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U4740 ( .A1(n3834), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U4741 ( .A1(n4258), .A2(n4257), .ZN(n4262) );
  OAI21_X1 U4742 ( .B1(n4258), .B2(n4257), .A(n4262), .ZN(n4844) );
  INV_X1 U4743 ( .A(n4844), .ZN(n4264) );
  NAND2_X1 U4744 ( .A1(n4290), .A2(n4264), .ZN(n4260) );
  INV_X1 U4745 ( .A(n4265), .ZN(n4259) );
  OAI211_X1 U4746 ( .C1(n4274), .C2(n4264), .A(n4260), .B(n4259), .ZN(n4269)
         );
  NAND2_X1 U4747 ( .A1(n4262), .A2(n4261), .ZN(n4273) );
  XNOR2_X1 U4748 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4263) );
  XNOR2_X1 U4749 ( .A(n4273), .B(n4263), .ZN(n4846) );
  INV_X1 U4750 ( .A(n4846), .ZN(n4267) );
  NAND3_X1 U4751 ( .A1(n4265), .A2(n4264), .A3(n4290), .ZN(n4266) );
  OAI21_X1 U4752 ( .B1(n4276), .B2(n4267), .A(n4266), .ZN(n4268) );
  AOI21_X1 U4753 ( .B1(n4270), .B2(n4269), .A(n4268), .ZN(n4279) );
  OR2_X1 U4754 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n7506), .ZN(n4272)
         );
  NOR2_X1 U4755 ( .A1(n5116), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4271)
         );
  AOI21_X1 U4756 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4280) );
  AND2_X1 U4757 ( .A1(n4280), .A2(n4281), .ZN(n4849) );
  OAI21_X1 U4758 ( .B1(n4849), .B2(n4846), .A(n4274), .ZN(n4275) );
  INV_X1 U4759 ( .A(n4275), .ZN(n4278) );
  AOI22_X1 U4760 ( .A1(n4287), .A2(n4849), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n3966), .ZN(n4277) );
  OAI21_X1 U4761 ( .B1(n4279), .B2(n4278), .A(n4277), .ZN(n4289) );
  INV_X1 U4762 ( .A(n4280), .ZN(n4283) );
  INV_X1 U4763 ( .A(n4281), .ZN(n4282) );
  NAND2_X1 U4764 ( .A1(n4283), .A2(n4282), .ZN(n4286) );
  INV_X1 U4765 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U4766 ( .A1(n4284), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U4767 ( .A1(n4286), .A2(n4285), .ZN(n4848) );
  NAND2_X1 U4768 ( .A1(n4287), .A2(n4848), .ZN(n4288) );
  NAND2_X1 U4769 ( .A1(n4289), .A2(n4288), .ZN(n4292) );
  NAND2_X1 U4770 ( .A1(n4290), .A2(n4848), .ZN(n4291) );
  NAND2_X1 U4771 ( .A1(n4293), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U4772 ( .A1(n5165), .A2(n3899), .ZN(n4296) );
  INV_X1 U4773 ( .A(n4960), .ZN(n4297) );
  AND2_X1 U4774 ( .A1(n4297), .A2(n3971), .ZN(n4298) );
  NOR2_X1 U4775 ( .A1(n4294), .A2(n4298), .ZN(n4879) );
  NAND2_X1 U4776 ( .A1(n4879), .A2(n4299), .ZN(n7509) );
  OR2_X1 U4777 ( .A1(n6583), .A2(n7482), .ZN(n4812) );
  NAND2_X1 U4778 ( .A1(n7522), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4498) );
  NAND2_X1 U4779 ( .A1(n3689), .A2(n4480), .ZN(n4307) );
  OR2_X1 U4780 ( .A1(n4039), .A2(n7522), .ZN(n4336) );
  NAND2_X1 U4781 ( .A1(n4312), .A2(EAX_REG_1__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U4782 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4303)
         );
  OAI211_X1 U4783 ( .C1(n4336), .C2(n4914), .A(n4304), .B(n4303), .ZN(n4305)
         );
  INV_X1 U4784 ( .A(n4305), .ZN(n4306) );
  NAND2_X1 U4785 ( .A1(n4307), .A2(n4306), .ZN(n5060) );
  NAND2_X1 U4786 ( .A1(n4308), .A2(n3671), .ZN(n4944) );
  NAND2_X1 U4787 ( .A1(n4310), .A2(n4480), .ZN(n4317) );
  NAND2_X1 U4788 ( .A1(n4312), .A2(EAX_REG_0__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U4789 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4313)
         );
  OAI211_X1 U4790 ( .C1(n4336), .C2(n4311), .A(n4314), .B(n4313), .ZN(n4315)
         );
  INV_X1 U4791 ( .A(n4315), .ZN(n4316) );
  NAND2_X1 U4792 ( .A1(n4317), .A2(n4316), .ZN(n4943) );
  AND2_X1 U4793 ( .A1(n4943), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U4794 ( .A1(n4944), .A2(n4318), .ZN(n4942) );
  OR2_X1 U4795 ( .A1(n4943), .A2(n5704), .ZN(n4319) );
  NAND2_X1 U4796 ( .A1(n4942), .A2(n4319), .ZN(n5059) );
  AND2_X2 U4797 ( .A1(n5060), .A2(n5059), .ZN(n5076) );
  NAND2_X1 U4798 ( .A1(n5077), .A2(n5076), .ZN(n4323) );
  NAND2_X1 U4799 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4326) );
  OAI21_X1 U4800 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4326), .ZN(n6292) );
  AOI22_X1 U4801 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4798), 
        .B2(n6292), .ZN(n4321) );
  NAND2_X1 U4802 ( .A1(n4766), .A2(EAX_REG_2__SCAN_IN), .ZN(n4320) );
  OAI211_X1 U4803 ( .C1(n4336), .C2(n3834), .A(n4321), .B(n4320), .ZN(n5075)
         );
  INV_X1 U4804 ( .A(n5075), .ZN(n4322) );
  NAND2_X1 U4805 ( .A1(n4323), .A2(n4322), .ZN(n4325) );
  NAND2_X1 U4806 ( .A1(n4766), .A2(EAX_REG_3__SCAN_IN), .ZN(n4330) );
  INV_X1 U4807 ( .A(n4326), .ZN(n4328) );
  INV_X1 U4808 ( .A(n4333), .ZN(n4327) );
  OAI21_X1 U4809 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4328), .A(n4327), 
        .ZN(n5844) );
  AOI22_X1 U4810 ( .A1(n4798), .A2(n5844), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4329) );
  OAI211_X1 U4811 ( .C1(n4336), .C2(n5116), .A(n4330), .B(n4329), .ZN(n4331)
         );
  AOI21_X1 U4812 ( .B1(n3664), .B2(n4480), .A(n4331), .ZN(n5111) );
  OAI21_X1 U4813 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4333), .A(n4342), 
        .ZN(n5644) );
  NAND2_X1 U4814 ( .A1(n4766), .A2(EAX_REG_4__SCAN_IN), .ZN(n4335) );
  OAI21_X1 U4815 ( .B1(n7303), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7522), 
        .ZN(n4334) );
  OAI211_X1 U4816 ( .C1(n4336), .C2(n7490), .A(n4335), .B(n4334), .ZN(n4337)
         );
  OAI21_X1 U4817 ( .B1(n5704), .B2(n5644), .A(n4337), .ZN(n4338) );
  NAND2_X1 U4818 ( .A1(n5113), .A2(n5156), .ZN(n5155) );
  INV_X1 U4819 ( .A(n4340), .ZN(n4347) );
  INV_X1 U4820 ( .A(n4349), .ZN(n4350) );
  INV_X1 U4821 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U4822 ( .A1(n4343), .A2(n4342), .ZN(n4344) );
  NAND2_X1 U4823 ( .A1(n4350), .A2(n4344), .ZN(n7374) );
  AOI22_X1 U4824 ( .A1(n7374), .A2(n4798), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4345) );
  OAI21_X1 U4825 ( .B1(n4348), .B2(n7181), .A(n4345), .ZN(n4346) );
  INV_X1 U4826 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4864) );
  INV_X1 U4827 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7379) );
  OAI22_X1 U4828 ( .A1(n4348), .A2(n4864), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7379), .ZN(n4354) );
  INV_X1 U4829 ( .A(n4359), .ZN(n4352) );
  NAND2_X1 U4830 ( .A1(n4350), .A2(n7379), .ZN(n4351) );
  NAND2_X1 U4831 ( .A1(n4352), .A2(n4351), .ZN(n7384) );
  AND2_X1 U4832 ( .A1(n7384), .A2(n4798), .ZN(n4353) );
  AOI21_X1 U4833 ( .B1(n4354), .B2(n5704), .A(n4353), .ZN(n4355) );
  OAI21_X1 U4834 ( .B1(n4359), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4380), 
        .ZN(n7397) );
  NAND2_X1 U4835 ( .A1(n7397), .A2(n4798), .ZN(n4361) );
  NAND2_X1 U4836 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4360)
         );
  NAND2_X1 U4837 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  AOI21_X1 U4838 ( .B1(n4766), .B2(EAX_REG_7__SCAN_IN), .A(n4362), .ZN(n4363)
         );
  AOI21_X2 U4839 ( .B1(n4365), .B2(n4480), .A(n4364), .ZN(n5557) );
  AOI22_X1 U4840 ( .A1(n4710), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4841 ( .A1(n4779), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4842 ( .A1(n3992), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U4843 ( .A1(n4752), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4366) );
  NAND4_X1 U4844 ( .A1(n4369), .A2(n4368), .A3(n4367), .A4(n4366), .ZN(n4375)
         );
  AOI22_X1 U4845 ( .A1(n4000), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4846 ( .A1(n4569), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U4847 ( .A1(n4730), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U4848 ( .A1(n3705), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4370) );
  NAND4_X1 U4849 ( .A1(n4373), .A2(n4372), .A3(n4371), .A4(n4370), .ZN(n4374)
         );
  OAI21_X1 U4850 ( .B1(n4375), .B2(n4374), .A(n4480), .ZN(n4379) );
  NAND2_X1 U4851 ( .A1(n4766), .A2(EAX_REG_8__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U4852 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4377)
         );
  XNOR2_X1 U4853 ( .A(n4380), .B(n5952), .ZN(n5714) );
  NAND2_X1 U4854 ( .A1(n5714), .A2(n4798), .ZN(n4376) );
  NAND4_X1 U4855 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(n5698)
         );
  XOR2_X1 U4856 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4394), .Z(n5968) );
  AOI22_X1 U4857 ( .A1(n4766), .A2(EAX_REG_9__SCAN_IN), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4858 ( .A1(n4779), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4859 ( .A1(n3992), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4860 ( .A1(n4710), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4861 ( .A1(n4730), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4381) );
  NAND4_X1 U4862 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4390)
         );
  AOI22_X1 U4863 ( .A1(n4000), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4864 ( .A1(n4569), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4865 ( .A1(n3674), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U4866 ( .A1(n4711), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4385) );
  NAND4_X1 U4867 ( .A1(n4388), .A2(n4387), .A3(n4386), .A4(n4385), .ZN(n4389)
         );
  OAI21_X1 U4868 ( .B1(n4390), .B2(n4389), .A(n4480), .ZN(n4391) );
  OAI211_X1 U4869 ( .C1(n5968), .C2(n5704), .A(n4392), .B(n4391), .ZN(n4393)
         );
  INV_X1 U4870 ( .A(n4393), .ZN(n5827) );
  XNOR2_X1 U4871 ( .A(n4410), .B(n4409), .ZN(n5992) );
  AOI22_X1 U4872 ( .A1(n4779), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U4873 ( .A1(n4730), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4874 ( .A1(n4757), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4875 ( .A1(n4752), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4395) );
  NAND4_X1 U4876 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(n4404)
         );
  AOI22_X1 U4877 ( .A1(n4569), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U4878 ( .A1(n4710), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4879 ( .A1(n4000), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4880 ( .A1(n3986), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4399) );
  NAND4_X1 U4881 ( .A1(n4402), .A2(n4401), .A3(n4400), .A4(n4399), .ZN(n4403)
         );
  OAI21_X1 U4882 ( .B1(n4404), .B2(n4403), .A(n4480), .ZN(n4407) );
  NAND2_X1 U4883 ( .A1(n4766), .A2(EAX_REG_10__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U4884 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4405)
         );
  NAND3_X1 U4885 ( .A1(n4407), .A2(n4406), .A3(n4405), .ZN(n4408) );
  XOR2_X1 U4886 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4424), .Z(n6545) );
  AOI22_X1 U4887 ( .A1(n4766), .A2(EAX_REG_11__SCAN_IN), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4423) );
  AOI22_X1 U4888 ( .A1(n4000), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4889 ( .A1(n4757), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4890 ( .A1(n4569), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4891 ( .A1(n3891), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U4892 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4421)
         );
  AOI22_X1 U4893 ( .A1(n4779), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U4894 ( .A1(n4564), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U4895 ( .A1(n4710), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4896 ( .A1(n3986), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4416) );
  NAND4_X1 U4897 ( .A1(n4419), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n4420)
         );
  OAI21_X1 U4898 ( .B1(n4421), .B2(n4420), .A(n4480), .ZN(n4422) );
  OAI211_X1 U4899 ( .C1(n6545), .C2(n5704), .A(n4423), .B(n4422), .ZN(n5958)
         );
  XNOR2_X1 U4900 ( .A(n4451), .B(n7413), .ZN(n7408) );
  NAND2_X1 U4901 ( .A1(n7408), .A2(n4798), .ZN(n4439) );
  AOI22_X1 U4902 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4000), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4903 ( .A1(n4757), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U4904 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4569), .B1(n4784), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U4905 ( .A1(n4730), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4425) );
  NAND4_X1 U4906 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), .ZN(n4434)
         );
  AOI22_X1 U4907 ( .A1(n4779), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4908 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3891), .B1(n3698), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U4909 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4710), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U4910 ( .A1(n3674), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4429) );
  NAND4_X1 U4911 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), .ZN(n4433)
         );
  OAI21_X1 U4912 ( .B1(n4434), .B2(n4433), .A(n4480), .ZN(n4437) );
  NAND2_X1 U4913 ( .A1(n4766), .A2(EAX_REG_12__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U4914 ( .A1(n6119), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4435)
         );
  AND3_X1 U4915 ( .A1(n4437), .A2(n4436), .A3(n4435), .ZN(n4438) );
  NAND2_X1 U4916 ( .A1(n4439), .A2(n4438), .ZN(n5976) );
  AOI22_X1 U4917 ( .A1(n4779), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4443) );
  AOI22_X1 U4918 ( .A1(n3992), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U4919 ( .A1(n3891), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U4920 ( .A1(n3986), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4440) );
  NAND4_X1 U4921 ( .A1(n4443), .A2(n4442), .A3(n4441), .A4(n4440), .ZN(n4449)
         );
  AOI22_X1 U4922 ( .A1(n4730), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U4923 ( .A1(n4587), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U4924 ( .A1(n4569), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4925 ( .A1(n4752), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4444) );
  NAND4_X1 U4926 ( .A1(n4447), .A2(n4446), .A3(n4445), .A4(n4444), .ZN(n4448)
         );
  OR2_X1 U4927 ( .A1(n4449), .A2(n4448), .ZN(n4450) );
  NAND2_X1 U4928 ( .A1(n4766), .A2(EAX_REG_13__SCAN_IN), .ZN(n4453) );
  XNOR2_X1 U4929 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4465), .ZN(n6532)
         );
  AOI22_X1 U4930 ( .A1(n4798), .A2(n6532), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U4931 ( .A1(n4453), .A2(n4452), .ZN(n6274) );
  AOI22_X1 U4932 ( .A1(n4757), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4933 ( .A1(n4730), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U4934 ( .A1(n3992), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U4935 ( .A1(n3697), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4455) );
  NAND4_X1 U4936 ( .A1(n4458), .A2(n4457), .A3(n4456), .A4(n4455), .ZN(n4464)
         );
  AOI22_X1 U4937 ( .A1(n4779), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U4938 ( .A1(n3891), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U4939 ( .A1(n4569), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U4940 ( .A1(n3705), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4459) );
  NAND4_X1 U4941 ( .A1(n4462), .A2(n4461), .A3(n4460), .A4(n4459), .ZN(n4463)
         );
  NOR2_X1 U4942 ( .A1(n4464), .A2(n4463), .ZN(n4469) );
  INV_X1 U4943 ( .A(n4471), .ZN(n4466) );
  XNOR2_X1 U4944 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4466), .ZN(n6525)
         );
  AOI22_X1 U4945 ( .A1(n4798), .A2(n6525), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U4946 ( .A1(n4766), .A2(EAX_REG_14__SCAN_IN), .ZN(n4467) );
  OAI211_X1 U4947 ( .C1(n4470), .C2(n4469), .A(n4468), .B(n4467), .ZN(n6256)
         );
  INV_X1 U4948 ( .A(n6248), .ZN(n4486) );
  XOR2_X1 U4949 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4487), .Z(n6512) );
  AOI22_X1 U4950 ( .A1(n4766), .A2(EAX_REG_15__SCAN_IN), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U4951 ( .A1(n4000), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4475) );
  AOI22_X1 U4952 ( .A1(n3891), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4752), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U4953 ( .A1(n3705), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U4954 ( .A1(n4784), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4472) );
  NAND4_X1 U4955 ( .A1(n4475), .A2(n4474), .A3(n4473), .A4(n4472), .ZN(n4482)
         );
  AOI22_X1 U4956 ( .A1(n4779), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4479) );
  AOI22_X1 U4957 ( .A1(n4569), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U4958 ( .A1(n4710), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U4959 ( .A1(n4730), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4476) );
  NAND4_X1 U4960 ( .A1(n4479), .A2(n4478), .A3(n4477), .A4(n4476), .ZN(n4481)
         );
  OAI21_X1 U4961 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n4483) );
  OAI211_X1 U4962 ( .C1(n6512), .C2(n5704), .A(n4484), .B(n4483), .ZN(n4485)
         );
  INV_X1 U4963 ( .A(n4485), .ZN(n6249) );
  XNOR2_X1 U4964 ( .A(n4518), .B(n6503), .ZN(n6242) );
  AOI22_X1 U4965 ( .A1(n4779), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U4966 ( .A1(n3992), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U4967 ( .A1(n3891), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U4968 ( .A1(n4569), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4488) );
  NAND4_X1 U4969 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(n4497)
         );
  AOI22_X1 U4970 ( .A1(n4757), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U4971 ( .A1(n4730), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U4972 ( .A1(n4784), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U4973 ( .A1(n4752), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4492) );
  NAND4_X1 U4974 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4496)
         );
  NOR2_X1 U4975 ( .A1(n4497), .A2(n4496), .ZN(n4501) );
  NOR2_X1 U4976 ( .A1(n4498), .A2(n6503), .ZN(n4499) );
  AOI21_X1 U4977 ( .B1(n4766), .B2(EAX_REG_16__SCAN_IN), .A(n4499), .ZN(n4500)
         );
  OAI21_X1 U4978 ( .B1(n4768), .B2(n4501), .A(n4500), .ZN(n4502) );
  AOI21_X1 U4979 ( .B1(n6242), .B2(n4798), .A(n4502), .ZN(n6233) );
  AOI22_X1 U4980 ( .A1(n4000), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U4981 ( .A1(n4569), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U4982 ( .A1(n4564), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U4983 ( .A1(n4784), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4504) );
  NAND4_X1 U4984 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(n4513)
         );
  AOI22_X1 U4985 ( .A1(n4757), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U4986 ( .A1(n3891), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U4987 ( .A1(n4779), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U4988 ( .A1(n3697), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4508) );
  NAND4_X1 U4989 ( .A1(n4511), .A2(n4510), .A3(n4509), .A4(n4508), .ZN(n4512)
         );
  NOR2_X1 U4990 ( .A1(n4513), .A2(n4512), .ZN(n4517) );
  OAI21_X1 U4991 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n7303), .A(n7522), 
        .ZN(n4514) );
  INV_X1 U4992 ( .A(n4514), .ZN(n4515) );
  AOI21_X1 U4993 ( .B1(n4766), .B2(EAX_REG_17__SCAN_IN), .A(n4515), .ZN(n4516)
         );
  OAI21_X1 U4994 ( .B1(n4768), .B2(n4517), .A(n4516), .ZN(n4525) );
  INV_X1 U4995 ( .A(n4556), .ZN(n4523) );
  INV_X1 U4996 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4521) );
  INV_X1 U4997 ( .A(n4519), .ZN(n4520) );
  NAND2_X1 U4998 ( .A1(n4521), .A2(n4520), .ZN(n4522) );
  NAND2_X1 U4999 ( .A1(n4523), .A2(n4522), .ZN(n7421) );
  NAND2_X1 U5000 ( .A1(n4525), .A2(n4524), .ZN(n6348) );
  NAND2_X1 U5001 ( .A1(n4768), .A2(n5704), .ZN(n4619) );
  AOI22_X1 U5002 ( .A1(n4779), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U5003 ( .A1(n4730), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3697), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U5004 ( .A1(n4711), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4527) );
  NAND2_X1 U5005 ( .A1(n4000), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4526)
         );
  AND3_X1 U5006 ( .A1(n4527), .A2(n4526), .A3(n5704), .ZN(n4529) );
  AOI22_X1 U5007 ( .A1(n3992), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4528) );
  NAND4_X1 U5008 ( .A1(n4531), .A2(n4530), .A3(n4529), .A4(n4528), .ZN(n4537)
         );
  AOI22_X1 U5009 ( .A1(n4757), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5010 ( .A1(n4569), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5011 ( .A1(n3925), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4533) );
  AOI22_X1 U5012 ( .A1(n4710), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4532) );
  NAND4_X1 U5013 ( .A1(n4535), .A2(n4534), .A3(n4533), .A4(n4532), .ZN(n4536)
         );
  OR2_X1 U5014 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  NAND2_X1 U5015 ( .A1(n4619), .A2(n4538), .ZN(n4541) );
  AOI22_X1 U5016 ( .A1(n4766), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n7522), .ZN(n4540) );
  INV_X1 U5017 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n7434) );
  XNOR2_X1 U5018 ( .A(n4556), .B(n7434), .ZN(n7440) );
  AND2_X1 U5019 ( .A1(n7440), .A2(n4798), .ZN(n4539) );
  AOI21_X1 U5020 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n6338) );
  AOI22_X1 U5021 ( .A1(n4000), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5022 ( .A1(n3697), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5023 ( .A1(n4779), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5024 ( .A1(n4569), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4542) );
  NAND4_X1 U5025 ( .A1(n4545), .A2(n4544), .A3(n4543), .A4(n4542), .ZN(n4551)
         );
  AOI22_X1 U5026 ( .A1(n3992), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5027 ( .A1(n4710), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5028 ( .A1(n3674), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4547) );
  AOI22_X1 U5029 ( .A1(n4730), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4546) );
  NAND4_X1 U5030 ( .A1(n4549), .A2(n4548), .A3(n4547), .A4(n4546), .ZN(n4550)
         );
  NOR2_X1 U5031 ( .A1(n4551), .A2(n4550), .ZN(n4555) );
  NAND2_X1 U5032 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4552)
         );
  NAND2_X1 U5033 ( .A1(n5704), .A2(n4552), .ZN(n4553) );
  AOI21_X1 U5034 ( .B1(n4766), .B2(EAX_REG_19__SCAN_IN), .A(n4553), .ZN(n4554)
         );
  OAI21_X1 U5035 ( .B1(n4768), .B2(n4555), .A(n4554), .ZN(n4562) );
  INV_X1 U5036 ( .A(n4557), .ZN(n4559) );
  INV_X1 U5037 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U5038 ( .A1(n4559), .A2(n4558), .ZN(n4560) );
  AND2_X1 U5039 ( .A1(n4597), .A2(n4560), .ZN(n7447) );
  NAND2_X1 U5040 ( .A1(n7447), .A2(n4798), .ZN(n4561) );
  NAND2_X1 U5041 ( .A1(n4562), .A2(n4561), .ZN(n6332) );
  AOI22_X1 U5042 ( .A1(n4710), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4752), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5043 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4779), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5044 ( .A1(n3696), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5045 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4564), .B1(n4784), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4565) );
  NAND4_X1 U5046 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(n4577)
         );
  AOI22_X1 U5047 ( .A1(n4757), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5048 ( .A1(n4569), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4571)
         );
  NAND2_X1 U5049 ( .A1(n4001), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4570) );
  AND3_X1 U5050 ( .A1(n4571), .A2(n4570), .A3(n5704), .ZN(n4574) );
  AOI22_X1 U5051 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3674), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5052 ( .A1(n3992), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4572) );
  NAND4_X1 U5053 ( .A1(n4575), .A2(n4574), .A3(n4573), .A4(n4572), .ZN(n4576)
         );
  OAI21_X1 U5054 ( .B1(n4577), .B2(n4576), .A(n4619), .ZN(n4579) );
  AOI22_X1 U5055 ( .A1(n4766), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n7522), .ZN(n4578) );
  NAND2_X1 U5056 ( .A1(n4579), .A2(n4578), .ZN(n4581) );
  XNOR2_X1 U5057 ( .A(n4597), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6485)
         );
  NAND2_X1 U5058 ( .A1(n6485), .A2(n4798), .ZN(n4580) );
  NAND2_X1 U5059 ( .A1(n4581), .A2(n4580), .ZN(n6219) );
  AOI22_X1 U5060 ( .A1(n4757), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5061 ( .A1(n3992), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5062 ( .A1(n4730), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5063 ( .A1(n4751), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4583) );
  NAND4_X1 U5064 ( .A1(n4586), .A2(n4585), .A3(n4584), .A4(n4583), .ZN(n4593)
         );
  AOI22_X1 U5065 ( .A1(n4779), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5066 ( .A1(n4710), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U5067 ( .A1(n4569), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5068 ( .A1(n4752), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4588) );
  NAND4_X1 U5069 ( .A1(n4591), .A2(n4590), .A3(n4589), .A4(n4588), .ZN(n4592)
         );
  NOR2_X1 U5070 ( .A1(n4593), .A2(n4592), .ZN(n4594) );
  OR2_X1 U5071 ( .A1(n4768), .A2(n4594), .ZN(n4603) );
  NAND2_X1 U5072 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4595)
         );
  NAND2_X1 U5073 ( .A1(n5704), .A2(n4595), .ZN(n4596) );
  AOI21_X1 U5074 ( .B1(n4766), .B2(EAX_REG_21__SCAN_IN), .A(n4596), .ZN(n4602)
         );
  INV_X1 U5075 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U5076 ( .A1(n4599), .A2(n6475), .ZN(n4600) );
  NAND2_X1 U5077 ( .A1(n4649), .A2(n4600), .ZN(n6474) );
  NOR2_X1 U5078 ( .A1(n6474), .A2(n5704), .ZN(n4601) );
  AOI21_X1 U5079 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n6320) );
  AOI22_X1 U5080 ( .A1(n4757), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3697), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5081 ( .A1(n4711), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5082 ( .A1(n3696), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4604)
         );
  AND3_X1 U5083 ( .A1(n4605), .A2(n4604), .A3(n5704), .ZN(n4608) );
  AOI22_X1 U5084 ( .A1(n4730), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4784), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5085 ( .A1(n4001), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4606) );
  NAND4_X1 U5086 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4617)
         );
  AOI22_X1 U5087 ( .A1(n4779), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5088 ( .A1(n4569), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5089 ( .A1(n4587), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5090 ( .A1(n3705), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4612) );
  NAND4_X1 U5091 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4616)
         );
  OR2_X1 U5092 ( .A1(n4617), .A2(n4616), .ZN(n4618) );
  NAND2_X1 U5093 ( .A1(n4619), .A2(n4618), .ZN(n4622) );
  AOI22_X1 U5094 ( .A1(n4766), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n7522), .ZN(n4621) );
  XNOR2_X1 U5095 ( .A(n4649), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6469)
         );
  AOI21_X1 U5096 ( .B1(n4622), .B2(n4621), .A(n4620), .ZN(n6209) );
  AOI22_X1 U5097 ( .A1(n4000), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4626) );
  AOI22_X1 U5098 ( .A1(n4569), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5099 ( .A1(n3992), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5100 ( .A1(n4779), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4623) );
  NAND4_X1 U5101 ( .A1(n4626), .A2(n4625), .A3(n4624), .A4(n4623), .ZN(n4632)
         );
  AOI22_X1 U5102 ( .A1(n4730), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5103 ( .A1(n4710), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5104 ( .A1(n4784), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5105 ( .A1(n3698), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4627) );
  NAND4_X1 U5106 ( .A1(n4630), .A2(n4629), .A3(n4628), .A4(n4627), .ZN(n4631)
         );
  OR2_X1 U5107 ( .A1(n4632), .A2(n4631), .ZN(n4644) );
  AOI22_X1 U5108 ( .A1(n4000), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5109 ( .A1(n4569), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5110 ( .A1(n3992), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3986), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5111 ( .A1(n4779), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4633) );
  NAND4_X1 U5112 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4642)
         );
  AOI22_X1 U5113 ( .A1(n4730), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5114 ( .A1(n4710), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5115 ( .A1(n4751), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5116 ( .A1(n3697), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4637) );
  NAND4_X1 U5117 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641)
         );
  OR2_X1 U5118 ( .A1(n4642), .A2(n4641), .ZN(n4643) );
  NAND2_X1 U5119 ( .A1(n4643), .A2(n4644), .ZN(n4680) );
  OAI21_X1 U5120 ( .B1(n4644), .B2(n4643), .A(n4680), .ZN(n4648) );
  NAND2_X1 U5121 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4645)
         );
  NAND2_X1 U5122 ( .A1(n5704), .A2(n4645), .ZN(n4646) );
  AOI21_X1 U5123 ( .B1(n4766), .B2(EAX_REG_23__SCAN_IN), .A(n4646), .ZN(n4647)
         );
  OAI21_X1 U5124 ( .B1(n4768), .B2(n4648), .A(n4647), .ZN(n4654) );
  INV_X1 U5125 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U5126 ( .A1(n4651), .A2(n6460), .ZN(n4652) );
  AND2_X1 U5127 ( .A1(n4685), .A2(n4652), .ZN(n7476) );
  NAND2_X1 U5128 ( .A1(n7476), .A2(n4798), .ZN(n4653) );
  NAND2_X1 U5129 ( .A1(n4654), .A2(n4653), .ZN(n6309) );
  AOI22_X1 U5130 ( .A1(n4779), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5131 ( .A1(n3992), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5132 ( .A1(n4001), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5133 ( .A1(n3698), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4655) );
  NAND4_X1 U5134 ( .A1(n4658), .A2(n4657), .A3(n4656), .A4(n4655), .ZN(n4664)
         );
  AOI22_X1 U5135 ( .A1(n4569), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5136 ( .A1(n4730), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5137 ( .A1(n4000), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5138 ( .A1(n4751), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4659) );
  NAND4_X1 U5139 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4663)
         );
  NOR2_X1 U5140 ( .A1(n4664), .A2(n4663), .ZN(n4681) );
  XNOR2_X1 U5141 ( .A(n4680), .B(n4681), .ZN(n4665) );
  OR2_X1 U5142 ( .A1(n4768), .A2(n4665), .ZN(n4668) );
  AOI22_X1 U5143 ( .A1(n4766), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6119), .ZN(n4667) );
  INV_X1 U5144 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6198) );
  XNOR2_X1 U5145 ( .A(n4685), .B(n6198), .ZN(n6451) );
  NAND2_X1 U5146 ( .A1(n6451), .A2(n4798), .ZN(n4666) );
  AOI22_X1 U5147 ( .A1(n4000), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5148 ( .A1(n4569), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5149 ( .A1(n3992), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3705), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U5150 ( .A1(n4779), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4670) );
  NAND4_X1 U5151 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4679)
         );
  AOI22_X1 U5152 ( .A1(n4730), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5153 ( .A1(n4710), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5154 ( .A1(n4784), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5155 ( .A1(n3698), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4674) );
  NAND4_X1 U5156 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4678)
         );
  OR2_X1 U5157 ( .A1(n4679), .A2(n4678), .ZN(n4701) );
  NOR2_X1 U5158 ( .A1(n4681), .A2(n4680), .ZN(n4702) );
  XNOR2_X1 U5159 ( .A(n4701), .B(n4702), .ZN(n4684) );
  INV_X1 U5160 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6180) );
  AOI21_X1 U5161 ( .B1(n6180), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4682) );
  AOI21_X1 U5162 ( .B1(n4766), .B2(EAX_REG_25__SCAN_IN), .A(n4682), .ZN(n4683)
         );
  OAI21_X1 U5163 ( .B1(n4768), .B2(n4684), .A(n4683), .ZN(n4690) );
  NAND2_X1 U5164 ( .A1(n4687), .A2(n6180), .ZN(n4688) );
  NAND2_X1 U5165 ( .A1(n4724), .A2(n4688), .ZN(n6437) );
  AOI22_X1 U5166 ( .A1(n4569), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5167 ( .A1(n4710), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5168 ( .A1(n3696), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5169 ( .A1(n3986), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4691) );
  NAND4_X1 U5170 ( .A1(n4694), .A2(n4693), .A3(n4692), .A4(n4691), .ZN(n4700)
         );
  AOI22_X1 U5171 ( .A1(n4779), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5172 ( .A1(n4730), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5173 ( .A1(n3992), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5174 ( .A1(n4752), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4695) );
  NAND4_X1 U5175 ( .A1(n4698), .A2(n4697), .A3(n4696), .A4(n4695), .ZN(n4699)
         );
  NOR2_X1 U5176 ( .A1(n4700), .A2(n4699), .ZN(n4709) );
  NAND2_X1 U5177 ( .A1(n4702), .A2(n4701), .ZN(n4708) );
  XOR2_X1 U5178 ( .A(n4709), .B(n4708), .Z(n4703) );
  INV_X1 U5179 ( .A(n4768), .ZN(n4794) );
  NAND2_X1 U5180 ( .A1(n4703), .A2(n4794), .ZN(n4707) );
  INV_X1 U5181 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6425) );
  AOI21_X1 U5182 ( .B1(n6425), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4704) );
  AOI21_X1 U5183 ( .B1(n4766), .B2(EAX_REG_26__SCAN_IN), .A(n4704), .ZN(n4706)
         );
  XNOR2_X1 U5184 ( .A(n4724), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6429)
         );
  AOI21_X1 U5185 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(n6167) );
  OR2_X1 U5186 ( .A1(n4709), .A2(n4708), .ZN(n4743) );
  AOI22_X1 U5187 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4730), .B1(n3891), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5188 ( .A1(n4779), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4710), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5189 ( .A1(n4569), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5190 ( .A1(n3925), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4712) );
  NAND4_X1 U5191 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4721)
         );
  AOI22_X1 U5192 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3992), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5193 ( .A1(n4757), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4718) );
  AOI22_X1 U5194 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3696), .B1(n4751), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5195 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3698), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4716) );
  NAND4_X1 U5196 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4720)
         );
  OR2_X1 U5197 ( .A1(n4721), .A2(n4720), .ZN(n4741) );
  XNOR2_X1 U5198 ( .A(n4743), .B(n4741), .ZN(n4722) );
  NAND2_X1 U5199 ( .A1(n4722), .A2(n4794), .ZN(n4729) );
  INV_X1 U5200 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6418) );
  AOI21_X1 U5201 ( .B1(n6418), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4723) );
  AOI21_X1 U5202 ( .B1(n4766), .B2(EAX_REG_27__SCAN_IN), .A(n4723), .ZN(n4728)
         );
  INV_X1 U5203 ( .A(n4725), .ZN(n4726) );
  NAND2_X1 U5204 ( .A1(n4726), .A2(n6418), .ZN(n4727) );
  AOI22_X1 U5205 ( .A1(n4729), .A2(n4728), .B1(n4798), .B2(n6422), .ZN(n6155)
         );
  AOI22_X1 U5206 ( .A1(n3696), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5207 ( .A1(n4757), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5208 ( .A1(n4710), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5209 ( .A1(n4730), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4731) );
  NAND4_X1 U5210 ( .A1(n4734), .A2(n4733), .A3(n4732), .A4(n4731), .ZN(n4740)
         );
  AOI22_X1 U5211 ( .A1(n4569), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5212 ( .A1(n4779), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U5213 ( .A1(n3697), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5214 ( .A1(n4001), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4735) );
  NAND4_X1 U5215 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4739)
         );
  OR2_X1 U5216 ( .A1(n4740), .A2(n4739), .ZN(n4750) );
  INV_X1 U5217 ( .A(n4741), .ZN(n4742) );
  NOR2_X1 U5218 ( .A1(n4743), .A2(n4742), .ZN(n4749) );
  XOR2_X1 U5219 ( .A(n4750), .B(n4749), .Z(n4744) );
  NAND2_X1 U5220 ( .A1(n4744), .A2(n4794), .ZN(n4748) );
  INV_X1 U5221 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4770) );
  AOI21_X1 U5222 ( .B1(n4770), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4745) );
  AOI21_X1 U5223 ( .B1(n4766), .B2(EAX_REG_28__SCAN_IN), .A(n4745), .ZN(n4747)
         );
  XNOR2_X1 U5224 ( .A(n4771), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6408)
         );
  AOI21_X1 U5225 ( .B1(n4748), .B2(n4747), .A(n4746), .ZN(n6143) );
  NAND2_X1 U5226 ( .A1(n4750), .A2(n4749), .ZN(n4777) );
  AOI22_X1 U5227 ( .A1(n4730), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5228 ( .A1(n4779), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4755) );
  AOI22_X1 U5229 ( .A1(n3986), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4751), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4754) );
  AOI22_X1 U5230 ( .A1(n4752), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4753) );
  NAND4_X1 U5231 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4763)
         );
  AOI22_X1 U5232 ( .A1(n3696), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5233 ( .A1(n4569), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5234 ( .A1(n4710), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3891), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5235 ( .A1(n3992), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4758) );
  NAND4_X1 U5236 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), .ZN(n4762)
         );
  NOR2_X1 U5237 ( .A1(n4763), .A2(n4762), .ZN(n4776) );
  XNOR2_X1 U5238 ( .A(n4777), .B(n4776), .ZN(n4769) );
  NAND2_X1 U5239 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4764)
         );
  NAND2_X1 U5240 ( .A1(n5704), .A2(n4764), .ZN(n4765) );
  AOI21_X1 U5241 ( .B1(n4766), .B2(EAX_REG_29__SCAN_IN), .A(n4765), .ZN(n4767)
         );
  OAI21_X1 U5242 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(n4775) );
  INV_X1 U5243 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U5244 ( .A1(n4772), .A2(n6134), .ZN(n4773) );
  NAND2_X1 U5245 ( .A1(n6132), .A2(n4798), .ZN(n4774) );
  NAND2_X1 U5246 ( .A1(n4775), .A2(n4774), .ZN(n4818) );
  NOR2_X1 U5247 ( .A1(n4777), .A2(n4776), .ZN(n4793) );
  AOI22_X1 U5248 ( .A1(n3696), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4587), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5249 ( .A1(n4569), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4757), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5250 ( .A1(n3992), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5251 ( .A1(n4779), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4778), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4780) );
  NAND4_X1 U5252 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4791)
         );
  AOI22_X1 U5253 ( .A1(n4730), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4001), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5254 ( .A1(n4710), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4711), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5255 ( .A1(n4784), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5256 ( .A1(n3697), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4785), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4786) );
  NAND4_X1 U5257 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4790)
         );
  NOR2_X1 U5258 ( .A1(n4791), .A2(n4790), .ZN(n4792) );
  XNOR2_X1 U5259 ( .A(n4793), .B(n4792), .ZN(n4795) );
  NAND2_X1 U5260 ( .A1(n4795), .A2(n4794), .ZN(n4801) );
  NAND2_X1 U5261 ( .A1(n7522), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4796)
         );
  NAND2_X1 U5262 ( .A1(n5704), .A2(n4796), .ZN(n4797) );
  AOI21_X1 U5263 ( .B1(n4766), .B2(EAX_REG_30__SCAN_IN), .A(n4797), .ZN(n4800)
         );
  XNOR2_X1 U5264 ( .A(n5709), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6074)
         );
  AOI21_X1 U5265 ( .B1(n4801), .B2(n4800), .A(n4799), .ZN(n6117) );
  NAND2_X1 U5266 ( .A1(n3966), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5703) );
  NOR2_X1 U5267 ( .A1(n5703), .A2(n7303), .ZN(n4832) );
  NOR2_X1 U5268 ( .A1(n6005), .A2(n6509), .ZN(n4810) );
  AND2_X1 U5269 ( .A1(n4802), .A2(n5456), .ZN(n7307) );
  OR2_X1 U5270 ( .A1(n7307), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U5271 ( .A1(n3966), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U5272 ( .A1(n7303), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4804) );
  AND2_X1 U5273 ( .A1(n4805), .A2(n4804), .ZN(n4947) );
  NAND2_X1 U5274 ( .A1(n6074), .A2(n6513), .ZN(n4808) );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5276 ( .A1(n6546), .A2(REIP_REG_30__SCAN_IN), .ZN(n6587) );
  OAI21_X1 U5277 ( .B1(n6516), .B2(n5708), .A(n6587), .ZN(n4806) );
  INV_X1 U5278 ( .A(n4806), .ZN(n4807) );
  NAND2_X1 U5279 ( .A1(n4812), .A2(n4811), .ZN(U2956) );
  NAND2_X1 U5280 ( .A1(n6399), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4814) );
  NOR2_X1 U5281 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4813) );
  INV_X1 U5282 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6584) );
  OAI21_X1 U5283 ( .B1(n3783), .B2(n6584), .A(n6395), .ZN(n4816) );
  AOI21_X1 U5284 ( .B1(n4818), .B2(n4817), .A(n6118), .ZN(n6131) );
  NAND2_X1 U5285 ( .A1(n6513), .A2(n6132), .ZN(n4819) );
  NAND2_X1 U5286 ( .A1(n7330), .A2(REIP_REG_29__SCAN_IN), .ZN(n6594) );
  OAI211_X1 U5287 ( .C1(n6134), .C2(n6516), .A(n4819), .B(n6594), .ZN(n4820)
         );
  AOI21_X1 U5288 ( .B1(n6131), .B2(n6534), .A(n4820), .ZN(n4821) );
  OAI21_X1 U5289 ( .B1(n6600), .B2(n7482), .A(n4821), .ZN(U2957) );
  AND2_X1 U5290 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7558) );
  INV_X1 U5291 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7559) );
  INV_X1 U5292 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7298) );
  NOR2_X1 U5293 ( .A1(n7559), .A2(n7298), .ZN(n4828) );
  AOI21_X1 U5294 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n4828), .ZN(n4823)
         );
  NAND2_X1 U5295 ( .A1(n4822), .A2(n7298), .ZN(n6105) );
  NAND2_X1 U5296 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n7560) );
  OAI211_X1 U5297 ( .C1(n7558), .C2(n4823), .A(n6105), .B(n7560), .ZN(U3182)
         );
  INV_X1 U5298 ( .A(HOLD), .ZN(n4824) );
  NOR2_X1 U5299 ( .A1(n4824), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n4826) );
  INV_X1 U5300 ( .A(READY_N), .ZN(n7516) );
  OAI21_X1 U5301 ( .B1(n7516), .B2(NA_N), .A(STATE_REG_1__SCAN_IN), .ZN(n4825)
         );
  AOI211_X1 U5302 ( .C1(n4826), .C2(n4825), .A(n7298), .B(n7558), .ZN(n4831)
         );
  INV_X1 U5303 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7562) );
  AOI21_X1 U5304 ( .B1(NA_N), .B2(n7098), .A(n7562), .ZN(n4827) );
  NOR2_X1 U5305 ( .A1(n4827), .A2(STATE_REG_0__SCAN_IN), .ZN(n7561) );
  INV_X1 U5306 ( .A(NA_N), .ZN(n4829) );
  AOI21_X1 U5307 ( .B1(n4829), .B2(n4828), .A(STATE_REG_2__SCAN_IN), .ZN(n4830) );
  OAI22_X1 U5308 ( .A1(n4831), .A2(n7561), .B1(n4830), .B2(n7560), .ZN(U3183)
         );
  NAND2_X1 U5309 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n7536) );
  NOR2_X1 U5310 ( .A1(n3966), .A2(n7536), .ZN(n7531) );
  NOR2_X1 U5311 ( .A1(n3966), .A2(n5711), .ZN(n7525) );
  AOI21_X1 U5312 ( .B1(n7516), .B2(n7525), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4834) );
  INV_X1 U5313 ( .A(n4832), .ZN(n4833) );
  OAI21_X1 U5314 ( .B1(n7531), .B2(n4834), .A(n4833), .ZN(U3150) );
  INV_X1 U5315 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4835) );
  AOI21_X1 U5316 ( .B1(n7562), .B2(STATE_REG_1__SCAN_IN), .A(n7298), .ZN(n4837) );
  OR2_X1 U5317 ( .A1(n7098), .A2(STATE_REG_0__SCAN_IN), .ZN(n7566) );
  INV_X2 U5318 ( .A(n7566), .ZN(n7569) );
  AOI21_X1 U5319 ( .B1(n4835), .B2(n4837), .A(n7569), .ZN(U2789) );
  INV_X1 U5320 ( .A(W_R_N_REG_SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5321 ( .A1(n4836), .A2(n7566), .B1(READREQUEST_REG_SCAN_IN), .B2(
        n7569), .ZN(U3470) );
  NOR2_X2 U5322 ( .A1(n7569), .A2(n4837), .ZN(n7170) );
  INV_X1 U5323 ( .A(n7170), .ZN(n7171) );
  INV_X1 U5324 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7103) );
  INV_X1 U5325 ( .A(BS16_N), .ZN(n4839) );
  NAND2_X1 U5326 ( .A1(n7562), .A2(n7298), .ZN(n4838) );
  AOI21_X1 U5327 ( .B1(n4839), .B2(n4838), .A(n7171), .ZN(n4840) );
  AOI21_X1 U5328 ( .B1(n7171), .B2(n7103), .A(n4840), .ZN(U3451) );
  INV_X1 U5329 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n4841) );
  INV_X1 U5330 ( .A(n4840), .ZN(n4842) );
  OAI21_X1 U5331 ( .B1(n7170), .B2(n4841), .A(n4842), .ZN(U3452) );
  OAI21_X1 U5332 ( .B1(n7170), .B2(n7303), .A(n4842), .ZN(U2792) );
  NOR3_X1 U5333 ( .A1(n4846), .A2(n4845), .A3(n4844), .ZN(n4847) );
  OR2_X1 U5334 ( .A1(n4848), .A2(n4847), .ZN(n4851) );
  INV_X1 U5335 ( .A(n4849), .ZN(n4850) );
  NAND2_X1 U5336 ( .A1(n4851), .A2(n4850), .ZN(n6096) );
  AND2_X1 U5337 ( .A1(n6096), .A2(n5175), .ZN(n4852) );
  NAND2_X1 U5338 ( .A1(n4843), .A2(n4852), .ZN(n4855) );
  INV_X1 U5339 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5340 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7568) );
  OAI211_X1 U5341 ( .C1(n4854), .C2(n7568), .A(n4861), .B(n5718), .ZN(U2788)
         );
  NAND2_X1 U5342 ( .A1(n4065), .A2(n5752), .ZN(n6106) );
  INV_X1 U5343 ( .A(n5718), .ZN(n4856) );
  OAI21_X1 U5344 ( .B1(n4856), .B2(READREQUEST_REG_SCAN_IN), .A(n7306), .ZN(
        n4857) );
  OAI21_X1 U5345 ( .B1(n7306), .B2(n6106), .A(n4857), .ZN(U3474) );
  INV_X1 U5346 ( .A(n4920), .ZN(n4860) );
  NAND2_X1 U5347 ( .A1(n3675), .A2(n7304), .ZN(n7519) );
  INV_X1 U5348 ( .A(n7519), .ZN(n4859) );
  INV_X1 U5349 ( .A(n4861), .ZN(n4862) );
  NAND2_X1 U5350 ( .A1(n5042), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5351 ( .A1(n3675), .A2(n6018), .ZN(n4967) );
  NOR2_X2 U5352 ( .A1(n4920), .A2(n4881), .ZN(n5062) );
  NAND2_X1 U5353 ( .A1(n5062), .A2(DATAI_6_), .ZN(n5007) );
  OAI211_X1 U5354 ( .C1(n5014), .C2(n4864), .A(n4863), .B(n5007), .ZN(U2945)
         );
  MUX2_X1 U5355 ( .A(n5206), .B(n4866), .S(n4865), .Z(n4867) );
  OR2_X1 U5356 ( .A1(n4867), .A2(n3971), .ZN(n4878) );
  NAND2_X2 U5357 ( .A1(n4868), .A2(n5721), .ZN(n6054) );
  INV_X1 U5358 ( .A(n5093), .ZN(n6049) );
  NOR2_X1 U5359 ( .A1(n4039), .A2(n5721), .ZN(n4869) );
  MUX2_X1 U5360 ( .A(n4869), .B(n5752), .S(n4957), .Z(n4870) );
  INV_X1 U5361 ( .A(n4870), .ZN(n4871) );
  AOI21_X1 U5362 ( .B1(n4294), .B2(n6114), .A(n4871), .ZN(n4872) );
  AND2_X1 U5363 ( .A1(n4878), .A2(n4872), .ZN(n4873) );
  NAND2_X1 U5364 ( .A1(n4874), .A2(n4873), .ZN(n4981) );
  INV_X1 U5365 ( .A(n4981), .ZN(n4877) );
  NAND2_X1 U5366 ( .A1(n3969), .A2(n5052), .ZN(n4875) );
  NOR2_X1 U5367 ( .A1(n3675), .A2(n4875), .ZN(n4876) );
  NAND2_X1 U5368 ( .A1(n4877), .A2(n4876), .ZN(n4896) );
  NAND2_X1 U5369 ( .A1(n3672), .A2(n5721), .ZN(n4956) );
  INV_X1 U5370 ( .A(n6099), .ZN(n6104) );
  NAND2_X1 U5371 ( .A1(n4879), .A2(n4878), .ZN(n4888) );
  INV_X1 U5372 ( .A(n4888), .ZN(n4880) );
  NAND2_X1 U5373 ( .A1(n4880), .A2(n6103), .ZN(n6095) );
  AND2_X1 U5374 ( .A1(n6095), .A2(n4881), .ZN(n4884) );
  NAND2_X1 U5375 ( .A1(n6096), .A2(n7516), .ZN(n4883) );
  OAI22_X1 U5376 ( .A1(n6099), .A2(n4884), .B1(n3692), .B2(n4883), .ZN(n5048)
         );
  INV_X1 U5377 ( .A(n5048), .ZN(n4892) );
  NAND2_X1 U5378 ( .A1(n4843), .A2(n5206), .ZN(n5134) );
  INV_X1 U5379 ( .A(n3675), .ZN(n4886) );
  OR2_X1 U5380 ( .A1(n6105), .A2(READY_N), .ZN(n4885) );
  AOI21_X1 U5381 ( .B1(n5134), .B2(n4886), .A(n4885), .ZN(n4890) );
  NAND2_X1 U5382 ( .A1(n4887), .A2(n4888), .ZN(n4963) );
  OAI21_X1 U5383 ( .B1(n5752), .B2(n5214), .A(n4963), .ZN(n4889) );
  AOI21_X1 U5384 ( .B1(n6104), .B2(n4890), .A(n4889), .ZN(n4891) );
  OAI211_X1 U5385 ( .C1(n6100), .C2(n6104), .A(n4892), .B(n4891), .ZN(n7495)
         );
  NAND2_X1 U5386 ( .A1(n7495), .A2(n5175), .ZN(n7485) );
  NAND2_X1 U5387 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7531), .ZN(n4893) );
  NAND2_X1 U5388 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n3966), .ZN(n7533) );
  AND2_X1 U5389 ( .A1(n4893), .A2(n7533), .ZN(n4894) );
  NAND2_X1 U5390 ( .A1(n7485), .A2(n4894), .ZN(n7491) );
  INV_X1 U5391 ( .A(n4882), .ZN(n4895) );
  OR2_X1 U5392 ( .A1(n4896), .A2(n4895), .ZN(n5130) );
  NAND2_X1 U5393 ( .A1(n4310), .A2(n5130), .ZN(n4898) );
  NAND2_X1 U5394 ( .A1(n4960), .A2(n3669), .ZN(n4897) );
  NAND2_X1 U5395 ( .A1(n4898), .A2(n4897), .ZN(n7494) );
  NOR2_X1 U5396 ( .A1(n5134), .A2(n3669), .ZN(n7493) );
  AOI21_X1 U5397 ( .B1(n7491), .B2(n7494), .A(n7493), .ZN(n4902) );
  INV_X1 U5398 ( .A(n6081), .ZN(n7486) );
  OAI22_X1 U5399 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7543), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5711), .ZN(n4900) );
  NOR2_X1 U5400 ( .A1(n7491), .A2(n3669), .ZN(n4899) );
  AOI21_X1 U5401 ( .B1(n4900), .B2(n7491), .A(n4899), .ZN(n4901) );
  OAI21_X1 U5402 ( .B1(n4902), .B2(n7486), .A(n4901), .ZN(U3461) );
  INV_X1 U5403 ( .A(n4905), .ZN(n5145) );
  INV_X1 U5404 ( .A(n4906), .ZN(n6086) );
  NAND3_X1 U5405 ( .A1(n4960), .A2(n5145), .A3(n6086), .ZN(n4907) );
  OAI21_X1 U5406 ( .B1(n5134), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4907), 
        .ZN(n4908) );
  AOI21_X1 U5407 ( .B1(n4054), .B2(n5130), .A(n4908), .ZN(n7496) );
  INV_X1 U5408 ( .A(n7496), .ZN(n4911) );
  AND2_X1 U5409 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6085) );
  INV_X1 U5410 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4909) );
  INV_X1 U5411 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5936) );
  AOI22_X1 U5412 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4909), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5936), .ZN(n6080) );
  AOI222_X1 U5413 ( .A1(n4911), .A2(n6081), .B1(n6085), .B2(n6080), .C1(n3670), 
        .C2(n6087), .ZN(n4917) );
  INV_X1 U5414 ( .A(n7491), .ZN(n6089) );
  INV_X1 U5415 ( .A(n4912), .ZN(n4913) );
  OAI22_X1 U5416 ( .A1(n7491), .A2(n4914), .B1(n4913), .B2(n7543), .ZN(n4915)
         );
  INV_X1 U5417 ( .A(n4915), .ZN(n4916) );
  OAI21_X1 U5418 ( .B1(n4917), .B2(n6089), .A(n4916), .ZN(U3460) );
  INV_X1 U5419 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5420 ( .A1(n5134), .A2(n7519), .ZN(n4918) );
  INV_X1 U5421 ( .A(n6105), .ZN(n5720) );
  NAND2_X1 U5422 ( .A1(n4918), .A2(n5720), .ZN(n4919) );
  NAND2_X1 U5423 ( .A1(n4921), .A2(n5721), .ZN(n5110) );
  OR2_X1 U5424 ( .A1(n7536), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7517) );
  AOI22_X1 U5427 ( .A1(n7182), .A2(UWORD_REG_8__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4922) );
  OAI21_X1 U5428 ( .B1(n4923), .B2(n5110), .A(n4922), .ZN(U2899) );
  INV_X1 U5429 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4925) );
  AOI22_X1 U5430 ( .A1(n7182), .A2(UWORD_REG_13__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4924) );
  OAI21_X1 U5431 ( .B1(n4925), .B2(n5110), .A(n4924), .ZN(U2894) );
  INV_X1 U5432 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U5433 ( .A1(n7182), .A2(UWORD_REG_12__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4926) );
  OAI21_X1 U5434 ( .B1(n4927), .B2(n5110), .A(n4926), .ZN(U2895) );
  INV_X1 U5435 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U5436 ( .A1(n7182), .A2(UWORD_REG_7__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4928) );
  OAI21_X1 U5437 ( .B1(n4929), .B2(n5110), .A(n4928), .ZN(U2900) );
  INV_X1 U5438 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4931) );
  AOI22_X1 U5439 ( .A1(n7182), .A2(UWORD_REG_10__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4930) );
  OAI21_X1 U5440 ( .B1(n4931), .B2(n5110), .A(n4930), .ZN(U2897) );
  INV_X1 U5441 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U5442 ( .A1(n7182), .A2(UWORD_REG_9__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4932) );
  OAI21_X1 U5443 ( .B1(n4996), .B2(n5110), .A(n4932), .ZN(U2898) );
  INV_X1 U5444 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U5445 ( .A1(n7182), .A2(UWORD_REG_5__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4933) );
  OAI21_X1 U5446 ( .B1(n4934), .B2(n5110), .A(n4933), .ZN(U2902) );
  INV_X1 U5447 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U5448 ( .A1(n7182), .A2(UWORD_REG_11__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4935) );
  OAI21_X1 U5449 ( .B1(n5010), .B2(n5110), .A(n4935), .ZN(U2896) );
  INV_X1 U5450 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U5451 ( .A1(n7182), .A2(UWORD_REG_6__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U5452 ( .B1(n4937), .B2(n5110), .A(n4936), .ZN(U2901) );
  INV_X1 U5453 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4939) );
  AOI22_X1 U5454 ( .A1(n7182), .A2(UWORD_REG_4__SCAN_IN), .B1(n7172), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U5455 ( .B1(n4939), .B2(n5110), .A(n4938), .ZN(U2903) );
  NOR2_X1 U5456 ( .A1(n4940), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4941)
         );
  NOR2_X1 U5457 ( .A1(n4954), .A2(n4941), .ZN(n7345) );
  INV_X1 U5458 ( .A(n7345), .ZN(n4951) );
  INV_X1 U5459 ( .A(n4942), .ZN(n4946) );
  AOI21_X1 U5460 ( .B1(n4944), .B2(STATE2_REG_2__SCAN_IN), .A(n4943), .ZN(
        n4945) );
  NOR2_X1 U5461 ( .A1(n4946), .A2(n4945), .ZN(n5058) );
  INV_X2 U5462 ( .A(n6509), .ZN(n6534) );
  NAND2_X1 U5463 ( .A1(n6546), .A2(REIP_REG_0__SCAN_IN), .ZN(n7339) );
  INV_X1 U5464 ( .A(n7339), .ZN(n4949) );
  INV_X1 U5465 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5858) );
  AOI21_X1 U5466 ( .B1(n6516), .B2(n4947), .A(n5858), .ZN(n4948) );
  AOI211_X1 U5467 ( .C1(n5058), .C2(n6534), .A(n4949), .B(n4948), .ZN(n4950)
         );
  OAI21_X1 U5468 ( .B1(n4951), .B2(n7482), .A(n4950), .ZN(U2986) );
  AOI222_X1 U5469 ( .A1(n5065), .A2(LWORD_REG_15__SCAN_IN), .B1(DATAI_15_), 
        .B2(n5062), .C1(EAX_REG_15__SCAN_IN), .C2(n5015), .ZN(n4952) );
  INV_X1 U5470 ( .A(n4952), .ZN(U2954) );
  XNOR2_X1 U5471 ( .A(n4953), .B(n4954), .ZN(n5074) );
  AOI21_X1 U5472 ( .B1(n4955), .B2(n6105), .A(READY_N), .ZN(n4958) );
  AOI22_X1 U5473 ( .A1(n3675), .A2(n4958), .B1(n4957), .B2(n4956), .ZN(n4959)
         );
  OR2_X1 U5474 ( .A1(n6099), .A2(n4959), .ZN(n4965) );
  NAND3_X1 U5475 ( .A1(n6099), .A2(n4960), .A3(n5206), .ZN(n4964) );
  NAND2_X1 U5476 ( .A1(n5206), .A2(n6105), .ZN(n4961) );
  NAND4_X1 U5477 ( .A1(n6096), .A2(n5214), .A3(n7516), .A4(n4961), .ZN(n4962)
         );
  NAND4_X1 U5478 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n4966)
         );
  OAI211_X1 U5479 ( .C1(n5050), .C2(n4971), .A(n7509), .B(n4967), .ZN(n4968)
         );
  INV_X1 U5480 ( .A(n4968), .ZN(n4969) );
  AND3_X1 U5481 ( .A1(n3692), .A2(n4969), .A3(n6095), .ZN(n4970) );
  OR2_X2 U5482 ( .A1(n4986), .A2(n4970), .ZN(n6765) );
  OR2_X1 U5483 ( .A1(n4971), .A2(n3899), .ZN(n4972) );
  AND2_X1 U5484 ( .A1(n7519), .A2(n4972), .ZN(n4973) );
  INV_X1 U5485 ( .A(n5093), .ZN(n5523) );
  INV_X1 U5486 ( .A(EBX_REG_1__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U5487 ( .A1(n6029), .A2(n7361), .ZN(n4976) );
  NAND2_X1 U5489 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4974)
         );
  OAI211_X1 U5490 ( .C1(n6113), .C2(EBX_REG_1__SCAN_IN), .A(n6054), .B(n4974), 
        .ZN(n4975) );
  NAND2_X1 U5491 ( .A1(n4976), .A2(n4975), .ZN(n5090) );
  INV_X1 U5492 ( .A(n6054), .ZN(n4977) );
  NAND2_X1 U5493 ( .A1(n4977), .A2(EBX_REG_0__SCAN_IN), .ZN(n4979) );
  INV_X1 U5494 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U5495 ( .A1(n5093), .A2(n5857), .ZN(n4978) );
  NAND2_X1 U5496 ( .A1(n4979), .A2(n4978), .ZN(n5483) );
  XNOR2_X1 U5497 ( .A(n5090), .B(n5483), .ZN(n7351) );
  XNOR2_X1 U5498 ( .A(n7351), .B(n6018), .ZN(n7278) );
  NAND2_X1 U5499 ( .A1(n6759), .A2(n4986), .ZN(n7347) );
  INV_X1 U5500 ( .A(n6683), .ZN(n6731) );
  NOR2_X1 U5501 ( .A1(n4981), .A2(n4980), .ZN(n4982) );
  INV_X1 U5502 ( .A(n6732), .ZN(n4983) );
  INV_X1 U5503 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7349) );
  OAI21_X1 U5504 ( .B1(n6731), .B2(n4983), .A(n7349), .ZN(n7340) );
  AOI21_X1 U5505 ( .B1(n7347), .B2(n7340), .A(n5936), .ZN(n4985) );
  INV_X1 U5506 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7350) );
  NOR2_X1 U5507 ( .A1(n6759), .A2(n7350), .ZN(n4984) );
  AOI211_X1 U5508 ( .C1(n7332), .C2(n7278), .A(n4985), .B(n4984), .ZN(n4988)
         );
  NAND2_X1 U5509 ( .A1(n6727), .A2(n6683), .ZN(n6687) );
  INV_X1 U5510 ( .A(n6687), .ZN(n6710) );
  OR3_X1 U5511 ( .A1(n6710), .A2(n5087), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4987) );
  OAI211_X1 U5512 ( .C1(n5074), .C2(n6765), .A(n4988), .B(n4987), .ZN(U3017)
         );
  NAND2_X1 U5513 ( .A1(n5065), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U5514 ( .A1(n5062), .A2(DATAI_7_), .ZN(n5026) );
  OAI211_X1 U5515 ( .C1(n5014), .C2(n4929), .A(n4989), .B(n5026), .ZN(U2931)
         );
  INV_X1 U5516 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5517 ( .A1(n5065), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U5518 ( .A1(n5062), .A2(DATAI_1_), .ZN(n5046) );
  OAI211_X1 U5519 ( .C1(n5014), .C2(n4991), .A(n4990), .B(n5046), .ZN(U2940)
         );
  INV_X1 U5520 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U5521 ( .A1(n5065), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U5522 ( .A1(n5062), .A2(DATAI_14_), .ZN(n4997) );
  OAI211_X1 U5523 ( .C1(n5014), .C2(n4993), .A(n4992), .B(n4997), .ZN(U2953)
         );
  NAND2_X1 U5524 ( .A1(n5065), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U5525 ( .A1(n5062), .A2(DATAI_8_), .ZN(n5043) );
  OAI211_X1 U5526 ( .C1(n5014), .C2(n4923), .A(n4994), .B(n5043), .ZN(U2932)
         );
  NAND2_X1 U5527 ( .A1(n5065), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U5528 ( .A1(n5062), .A2(DATAI_9_), .ZN(n5016) );
  OAI211_X1 U5529 ( .C1(n5014), .C2(n4996), .A(n4995), .B(n5016), .ZN(U2933)
         );
  INV_X1 U5530 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U5531 ( .A1(n5065), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4998) );
  OAI211_X1 U5532 ( .C1(n5014), .C2(n4999), .A(n4998), .B(n4997), .ZN(U2938)
         );
  INV_X1 U5533 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5534 ( .A1(n5065), .A2(UWORD_REG_3__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5535 ( .A1(n5062), .A2(DATAI_3_), .ZN(n5031) );
  OAI211_X1 U5536 ( .C1(n5014), .C2(n5001), .A(n5000), .B(n5031), .ZN(U2927)
         );
  INV_X1 U5537 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5538 ( .A1(n5065), .A2(LWORD_REG_2__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U5539 ( .A1(n5062), .A2(DATAI_2_), .ZN(n5004) );
  OAI211_X1 U5540 ( .C1(n5014), .C2(n5003), .A(n5002), .B(n5004), .ZN(U2941)
         );
  INV_X1 U5541 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U5542 ( .A1(n5065), .A2(UWORD_REG_2__SCAN_IN), .ZN(n5005) );
  OAI211_X1 U5543 ( .C1(n5014), .C2(n5006), .A(n5005), .B(n5004), .ZN(U2926)
         );
  NAND2_X1 U5544 ( .A1(n5065), .A2(UWORD_REG_6__SCAN_IN), .ZN(n5008) );
  OAI211_X1 U5545 ( .C1(n5014), .C2(n4937), .A(n5008), .B(n5007), .ZN(U2930)
         );
  NAND2_X1 U5546 ( .A1(n5065), .A2(UWORD_REG_11__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U5547 ( .A1(n5062), .A2(DATAI_11_), .ZN(n5020) );
  OAI211_X1 U5548 ( .C1(n5014), .C2(n5010), .A(n5009), .B(n5020), .ZN(U2935)
         );
  NAND2_X1 U5549 ( .A1(n5065), .A2(UWORD_REG_12__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U5550 ( .A1(n5062), .A2(DATAI_12_), .ZN(n5037) );
  OAI211_X1 U5551 ( .C1(n5014), .C2(n4927), .A(n5011), .B(n5037), .ZN(U2936)
         );
  NAND2_X1 U5552 ( .A1(n5065), .A2(UWORD_REG_13__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U5553 ( .A1(n5062), .A2(DATAI_13_), .ZN(n5040) );
  OAI211_X1 U5554 ( .C1(n5014), .C2(n4925), .A(n5012), .B(n5040), .ZN(U2937)
         );
  NAND2_X1 U5555 ( .A1(n5065), .A2(UWORD_REG_10__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U5556 ( .A1(n5062), .A2(DATAI_10_), .ZN(n5023) );
  OAI211_X1 U5557 ( .C1(n5014), .C2(n4931), .A(n5013), .B(n5023), .ZN(U2934)
         );
  INV_X1 U5558 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U5559 ( .A1(n5042), .A2(LWORD_REG_9__SCAN_IN), .ZN(n5017) );
  OAI211_X1 U5560 ( .C1(n5068), .C2(n5018), .A(n5017), .B(n5016), .ZN(U2948)
         );
  NAND2_X1 U5561 ( .A1(n5065), .A2(UWORD_REG_5__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U5562 ( .A1(n5062), .A2(DATAI_5_), .ZN(n5029) );
  OAI211_X1 U5563 ( .C1(n5068), .C2(n4934), .A(n5019), .B(n5029), .ZN(U2929)
         );
  INV_X1 U5564 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U5565 ( .A1(n5065), .A2(LWORD_REG_11__SCAN_IN), .ZN(n5021) );
  OAI211_X1 U5566 ( .C1(n5068), .C2(n5022), .A(n5021), .B(n5020), .ZN(U2950)
         );
  INV_X1 U5567 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U5568 ( .A1(n5065), .A2(LWORD_REG_10__SCAN_IN), .ZN(n5024) );
  OAI211_X1 U5569 ( .C1(n5068), .C2(n5025), .A(n5024), .B(n5023), .ZN(U2949)
         );
  INV_X1 U5570 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U5571 ( .A1(n5042), .A2(LWORD_REG_7__SCAN_IN), .ZN(n5027) );
  OAI211_X1 U5572 ( .C1(n5068), .C2(n5028), .A(n5027), .B(n5026), .ZN(U2946)
         );
  NAND2_X1 U5573 ( .A1(n5042), .A2(LWORD_REG_5__SCAN_IN), .ZN(n5030) );
  OAI211_X1 U5574 ( .C1(n5068), .C2(n7181), .A(n5030), .B(n5029), .ZN(U2944)
         );
  INV_X1 U5575 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U5576 ( .A1(n5065), .A2(LWORD_REG_3__SCAN_IN), .ZN(n5032) );
  OAI211_X1 U5577 ( .C1(n5068), .C2(n5033), .A(n5032), .B(n5031), .ZN(U2942)
         );
  INV_X1 U5578 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U5579 ( .A1(n5042), .A2(LWORD_REG_4__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U5580 ( .A1(n5062), .A2(DATAI_4_), .ZN(n5035) );
  OAI211_X1 U5581 ( .C1(n5068), .C2(n7179), .A(n5034), .B(n5035), .ZN(U2943)
         );
  NAND2_X1 U5582 ( .A1(n5065), .A2(UWORD_REG_4__SCAN_IN), .ZN(n5036) );
  OAI211_X1 U5583 ( .C1(n5068), .C2(n4939), .A(n5036), .B(n5035), .ZN(U2928)
         );
  INV_X1 U5584 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U5585 ( .A1(n5065), .A2(LWORD_REG_12__SCAN_IN), .ZN(n5038) );
  OAI211_X1 U5586 ( .C1(n5068), .C2(n5039), .A(n5038), .B(n5037), .ZN(U2951)
         );
  INV_X1 U5587 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U5588 ( .A1(n5065), .A2(LWORD_REG_13__SCAN_IN), .ZN(n5041) );
  OAI211_X1 U5589 ( .C1(n5068), .C2(n7191), .A(n5041), .B(n5040), .ZN(U2952)
         );
  INV_X1 U5590 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U5591 ( .A1(n5042), .A2(LWORD_REG_8__SCAN_IN), .ZN(n5044) );
  OAI211_X1 U5592 ( .C1(n5068), .C2(n5045), .A(n5044), .B(n5043), .ZN(U2947)
         );
  INV_X1 U5593 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U5594 ( .A1(n5065), .A2(UWORD_REG_1__SCAN_IN), .ZN(n5047) );
  OAI211_X1 U5595 ( .C1(n5068), .C2(n5107), .A(n5047), .B(n5046), .ZN(U2925)
         );
  NAND2_X1 U5596 ( .A1(n5048), .A2(n5175), .ZN(n5054) );
  NAND4_X1 U5597 ( .A1(n3901), .A2(n5050), .A3(n5175), .A4(n5049), .ZN(n5051)
         );
  NOR2_X1 U5598 ( .A1(n5052), .A2(n5051), .ZN(n5176) );
  NAND2_X1 U5599 ( .A1(n5176), .A2(n6103), .ZN(n5053) );
  AND2_X1 U5600 ( .A1(n3900), .A2(n5219), .ZN(n6006) );
  INV_X1 U5601 ( .A(n6006), .ZN(n5055) );
  AND2_X1 U5602 ( .A1(n5055), .A2(n3672), .ZN(n5057) );
  INV_X1 U5603 ( .A(n5057), .ZN(n5056) );
  INV_X1 U5604 ( .A(DATAI_0_), .ZN(n5199) );
  INV_X1 U5605 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7174) );
  INV_X1 U5606 ( .A(n5058), .ZN(n5863) );
  OAI222_X1 U5607 ( .A1(n6394), .A2(n5199), .B1(n6391), .B2(n7174), .C1(n7570), 
        .C2(n5863), .ZN(U2891) );
  INV_X1 U5608 ( .A(DATAI_1_), .ZN(n5207) );
  NOR2_X1 U5609 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  OR2_X1 U5610 ( .A1(n5076), .A2(n5061), .ZN(n7355) );
  OAI222_X1 U5611 ( .A1(n5207), .A2(n6394), .B1(n6391), .B2(n4991), .C1(n7570), 
        .C2(n7355), .ZN(U2890) );
  INV_X1 U5612 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U5613 ( .A1(n5065), .A2(UWORD_REG_0__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U5614 ( .A1(n5062), .A2(DATAI_0_), .ZN(n5066) );
  OAI211_X1 U5615 ( .C1(n5064), .C2(n5068), .A(n5063), .B(n5066), .ZN(U2924)
         );
  NAND2_X1 U5616 ( .A1(n5065), .A2(LWORD_REG_0__SCAN_IN), .ZN(n5067) );
  OAI211_X1 U5617 ( .C1(n7174), .C2(n5068), .A(n5067), .B(n5066), .ZN(U2939)
         );
  AOI22_X1 U5618 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7330), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5071) );
  INV_X1 U5619 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U5620 ( .A1(n6513), .A2(n5069), .ZN(n5070) );
  OAI211_X1 U5621 ( .C1(n7355), .C2(n6509), .A(n5071), .B(n5070), .ZN(n5072)
         );
  INV_X1 U5622 ( .A(n5072), .ZN(n5073) );
  OAI21_X1 U5623 ( .B1(n5074), .B2(n7482), .A(n5073), .ZN(U2985) );
  INV_X1 U5624 ( .A(DATAI_2_), .ZN(n5215) );
  INV_X1 U5625 ( .A(n5112), .ZN(n5079) );
  NOR3_X1 U5626 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(n5078) );
  NOR2_X1 U5627 ( .A1(n5079), .A2(n5078), .ZN(n6289) );
  INV_X1 U5628 ( .A(n6289), .ZN(n5181) );
  OAI222_X1 U5629 ( .A1(n6394), .A2(n5215), .B1(n6391), .B2(n5003), .C1(n7570), 
        .C2(n5181), .ZN(U2889) );
  XNOR2_X1 U5630 ( .A(n3691), .B(n5081), .ZN(n5103) );
  INV_X1 U5631 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7199) );
  NOR2_X1 U5632 ( .A1(n6759), .A2(n7199), .ZN(n5099) );
  AOI21_X1 U5633 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5099), 
        .ZN(n5082) );
  OAI21_X1 U5634 ( .B1(n7294), .B2(n6292), .A(n5082), .ZN(n5083) );
  AOI21_X1 U5635 ( .B1(n6289), .B2(n6534), .A(n5083), .ZN(n5084) );
  OAI21_X1 U5636 ( .B1(n5103), .B2(n7482), .A(n5084), .ZN(U2984) );
  NOR2_X1 U5637 ( .A1(n5937), .A2(n5936), .ZN(n5086) );
  OR2_X1 U5638 ( .A1(n6732), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5085)
         );
  AND2_X1 U5639 ( .A1(n5085), .A2(n7347), .ZN(n6563) );
  OAI21_X1 U5640 ( .B1(n6727), .B2(n5086), .A(n6563), .ZN(n5511) );
  NOR2_X1 U5641 ( .A1(n5936), .A2(n6741), .ZN(n5088) );
  AOI22_X1 U5642 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5511), .B1(n5088), 
        .B2(n5937), .ZN(n5102) );
  NAND2_X1 U5643 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5089) );
  OAI21_X1 U5644 ( .B1(n5936), .B2(n7349), .A(n5937), .ZN(n5631) );
  OAI21_X1 U5645 ( .B1(n5937), .B2(n5089), .A(n5631), .ZN(n5100) );
  NAND2_X1 U5646 ( .A1(n7351), .A2(n6018), .ZN(n5092) );
  INV_X1 U5647 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U5648 ( .A1(n5092), .A2(n5091), .ZN(n5097) );
  MUX2_X1 U5649 ( .A(n6058), .B(n5523), .S(EBX_REG_2__SCAN_IN), .Z(n5094) );
  OAI21_X1 U5650 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6114), .A(n5094), 
        .ZN(n5096) );
  INV_X1 U5651 ( .A(n5293), .ZN(n5095) );
  AOI21_X1 U5652 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n6290) );
  INV_X1 U5653 ( .A(n6290), .ZN(n5179) );
  NOR2_X1 U5654 ( .A1(n7342), .A2(n5179), .ZN(n5098) );
  AOI211_X1 U5655 ( .C1(n6731), .C2(n5100), .A(n5099), .B(n5098), .ZN(n5101)
         );
  OAI211_X1 U5656 ( .C1(n5103), .C2(n6765), .A(n5102), .B(n5101), .ZN(U3016)
         );
  AOI22_X1 U5657 ( .A1(n7182), .A2(UWORD_REG_14__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5104) );
  OAI21_X1 U5658 ( .B1(n4999), .B2(n5110), .A(n5104), .ZN(U2893) );
  AOI22_X1 U5659 ( .A1(n7182), .A2(UWORD_REG_0__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5105) );
  OAI21_X1 U5660 ( .B1(n5064), .B2(n5110), .A(n5105), .ZN(U2907) );
  AOI22_X1 U5661 ( .A1(n7182), .A2(UWORD_REG_1__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5106) );
  OAI21_X1 U5662 ( .B1(n5107), .B2(n5110), .A(n5106), .ZN(U2906) );
  AOI22_X1 U5663 ( .A1(n7182), .A2(UWORD_REG_2__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5108) );
  OAI21_X1 U5664 ( .B1(n5006), .B2(n5110), .A(n5108), .ZN(U2905) );
  AOI22_X1 U5665 ( .A1(n7182), .A2(UWORD_REG_3__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5109) );
  OAI21_X1 U5666 ( .B1(n5001), .B2(n5110), .A(n5109), .ZN(U2904) );
  INV_X1 U5667 ( .A(DATAI_3_), .ZN(n5115) );
  AND2_X1 U5668 ( .A1(n5112), .A2(n5111), .ZN(n5114) );
  OR2_X1 U5669 ( .A1(n5114), .A2(n5113), .ZN(n5856) );
  OAI222_X1 U5670 ( .A1(n5115), .A2(n6394), .B1(n6391), .B2(n5033), .C1(n7570), 
        .C2(n5856), .ZN(U2888) );
  NAND2_X1 U5671 ( .A1(n5854), .A2(n5130), .ZN(n5128) );
  AOI21_X1 U5672 ( .B1(n4906), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n5116), 
        .ZN(n5117) );
  NOR2_X1 U5673 ( .A1(n3674), .A2(n5117), .ZN(n6768) );
  NAND2_X1 U5674 ( .A1(n6100), .A2(n6095), .ZN(n5137) );
  NAND2_X1 U5675 ( .A1(n6086), .A2(n3834), .ZN(n5119) );
  INV_X1 U5676 ( .A(n5134), .ZN(n5118) );
  AND2_X1 U5677 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U5678 ( .A1(n5137), .A2(n5119), .B1(n5118), .B2(n5120), .ZN(n5122)
         );
  OR2_X1 U5679 ( .A1(n5134), .A2(n5120), .ZN(n5121) );
  MUX2_X1 U5680 ( .A(n5122), .B(n5121), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5125) );
  NAND2_X1 U5681 ( .A1(n6086), .A2(n5123), .ZN(n5124) );
  OAI211_X1 U5682 ( .C1(n6768), .C2(n5132), .A(n5125), .B(n5124), .ZN(n5126)
         );
  INV_X1 U5683 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U5684 ( .A1(n5128), .A2(n5127), .ZN(n6767) );
  MUX2_X1 U5685 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6767), .S(n7495), 
        .Z(n7505) );
  INV_X1 U5686 ( .A(n5130), .ZN(n5131) );
  OR2_X1 U5687 ( .A1(n5129), .A2(n5131), .ZN(n5139) );
  XNOR2_X1 U5688 ( .A(n4906), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5136)
         );
  XNOR2_X1 U5689 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5133) );
  OAI22_X1 U5690 ( .A1(n5134), .A2(n5133), .B1(n5132), .B2(n5136), .ZN(n5135)
         );
  AOI21_X1 U5691 ( .B1(n5137), .B2(n5136), .A(n5135), .ZN(n5138) );
  NAND2_X1 U5692 ( .A1(n5139), .A2(n5138), .ZN(n6082) );
  NAND2_X1 U5693 ( .A1(n6082), .A2(n7495), .ZN(n5141) );
  OR2_X1 U5694 ( .A1(n7495), .A2(n3834), .ZN(n5140) );
  NAND2_X1 U5695 ( .A1(n5141), .A2(n5140), .ZN(n7502) );
  NAND3_X1 U5696 ( .A1(n7505), .A2(n5711), .A3(n7502), .ZN(n5144) );
  INV_X1 U5697 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7483) );
  AND2_X1 U5698 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7483), .ZN(n5142) );
  NAND2_X1 U5699 ( .A1(n5144), .A2(n5143), .ZN(n7515) );
  NAND2_X1 U5700 ( .A1(n7515), .A2(n5145), .ZN(n5152) );
  OR2_X1 U5701 ( .A1(n5147), .A2(n3802), .ZN(n5148) );
  XNOR2_X1 U5702 ( .A(n5148), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7488)
         );
  NOR2_X1 U5703 ( .A1(n3692), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5151) );
  MUX2_X1 U5704 ( .A(n7495), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5149) );
  NOR2_X1 U5705 ( .A1(n5149), .A2(n7490), .ZN(n5150) );
  AOI21_X1 U5706 ( .B1(n7488), .B2(n5151), .A(n5150), .ZN(n7492) );
  NAND2_X1 U5707 ( .A1(n5152), .A2(n7492), .ZN(n7537) );
  OAI21_X1 U5708 ( .B1(n7537), .B2(FLUSH_REG_SCAN_IN), .A(n7531), .ZN(n5153)
         );
  NAND2_X1 U5709 ( .A1(n7522), .A2(n5711), .ZN(n7542) );
  NAND2_X1 U5710 ( .A1(n5153), .A2(n5227), .ZN(n7556) );
  NAND2_X1 U5711 ( .A1(n7556), .A2(n5575), .ZN(n5182) );
  XNOR2_X1 U5712 ( .A(n3689), .B(STATEBS16_REG_SCAN_IN), .ZN(n5154) );
  OAI21_X1 U5713 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5711), .A(n7556), .ZN(
        n7549) );
  OAI222_X1 U5714 ( .A1(n7556), .A2(n5348), .B1(n5182), .B2(n5154), .C1(n4904), 
        .C2(n7549), .ZN(U3464) );
  OAI21_X1 U5715 ( .B1(n5113), .B2(n5156), .A(n5333), .ZN(n5763) );
  INV_X1 U5716 ( .A(DATAI_4_), .ZN(n5195) );
  OAI222_X1 U5717 ( .A1(n5763), .A2(n7570), .B1(n6391), .B2(n7179), .C1(n6394), 
        .C2(n5195), .ZN(U2887) );
  AND2_X1 U5718 ( .A1(n4137), .A2(n3688), .ZN(n5158) );
  OR2_X1 U5719 ( .A1(n5456), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5577) );
  OAI21_X1 U5720 ( .B1(n5163), .B2(n5456), .A(n5577), .ZN(n5160) );
  INV_X1 U5721 ( .A(n5160), .ZN(n5159) );
  AND2_X1 U5722 ( .A1(n5854), .A2(n4310), .ZN(n5310) );
  NOR2_X1 U5723 ( .A1(n5129), .A2(n4054), .ZN(n5657) );
  NAND3_X1 U5724 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5348), .ZN(n5651) );
  NOR2_X1 U5725 ( .A1(n7557), .A2(n5651), .ZN(n5166) );
  AOI21_X1 U5726 ( .B1(n5310), .B2(n5657), .A(n5166), .ZN(n5161) );
  OAI22_X1 U5727 ( .A1(n5159), .A2(n5161), .B1(n5651), .B2(n7522), .ZN(n5531)
         );
  INV_X1 U5728 ( .A(n5531), .ZN(n5174) );
  NAND2_X1 U5729 ( .A1(n5396), .A2(DATAI_5_), .ZN(n5888) );
  AOI22_X1 U5730 ( .A1(n5161), .A2(n5160), .B1(n5456), .B2(n5651), .ZN(n5162)
         );
  NAND2_X1 U5731 ( .A1(n5461), .A2(n5162), .ZN(n5532) );
  NAND2_X1 U5732 ( .A1(n5532), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5169)
         );
  AND2_X1 U5733 ( .A1(n6534), .A2(DATAI_29_), .ZN(n5890) );
  NAND2_X1 U5734 ( .A1(n6534), .A2(DATAI_21_), .ZN(n5893) );
  OR2_X1 U5735 ( .A1(n5164), .A2(n7533), .ZN(n5226) );
  NAND2_X1 U5736 ( .A1(n5220), .A2(n5165), .ZN(n5887) );
  INV_X1 U5737 ( .A(n5166), .ZN(n5534) );
  OAI22_X1 U5738 ( .A1(n5537), .A2(n5893), .B1(n5887), .B2(n5534), .ZN(n5167)
         );
  AOI21_X1 U5739 ( .B1(n5890), .B2(n5822), .A(n5167), .ZN(n5168) );
  OAI211_X1 U5740 ( .C1(n5174), .C2(n5888), .A(n5169), .B(n5168), .ZN(U3129)
         );
  NAND2_X1 U5741 ( .A1(n5396), .A2(DATAI_3_), .ZN(n5901) );
  NAND2_X1 U5742 ( .A1(n5532), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5173)
         );
  AND2_X1 U5743 ( .A1(n6534), .A2(DATAI_27_), .ZN(n5903) );
  NAND2_X1 U5744 ( .A1(n6534), .A2(DATAI_19_), .ZN(n5906) );
  NAND2_X1 U5745 ( .A1(n5220), .A2(n5170), .ZN(n5900) );
  OAI22_X1 U5746 ( .A1(n5537), .A2(n5906), .B1(n5900), .B2(n5534), .ZN(n5171)
         );
  AOI21_X1 U5747 ( .B1(n5903), .B2(n5822), .A(n5171), .ZN(n5172) );
  OAI211_X1 U5748 ( .C1(n5174), .C2(n5901), .A(n5173), .B(n5172), .ZN(U3127)
         );
  NAND2_X1 U5749 ( .A1(n6099), .A2(n5175), .ZN(n5178) );
  NAND2_X1 U5750 ( .A1(n5176), .A2(n6018), .ZN(n5177) );
  OAI21_X4 U5751 ( .B1(n6100), .B2(n5178), .A(n5177), .ZN(n6352) );
  INV_X1 U5752 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5180) );
  OAI222_X1 U5753 ( .A1(n5181), .A2(n6355), .B1(n6352), .B2(n5180), .C1(n5179), 
        .C2(n6359), .ZN(U2857) );
  INV_X1 U5754 ( .A(n5854), .ZN(n5186) );
  INV_X1 U5755 ( .A(n4137), .ZN(n5441) );
  NOR2_X1 U5756 ( .A1(n3688), .A2(n7303), .ZN(n6092) );
  NAND2_X1 U5757 ( .A1(n6092), .A2(n3706), .ZN(n6091) );
  INV_X1 U5758 ( .A(n5182), .ZN(n7553) );
  INV_X1 U5759 ( .A(n3664), .ZN(n5346) );
  NAND2_X1 U5760 ( .A1(n5346), .A2(n6091), .ZN(n5183) );
  OAI211_X1 U5761 ( .C1(n5441), .C2(n6091), .A(n7553), .B(n5183), .ZN(n5185)
         );
  INV_X1 U5762 ( .A(n7556), .ZN(n7551) );
  NAND2_X1 U5763 ( .A1(n7551), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5184) );
  OAI211_X1 U5764 ( .C1(n5186), .C2(n7549), .A(n5185), .B(n5184), .ZN(U3462)
         );
  AND2_X1 U5765 ( .A1(n4137), .A2(n4301), .ZN(n5187) );
  NAND2_X1 U5766 ( .A1(n3706), .A2(n5187), .ZN(n5238) );
  NAND2_X1 U5767 ( .A1(n6534), .A2(DATAI_20_), .ZN(n7653) );
  NAND3_X1 U5768 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5240) );
  OR2_X1 U5769 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5240), .ZN(n5229)
         );
  OR2_X1 U5770 ( .A1(n5652), .A2(n7506), .ZN(n5194) );
  AND2_X1 U5771 ( .A1(n5194), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5582) );
  AND2_X1 U5772 ( .A1(n5193), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5874) );
  NOR2_X1 U5773 ( .A1(n5227), .A2(n5874), .ZN(n5363) );
  INV_X1 U5774 ( .A(n5363), .ZN(n5543) );
  AOI211_X1 U5775 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5229), .A(n5582), .B(
        n5543), .ZN(n5192) );
  NOR2_X1 U5776 ( .A1(n5129), .A2(n4904), .ZN(n5550) );
  INV_X1 U5777 ( .A(n5550), .ZN(n5189) );
  INV_X1 U5778 ( .A(n5577), .ZN(n5188) );
  NAND2_X1 U5779 ( .A1(n5189), .A2(n5188), .ZN(n5191) );
  OR2_X1 U5780 ( .A1(n5854), .A2(n5456), .ZN(n5650) );
  INV_X1 U5781 ( .A(n5650), .ZN(n5866) );
  NOR2_X1 U5782 ( .A1(n5550), .A2(n5456), .ZN(n5539) );
  OAI211_X1 U5783 ( .C1(n5866), .C2(n5539), .A(n5537), .B(n5271), .ZN(n5190)
         );
  NAND3_X1 U5784 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(n5224) );
  NAND2_X1 U5785 ( .A1(n5224), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5198)
         );
  AND2_X1 U5786 ( .A1(n6534), .A2(DATAI_28_), .ZN(n7670) );
  NAND2_X1 U5787 ( .A1(n5220), .A2(n3899), .ZN(n7667) );
  AND2_X1 U5788 ( .A1(n5854), .A2(n5575), .ZN(n5876) );
  OR2_X1 U5789 ( .A1(n5193), .A2(n7522), .ZN(n5548) );
  INV_X1 U5790 ( .A(n5548), .ZN(n5659) );
  INV_X1 U5791 ( .A(n5194), .ZN(n5579) );
  AOI22_X1 U5792 ( .A1(n5876), .A2(n5550), .B1(n5659), .B2(n5579), .ZN(n5228)
         );
  NOR2_X1 U5793 ( .A1(n5195), .A2(n5227), .ZN(n5773) );
  OAI22_X1 U5794 ( .A1(n7667), .A2(n5229), .B1(n5228), .B2(n7673), .ZN(n5196)
         );
  AOI21_X1 U5795 ( .B1(n7670), .B2(n5231), .A(n5196), .ZN(n5197) );
  OAI211_X1 U5796 ( .C1(n5271), .C2(n7653), .A(n5198), .B(n5197), .ZN(U3136)
         );
  NAND2_X1 U5797 ( .A1(n6534), .A2(DATAI_16_), .ZN(n7597) );
  NAND2_X1 U5798 ( .A1(n5224), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5202)
         );
  AND2_X1 U5799 ( .A1(n6534), .A2(DATAI_24_), .ZN(n7605) );
  NAND2_X1 U5800 ( .A1(n5220), .A2(n5721), .ZN(n7601) );
  NOR2_X1 U5801 ( .A1(n5199), .A2(n5227), .ZN(n5498) );
  OAI22_X1 U5802 ( .A1(n7601), .A2(n5229), .B1(n5228), .B2(n7608), .ZN(n5200)
         );
  AOI21_X1 U5803 ( .B1(n7605), .B2(n5231), .A(n5200), .ZN(n5201) );
  OAI211_X1 U5804 ( .C1(n5271), .C2(n7597), .A(n5202), .B(n5201), .ZN(U3132)
         );
  NAND2_X1 U5805 ( .A1(n5224), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5205)
         );
  OAI22_X1 U5806 ( .A1(n5888), .A2(n5228), .B1(n5887), .B2(n5229), .ZN(n5203)
         );
  AOI21_X1 U5807 ( .B1(n5890), .B2(n5231), .A(n5203), .ZN(n5204) );
  OAI211_X1 U5808 ( .C1(n5271), .C2(n5893), .A(n5205), .B(n5204), .ZN(U3137)
         );
  NAND2_X1 U5809 ( .A1(n6534), .A2(DATAI_17_), .ZN(n7620) );
  NAND2_X1 U5810 ( .A1(n5224), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5210)
         );
  AND2_X1 U5811 ( .A1(n6534), .A2(DATAI_25_), .ZN(n7622) );
  NAND2_X1 U5812 ( .A1(n5220), .A2(n5206), .ZN(n7625) );
  NOR2_X1 U5813 ( .A1(n5207), .A2(n5227), .ZN(n5790) );
  OAI22_X1 U5814 ( .A1(n7625), .A2(n5229), .B1(n5228), .B2(n7631), .ZN(n5208)
         );
  AOI21_X1 U5815 ( .B1(n7622), .B2(n5231), .A(n5208), .ZN(n5209) );
  OAI211_X1 U5816 ( .C1(n5271), .C2(n7620), .A(n5210), .B(n5209), .ZN(U3133)
         );
  NAND2_X1 U5817 ( .A1(n5224), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5213)
         );
  OAI22_X1 U5818 ( .A1(n5901), .A2(n5228), .B1(n5900), .B2(n5229), .ZN(n5211)
         );
  AOI21_X1 U5819 ( .B1(n5903), .B2(n5231), .A(n5211), .ZN(n5212) );
  OAI211_X1 U5820 ( .C1(n5271), .C2(n5906), .A(n5213), .B(n5212), .ZN(U3135)
         );
  NAND2_X1 U5821 ( .A1(n6534), .A2(DATAI_18_), .ZN(n5886) );
  NAND2_X1 U5822 ( .A1(n5224), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5218)
         );
  AND2_X1 U5823 ( .A1(n6534), .A2(DATAI_26_), .ZN(n7649) );
  NAND2_X1 U5824 ( .A1(n5220), .A2(n5214), .ZN(n7646) );
  NOR2_X1 U5825 ( .A1(n5215), .A2(n5227), .ZN(n5785) );
  OAI22_X1 U5826 ( .A1(n7646), .A2(n5229), .B1(n5228), .B2(n7652), .ZN(n5216)
         );
  AOI21_X1 U5827 ( .B1(n7649), .B2(n5231), .A(n5216), .ZN(n5217) );
  OAI211_X1 U5828 ( .C1(n5271), .C2(n5886), .A(n5218), .B(n5217), .ZN(U3134)
         );
  NAND2_X1 U5829 ( .A1(n6534), .A2(DATAI_23_), .ZN(n7707) );
  NAND2_X1 U5830 ( .A1(n5224), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5223)
         );
  AND2_X1 U5831 ( .A1(n6534), .A2(DATAI_31_), .ZN(n7730) );
  NAND2_X1 U5832 ( .A1(n5220), .A2(n5219), .ZN(n7738) );
  INV_X1 U5833 ( .A(DATAI_7_), .ZN(n5628) );
  NOR2_X1 U5834 ( .A1(n5628), .A2(n5227), .ZN(n5768) );
  OAI22_X1 U5835 ( .A1(n7738), .A2(n5229), .B1(n5228), .B2(n7747), .ZN(n5221)
         );
  AOI21_X1 U5836 ( .B1(n7730), .B2(n5231), .A(n5221), .ZN(n5222) );
  OAI211_X1 U5837 ( .C1(n5271), .C2(n7707), .A(n5223), .B(n5222), .ZN(U3139)
         );
  NAND2_X1 U5838 ( .A1(n6534), .A2(DATAI_22_), .ZN(n7680) );
  NAND2_X1 U5839 ( .A1(n5224), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5233)
         );
  NAND2_X1 U5840 ( .A1(n6534), .A2(DATAI_30_), .ZN(n7674) );
  INV_X1 U5841 ( .A(n7674), .ZN(n7693) );
  NOR2_X1 U5842 ( .A1(n5226), .A2(n5225), .ZN(n7691) );
  INV_X1 U5843 ( .A(n7691), .ZN(n7679) );
  INV_X1 U5844 ( .A(DATAI_6_), .ZN(n5696) );
  NOR2_X1 U5845 ( .A1(n5696), .A2(n5227), .ZN(n7144) );
  OAI22_X1 U5846 ( .A1(n7679), .A2(n5229), .B1(n5228), .B2(n7697), .ZN(n5230)
         );
  AOI21_X1 U5847 ( .B1(n7693), .B2(n5231), .A(n5230), .ZN(n5232) );
  OAI211_X1 U5848 ( .C1(n5271), .C2(n7680), .A(n5233), .B(n5232), .ZN(U3138)
         );
  INV_X1 U5849 ( .A(n5903), .ZN(n5610) );
  NOR2_X1 U5850 ( .A1(n5234), .A2(n7506), .ZN(n5243) );
  AOI21_X1 U5851 ( .B1(n5310), .B2(n5550), .A(n5243), .ZN(n5239) );
  INV_X1 U5852 ( .A(n5238), .ZN(n5235) );
  OAI21_X1 U5853 ( .B1(n5235), .B2(n6509), .A(n5577), .ZN(n5236) );
  AOI22_X1 U5854 ( .A1(n5239), .A2(n5236), .B1(n5456), .B2(n5240), .ZN(n5237)
         );
  NAND2_X1 U5855 ( .A1(n5461), .A2(n5237), .ZN(n5265) );
  NAND2_X1 U5856 ( .A1(n5265), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5246)
         );
  OR2_X1 U5857 ( .A1(n5238), .A2(n4308), .ZN(n7147) );
  INV_X1 U5858 ( .A(n5906), .ZN(n5607) );
  INV_X1 U5859 ( .A(n5239), .ZN(n5242) );
  INV_X1 U5860 ( .A(n5240), .ZN(n5241) );
  AOI22_X1 U5861 ( .A1(n5242), .A2(n5575), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5241), .ZN(n5267) );
  INV_X1 U5862 ( .A(n5243), .ZN(n5266) );
  OAI22_X1 U5863 ( .A1(n5267), .A2(n5901), .B1(n5900), .B2(n5266), .ZN(n5244)
         );
  AOI21_X1 U5864 ( .B1(n5432), .B2(n5607), .A(n5244), .ZN(n5245) );
  OAI211_X1 U5865 ( .C1(n5271), .C2(n5610), .A(n5246), .B(n5245), .ZN(U3143)
         );
  INV_X1 U5866 ( .A(n5890), .ZN(n5601) );
  NAND2_X1 U5867 ( .A1(n5265), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5249)
         );
  INV_X1 U5868 ( .A(n5893), .ZN(n5598) );
  OAI22_X1 U5869 ( .A1(n5267), .A2(n5888), .B1(n5887), .B2(n5266), .ZN(n5247)
         );
  AOI21_X1 U5870 ( .B1(n5432), .B2(n5598), .A(n5247), .ZN(n5248) );
  OAI211_X1 U5871 ( .C1(n5271), .C2(n5601), .A(n5249), .B(n5248), .ZN(U3145)
         );
  INV_X1 U5872 ( .A(n7670), .ZN(n5778) );
  NAND2_X1 U5873 ( .A1(n5265), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5252)
         );
  INV_X1 U5874 ( .A(n7653), .ZN(n7669) );
  OAI22_X1 U5875 ( .A1(n5267), .A2(n7673), .B1(n7667), .B2(n5266), .ZN(n5250)
         );
  AOI21_X1 U5876 ( .B1(n5432), .B2(n7669), .A(n5250), .ZN(n5251) );
  OAI211_X1 U5877 ( .C1(n5271), .C2(n5778), .A(n5252), .B(n5251), .ZN(U3144)
         );
  INV_X1 U5878 ( .A(n7730), .ZN(n7739) );
  NAND2_X1 U5879 ( .A1(n5265), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5255)
         );
  INV_X1 U5880 ( .A(n7707), .ZN(n7743) );
  OAI22_X1 U5881 ( .A1(n5267), .A2(n7747), .B1(n7738), .B2(n5266), .ZN(n5253)
         );
  AOI21_X1 U5882 ( .B1(n5432), .B2(n7743), .A(n5253), .ZN(n5254) );
  OAI211_X1 U5883 ( .C1(n5271), .C2(n7739), .A(n5255), .B(n5254), .ZN(U3147)
         );
  NAND2_X1 U5884 ( .A1(n5265), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5258)
         );
  INV_X1 U5885 ( .A(n7680), .ZN(n7692) );
  OAI22_X1 U5886 ( .A1(n5267), .A2(n7697), .B1(n7679), .B2(n5266), .ZN(n5256)
         );
  AOI21_X1 U5887 ( .B1(n5432), .B2(n7692), .A(n5256), .ZN(n5257) );
  OAI211_X1 U5888 ( .C1(n5271), .C2(n7674), .A(n5258), .B(n5257), .ZN(U3146)
         );
  INV_X1 U5889 ( .A(n7605), .ZN(n5825) );
  NAND2_X1 U5890 ( .A1(n5265), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5261)
         );
  INV_X1 U5891 ( .A(n7597), .ZN(n7603) );
  OAI22_X1 U5892 ( .A1(n5267), .A2(n7608), .B1(n7601), .B2(n5266), .ZN(n5259)
         );
  AOI21_X1 U5893 ( .B1(n5432), .B2(n7603), .A(n5259), .ZN(n5260) );
  OAI211_X1 U5894 ( .C1(n5825), .C2(n5271), .A(n5261), .B(n5260), .ZN(U3140)
         );
  INV_X1 U5895 ( .A(n7649), .ZN(n7632) );
  NAND2_X1 U5896 ( .A1(n5265), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5264)
         );
  INV_X1 U5897 ( .A(n5886), .ZN(n7648) );
  OAI22_X1 U5898 ( .A1(n5267), .A2(n7652), .B1(n7646), .B2(n5266), .ZN(n5262)
         );
  AOI21_X1 U5899 ( .B1(n5432), .B2(n7648), .A(n5262), .ZN(n5263) );
  OAI211_X1 U5900 ( .C1(n5271), .C2(n7632), .A(n5264), .B(n5263), .ZN(U3142)
         );
  INV_X1 U5901 ( .A(n7622), .ZN(n7626) );
  NAND2_X1 U5902 ( .A1(n5265), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5270)
         );
  INV_X1 U5903 ( .A(n7620), .ZN(n7628) );
  OAI22_X1 U5904 ( .A1(n5267), .A2(n7631), .B1(n7625), .B2(n5266), .ZN(n5268)
         );
  AOI21_X1 U5905 ( .B1(n5432), .B2(n7628), .A(n5268), .ZN(n5269) );
  OAI211_X1 U5906 ( .C1(n5271), .C2(n7626), .A(n5270), .B(n5269), .ZN(U3141)
         );
  NOR2_X1 U5907 ( .A1(n4137), .A2(n3689), .ZN(n5272) );
  NAND2_X1 U5908 ( .A1(n3706), .A2(n5272), .ZN(n5280) );
  INV_X1 U5909 ( .A(n5280), .ZN(n5273) );
  OAI21_X1 U5910 ( .B1(n5273), .B2(n5456), .A(n5577), .ZN(n5277) );
  INV_X1 U5911 ( .A(n4310), .ZN(n7548) );
  OR2_X1 U5912 ( .A1(n5854), .A2(n7548), .ZN(n5458) );
  INV_X1 U5913 ( .A(n5458), .ZN(n5438) );
  NAND2_X1 U5914 ( .A1(n5438), .A2(n5657), .ZN(n5274) );
  NAND3_X1 U5915 ( .A1(n5348), .A2(n7506), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5361) );
  NOR2_X1 U5916 ( .A1(n7557), .A2(n5361), .ZN(n7721) );
  INV_X1 U5917 ( .A(n7721), .ZN(n5284) );
  NAND2_X1 U5918 ( .A1(n5274), .A2(n5284), .ZN(n5275) );
  INV_X1 U5919 ( .A(n5361), .ZN(n5279) );
  AOI22_X1 U5920 ( .A1(n5277), .A2(n5275), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5279), .ZN(n7727) );
  INV_X1 U5921 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U5922 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  OAI211_X1 U5923 ( .C1(n5575), .C2(n5279), .A(n5278), .B(n5461), .ZN(n7724)
         );
  NOR2_X1 U5924 ( .A1(n5627), .A2(n5893), .ZN(n5282) );
  OAI22_X1 U5925 ( .A1(n5367), .A2(n5601), .B1(n5887), .B2(n5284), .ZN(n5281)
         );
  AOI211_X1 U5926 ( .C1(n7724), .C2(INSTQUEUE_REG_5__5__SCAN_IN), .A(n5282), 
        .B(n5281), .ZN(n5283) );
  OAI21_X1 U5927 ( .B1(n7727), .B2(n5888), .A(n5283), .ZN(U3065) );
  NOR2_X1 U5928 ( .A1(n5627), .A2(n5906), .ZN(n5286) );
  OAI22_X1 U5929 ( .A1(n5367), .A2(n5610), .B1(n5900), .B2(n5284), .ZN(n5285)
         );
  AOI211_X1 U5930 ( .C1(n7724), .C2(INSTQUEUE_REG_5__3__SCAN_IN), .A(n5286), 
        .B(n5285), .ZN(n5287) );
  OAI21_X1 U5931 ( .B1(n7727), .B2(n5901), .A(n5287), .ZN(U3063) );
  INV_X1 U5932 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5933 ( .A1(n6052), .A2(n5849), .ZN(n5291) );
  NAND2_X1 U5934 ( .A1(n6054), .A2(n5515), .ZN(n5289) );
  NAND2_X1 U5935 ( .A1(n6018), .A2(n5849), .ZN(n5288) );
  NAND3_X1 U5936 ( .A1(n5289), .A2(n6049), .A3(n5288), .ZN(n5290) );
  AND2_X1 U5937 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  NOR2_X1 U5938 ( .A1(n5478), .A2(n5294), .ZN(n5846) );
  AOI22_X1 U5939 ( .A1(n7284), .A2(n5846), .B1(n6353), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5295) );
  OAI21_X1 U5940 ( .B1(n5856), .B2(n6355), .A(n5295), .ZN(U2856) );
  NOR2_X1 U5941 ( .A1(n3706), .A2(n3688), .ZN(n5345) );
  AOI21_X1 U5942 ( .B1(n5302), .B2(STATEBS16_REG_SCAN_IN), .A(n5456), .ZN(
        n5299) );
  AND2_X1 U5943 ( .A1(n5129), .A2(n4054), .ZN(n5347) );
  AND2_X1 U5944 ( .A1(n5347), .A2(n5854), .ZN(n5584) );
  NAND2_X1 U5945 ( .A1(n5584), .A2(n4310), .ZN(n5296) );
  NAND3_X1 U5946 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n7501), .ZN(n5581) );
  NOR2_X1 U5947 ( .A1(n7557), .A2(n5581), .ZN(n5306) );
  INV_X1 U5948 ( .A(n5306), .ZN(n7698) );
  NAND2_X1 U5949 ( .A1(n5296), .A2(n7698), .ZN(n5297) );
  INV_X1 U5950 ( .A(n5581), .ZN(n5301) );
  AOI22_X1 U5951 ( .A1(n5299), .A2(n5297), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5301), .ZN(n7705) );
  INV_X1 U5952 ( .A(n5297), .ZN(n5298) );
  NAND2_X1 U5953 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  OAI211_X1 U5954 ( .C1(n5575), .C2(n5301), .A(n5300), .B(n5461), .ZN(n7702)
         );
  NAND2_X1 U5955 ( .A1(n5302), .A2(n7554), .ZN(n7699) );
  NAND2_X1 U5956 ( .A1(n5302), .A2(n4308), .ZN(n7708) );
  INV_X1 U5957 ( .A(n5887), .ZN(n5674) );
  AOI22_X1 U5958 ( .A1(n7701), .A2(n5890), .B1(n5674), .B2(n5306), .ZN(n5303)
         );
  OAI21_X1 U5959 ( .B1(n5893), .B2(n7699), .A(n5303), .ZN(n5304) );
  AOI21_X1 U5960 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n7702), .A(n5304), 
        .ZN(n5305) );
  OAI21_X1 U5961 ( .B1(n7705), .B2(n5888), .A(n5305), .ZN(U3113) );
  INV_X1 U5962 ( .A(n5900), .ZN(n5688) );
  AOI22_X1 U5963 ( .A1(n7701), .A2(n5903), .B1(n5688), .B2(n5306), .ZN(n5307)
         );
  OAI21_X1 U5964 ( .B1(n5906), .B2(n7699), .A(n5307), .ZN(n5308) );
  AOI21_X1 U5965 ( .B1(INSTQUEUE_REG_11__3__SCAN_IN), .B2(n7702), .A(n5308), 
        .ZN(n5309) );
  OAI21_X1 U5966 ( .B1(n7705), .B2(n5901), .A(n5309), .ZN(U3111) );
  AND2_X1 U5967 ( .A1(n5129), .A2(n4904), .ZN(n5875) );
  NAND3_X1 U5968 ( .A1(n7501), .A2(n5348), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5864) );
  NOR2_X1 U5969 ( .A1(n7557), .A2(n5864), .ZN(n7714) );
  AOI21_X1 U5970 ( .B1(n5310), .B2(n5875), .A(n7714), .ZN(n5313) );
  INV_X1 U5971 ( .A(n5395), .ZN(n5311) );
  OAI21_X1 U5972 ( .B1(n5319), .B2(n5456), .A(n5577), .ZN(n5315) );
  AOI22_X1 U5973 ( .A1(n5313), .A2(n5315), .B1(n5456), .B2(n5864), .ZN(n5312)
         );
  NAND2_X1 U5974 ( .A1(n5461), .A2(n5312), .ZN(n7717) );
  INV_X1 U5975 ( .A(n7717), .ZN(n5331) );
  INV_X1 U5976 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5324) );
  INV_X1 U5977 ( .A(n5313), .ZN(n5314) );
  NAND2_X1 U5978 ( .A1(n5315), .A2(n5314), .ZN(n5318) );
  INV_X1 U5979 ( .A(n5864), .ZN(n5316) );
  NAND2_X1 U5980 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5316), .ZN(n5317) );
  INV_X1 U5981 ( .A(n7720), .ZN(n5328) );
  INV_X1 U5982 ( .A(n5901), .ZN(n5689) );
  NAND2_X1 U5983 ( .A1(n7716), .A2(n5607), .ZN(n5321) );
  NAND2_X1 U5984 ( .A1(n5688), .A2(n7714), .ZN(n5320) );
  OAI211_X1 U5985 ( .C1(n5610), .C2(n5914), .A(n5321), .B(n5320), .ZN(n5322)
         );
  AOI21_X1 U5986 ( .B1(n5328), .B2(n5689), .A(n5322), .ZN(n5323) );
  OAI21_X1 U5987 ( .B1(n5331), .B2(n5324), .A(n5323), .ZN(U3095) );
  INV_X1 U5988 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5330) );
  INV_X1 U5989 ( .A(n5888), .ZN(n5675) );
  NAND2_X1 U5990 ( .A1(n7716), .A2(n5598), .ZN(n5326) );
  NAND2_X1 U5991 ( .A1(n5674), .A2(n7714), .ZN(n5325) );
  OAI211_X1 U5992 ( .C1(n5601), .C2(n5914), .A(n5326), .B(n5325), .ZN(n5327)
         );
  AOI21_X1 U5993 ( .B1(n5328), .B2(n5675), .A(n5327), .ZN(n5329) );
  OAI21_X1 U5994 ( .B1(n5331), .B2(n5330), .A(n5329), .ZN(U3097) );
  AOI21_X1 U5995 ( .B1(n5334), .B2(n5333), .A(n3683), .ZN(n7371) );
  INV_X1 U5996 ( .A(n7371), .ZN(n5484) );
  MUX2_X1 U5997 ( .A(n6058), .B(n6049), .S(EBX_REG_4__SCAN_IN), .Z(n5336) );
  OR2_X1 U5998 ( .A1(n6114), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5335)
         );
  NAND2_X1 U5999 ( .A1(n6054), .A2(n5337), .ZN(n5339) );
  INV_X1 U6000 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U6001 ( .A1(n6018), .A2(n7363), .ZN(n5338) );
  NAND3_X1 U6002 ( .A1(n5339), .A2(n5523), .A3(n5338), .ZN(n5340) );
  OAI21_X1 U6003 ( .B1(n6107), .B2(EBX_REG_5__SCAN_IN), .A(n5340), .ZN(n5341)
         );
  OR2_X1 U6004 ( .A1(n5480), .A2(n5341), .ZN(n5342) );
  NAND2_X1 U6005 ( .A1(n5525), .A2(n5342), .ZN(n7362) );
  INV_X1 U6006 ( .A(n7362), .ZN(n5343) );
  AOI22_X1 U6007 ( .A1(n7284), .A2(n5343), .B1(n6353), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5344) );
  OAI21_X1 U6008 ( .B1(n5484), .B2(n6355), .A(n5344), .ZN(U2854) );
  OAI21_X1 U6009 ( .B1(n5354), .B2(n5456), .A(n5577), .ZN(n5350) );
  INV_X1 U6010 ( .A(n5347), .ZN(n5493) );
  NOR3_X1 U6011 ( .A1(n5348), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5349) );
  INV_X1 U6012 ( .A(n5349), .ZN(n5487) );
  NOR2_X1 U6013 ( .A1(n7557), .A2(n5487), .ZN(n7728) );
  INV_X1 U6014 ( .A(n7728), .ZN(n7619) );
  OAI21_X1 U6015 ( .B1(n5458), .B2(n5493), .A(n7619), .ZN(n5352) );
  AOI22_X1 U6016 ( .A1(n5350), .A2(n5352), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5349), .ZN(n7736) );
  INV_X1 U6017 ( .A(n5350), .ZN(n5353) );
  NAND2_X1 U6018 ( .A1(n5456), .A2(n5487), .ZN(n5351) );
  OAI211_X1 U6019 ( .C1(n5353), .C2(n5352), .A(n5461), .B(n5351), .ZN(n7733)
         );
  AOI22_X1 U6020 ( .A1(n7731), .A2(n5890), .B1(n5674), .B2(n7728), .ZN(n5355)
         );
  OAI21_X1 U6021 ( .B1(n5893), .B2(n7643), .A(n5355), .ZN(n5356) );
  AOI21_X1 U6022 ( .B1(n7733), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n5356), 
        .ZN(n5357) );
  OAI21_X1 U6023 ( .B1(n7736), .B2(n5888), .A(n5357), .ZN(U3049) );
  AOI22_X1 U6024 ( .A1(n7731), .A2(n5903), .B1(n5688), .B2(n7728), .ZN(n5358)
         );
  OAI21_X1 U6025 ( .B1(n5906), .B2(n7643), .A(n5358), .ZN(n5359) );
  AOI21_X1 U6026 ( .B1(n7733), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n5359), 
        .ZN(n5360) );
  OAI21_X1 U6027 ( .B1(n7736), .B2(n5901), .A(n5360), .ZN(U3047) );
  NOR2_X1 U6028 ( .A1(n5657), .A2(n5456), .ZN(n5648) );
  OAI211_X1 U6029 ( .C1(n5876), .C2(n5648), .A(n7643), .B(n5367), .ZN(n5366)
         );
  OR2_X1 U6030 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5361), .ZN(n5390)
         );
  INV_X1 U6031 ( .A(n5652), .ZN(n5362) );
  NOR2_X1 U6032 ( .A1(n5653), .A2(n5362), .ZN(n5401) );
  NOR2_X1 U6033 ( .A1(n5401), .A2(n7522), .ZN(n5397) );
  AOI21_X1 U6034 ( .B1(n5390), .B2(STATE2_REG_3__SCAN_IN), .A(n5397), .ZN(
        n5365) );
  OR2_X1 U6035 ( .A1(n5657), .A2(n5577), .ZN(n5364) );
  AND2_X1 U6036 ( .A1(n5364), .A2(n5363), .ZN(n5654) );
  NAND3_X1 U6037 ( .A1(n5366), .A2(n5365), .A3(n5654), .ZN(n5389) );
  NAND2_X1 U6038 ( .A1(n5389), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5370) );
  AOI22_X1 U6039 ( .A1(n5866), .A2(n5657), .B1(n5401), .B2(n5659), .ZN(n5391)
         );
  OAI22_X1 U6040 ( .A1(n5391), .A2(n7673), .B1(n7667), .B2(n5390), .ZN(n5368)
         );
  AOI21_X1 U6041 ( .B1(n7669), .B2(n7722), .A(n5368), .ZN(n5369) );
  OAI211_X1 U6042 ( .C1(n7643), .C2(n5778), .A(n5370), .B(n5369), .ZN(U3056)
         );
  NAND2_X1 U6043 ( .A1(n5389), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5373) );
  OAI22_X1 U6044 ( .A1(n5391), .A2(n7608), .B1(n7601), .B2(n5390), .ZN(n5371)
         );
  AOI21_X1 U6045 ( .B1(n7603), .B2(n7722), .A(n5371), .ZN(n5372) );
  OAI211_X1 U6046 ( .C1(n7643), .C2(n5825), .A(n5373), .B(n5372), .ZN(U3052)
         );
  NAND2_X1 U6047 ( .A1(n5389), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5376) );
  OAI22_X1 U6048 ( .A1(n5391), .A2(n7747), .B1(n7738), .B2(n5390), .ZN(n5374)
         );
  AOI21_X1 U6049 ( .B1(n7743), .B2(n7722), .A(n5374), .ZN(n5375) );
  OAI211_X1 U6050 ( .C1(n7643), .C2(n7739), .A(n5376), .B(n5375), .ZN(U3059)
         );
  NAND2_X1 U6051 ( .A1(n5389), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5379) );
  OAI22_X1 U6052 ( .A1(n5391), .A2(n7652), .B1(n7646), .B2(n5390), .ZN(n5377)
         );
  AOI21_X1 U6053 ( .B1(n7648), .B2(n7722), .A(n5377), .ZN(n5378) );
  OAI211_X1 U6054 ( .C1(n7643), .C2(n7632), .A(n5379), .B(n5378), .ZN(U3054)
         );
  NAND2_X1 U6055 ( .A1(n5389), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5382) );
  OAI22_X1 U6056 ( .A1(n5888), .A2(n5391), .B1(n5887), .B2(n5390), .ZN(n5380)
         );
  AOI21_X1 U6057 ( .B1(n5598), .B2(n7722), .A(n5380), .ZN(n5381) );
  OAI211_X1 U6058 ( .C1(n7643), .C2(n5601), .A(n5382), .B(n5381), .ZN(U3057)
         );
  NAND2_X1 U6059 ( .A1(n5389), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5385) );
  OAI22_X1 U6060 ( .A1(n7679), .A2(n5390), .B1(n5391), .B2(n7697), .ZN(n5383)
         );
  AOI21_X1 U6061 ( .B1(n7692), .B2(n7722), .A(n5383), .ZN(n5384) );
  OAI211_X1 U6062 ( .C1(n7643), .C2(n7674), .A(n5385), .B(n5384), .ZN(U3058)
         );
  NAND2_X1 U6063 ( .A1(n5389), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5388) );
  OAI22_X1 U6064 ( .A1(n5901), .A2(n5391), .B1(n5900), .B2(n5390), .ZN(n5386)
         );
  AOI21_X1 U6065 ( .B1(n5607), .B2(n7722), .A(n5386), .ZN(n5387) );
  OAI211_X1 U6066 ( .C1(n7643), .C2(n5610), .A(n5388), .B(n5387), .ZN(U3055)
         );
  NAND2_X1 U6067 ( .A1(n5389), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5394) );
  OAI22_X1 U6068 ( .A1(n5391), .A2(n7631), .B1(n7625), .B2(n5390), .ZN(n5392)
         );
  AOI21_X1 U6069 ( .B1(n7628), .B2(n7722), .A(n5392), .ZN(n5393) );
  OAI211_X1 U6070 ( .C1(n7643), .C2(n7626), .A(n5394), .B(n5393), .ZN(U3053)
         );
  NOR2_X1 U6071 ( .A1(n5875), .A2(n5456), .ZN(n5865) );
  NAND2_X1 U6072 ( .A1(n5459), .A2(n4308), .ZN(n7740) );
  OAI211_X1 U6073 ( .C1(n5876), .C2(n5865), .A(n7740), .B(n7147), .ZN(n5400)
         );
  INV_X1 U6074 ( .A(n5876), .ZN(n5542) );
  NOR3_X1 U6075 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5462) );
  NAND2_X1 U6076 ( .A1(n5462), .A2(n7557), .ZN(n5403) );
  NAND2_X1 U6077 ( .A1(n5396), .A2(n5548), .ZN(n5867) );
  AOI211_X1 U6078 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5403), .A(n5397), .B(
        n5867), .ZN(n5398) );
  NAND3_X1 U6079 ( .A1(n5400), .A2(n5399), .A3(n5398), .ZN(n7150) );
  INV_X1 U6080 ( .A(n7150), .ZN(n5415) );
  INV_X1 U6081 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5408) );
  INV_X1 U6082 ( .A(n5875), .ZN(n5457) );
  NAND2_X1 U6083 ( .A1(n5401), .A2(n5874), .ZN(n5402) );
  OAI21_X1 U6084 ( .B1(n5650), .B2(n5457), .A(n5402), .ZN(n7143) );
  INV_X1 U6085 ( .A(n7143), .ZN(n5411) );
  NAND2_X1 U6086 ( .A1(n5432), .A2(n5903), .ZN(n5405) );
  INV_X1 U6087 ( .A(n5403), .ZN(n7145) );
  NAND2_X1 U6088 ( .A1(n5688), .A2(n7145), .ZN(n5404) );
  OAI211_X1 U6089 ( .C1(n5901), .C2(n5411), .A(n5405), .B(n5404), .ZN(n5406)
         );
  AOI21_X1 U6090 ( .B1(n7694), .B2(n5607), .A(n5406), .ZN(n5407) );
  OAI21_X1 U6091 ( .B1(n5415), .B2(n5408), .A(n5407), .ZN(U3023) );
  INV_X1 U6092 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6093 ( .A1(n5432), .A2(n5890), .ZN(n5410) );
  NAND2_X1 U6094 ( .A1(n5674), .A2(n7145), .ZN(n5409) );
  OAI211_X1 U6095 ( .C1(n5888), .C2(n5411), .A(n5410), .B(n5409), .ZN(n5412)
         );
  AOI21_X1 U6096 ( .B1(n7694), .B2(n5598), .A(n5412), .ZN(n5413) );
  OAI21_X1 U6097 ( .B1(n5415), .B2(n5414), .A(n5413), .ZN(U3025) );
  INV_X1 U6098 ( .A(n7667), .ZN(n7664) );
  AOI22_X1 U6099 ( .A1(n7664), .A2(n7145), .B1(n5773), .B2(n7143), .ZN(n5417)
         );
  NAND2_X1 U6100 ( .A1(n5432), .A2(n7670), .ZN(n5416) );
  OAI211_X1 U6101 ( .C1(n7740), .C2(n7653), .A(n5417), .B(n5416), .ZN(n5418)
         );
  AOI21_X1 U6102 ( .B1(n7150), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n5418), 
        .ZN(n5419) );
  INV_X1 U6103 ( .A(n5419), .ZN(U3024) );
  INV_X1 U6104 ( .A(n7601), .ZN(n7594) );
  AOI22_X1 U6105 ( .A1(n7594), .A2(n7145), .B1(n5498), .B2(n7143), .ZN(n5421)
         );
  NAND2_X1 U6106 ( .A1(n5432), .A2(n7605), .ZN(n5420) );
  OAI211_X1 U6107 ( .C1(n7740), .C2(n7597), .A(n5421), .B(n5420), .ZN(n5422)
         );
  AOI21_X1 U6108 ( .B1(n7150), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n5422), 
        .ZN(n5423) );
  INV_X1 U6109 ( .A(n5423), .ZN(U3020) );
  INV_X1 U6110 ( .A(n7625), .ZN(n7616) );
  AOI22_X1 U6111 ( .A1(n7616), .A2(n7145), .B1(n5790), .B2(n7143), .ZN(n5425)
         );
  NAND2_X1 U6112 ( .A1(n5432), .A2(n7622), .ZN(n5424) );
  OAI211_X1 U6113 ( .C1(n7740), .C2(n7620), .A(n5425), .B(n5424), .ZN(n5426)
         );
  AOI21_X1 U6114 ( .B1(n7150), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n5426), 
        .ZN(n5427) );
  INV_X1 U6115 ( .A(n5427), .ZN(U3021) );
  AOI22_X1 U6116 ( .A1(n7642), .A2(n7145), .B1(n5785), .B2(n7143), .ZN(n5429)
         );
  NAND2_X1 U6117 ( .A1(n5432), .A2(n7649), .ZN(n5428) );
  OAI211_X1 U6118 ( .C1(n7740), .C2(n5886), .A(n5429), .B(n5428), .ZN(n5430)
         );
  AOI21_X1 U6119 ( .B1(n7150), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n5430), 
        .ZN(n5431) );
  INV_X1 U6120 ( .A(n5431), .ZN(U3022) );
  INV_X1 U6121 ( .A(n7738), .ZN(n7729) );
  AOI22_X1 U6122 ( .A1(n7729), .A2(n7145), .B1(n5768), .B2(n7143), .ZN(n5434)
         );
  NAND2_X1 U6123 ( .A1(n5432), .A2(n7730), .ZN(n5433) );
  OAI211_X1 U6124 ( .C1(n7740), .C2(n7707), .A(n5434), .B(n5433), .ZN(n5435)
         );
  AOI21_X1 U6125 ( .B1(n7150), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n5435), 
        .ZN(n5436) );
  INV_X1 U6126 ( .A(n5436), .ZN(U3027) );
  INV_X1 U6127 ( .A(n6091), .ZN(n5437) );
  AOI21_X1 U6128 ( .B1(n5437), .B2(n5441), .A(n5456), .ZN(n5444) );
  NAND2_X1 U6129 ( .A1(n5438), .A2(n5550), .ZN(n5439) );
  NAND2_X1 U6130 ( .A1(n5439), .A2(n5742), .ZN(n5446) );
  NAND3_X1 U6131 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(n7506), .ZN(n5538) );
  INV_X1 U6132 ( .A(n5538), .ZN(n5440) );
  AOI22_X1 U6133 ( .A1(n5444), .A2(n5446), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5440), .ZN(n5749) );
  NAND3_X1 U6134 ( .A1(n3706), .A2(n5441), .A3(n3689), .ZN(n5442) );
  NOR2_X2 U6135 ( .A1(n5442), .A2(n4308), .ZN(n5911) );
  OAI22_X1 U6136 ( .A1(n5620), .A2(n7632), .B1(n7646), .B2(n5742), .ZN(n5443)
         );
  AOI21_X1 U6137 ( .B1(n5911), .B2(n7648), .A(n5443), .ZN(n5449) );
  INV_X1 U6138 ( .A(n5444), .ZN(n5447) );
  NAND2_X1 U6139 ( .A1(n5456), .A2(n5538), .ZN(n5445) );
  OAI211_X1 U6140 ( .C1(n5447), .C2(n5446), .A(n5461), .B(n5445), .ZN(n5746)
         );
  NAND2_X1 U6141 ( .A1(n5746), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5448) );
  OAI211_X1 U6142 ( .C1(n5749), .C2(n7652), .A(n5449), .B(n5448), .ZN(U3078)
         );
  OAI22_X1 U6143 ( .A1(n5620), .A2(n5601), .B1(n5887), .B2(n5742), .ZN(n5450)
         );
  AOI21_X1 U6144 ( .B1(n5911), .B2(n5598), .A(n5450), .ZN(n5452) );
  NAND2_X1 U6145 ( .A1(n5746), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6146 ( .C1(n5749), .C2(n5888), .A(n5452), .B(n5451), .ZN(U3081)
         );
  OAI22_X1 U6147 ( .A1(n5620), .A2(n5610), .B1(n5900), .B2(n5742), .ZN(n5453)
         );
  AOI21_X1 U6148 ( .B1(n5911), .B2(n5607), .A(n5453), .ZN(n5455) );
  NAND2_X1 U6149 ( .A1(n5746), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6150 ( .C1(n5749), .C2(n5901), .A(n5455), .B(n5454), .ZN(U3079)
         );
  OAI21_X1 U6151 ( .B1(n5459), .B2(n5456), .A(n5577), .ZN(n5465) );
  NAND2_X1 U6152 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5462), .ZN(n7737) );
  OAI21_X1 U6153 ( .B1(n5458), .B2(n5457), .A(n7737), .ZN(n5460) );
  AOI22_X1 U6154 ( .A1(n5465), .A2(n5460), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5462), .ZN(n7748) );
  OAI22_X1 U6155 ( .A1(n7740), .A2(n5610), .B1(n5900), .B2(n7737), .ZN(n5468)
         );
  INV_X1 U6156 ( .A(n5460), .ZN(n5464) );
  OAI21_X1 U6157 ( .B1(n5575), .B2(n5462), .A(n5461), .ZN(n5463) );
  AOI21_X1 U6158 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n7604) );
  INV_X1 U6159 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5466) );
  NOR2_X1 U6160 ( .A1(n7604), .A2(n5466), .ZN(n5467) );
  AOI211_X1 U6161 ( .C1(n7742), .C2(n5607), .A(n5468), .B(n5467), .ZN(n5469)
         );
  OAI21_X1 U6162 ( .B1(n7748), .B2(n5901), .A(n5469), .ZN(U3031) );
  OAI22_X1 U6163 ( .A1(n7740), .A2(n5601), .B1(n5887), .B2(n7737), .ZN(n5472)
         );
  INV_X1 U6164 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5470) );
  NOR2_X1 U6165 ( .A1(n7604), .A2(n5470), .ZN(n5471) );
  AOI211_X1 U6166 ( .C1(n7742), .C2(n5598), .A(n5472), .B(n5471), .ZN(n5473)
         );
  OAI21_X1 U6167 ( .B1(n7748), .B2(n5888), .A(n5473), .ZN(U3033) );
  OAI22_X1 U6168 ( .A1(n5742), .A2(n7679), .B1(n5620), .B2(n7674), .ZN(n5474)
         );
  AOI21_X1 U6169 ( .B1(n7692), .B2(n5911), .A(n5474), .ZN(n5476) );
  NAND2_X1 U6170 ( .A1(n5746), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5475) );
  OAI211_X1 U6171 ( .C1(n5749), .C2(n7697), .A(n5476), .B(n5475), .ZN(U3082)
         );
  NOR2_X1 U6172 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  OR2_X1 U6173 ( .A1(n5480), .A2(n5479), .ZN(n7312) );
  INV_X1 U6174 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5481) );
  OAI222_X1 U6175 ( .A1(n7312), .A2(n6359), .B1(n5481), .B2(n6352), .C1(n5763), 
        .C2(n6355), .ZN(U2855) );
  NOR2_X1 U6176 ( .A1(n6114), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5482)
         );
  OR2_X1 U6177 ( .A1(n5483), .A2(n5482), .ZN(n7341) );
  OAI222_X1 U6178 ( .A1(n7341), .A2(n6359), .B1(n6352), .B2(n5857), .C1(n5863), 
        .C2(n6355), .ZN(U2859) );
  INV_X1 U6179 ( .A(DATAI_5_), .ZN(n5485) );
  INV_X1 U6180 ( .A(EAX_REG_5__SCAN_IN), .ZN(n7181) );
  OAI222_X1 U6181 ( .A1(n5485), .A2(n6394), .B1(n6391), .B2(n7181), .C1(n7570), 
        .C2(n5484), .ZN(U2886) );
  OAI21_X1 U6182 ( .B1(n7731), .B2(n7742), .A(n5577), .ZN(n5486) );
  OAI21_X1 U6183 ( .B1(n5493), .B2(n5854), .A(n5486), .ZN(n5488) );
  NOR2_X1 U6184 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5487), .ZN(n5797)
         );
  AOI21_X1 U6185 ( .B1(n5488), .B2(n7534), .A(n5797), .ZN(n5490) );
  OR2_X1 U6186 ( .A1(n5652), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5547)
         );
  NAND2_X1 U6187 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5547), .ZN(n5545) );
  INV_X1 U6188 ( .A(n5545), .ZN(n5489) );
  NOR3_X1 U6189 ( .A1(n5490), .A2(n5867), .A3(n5489), .ZN(n5764) );
  INV_X1 U6190 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5497) );
  INV_X1 U6191 ( .A(n5547), .ZN(n5491) );
  NAND2_X1 U6192 ( .A1(n5874), .A2(n5491), .ZN(n5492) );
  OAI21_X1 U6193 ( .B1(n5650), .B2(n5493), .A(n5492), .ZN(n5796) );
  AOI22_X1 U6194 ( .A1(n7594), .A2(n5797), .B1(n5498), .B2(n5796), .ZN(n5494)
         );
  OAI21_X1 U6195 ( .B1(n5793), .B2(n7597), .A(n5494), .ZN(n5495) );
  AOI21_X1 U6196 ( .B1(n7605), .B2(n7742), .A(n5495), .ZN(n5496) );
  OAI21_X1 U6197 ( .B1(n5764), .B2(n5497), .A(n5496), .ZN(U3036) );
  AOI22_X1 U6198 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5532), .B1(n5498), 
        .B2(n5531), .ZN(n5499) );
  OAI21_X1 U6199 ( .B1(n7601), .B2(n5534), .A(n5499), .ZN(n5500) );
  AOI21_X1 U6200 ( .B1(n7605), .B2(n5822), .A(n5500), .ZN(n5501) );
  OAI21_X1 U6201 ( .B1(n7597), .B2(n5537), .A(n5501), .ZN(U3124) );
  AOI22_X1 U6202 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5532), .B1(n7144), 
        .B2(n5531), .ZN(n5502) );
  OAI21_X1 U6203 ( .B1(n7679), .B2(n5534), .A(n5502), .ZN(n5503) );
  AOI21_X1 U6204 ( .B1(n7693), .B2(n5822), .A(n5503), .ZN(n5504) );
  OAI21_X1 U6205 ( .B1(n7680), .B2(n5537), .A(n5504), .ZN(U3130) );
  AOI22_X1 U6206 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5532), .B1(n5785), 
        .B2(n5531), .ZN(n5505) );
  OAI21_X1 U6207 ( .B1(n7646), .B2(n5534), .A(n5505), .ZN(n5506) );
  AOI21_X1 U6208 ( .B1(n7649), .B2(n5822), .A(n5506), .ZN(n5507) );
  OAI21_X1 U6209 ( .B1(n5886), .B2(n5537), .A(n5507), .ZN(U3126) );
  XOR2_X1 U6210 ( .A(n5508), .B(n5509), .Z(n5570) );
  NOR2_X1 U6211 ( .A1(n6683), .A2(n5631), .ZN(n5510) );
  NOR2_X1 U6212 ( .A1(n5511), .A2(n5510), .ZN(n7310) );
  INV_X1 U6213 ( .A(n5631), .ZN(n5939) );
  INV_X1 U6214 ( .A(n6741), .ZN(n5512) );
  NAND3_X1 U6215 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5512), .ZN(n5633) );
  OAI21_X1 U6216 ( .B1(n5939), .B2(n6683), .A(n5633), .ZN(n7317) );
  NAND2_X1 U6217 ( .A1(n7317), .A2(n5515), .ZN(n5514) );
  AND2_X1 U6218 ( .A1(n7330), .A2(REIP_REG_3__SCAN_IN), .ZN(n5572) );
  AOI21_X1 U6219 ( .B1(n7332), .B2(n5846), .A(n5572), .ZN(n5513) );
  OAI211_X1 U6220 ( .C1(n7310), .C2(n5515), .A(n5514), .B(n5513), .ZN(n5516)
         );
  AOI21_X1 U6221 ( .B1(n5570), .B2(n7344), .A(n5516), .ZN(n5517) );
  INV_X1 U6222 ( .A(n5517), .ZN(U3015) );
  AOI22_X1 U6223 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5532), .B1(n5773), 
        .B2(n5531), .ZN(n5518) );
  OAI21_X1 U6224 ( .B1(n7667), .B2(n5534), .A(n5518), .ZN(n5519) );
  AOI21_X1 U6225 ( .B1(n7670), .B2(n5822), .A(n5519), .ZN(n5520) );
  OAI21_X1 U6226 ( .B1(n7653), .B2(n5537), .A(n5520), .ZN(U3128) );
  AOI21_X1 U6227 ( .B1(n5522), .B2(n5332), .A(n3816), .ZN(n7382) );
  INV_X1 U6228 ( .A(n7382), .ZN(n5695) );
  MUX2_X1 U6229 ( .A(n6058), .B(n5523), .S(EBX_REG_6__SCAN_IN), .Z(n5524) );
  OAI21_X1 U6230 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6114), .A(n5524), 
        .ZN(n5526) );
  AOI21_X1 U6231 ( .B1(n5526), .B2(n5525), .A(n3757), .ZN(n7377) );
  AOI22_X1 U6232 ( .A1(n7377), .A2(n7284), .B1(EBX_REG_6__SCAN_IN), .B2(n6353), 
        .ZN(n5527) );
  OAI21_X1 U6233 ( .B1(n5695), .B2(n6355), .A(n5527), .ZN(U2853) );
  AOI22_X1 U6234 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5532), .B1(n5790), 
        .B2(n5531), .ZN(n5528) );
  OAI21_X1 U6235 ( .B1(n7625), .B2(n5534), .A(n5528), .ZN(n5529) );
  AOI21_X1 U6236 ( .B1(n7622), .B2(n5822), .A(n5529), .ZN(n5530) );
  OAI21_X1 U6237 ( .B1(n7620), .B2(n5537), .A(n5530), .ZN(U3125) );
  AOI22_X1 U6238 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5532), .B1(n5768), 
        .B2(n5531), .ZN(n5533) );
  OAI21_X1 U6239 ( .B1(n7738), .B2(n5534), .A(n5533), .ZN(n5535) );
  AOI21_X1 U6240 ( .B1(n7730), .B2(n5822), .A(n5535), .ZN(n5536) );
  OAI21_X1 U6241 ( .B1(n7707), .B2(n5537), .A(n5536), .ZN(U3131) );
  NOR2_X1 U6242 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5538), .ZN(n5592)
         );
  INV_X1 U6243 ( .A(n5539), .ZN(n5541) );
  AOI21_X1 U6244 ( .B1(n5620), .B2(n5627), .A(n7303), .ZN(n5540) );
  AOI21_X1 U6245 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5544) );
  NOR2_X1 U6246 ( .A1(n5544), .A2(n5543), .ZN(n5546) );
  NOR2_X1 U6247 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  AOI21_X1 U6248 ( .B1(n5866), .B2(n5550), .A(n5549), .ZN(n5621) );
  INV_X1 U6249 ( .A(n5621), .ZN(n5551) );
  AOI22_X1 U6250 ( .A1(n5551), .A2(n7144), .B1(n7691), .B2(n5592), .ZN(n5553)
         );
  NAND2_X1 U6251 ( .A1(n7723), .A2(n7693), .ZN(n5552) );
  OAI211_X1 U6252 ( .C1(n5620), .C2(n7680), .A(n5553), .B(n5552), .ZN(n5554)
         );
  AOI21_X1 U6253 ( .B1(n5619), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n5554), 
        .ZN(n5555) );
  INV_X1 U6254 ( .A(n5555), .ZN(U3074) );
  INV_X1 U6255 ( .A(n5556), .ZN(n5559) );
  NAND2_X1 U6256 ( .A1(n5521), .A2(n5557), .ZN(n5558) );
  NAND2_X1 U6257 ( .A1(n5559), .A2(n5558), .ZN(n7394) );
  INV_X1 U6258 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6259 ( .A1(n6052), .A2(n5561), .ZN(n5565) );
  NAND2_X1 U6260 ( .A1(n6054), .A2(n5560), .ZN(n5563) );
  NAND2_X1 U6261 ( .A1(n6018), .A2(n5561), .ZN(n5562) );
  NAND3_X1 U6262 ( .A1(n5563), .A2(n6049), .A3(n5562), .ZN(n5564) );
  NAND2_X1 U6263 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U6264 ( .A1(n5700), .A2(n5568), .ZN(n5941) );
  INV_X1 U6265 ( .A(n5941), .ZN(n7391) );
  AOI22_X1 U6266 ( .A1(n7284), .A2(n7391), .B1(n6353), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5569) );
  OAI21_X1 U6267 ( .B1(n7394), .B2(n6355), .A(n5569), .ZN(U2852) );
  INV_X1 U6268 ( .A(n7482), .ZN(n7290) );
  NAND2_X1 U6269 ( .A1(n5570), .A2(n7290), .ZN(n5574) );
  NOR2_X1 U6270 ( .A1(n7294), .A2(n5844), .ZN(n5571) );
  AOI211_X1 U6271 ( .C1(n7289), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5572), 
        .B(n5571), .ZN(n5573) );
  OAI211_X1 U6272 ( .C1(n6509), .C2(n5856), .A(n5574), .B(n5573), .ZN(U2983)
         );
  INV_X1 U6273 ( .A(n7716), .ZN(n5576) );
  NAND3_X1 U6274 ( .A1(n5576), .A2(n5575), .A3(n7708), .ZN(n5578) );
  NAND2_X1 U6275 ( .A1(n5578), .A2(n5577), .ZN(n5580) );
  INV_X1 U6276 ( .A(n5580), .ZN(n5585) );
  NOR2_X1 U6277 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5581), .ZN(n7657)
         );
  INV_X1 U6278 ( .A(n7657), .ZN(n7706) );
  AOI211_X1 U6279 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7706), .A(n5582), .B(
        n5867), .ZN(n5583) );
  AOI22_X1 U6280 ( .A1(n7716), .A2(n5890), .B1(n5674), .B2(n7657), .ZN(n5586)
         );
  OAI21_X1 U6281 ( .B1(n5893), .B2(n7708), .A(n5586), .ZN(n5587) );
  AOI21_X1 U6282 ( .B1(n7710), .B2(INSTQUEUE_REG_10__5__SCAN_IN), .A(n5587), 
        .ZN(n5588) );
  OAI21_X1 U6283 ( .B1(n7713), .B2(n5888), .A(n5588), .ZN(U3105) );
  AOI22_X1 U6284 ( .A1(n7716), .A2(n5903), .B1(n5688), .B2(n7657), .ZN(n5589)
         );
  OAI21_X1 U6285 ( .B1(n5906), .B2(n7708), .A(n5589), .ZN(n5590) );
  AOI21_X1 U6286 ( .B1(n7710), .B2(INSTQUEUE_REG_10__3__SCAN_IN), .A(n5590), 
        .ZN(n5591) );
  OAI21_X1 U6287 ( .B1(n7713), .B2(n5901), .A(n5591), .ZN(U3103) );
  NAND2_X1 U6288 ( .A1(n5619), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5596) );
  NOR2_X1 U6289 ( .A1(n5620), .A2(n5886), .ZN(n5594) );
  INV_X1 U6290 ( .A(n5592), .ZN(n5622) );
  OAI22_X1 U6291 ( .A1(n7646), .A2(n5622), .B1(n5621), .B2(n7652), .ZN(n5593)
         );
  NOR2_X1 U6292 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  OAI211_X1 U6293 ( .C1(n7632), .C2(n5627), .A(n5596), .B(n5595), .ZN(U3070)
         );
  NAND2_X1 U6294 ( .A1(n5619), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5600) );
  OAI22_X1 U6295 ( .A1(n5888), .A2(n5621), .B1(n5887), .B2(n5622), .ZN(n5597)
         );
  AOI21_X1 U6296 ( .B1(n5598), .B2(n5745), .A(n5597), .ZN(n5599) );
  OAI211_X1 U6297 ( .C1(n5627), .C2(n5601), .A(n5600), .B(n5599), .ZN(U3073)
         );
  NAND2_X1 U6298 ( .A1(n5619), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5605) );
  NOR2_X1 U6299 ( .A1(n5620), .A2(n7653), .ZN(n5603) );
  OAI22_X1 U6300 ( .A1(n7667), .A2(n5622), .B1(n5621), .B2(n7673), .ZN(n5602)
         );
  NOR2_X1 U6301 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  OAI211_X1 U6302 ( .C1(n5627), .C2(n5778), .A(n5605), .B(n5604), .ZN(U3072)
         );
  NAND2_X1 U6303 ( .A1(n5619), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5609) );
  OAI22_X1 U6304 ( .A1(n5901), .A2(n5621), .B1(n5900), .B2(n5622), .ZN(n5606)
         );
  AOI21_X1 U6305 ( .B1(n5607), .B2(n5745), .A(n5606), .ZN(n5608) );
  OAI211_X1 U6306 ( .C1(n5627), .C2(n5610), .A(n5609), .B(n5608), .ZN(U3071)
         );
  NAND2_X1 U6307 ( .A1(n5619), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5614) );
  NOR2_X1 U6308 ( .A1(n5620), .A2(n7707), .ZN(n5612) );
  OAI22_X1 U6309 ( .A1(n7738), .A2(n5622), .B1(n5621), .B2(n7747), .ZN(n5611)
         );
  NOR2_X1 U6310 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  OAI211_X1 U6311 ( .C1(n5627), .C2(n7739), .A(n5614), .B(n5613), .ZN(U3075)
         );
  NAND2_X1 U6312 ( .A1(n5619), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5618) );
  NOR2_X1 U6313 ( .A1(n5620), .A2(n7597), .ZN(n5616) );
  OAI22_X1 U6314 ( .A1(n7601), .A2(n5622), .B1(n5621), .B2(n7608), .ZN(n5615)
         );
  NOR2_X1 U6315 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  OAI211_X1 U6316 ( .C1(n5627), .C2(n5825), .A(n5618), .B(n5617), .ZN(U3068)
         );
  NAND2_X1 U6317 ( .A1(n5619), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5626) );
  NOR2_X1 U6318 ( .A1(n5620), .A2(n7620), .ZN(n5624) );
  OAI22_X1 U6319 ( .A1(n7625), .A2(n5622), .B1(n5621), .B2(n7631), .ZN(n5623)
         );
  NOR2_X1 U6320 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  OAI211_X1 U6321 ( .C1(n5627), .C2(n7626), .A(n5626), .B(n5625), .ZN(U3069)
         );
  OAI222_X1 U6322 ( .A1(n5628), .A2(n6394), .B1(n6391), .B2(n5028), .C1(n7570), 
        .C2(n7394), .ZN(U2884) );
  XNOR2_X1 U6323 ( .A(n5630), .B(n5629), .ZN(n5641) );
  NAND2_X1 U6324 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7316) );
  NOR2_X1 U6325 ( .A1(n5337), .A2(n7316), .ZN(n5932) );
  OAI21_X1 U6326 ( .B1(n5932), .B2(n6710), .A(n7310), .ZN(n5809) );
  NAND2_X1 U6327 ( .A1(n6731), .A2(n5631), .ZN(n5632) );
  OAI21_X1 U6328 ( .B1(n7316), .B2(n5632), .A(n5337), .ZN(n5636) );
  INV_X1 U6329 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7366) );
  OAI22_X1 U6330 ( .A1(n7342), .A2(n7362), .B1(n7366), .B2(n6759), .ZN(n5635)
         );
  NOR3_X1 U6331 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n7316), .A3(n5633), 
        .ZN(n5634) );
  AOI211_X1 U6332 ( .C1(n5809), .C2(n5636), .A(n5635), .B(n5634), .ZN(n5637)
         );
  OAI21_X1 U6333 ( .B1(n5641), .B2(n6765), .A(n5637), .ZN(U3013) );
  AOI22_X1 U6334 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6546), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5638) );
  OAI21_X1 U6335 ( .B1(n7294), .B2(n7374), .A(n5638), .ZN(n5639) );
  AOI21_X1 U6336 ( .B1(n7371), .B2(n6534), .A(n5639), .ZN(n5640) );
  OAI21_X1 U6337 ( .B1(n5641), .B2(n7482), .A(n5640), .ZN(U2981) );
  XOR2_X1 U6338 ( .A(n5642), .B(n5643), .Z(n7315) );
  NAND2_X1 U6339 ( .A1(n7315), .A2(n7290), .ZN(n5647) );
  INV_X1 U6340 ( .A(n5644), .ZN(n5757) );
  INV_X1 U6341 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6342 ( .A1(n7330), .A2(REIP_REG_4__SCAN_IN), .ZN(n7311) );
  OAI21_X1 U6343 ( .B1(n6516), .B2(n5755), .A(n7311), .ZN(n5645) );
  AOI21_X1 U6344 ( .B1(n5757), .B2(n6513), .A(n5645), .ZN(n5646) );
  OAI211_X1 U6345 ( .C1(n6509), .C2(n5763), .A(n5647), .B(n5646), .ZN(U2982)
         );
  INV_X1 U6346 ( .A(n5648), .ZN(n5649) );
  AOI211_X1 U6347 ( .C1(n5650), .C2(n5649), .A(n5822), .B(n7676), .ZN(n5656)
         );
  NOR2_X1 U6348 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5651), .ZN(n5817)
         );
  NAND2_X1 U6349 ( .A1(n5653), .A2(n5652), .ZN(n5658) );
  NAND2_X1 U6350 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5658), .ZN(n5870) );
  OAI211_X1 U6351 ( .C1(n5817), .C2(n7534), .A(n5654), .B(n5870), .ZN(n5655)
         );
  NOR2_X1 U6352 ( .A1(n5656), .A2(n5655), .ZN(n5815) );
  INV_X1 U6353 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6354 ( .A1(n5876), .A2(n5657), .ZN(n5661) );
  INV_X1 U6355 ( .A(n5658), .ZN(n5873) );
  NAND2_X1 U6356 ( .A1(n5873), .A2(n5659), .ZN(n5660) );
  NAND2_X1 U6357 ( .A1(n5661), .A2(n5660), .ZN(n5818) );
  AOI22_X1 U6358 ( .A1(n7729), .A2(n5817), .B1(n5768), .B2(n5818), .ZN(n5662)
         );
  OAI21_X1 U6359 ( .B1(n5691), .B2(n7707), .A(n5662), .ZN(n5663) );
  AOI21_X1 U6360 ( .B1(n7730), .B2(n7676), .A(n5663), .ZN(n5664) );
  OAI21_X1 U6361 ( .B1(n5815), .B2(n5665), .A(n5664), .ZN(U3123) );
  INV_X1 U6362 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5669) );
  AOI22_X1 U6363 ( .A1(n7691), .A2(n5817), .B1(n7144), .B2(n5818), .ZN(n5666)
         );
  OAI21_X1 U6364 ( .B1(n5691), .B2(n7680), .A(n5666), .ZN(n5667) );
  AOI21_X1 U6365 ( .B1(n7693), .B2(n7676), .A(n5667), .ZN(n5668) );
  OAI21_X1 U6366 ( .B1(n5815), .B2(n5669), .A(n5668), .ZN(U3122) );
  INV_X1 U6367 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5673) );
  AOI22_X1 U6368 ( .A1(n7642), .A2(n5817), .B1(n5785), .B2(n5818), .ZN(n5670)
         );
  OAI21_X1 U6369 ( .B1(n5691), .B2(n5886), .A(n5670), .ZN(n5671) );
  AOI21_X1 U6370 ( .B1(n7649), .B2(n7676), .A(n5671), .ZN(n5672) );
  OAI21_X1 U6371 ( .B1(n5815), .B2(n5673), .A(n5672), .ZN(U3118) );
  INV_X1 U6372 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5679) );
  AOI22_X1 U6373 ( .A1(n5675), .A2(n5818), .B1(n5674), .B2(n5817), .ZN(n5676)
         );
  OAI21_X1 U6374 ( .B1(n5893), .B2(n5691), .A(n5676), .ZN(n5677) );
  AOI21_X1 U6375 ( .B1(n5890), .B2(n7676), .A(n5677), .ZN(n5678) );
  OAI21_X1 U6376 ( .B1(n5815), .B2(n5679), .A(n5678), .ZN(U3121) );
  INV_X1 U6377 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5683) );
  AOI22_X1 U6378 ( .A1(n7664), .A2(n5817), .B1(n5773), .B2(n5818), .ZN(n5680)
         );
  OAI21_X1 U6379 ( .B1(n5691), .B2(n7653), .A(n5680), .ZN(n5681) );
  AOI21_X1 U6380 ( .B1(n7670), .B2(n7676), .A(n5681), .ZN(n5682) );
  OAI21_X1 U6381 ( .B1(n5815), .B2(n5683), .A(n5682), .ZN(U3120) );
  INV_X1 U6382 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5687) );
  AOI22_X1 U6383 ( .A1(n7616), .A2(n5817), .B1(n5790), .B2(n5818), .ZN(n5684)
         );
  OAI21_X1 U6384 ( .B1(n5691), .B2(n7620), .A(n5684), .ZN(n5685) );
  AOI21_X1 U6385 ( .B1(n7622), .B2(n7676), .A(n5685), .ZN(n5686) );
  OAI21_X1 U6386 ( .B1(n5815), .B2(n5687), .A(n5686), .ZN(U3117) );
  INV_X1 U6387 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5694) );
  AOI22_X1 U6388 ( .A1(n5689), .A2(n5818), .B1(n5688), .B2(n5817), .ZN(n5690)
         );
  OAI21_X1 U6389 ( .B1(n5906), .B2(n5691), .A(n5690), .ZN(n5692) );
  AOI21_X1 U6390 ( .B1(n5903), .B2(n7676), .A(n5692), .ZN(n5693) );
  OAI21_X1 U6391 ( .B1(n5815), .B2(n5694), .A(n5693), .ZN(U3119) );
  OAI222_X1 U6392 ( .A1(n6394), .A2(n5696), .B1(n6391), .B2(n4864), .C1(n7570), 
        .C2(n5695), .ZN(U2885) );
  OAI21_X1 U6393 ( .B1(n5556), .B2(n5698), .A(n5697), .ZN(n5957) );
  MUX2_X1 U6394 ( .A(n6058), .B(n5523), .S(EBX_REG_8__SCAN_IN), .Z(n5699) );
  OAI21_X1 U6395 ( .B1(n6114), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5699), 
        .ZN(n5701) );
  AOI21_X1 U6396 ( .B1(n5701), .B2(n5700), .A(n5832), .ZN(n7321) );
  AOI22_X1 U6397 ( .A1(n7321), .A2(n7284), .B1(EBX_REG_8__SCAN_IN), .B2(n6353), 
        .ZN(n5702) );
  OAI21_X1 U6398 ( .B1(n5957), .B2(n6355), .A(n5702), .ZN(U2851) );
  OR2_X1 U6399 ( .A1(n5704), .A2(n5703), .ZN(n7523) );
  NOR3_X1 U6400 ( .A1(n3966), .A2(n7534), .A3(n7542), .ZN(n7539) );
  INV_X1 U6401 ( .A(n7539), .ZN(n5705) );
  NAND2_X1 U6402 ( .A1(n7523), .A2(n5705), .ZN(n5706) );
  NOR2_X1 U6403 ( .A1(n7330), .A2(n5706), .ZN(n5707) );
  NOR2_X1 U6404 ( .A1(n6402), .A2(n5711), .ZN(n5712) );
  INV_X1 U6405 ( .A(n5714), .ZN(n5954) );
  NAND2_X1 U6406 ( .A1(n7516), .A2(n7303), .ZN(n5723) );
  OR2_X1 U6407 ( .A1(n6105), .A2(n5723), .ZN(n7520) );
  NAND2_X1 U6408 ( .A1(n7304), .A2(n7520), .ZN(n6123) );
  INV_X1 U6409 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6300) );
  NAND3_X1 U6410 ( .A1(n5721), .A2(n6300), .A3(n5723), .ZN(n5715) );
  AND2_X1 U6411 ( .A1(n6123), .A2(n5715), .ZN(n5716) );
  NAND2_X1 U6412 ( .A1(n5723), .A2(EBX_REG_31__SCAN_IN), .ZN(n5717) );
  AOI22_X1 U6413 ( .A1(EBX_REG_8__SCAN_IN), .A2(n7471), .B1(n7473), .B2(n7321), 
        .ZN(n5719) );
  INV_X1 U6414 ( .A(n7426), .ZN(n7352) );
  NOR2_X1 U6415 ( .A1(n5718), .A2(n7352), .ZN(n7423) );
  INV_X1 U6416 ( .A(n7423), .ZN(n7448) );
  OAI211_X1 U6417 ( .C1(n7450), .C2(n5952), .A(n5719), .B(n7448), .ZN(n5731)
         );
  NAND2_X1 U6418 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n5726) );
  AND2_X1 U6419 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NOR2_X1 U6420 ( .A1(n6018), .A2(n5722), .ZN(n5724) );
  NAND3_X1 U6421 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n5754) );
  INV_X1 U6422 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7203) );
  NOR2_X1 U6423 ( .A1(n5754), .A2(n7203), .ZN(n7365) );
  AND2_X1 U6424 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7365), .ZN(n5725) );
  NAND2_X1 U6425 ( .A1(n7470), .A2(n5725), .ZN(n7388) );
  NOR2_X1 U6426 ( .A1(n5726), .A2(n7388), .ZN(n5729) );
  INV_X1 U6427 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7209) );
  NOR2_X1 U6428 ( .A1(n5726), .A2(n7209), .ZN(n6063) );
  INV_X1 U6429 ( .A(n6063), .ZN(n5836) );
  NAND2_X1 U6430 ( .A1(n7365), .A2(REIP_REG_5__SCAN_IN), .ZN(n6064) );
  INV_X1 U6431 ( .A(n6064), .ZN(n5727) );
  NAND2_X1 U6432 ( .A1(n7426), .A2(n5727), .ZN(n7376) );
  NAND2_X1 U6433 ( .A1(n7446), .A2(n7426), .ZN(n7375) );
  OAI21_X1 U6434 ( .B1(n5836), .B2(n7376), .A(n7375), .ZN(n6278) );
  INV_X1 U6435 ( .A(n6278), .ZN(n5728) );
  MUX2_X1 U6436 ( .A(n5729), .B(n5728), .S(REIP_REG_8__SCAN_IN), .Z(n5730) );
  AOI211_X1 U6437 ( .C1(n7475), .C2(n5954), .A(n5731), .B(n5730), .ZN(n5732)
         );
  OAI21_X1 U6438 ( .B1(n7437), .B2(n5957), .A(n5732), .ZN(U2819) );
  INV_X1 U6439 ( .A(n5911), .ZN(n5743) );
  OAI22_X1 U6440 ( .A1(n5743), .A2(n7707), .B1(n5742), .B2(n7738), .ZN(n5733)
         );
  AOI21_X1 U6441 ( .B1(n7730), .B2(n5745), .A(n5733), .ZN(n5735) );
  NAND2_X1 U6442 ( .A1(n5746), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U6443 ( .C1(n5749), .C2(n7747), .A(n5735), .B(n5734), .ZN(U3083)
         );
  OAI22_X1 U6444 ( .A1(n5743), .A2(n7620), .B1(n5742), .B2(n7625), .ZN(n5736)
         );
  AOI21_X1 U6445 ( .B1(n7622), .B2(n5745), .A(n5736), .ZN(n5738) );
  NAND2_X1 U6446 ( .A1(n5746), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U6447 ( .C1(n5749), .C2(n7631), .A(n5738), .B(n5737), .ZN(U3077)
         );
  OAI22_X1 U6448 ( .A1(n5743), .A2(n7653), .B1(n5742), .B2(n7667), .ZN(n5739)
         );
  AOI21_X1 U6449 ( .B1(n7670), .B2(n5745), .A(n5739), .ZN(n5741) );
  NAND2_X1 U6450 ( .A1(n5746), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5740) );
  OAI211_X1 U6451 ( .C1(n5749), .C2(n7673), .A(n5741), .B(n5740), .ZN(U3080)
         );
  OAI22_X1 U6452 ( .A1(n5743), .A2(n7597), .B1(n5742), .B2(n7601), .ZN(n5744)
         );
  AOI21_X1 U6453 ( .B1(n7605), .B2(n5745), .A(n5744), .ZN(n5748) );
  NAND2_X1 U6454 ( .A1(n5746), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n5747) );
  OAI211_X1 U6455 ( .C1(n5749), .C2(n7608), .A(n5748), .B(n5747), .ZN(U3076)
         );
  INV_X1 U6456 ( .A(n6103), .ZN(n5750) );
  NOR2_X1 U6457 ( .A1(n6124), .A2(n5750), .ZN(n5751) );
  OR2_X1 U6458 ( .A1(n5751), .A2(n7477), .ZN(n7370) );
  NOR2_X1 U6459 ( .A1(n6124), .A2(n5752), .ZN(n7358) );
  OR3_X1 U6460 ( .A1(n7446), .A2(REIP_REG_4__SCAN_IN), .A3(n5754), .ZN(n5760)
         );
  INV_X1 U6461 ( .A(n7312), .ZN(n5753) );
  AOI22_X1 U6462 ( .A1(n7471), .A2(EBX_REG_4__SCAN_IN), .B1(n7473), .B2(n5753), 
        .ZN(n5759) );
  OAI21_X1 U6463 ( .B1(n7352), .B2(n5754), .A(n7375), .ZN(n5850) );
  OAI22_X1 U6464 ( .A1(n5755), .A2(n7450), .B1(n7203), .B2(n5850), .ZN(n5756)
         );
  AOI211_X1 U6465 ( .C1(n7475), .C2(n5757), .A(n7423), .B(n5756), .ZN(n5758)
         );
  NAND3_X1 U6466 ( .A1(n5760), .A2(n5759), .A3(n5758), .ZN(n5761) );
  AOI21_X1 U6467 ( .B1(n7488), .B2(n7358), .A(n5761), .ZN(n5762) );
  OAI21_X1 U6468 ( .B1(n5763), .B2(n7354), .A(n5762), .ZN(U2823) );
  INV_X1 U6469 ( .A(n5764), .ZN(n5802) );
  NAND2_X1 U6470 ( .A1(n5802), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5767) );
  INV_X1 U6471 ( .A(n5796), .ZN(n5780) );
  INV_X1 U6472 ( .A(n5797), .ZN(n5779) );
  OAI22_X1 U6473 ( .A1(n5888), .A2(n5780), .B1(n5887), .B2(n5779), .ZN(n5765)
         );
  AOI21_X1 U6474 ( .B1(n5890), .B2(n7742), .A(n5765), .ZN(n5766) );
  OAI211_X1 U6475 ( .C1(n5793), .C2(n5893), .A(n5767), .B(n5766), .ZN(U3041)
         );
  INV_X1 U6476 ( .A(n7742), .ZN(n5800) );
  NAND2_X1 U6477 ( .A1(n5802), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U6478 ( .A1(n5796), .A2(n5768), .ZN(n5769) );
  OAI21_X1 U6479 ( .B1(n7738), .B2(n5779), .A(n5769), .ZN(n5770) );
  AOI21_X1 U6480 ( .B1(n7731), .B2(n7743), .A(n5770), .ZN(n5771) );
  OAI211_X1 U6481 ( .C1(n5800), .C2(n7739), .A(n5772), .B(n5771), .ZN(U3043)
         );
  NAND2_X1 U6482 ( .A1(n5802), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U6483 ( .A1(n5796), .A2(n5773), .ZN(n5774) );
  OAI21_X1 U6484 ( .B1(n7667), .B2(n5779), .A(n5774), .ZN(n5775) );
  AOI21_X1 U6485 ( .B1(n7731), .B2(n7669), .A(n5775), .ZN(n5776) );
  OAI211_X1 U6486 ( .C1(n5800), .C2(n5778), .A(n5777), .B(n5776), .ZN(U3040)
         );
  NAND2_X1 U6487 ( .A1(n5802), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5783) );
  OAI22_X1 U6488 ( .A1(n5901), .A2(n5780), .B1(n5900), .B2(n5779), .ZN(n5781)
         );
  AOI21_X1 U6489 ( .B1(n5903), .B2(n7742), .A(n5781), .ZN(n5782) );
  OAI211_X1 U6490 ( .C1(n5793), .C2(n5906), .A(n5783), .B(n5782), .ZN(U3039)
         );
  INV_X1 U6491 ( .A(DATAI_8_), .ZN(n5784) );
  OAI222_X1 U6492 ( .A1(n5957), .A2(n7570), .B1(n6394), .B2(n5784), .C1(n6391), 
        .C2(n5045), .ZN(U2883) );
  AOI22_X1 U6493 ( .A1(n7642), .A2(n5797), .B1(n5785), .B2(n5796), .ZN(n5787)
         );
  NAND2_X1 U6494 ( .A1(n7742), .A2(n7649), .ZN(n5786) );
  OAI211_X1 U6495 ( .C1(n5793), .C2(n5886), .A(n5787), .B(n5786), .ZN(n5788)
         );
  AOI21_X1 U6496 ( .B1(n5802), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n5788), 
        .ZN(n5789) );
  INV_X1 U6497 ( .A(n5789), .ZN(U3038) );
  AOI22_X1 U6498 ( .A1(n7616), .A2(n5797), .B1(n5790), .B2(n5796), .ZN(n5792)
         );
  NAND2_X1 U6499 ( .A1(n7742), .A2(n7622), .ZN(n5791) );
  OAI211_X1 U6500 ( .C1(n5793), .C2(n7620), .A(n5792), .B(n5791), .ZN(n5794)
         );
  AOI21_X1 U6501 ( .B1(n5802), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n5794), 
        .ZN(n5795) );
  INV_X1 U6502 ( .A(n5795), .ZN(U3037) );
  AOI22_X1 U6503 ( .A1(n7691), .A2(n5797), .B1(n7144), .B2(n5796), .ZN(n5799)
         );
  NAND2_X1 U6504 ( .A1(n7731), .A2(n7692), .ZN(n5798) );
  OAI211_X1 U6505 ( .C1(n5800), .C2(n7674), .A(n5799), .B(n5798), .ZN(n5801)
         );
  AOI21_X1 U6506 ( .B1(n5802), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n5801), 
        .ZN(n5803) );
  INV_X1 U6507 ( .A(n5803), .ZN(U3042) );
  XNOR2_X1 U6508 ( .A(n3694), .B(n5804), .ZN(n5814) );
  INV_X1 U6509 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7387) );
  NOR2_X1 U6510 ( .A1(n6759), .A2(n7387), .ZN(n5811) );
  AOI21_X1 U6511 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5811), 
        .ZN(n5806) );
  OAI21_X1 U6512 ( .B1(n7294), .B2(n7384), .A(n5806), .ZN(n5807) );
  AOI21_X1 U6513 ( .B1(n7382), .B2(n6534), .A(n5807), .ZN(n5808) );
  OAI21_X1 U6514 ( .B1(n5814), .B2(n7482), .A(n5808), .ZN(U2980) );
  INV_X1 U6515 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5810) );
  OAI222_X1 U6516 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5932), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n7317), .C1(n5810), .C2(n5809), 
        .ZN(n5813) );
  AOI21_X1 U6517 ( .B1(n7377), .B2(n7332), .A(n5811), .ZN(n5812) );
  OAI211_X1 U6518 ( .C1(n5814), .C2(n6765), .A(n5813), .B(n5812), .ZN(U3012)
         );
  INV_X1 U6519 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U6520 ( .A1(n5816), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5824)
         );
  INV_X1 U6521 ( .A(n5817), .ZN(n5820) );
  INV_X1 U6522 ( .A(n5818), .ZN(n5819) );
  OAI22_X1 U6523 ( .A1(n7601), .A2(n5820), .B1(n5819), .B2(n7608), .ZN(n5821)
         );
  AOI21_X1 U6524 ( .B1(n7603), .B2(n5822), .A(n5821), .ZN(n5823) );
  OAI211_X1 U6525 ( .C1(n7699), .C2(n5825), .A(n5824), .B(n5823), .ZN(U3116)
         );
  AOI21_X1 U6526 ( .B1(n5827), .B2(n5697), .A(n5826), .ZN(n5972) );
  INV_X1 U6527 ( .A(n6355), .ZN(n7285) );
  NAND2_X1 U6528 ( .A1(n6054), .A2(n6551), .ZN(n5829) );
  INV_X1 U6529 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U6530 ( .A1(n6018), .A2(n5837), .ZN(n5828) );
  NAND3_X1 U6531 ( .A1(n5829), .A2(n6049), .A3(n5828), .ZN(n5830) );
  OAI21_X1 U6532 ( .B1(n6107), .B2(EBX_REG_9__SCAN_IN), .A(n5830), .ZN(n5831)
         );
  NOR2_X1 U6533 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  OR2_X1 U6534 ( .A1(n5920), .A2(n5833), .ZN(n5963) );
  OAI22_X1 U6535 ( .A1(n5963), .A2(n6359), .B1(n5837), .B2(n6352), .ZN(n5834)
         );
  AOI21_X1 U6536 ( .B1(n5972), .B2(n7285), .A(n5834), .ZN(n5835) );
  INV_X1 U6537 ( .A(n5835), .ZN(U2850) );
  INV_X1 U6538 ( .A(n5972), .ZN(n5843) );
  INV_X1 U6539 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7210) );
  OAI22_X1 U6540 ( .A1(n5837), .A2(n7443), .B1(n7467), .B2(n5963), .ZN(n5838)
         );
  AOI211_X1 U6541 ( .C1(n7472), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n7423), 
        .B(n5838), .ZN(n5839) );
  OAI221_X1 U6542 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6281), .C1(n7210), .C2(
        n6278), .A(n5839), .ZN(n5840) );
  AOI21_X1 U6543 ( .B1(n5968), .B2(n7475), .A(n5840), .ZN(n5841) );
  OAI21_X1 U6544 ( .B1(n5843), .B2(n7437), .A(n5841), .ZN(U2818) );
  INV_X1 U6545 ( .A(DATAI_9_), .ZN(n5842) );
  OAI222_X1 U6546 ( .A1(n5843), .A2(n7570), .B1(n6394), .B2(n5842), .C1(n6391), 
        .C2(n5018), .ZN(U2882) );
  INV_X1 U6547 ( .A(n5844), .ZN(n5845) );
  AOI22_X1 U6548 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7472), .B1(n7475), 
        .B2(n5845), .ZN(n5848) );
  NAND2_X1 U6549 ( .A1(n7473), .A2(n5846), .ZN(n5847) );
  OAI211_X1 U6550 ( .C1(n5849), .C2(n7443), .A(n5848), .B(n5847), .ZN(n5853)
         );
  INV_X1 U6551 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U6552 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6295) );
  OR2_X1 U6553 ( .A1(n7352), .A2(n6295), .ZN(n5851) );
  AOI21_X1 U6554 ( .B1(n7201), .B2(n5851), .A(n5850), .ZN(n5852) );
  AOI211_X1 U6555 ( .C1(n7358), .C2(n5854), .A(n5853), .B(n5852), .ZN(n5855)
         );
  OAI21_X1 U6556 ( .B1(n5856), .B2(n7354), .A(n5855), .ZN(U2824) );
  OAI22_X1 U6557 ( .A1(n5857), .A2(n7443), .B1(n7467), .B2(n7341), .ZN(n5860)
         );
  AOI21_X1 U6558 ( .B1(n7450), .B2(n7420), .A(n5858), .ZN(n5859) );
  AOI211_X1 U6559 ( .C1(n7358), .C2(n4310), .A(n5860), .B(n5859), .ZN(n5862)
         );
  NAND2_X1 U6560 ( .A1(n7375), .A2(REIP_REG_0__SCAN_IN), .ZN(n5861) );
  OAI211_X1 U6561 ( .C1(n7354), .C2(n5863), .A(n5862), .B(n5861), .ZN(U2827)
         );
  NOR2_X1 U6562 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5864), .ZN(n5872)
         );
  OAI21_X1 U6563 ( .B1(n7715), .B2(n5911), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5869) );
  OR2_X1 U6564 ( .A1(n5866), .A2(n5865), .ZN(n5868) );
  AOI21_X1 U6565 ( .B1(n5869), .B2(n5868), .A(n5867), .ZN(n5871) );
  NAND2_X1 U6566 ( .A1(n5907), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5879) );
  INV_X1 U6567 ( .A(n5872), .ZN(n5909) );
  AOI22_X1 U6568 ( .A1(n5876), .A2(n5875), .B1(n5874), .B2(n5873), .ZN(n5908)
         );
  OAI22_X1 U6569 ( .A1(n7679), .A2(n5909), .B1(n5908), .B2(n7697), .ZN(n5877)
         );
  AOI21_X1 U6570 ( .B1(n7693), .B2(n5911), .A(n5877), .ZN(n5878) );
  OAI211_X1 U6571 ( .C1(n5914), .C2(n7680), .A(n5879), .B(n5878), .ZN(U3090)
         );
  NAND2_X1 U6572 ( .A1(n5907), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5882) );
  OAI22_X1 U6573 ( .A1(n7625), .A2(n5909), .B1(n5908), .B2(n7631), .ZN(n5880)
         );
  AOI21_X1 U6574 ( .B1(n5911), .B2(n7622), .A(n5880), .ZN(n5881) );
  OAI211_X1 U6575 ( .C1(n5914), .C2(n7620), .A(n5882), .B(n5881), .ZN(U3085)
         );
  NAND2_X1 U6576 ( .A1(n5907), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5885) );
  OAI22_X1 U6577 ( .A1(n7646), .A2(n5909), .B1(n5908), .B2(n7652), .ZN(n5883)
         );
  AOI21_X1 U6578 ( .B1(n5911), .B2(n7649), .A(n5883), .ZN(n5884) );
  OAI211_X1 U6579 ( .C1(n5914), .C2(n5886), .A(n5885), .B(n5884), .ZN(U3086)
         );
  NAND2_X1 U6580 ( .A1(n5907), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5892) );
  OAI22_X1 U6581 ( .A1(n5888), .A2(n5908), .B1(n5909), .B2(n5887), .ZN(n5889)
         );
  AOI21_X1 U6582 ( .B1(n5911), .B2(n5890), .A(n5889), .ZN(n5891) );
  OAI211_X1 U6583 ( .C1(n5914), .C2(n5893), .A(n5892), .B(n5891), .ZN(U3089)
         );
  NAND2_X1 U6584 ( .A1(n5907), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5896) );
  OAI22_X1 U6585 ( .A1(n7667), .A2(n5909), .B1(n5908), .B2(n7673), .ZN(n5894)
         );
  AOI21_X1 U6586 ( .B1(n5911), .B2(n7670), .A(n5894), .ZN(n5895) );
  OAI211_X1 U6587 ( .C1(n5914), .C2(n7653), .A(n5896), .B(n5895), .ZN(U3088)
         );
  NAND2_X1 U6588 ( .A1(n5907), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5899) );
  OAI22_X1 U6589 ( .A1(n7601), .A2(n5909), .B1(n5908), .B2(n7608), .ZN(n5897)
         );
  AOI21_X1 U6590 ( .B1(n7605), .B2(n5911), .A(n5897), .ZN(n5898) );
  OAI211_X1 U6591 ( .C1(n7597), .C2(n5914), .A(n5899), .B(n5898), .ZN(U3084)
         );
  NAND2_X1 U6592 ( .A1(n5907), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5905) );
  OAI22_X1 U6593 ( .A1(n5901), .A2(n5908), .B1(n5909), .B2(n5900), .ZN(n5902)
         );
  AOI21_X1 U6594 ( .B1(n5911), .B2(n5903), .A(n5902), .ZN(n5904) );
  OAI211_X1 U6595 ( .C1(n5914), .C2(n5906), .A(n5905), .B(n5904), .ZN(U3087)
         );
  NAND2_X1 U6596 ( .A1(n5907), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5913) );
  OAI22_X1 U6597 ( .A1(n7738), .A2(n5909), .B1(n5908), .B2(n7747), .ZN(n5910)
         );
  AOI21_X1 U6598 ( .B1(n5911), .B2(n7730), .A(n5910), .ZN(n5912) );
  OAI211_X1 U6599 ( .C1(n5914), .C2(n7707), .A(n5913), .B(n5912), .ZN(U3091)
         );
  AND2_X1 U6600 ( .A1(n3819), .A2(n5916), .ZN(n5917) );
  NOR2_X1 U6601 ( .A1(n5915), .A2(n5917), .ZN(n5994) );
  INV_X1 U6602 ( .A(n5994), .ZN(n5931) );
  MUX2_X1 U6603 ( .A(n6058), .B(n5523), .S(EBX_REG_10__SCAN_IN), .Z(n5918) );
  OAI21_X1 U6604 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6114), .A(n5918), 
        .ZN(n5923) );
  INV_X1 U6605 ( .A(n5920), .ZN(n5922) );
  INV_X1 U6606 ( .A(n5923), .ZN(n5919) );
  INV_X1 U6607 ( .A(n5984), .ZN(n5921) );
  AOI21_X1 U6608 ( .B1(n5923), .B2(n5922), .A(n5921), .ZN(n6001) );
  AOI22_X1 U6609 ( .A1(n6001), .A2(n7284), .B1(n6353), .B2(EBX_REG_10__SCAN_IN), .ZN(n5924) );
  OAI21_X1 U6610 ( .B1(n5931), .B2(n6355), .A(n5924), .ZN(U2849) );
  AOI22_X1 U6611 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n7472), .B1(n7473), 
        .B2(n6001), .ZN(n5925) );
  OAI211_X1 U6612 ( .C1(n7420), .C2(n5992), .A(n5925), .B(n7448), .ZN(n5926)
         );
  AOI21_X1 U6613 ( .B1(n7471), .B2(EBX_REG_10__SCAN_IN), .A(n5926), .ZN(n5929)
         );
  OAI211_X1 U6614 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6281), .A(
        REIP_REG_10__SCAN_IN), .B(n6278), .ZN(n7406) );
  INV_X1 U6615 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U6616 ( .B1(n7210), .B2(n6281), .A(n7213), .ZN(n5927) );
  NAND2_X1 U6617 ( .A1(n7406), .A2(n5927), .ZN(n5928) );
  OAI211_X1 U6618 ( .C1(n5931), .C2(n7437), .A(n5929), .B(n5928), .ZN(U2817)
         );
  INV_X1 U6619 ( .A(DATAI_10_), .ZN(n5930) );
  OAI222_X1 U6620 ( .A1(n5931), .A2(n7570), .B1(n6394), .B2(n5930), .C1(n6391), 
        .C2(n5025), .ZN(U2881) );
  NAND2_X1 U6621 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5932), .ZN(n5938)
         );
  INV_X1 U6622 ( .A(n5938), .ZN(n5933) );
  NAND2_X1 U6623 ( .A1(n5933), .A2(n7317), .ZN(n7328) );
  XOR2_X1 U6624 ( .A(n5934), .B(n5935), .Z(n5945) );
  NAND2_X1 U6625 ( .A1(n5945), .A2(n7344), .ZN(n5944) );
  INV_X1 U6626 ( .A(n6563), .ZN(n6729) );
  NOR3_X1 U6627 ( .A1(n5937), .A2(n5936), .A3(n5938), .ZN(n6553) );
  NOR2_X1 U6628 ( .A1(n5939), .A2(n5938), .ZN(n6556) );
  OAI22_X1 U6629 ( .A1(n6727), .A2(n6553), .B1(n6556), .B2(n6683), .ZN(n5940)
         );
  NOR2_X1 U6630 ( .A1(n6729), .A2(n5940), .ZN(n7323) );
  INV_X1 U6631 ( .A(n7323), .ZN(n5964) );
  AND2_X1 U6632 ( .A1(n6546), .A2(REIP_REG_7__SCAN_IN), .ZN(n5947) );
  NOR2_X1 U6633 ( .A1(n5941), .A2(n7342), .ZN(n5942) );
  AOI211_X1 U6634 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n5964), .A(n5947), 
        .B(n5942), .ZN(n5943) );
  OAI211_X1 U6635 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n7328), .A(n5944), 
        .B(n5943), .ZN(U3011) );
  NAND2_X1 U6636 ( .A1(n5945), .A2(n7290), .ZN(n5949) );
  NOR2_X1 U6637 ( .A1(n7294), .A2(n7397), .ZN(n5946) );
  AOI211_X1 U6638 ( .C1(n7289), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5947), 
        .B(n5946), .ZN(n5948) );
  OAI211_X1 U6639 ( .C1(n6509), .C2(n7394), .A(n5949), .B(n5948), .ZN(U2979)
         );
  XOR2_X1 U6640 ( .A(n5951), .B(n5950), .Z(n7325) );
  NAND2_X1 U6641 ( .A1(n7325), .A2(n7290), .ZN(n5956) );
  OAI22_X1 U6642 ( .A1(n6516), .A2(n5952), .B1(n6759), .B2(n7209), .ZN(n5953)
         );
  AOI21_X1 U6643 ( .B1(n5954), .B2(n6513), .A(n5953), .ZN(n5955) );
  OAI211_X1 U6644 ( .C1(n6509), .C2(n5957), .A(n5956), .B(n5955), .ZN(U2978)
         );
  INV_X1 U6645 ( .A(DATAI_11_), .ZN(n5960) );
  NOR2_X1 U6646 ( .A1(n5915), .A2(n5958), .ZN(n5959) );
  OR2_X1 U6647 ( .A1(n5977), .A2(n5959), .ZN(n7402) );
  OAI222_X1 U6648 ( .A1(n6394), .A2(n5960), .B1(n6391), .B2(n5022), .C1(n7570), 
        .C2(n7402), .ZN(U2880) );
  XNOR2_X1 U6649 ( .A(n3690), .B(n5962), .ZN(n5974) );
  NAND2_X1 U6650 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7320) );
  NOR2_X1 U6651 ( .A1(n7320), .A2(n7328), .ZN(n5998) );
  OAI22_X1 U6652 ( .A1(n5963), .A2(n7342), .B1(n7210), .B2(n6759), .ZN(n5966)
         );
  AOI21_X1 U6653 ( .B1(n7320), .B2(n6687), .A(n5964), .ZN(n5996) );
  NOR2_X1 U6654 ( .A1(n5996), .A2(n6551), .ZN(n5965) );
  AOI211_X1 U6655 ( .C1(n5998), .C2(n6551), .A(n5966), .B(n5965), .ZN(n5967)
         );
  OAI21_X1 U6656 ( .B1(n5974), .B2(n6765), .A(n5967), .ZN(U3009) );
  INV_X1 U6657 ( .A(n5968), .ZN(n5970) );
  AOI22_X1 U6658 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6546), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5969) );
  OAI21_X1 U6659 ( .B1(n7294), .B2(n5970), .A(n5969), .ZN(n5971) );
  AOI21_X1 U6660 ( .B1(n5972), .B2(n6534), .A(n5971), .ZN(n5973) );
  OAI21_X1 U6661 ( .B1(n5974), .B2(n7482), .A(n5973), .ZN(U2977) );
  INV_X1 U6662 ( .A(DATAI_12_), .ZN(n5978) );
  OAI21_X1 U6663 ( .B1(n5977), .B2(n5976), .A(n5975), .ZN(n6539) );
  OAI222_X1 U6664 ( .A1(n6394), .A2(n5978), .B1(n6391), .B2(n5039), .C1(n7570), 
        .C2(n6539), .ZN(U2879) );
  INV_X1 U6665 ( .A(n7402), .ZN(n6549) );
  INV_X1 U6666 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U6667 ( .A1(n6052), .A2(n5986), .ZN(n5982) );
  NAND2_X1 U6668 ( .A1(n6054), .A2(n6752), .ZN(n5980) );
  NAND2_X1 U6669 ( .A1(n6018), .A2(n5986), .ZN(n5979) );
  NAND3_X1 U6670 ( .A1(n5980), .A2(n5523), .A3(n5979), .ZN(n5981) );
  NAND2_X1 U6671 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  NAND2_X1 U6672 ( .A1(n6749), .A2(n5985), .ZN(n7399) );
  OAI22_X1 U6673 ( .A1(n7399), .A2(n6359), .B1(n5986), .B2(n6352), .ZN(n5987)
         );
  AOI21_X1 U6674 ( .B1(n6549), .B2(n7285), .A(n5987), .ZN(n5988) );
  INV_X1 U6675 ( .A(n5988), .ZN(U2848) );
  XNOR2_X1 U6676 ( .A(n5990), .B(n5989), .ZN(n6004) );
  NOR2_X1 U6677 ( .A1(n6759), .A2(n7213), .ZN(n6000) );
  AOI21_X1 U6678 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6000), 
        .ZN(n5991) );
  OAI21_X1 U6679 ( .B1(n7294), .B2(n5992), .A(n5991), .ZN(n5993) );
  AOI21_X1 U6680 ( .B1(n5994), .B2(n6534), .A(n5993), .ZN(n5995) );
  OAI21_X1 U6681 ( .B1(n6004), .B2(n7482), .A(n5995), .ZN(U2976) );
  INV_X1 U6682 ( .A(n5996), .ZN(n5999) );
  INV_X1 U6683 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6552) );
  AOI22_X1 U6684 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6551), .B2(n6552), .ZN(n5997) );
  AOI22_X1 U6685 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5999), .B1(n5998), .B2(n5997), .ZN(n6003) );
  AOI21_X1 U6686 ( .B1(n6001), .B2(n7332), .A(n6000), .ZN(n6002) );
  OAI211_X1 U6687 ( .C1(n6004), .C2(n6765), .A(n6003), .B(n6002), .ZN(U3008)
         );
  NOR2_X2 U6688 ( .A1(n7583), .A2(n3672), .ZN(n7580) );
  AOI22_X1 U6689 ( .A1(n7580), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n7583), .ZN(n6008) );
  NAND2_X1 U6690 ( .A1(n7584), .A2(DATAI_14_), .ZN(n6007) );
  OAI211_X1 U6691 ( .C1(n6005), .C2(n7570), .A(n6008), .B(n6007), .ZN(U2861)
         );
  INV_X1 U6692 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6076) );
  OAI22_X1 U6693 ( .A1(n6114), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n6113), .ZN(n6108) );
  INV_X1 U6694 ( .A(n6108), .ZN(n6060) );
  NAND2_X1 U6695 ( .A1(n5523), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U6696 ( .C1(n6113), .C2(EBX_REG_12__SCAN_IN), .A(n6054), .B(n6009), 
        .ZN(n6010) );
  OAI21_X1 U6697 ( .B1(n6058), .B2(EBX_REG_12__SCAN_IN), .A(n6010), .ZN(n6750)
         );
  NAND2_X1 U6698 ( .A1(n6054), .A2(n6730), .ZN(n6012) );
  INV_X1 U6699 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U6700 ( .A1(n6018), .A2(n6358), .ZN(n6011) );
  NAND3_X1 U6701 ( .A1(n6012), .A2(n6049), .A3(n6011), .ZN(n6013) );
  OAI21_X1 U6702 ( .B1(n6107), .B2(EBX_REG_13__SCAN_IN), .A(n6013), .ZN(n6275)
         );
  MUX2_X1 U6703 ( .A(n6058), .B(n5523), .S(EBX_REG_14__SCAN_IN), .Z(n6015) );
  OR2_X1 U6704 ( .A1(n6114), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6014)
         );
  MUX2_X1 U6705 ( .A(n6058), .B(n6049), .S(EBX_REG_16__SCAN_IN), .Z(n6017) );
  OR2_X1 U6706 ( .A1(n6114), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6016)
         );
  NAND2_X1 U6707 ( .A1(n6017), .A2(n6016), .ZN(n6239) );
  INV_X1 U6708 ( .A(n6239), .ZN(n6023) );
  INV_X1 U6709 ( .A(EBX_REG_15__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U6710 ( .A1(n6052), .A2(n7288), .ZN(n6022) );
  NAND2_X1 U6711 ( .A1(n6054), .A2(n4223), .ZN(n6020) );
  NAND2_X1 U6712 ( .A1(n6018), .A2(n7288), .ZN(n6019) );
  NAND3_X1 U6713 ( .A1(n6020), .A2(n5523), .A3(n6019), .ZN(n6021) );
  NAND2_X1 U6714 ( .A1(n6022), .A2(n6021), .ZN(n6250) );
  NAND2_X1 U6715 ( .A1(n6023), .A2(n6250), .ZN(n6024) );
  INV_X1 U6716 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U6717 ( .A1(n6052), .A2(n6351), .ZN(n6028) );
  NAND2_X1 U6718 ( .A1(n5523), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U6719 ( .A1(n6054), .A2(n6025), .ZN(n6026) );
  OAI21_X1 U6720 ( .B1(EBX_REG_17__SCAN_IN), .B2(n6113), .A(n6026), .ZN(n6027)
         );
  INV_X1 U6721 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U6722 ( .A1(n6029), .A2(n7444), .ZN(n6032) );
  NAND2_X1 U6723 ( .A1(n5523), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6030) );
  OAI211_X1 U6724 ( .C1(n6113), .C2(EBX_REG_18__SCAN_IN), .A(n6054), .B(n6030), 
        .ZN(n6031) );
  NAND2_X1 U6725 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U6726 ( .A1(n6054), .A2(n6033), .ZN(n6034) );
  OAI21_X1 U6727 ( .B1(EBX_REG_19__SCAN_IN), .B2(n6113), .A(n6034), .ZN(n6035)
         );
  OAI21_X1 U6728 ( .B1(n6107), .B2(EBX_REG_19__SCAN_IN), .A(n6035), .ZN(n6333)
         );
  NAND2_X1 U6729 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U6730 ( .C1(n6113), .C2(EBX_REG_20__SCAN_IN), .A(n6054), .B(n6036), 
        .ZN(n6037) );
  OAI21_X1 U6731 ( .B1(n6058), .B2(EBX_REG_20__SCAN_IN), .A(n6037), .ZN(n6222)
         );
  NAND2_X1 U6732 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U6733 ( .A1(n6054), .A2(n6038), .ZN(n6039) );
  OAI21_X1 U6734 ( .B1(EBX_REG_21__SCAN_IN), .B2(n6113), .A(n6039), .ZN(n6040)
         );
  OAI21_X1 U6735 ( .B1(n6107), .B2(EBX_REG_21__SCAN_IN), .A(n6040), .ZN(n6321)
         );
  MUX2_X1 U6736 ( .A(n6058), .B(n5523), .S(EBX_REG_22__SCAN_IN), .Z(n6041) );
  OAI21_X1 U6737 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6114), .A(n6041), 
        .ZN(n6210) );
  INV_X1 U6738 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U6739 ( .A1(n6052), .A2(n6315), .ZN(n6045) );
  NAND2_X1 U6740 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U6741 ( .A1(n6054), .A2(n6042), .ZN(n6043) );
  OAI21_X1 U6742 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6113), .A(n6043), .ZN(n6044)
         );
  AND2_X1 U6743 ( .A1(n6045), .A2(n6044), .ZN(n6313) );
  MUX2_X1 U6744 ( .A(n6058), .B(n5523), .S(EBX_REG_24__SCAN_IN), .Z(n6046) );
  OAI21_X1 U6745 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n6114), .A(n6046), 
        .ZN(n6204) );
  INV_X1 U6746 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U6747 ( .A1(n6054), .A2(n6630), .ZN(n6047) );
  OAI211_X1 U6748 ( .C1(EBX_REG_25__SCAN_IN), .C2(n6113), .A(n6047), .B(n6049), 
        .ZN(n6048) );
  OAI21_X1 U6749 ( .B1(n6107), .B2(EBX_REG_25__SCAN_IN), .A(n6048), .ZN(n6188)
         );
  NAND2_X1 U6750 ( .A1(n6049), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U6751 ( .C1(n6113), .C2(EBX_REG_26__SCAN_IN), .A(n6054), .B(n6050), 
        .ZN(n6051) );
  OAI21_X1 U6752 ( .B1(n6058), .B2(EBX_REG_26__SCAN_IN), .A(n6051), .ZN(n6168)
         );
  INV_X1 U6753 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U6754 ( .A1(n6052), .A2(n6303), .ZN(n6057) );
  NAND2_X1 U6755 ( .A1(n5523), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U6756 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  OAI21_X1 U6757 ( .B1(EBX_REG_27__SCAN_IN), .B2(n6113), .A(n6055), .ZN(n6056)
         );
  AND2_X1 U6758 ( .A1(n6057), .A2(n6056), .ZN(n6157) );
  MUX2_X1 U6759 ( .A(n6058), .B(n6049), .S(EBX_REG_28__SCAN_IN), .Z(n6059) );
  OAI21_X1 U6760 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n6114), .A(n6059), 
        .ZN(n6146) );
  AOI22_X1 U6761 ( .A1(n6114), .A2(EBX_REG_30__SCAN_IN), .B1(n6113), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6109) );
  XNOR2_X1 U6762 ( .A(n6061), .B(n6109), .ZN(n6062) );
  OAI222_X1 U6763 ( .A1(n6355), .A2(n6005), .B1(n6352), .B2(n6076), .C1(n6062), 
        .C2(n6359), .ZN(U2829) );
  INV_X1 U6764 ( .A(n6062), .ZN(n6591) );
  INV_X1 U6765 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7232) );
  INV_X1 U6766 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7461) );
  INV_X1 U6767 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7228) );
  INV_X1 U6768 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7433) );
  INV_X1 U6769 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7223) );
  INV_X1 U6770 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7221) );
  NOR2_X1 U6771 ( .A1(n7223), .A2(n7221), .ZN(n7425) );
  INV_X1 U6772 ( .A(n7425), .ZN(n6236) );
  NAND2_X1 U6773 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n6283) );
  NAND3_X1 U6774 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n6282) );
  NOR2_X1 U6775 ( .A1(n6283), .A2(n6282), .ZN(n6265) );
  NAND3_X1 U6776 ( .A1(n6265), .A2(n6063), .A3(REIP_REG_14__SCAN_IN), .ZN(
        n6235) );
  NOR4_X1 U6777 ( .A1(n7433), .A2(n6064), .A3(n6236), .A4(n6235), .ZN(n7427)
         );
  NAND2_X1 U6778 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7427), .ZN(n7445) );
  NOR2_X1 U6779 ( .A1(n7228), .A2(n7445), .ZN(n6213) );
  NAND2_X1 U6780 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6213), .ZN(n6225) );
  NOR3_X1 U6781 ( .A1(n7232), .A2(n7461), .A3(n6225), .ZN(n7469) );
  NAND2_X1 U6782 ( .A1(REIP_REG_23__SCAN_IN), .A2(n7469), .ZN(n6196) );
  INV_X1 U6783 ( .A(n6196), .ZN(n6182) );
  NAND2_X1 U6784 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6182), .ZN(n6181) );
  INV_X1 U6785 ( .A(n6181), .ZN(n6065) );
  NAND2_X1 U6786 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6065), .ZN(n6066) );
  NOR2_X1 U6787 ( .A1(n7446), .A2(n6066), .ZN(n6173) );
  NAND2_X1 U6788 ( .A1(n6173), .A2(REIP_REG_26__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U6789 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n6069) );
  OR2_X1 U6790 ( .A1(n6159), .A2(n6069), .ZN(n6135) );
  INV_X1 U6791 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7248) );
  NOR2_X1 U6792 ( .A1(n6135), .A2(n7248), .ZN(n6073) );
  NAND2_X1 U6793 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n6071) );
  INV_X1 U6794 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7240) );
  INV_X1 U6795 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7239) );
  NOR3_X1 U6796 ( .A1(n7240), .A2(n7239), .A3(n6181), .ZN(n6067) );
  NAND2_X1 U6797 ( .A1(n7426), .A2(n6067), .ZN(n6068) );
  NAND2_X1 U6798 ( .A1(n7375), .A2(n6068), .ZN(n6171) );
  NAND2_X1 U6799 ( .A1(n7375), .A2(n6069), .ZN(n6070) );
  NAND2_X1 U6800 ( .A1(n6171), .A2(n6070), .ZN(n6147) );
  AOI21_X1 U6801 ( .B1(n7470), .B2(n6071), .A(n6147), .ZN(n6072) );
  INV_X1 U6802 ( .A(n6072), .ZN(n6125) );
  MUX2_X1 U6803 ( .A(n6073), .B(n6125), .S(REIP_REG_30__SCAN_IN), .Z(n6078) );
  AOI22_X1 U6804 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7472), .B1(n7475), 
        .B2(n6074), .ZN(n6075) );
  OAI21_X1 U6805 ( .B1(n6076), .B2(n7443), .A(n6075), .ZN(n6077) );
  AOI211_X1 U6806 ( .C1(n6591), .C2(n7473), .A(n6078), .B(n6077), .ZN(n6079)
         );
  OAI21_X1 U6807 ( .B1(n6005), .B2(n7437), .A(n6079), .ZN(U2797) );
  INV_X1 U6808 ( .A(n6080), .ZN(n6084) );
  NOR2_X1 U6809 ( .A1(n7543), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6083)
         );
  AOI222_X1 U6810 ( .A1(n6085), .A2(n6084), .B1(n4906), .B2(n6083), .C1(n6082), 
        .C2(n6081), .ZN(n6090) );
  AOI21_X1 U6811 ( .B1(n6087), .B2(n6086), .A(n6089), .ZN(n6088) );
  OAI22_X1 U6812 ( .A1(n6090), .A2(n6089), .B1(n6088), .B2(n3834), .ZN(U3459)
         );
  OAI211_X1 U6813 ( .C1(n6092), .C2(n3706), .A(n7553), .B(n6091), .ZN(n6094)
         );
  NAND2_X1 U6814 ( .A1(n7551), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6093) );
  OAI211_X1 U6815 ( .C1(n7549), .C2(n5129), .A(n6094), .B(n6093), .ZN(U3463)
         );
  NAND3_X1 U6816 ( .A1(n6095), .A2(n4853), .A3(n7509), .ZN(n6097) );
  INV_X1 U6817 ( .A(n6096), .ZN(n6101) );
  AOI22_X1 U6818 ( .A1(n6099), .A2(n6097), .B1(n4843), .B2(n6101), .ZN(n6098)
         );
  OAI21_X1 U6819 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n7513) );
  OAI21_X1 U6820 ( .B1(n4887), .B2(n6101), .A(n4853), .ZN(n6102) );
  OAI21_X1 U6821 ( .B1(n6104), .B2(n6103), .A(n6102), .ZN(n7295) );
  AOI21_X1 U6822 ( .B1(n6106), .B2(n6105), .A(READY_N), .ZN(n7301) );
  NOR2_X1 U6823 ( .A1(n7295), .A2(n7301), .ZN(n7508) );
  NOR2_X1 U6824 ( .A1(n7508), .A2(n7546), .ZN(n7484) );
  MUX2_X1 U6825 ( .A(MORE_REG_SCAN_IN), .B(n7513), .S(n7484), .Z(U3471) );
  OAI22_X1 U6826 ( .A1(n6108), .A2(n5093), .B1(EBX_REG_29__SCAN_IN), .B2(n6107), .ZN(n6139) );
  INV_X1 U6827 ( .A(n6139), .ZN(n6110) );
  NOR2_X1 U6828 ( .A1(n6110), .A2(n6109), .ZN(n6112) );
  AOI21_X1 U6829 ( .B1(n6145), .B2(n6112), .A(n6111), .ZN(n6116) );
  AOI22_X1 U6830 ( .A1(n6114), .A2(EBX_REG_31__SCAN_IN), .B1(n6113), .B2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U6831 ( .A(n6116), .B(n6115), .ZN(n6578) );
  NAND2_X1 U6832 ( .A1(n6118), .A2(n6117), .ZN(n6122) );
  AOI22_X1 U6833 ( .A1(n4766), .A2(EAX_REG_31__SCAN_IN), .B1(n6119), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6120) );
  INV_X1 U6834 ( .A(n6120), .ZN(n6121) );
  XNOR2_X2 U6835 ( .A(n6122), .B(n6121), .ZN(n6404) );
  NAND2_X1 U6836 ( .A1(n6404), .A2(n7477), .ZN(n6130) );
  NOR3_X1 U6837 ( .A1(n6124), .A2(n6300), .A3(n6123), .ZN(n6128) );
  INV_X1 U6838 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7251) );
  NOR3_X1 U6839 ( .A1(n6135), .A2(n7248), .A3(n7251), .ZN(n6126) );
  MUX2_X1 U6840 ( .A(n6126), .B(n6125), .S(REIP_REG_31__SCAN_IN), .Z(n6127) );
  AOI211_X1 U6841 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n7472), .A(n6128), 
        .B(n6127), .ZN(n6129) );
  OAI211_X1 U6842 ( .C1(n6578), .C2(n7467), .A(n6130), .B(n6129), .ZN(U2796)
         );
  INV_X1 U6843 ( .A(n6131), .ZN(n6366) );
  INV_X1 U6844 ( .A(n6132), .ZN(n6133) );
  OAI22_X1 U6845 ( .A1(n6134), .A2(n7450), .B1(n7420), .B2(n6133), .ZN(n6138)
         );
  INV_X1 U6846 ( .A(n6135), .ZN(n6136) );
  MUX2_X1 U6847 ( .A(n6136), .B(n6147), .S(REIP_REG_29__SCAN_IN), .Z(n6137) );
  AOI211_X1 U6848 ( .C1(EBX_REG_29__SCAN_IN), .C2(n7471), .A(n6138), .B(n6137), 
        .ZN(n6141) );
  XOR2_X1 U6849 ( .A(n6139), .B(n6145), .Z(n6598) );
  NAND2_X1 U6850 ( .A1(n6598), .A2(n7473), .ZN(n6140) );
  OAI211_X1 U6851 ( .C1(n6366), .C2(n7437), .A(n6141), .B(n6140), .ZN(U2798)
         );
  OR2_X1 U6852 ( .A1(n6142), .A2(n6143), .ZN(n6144) );
  AOI21_X1 U6853 ( .B1(n6146), .B2(n3714), .A(n6145), .ZN(n6606) );
  INV_X1 U6854 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6151) );
  INV_X1 U6855 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7244) );
  NOR2_X1 U6856 ( .A1(n6159), .A2(n7244), .ZN(n6148) );
  OAI21_X1 U6857 ( .B1(n6148), .B2(REIP_REG_28__SCAN_IN), .A(n6147), .ZN(n6150) );
  AOI22_X1 U6858 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7472), .B1(n7475), 
        .B2(n6408), .ZN(n6149) );
  OAI211_X1 U6859 ( .C1(n6151), .C2(n7443), .A(n6150), .B(n6149), .ZN(n6152)
         );
  AOI21_X1 U6860 ( .B1(n6606), .B2(n7473), .A(n6152), .ZN(n6153) );
  OAI21_X1 U6861 ( .B1(n6369), .B2(n7437), .A(n6153), .ZN(U2799) );
  NOR2_X1 U6862 ( .A1(n6154), .A2(n6155), .ZN(n6156) );
  NAND2_X1 U6863 ( .A1(n6170), .A2(n6157), .ZN(n6158) );
  NAND2_X1 U6864 ( .A1(n3714), .A2(n6158), .ZN(n6612) );
  INV_X1 U6865 ( .A(n6612), .ZN(n6163) );
  MUX2_X1 U6866 ( .A(n6159), .B(n6171), .S(REIP_REG_27__SCAN_IN), .Z(n6161) );
  AOI22_X1 U6867 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n7472), .B1(n7475), 
        .B2(n6422), .ZN(n6160) );
  OAI211_X1 U6868 ( .C1(n6303), .C2(n7443), .A(n6161), .B(n6160), .ZN(n6162)
         );
  AOI21_X1 U6869 ( .B1(n6163), .B2(n7473), .A(n6162), .ZN(n6164) );
  OAI21_X1 U6870 ( .B1(n6419), .B2(n7437), .A(n6164), .ZN(U2800) );
  INV_X1 U6871 ( .A(n6154), .ZN(n6166) );
  OAI21_X1 U6872 ( .B1(n6167), .B2(n6165), .A(n6166), .ZN(n6426) );
  NAND2_X1 U6873 ( .A1(n6190), .A2(n6168), .ZN(n6169) );
  AND2_X1 U6874 ( .A1(n6170), .A2(n6169), .ZN(n6624) );
  INV_X1 U6875 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6305) );
  INV_X1 U6876 ( .A(n6171), .ZN(n6172) );
  OAI21_X1 U6877 ( .B1(REIP_REG_26__SCAN_IN), .B2(n6173), .A(n6172), .ZN(n6175) );
  AOI22_X1 U6878 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n7472), .B1(n7475), 
        .B2(n6429), .ZN(n6174) );
  OAI211_X1 U6879 ( .C1(n7443), .C2(n6305), .A(n6175), .B(n6174), .ZN(n6176)
         );
  AOI21_X1 U6880 ( .B1(n6624), .B2(n7473), .A(n6176), .ZN(n6177) );
  OAI21_X1 U6881 ( .B1(n6426), .B2(n7437), .A(n6177), .ZN(U2801) );
  AOI21_X1 U6882 ( .B1(n6179), .B2(n6178), .A(n6165), .ZN(n6439) );
  INV_X1 U6883 ( .A(n6439), .ZN(n6376) );
  OAI22_X1 U6884 ( .A1(n6180), .A2(n7450), .B1(n7420), .B2(n6437), .ZN(n6187)
         );
  NOR2_X1 U6885 ( .A1(n7446), .A2(n6181), .ZN(n6185) );
  NAND2_X1 U6886 ( .A1(n7426), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U6887 ( .A1(n7375), .A2(n6183), .ZN(n7481) );
  INV_X1 U6888 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U6889 ( .A1(n7470), .A2(n7237), .ZN(n6184) );
  NAND2_X1 U6890 ( .A1(n7481), .A2(n6184), .ZN(n6202) );
  MUX2_X1 U6891 ( .A(n6185), .B(n6202), .S(REIP_REG_25__SCAN_IN), .Z(n6186) );
  AOI211_X1 U6892 ( .C1(EBX_REG_25__SCAN_IN), .C2(n7471), .A(n6187), .B(n6186), 
        .ZN(n6192) );
  OR2_X1 U6893 ( .A1(n6203), .A2(n6188), .ZN(n6189) );
  AND2_X1 U6894 ( .A1(n6190), .A2(n6189), .ZN(n6632) );
  NAND2_X1 U6895 ( .A1(n6632), .A2(n7473), .ZN(n6191) );
  OAI211_X1 U6896 ( .C1(n6376), .C2(n7437), .A(n6192), .B(n6191), .ZN(U2802)
         );
  INV_X1 U6897 ( .A(n6178), .ZN(n6194) );
  AOI21_X1 U6898 ( .B1(n6195), .B2(n6308), .A(n6194), .ZN(n6453) );
  INV_X1 U6899 ( .A(n6453), .ZN(n6379) );
  OAI21_X1 U6900 ( .B1(n7446), .B2(n6196), .A(n7237), .ZN(n6201) );
  INV_X1 U6901 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6197) );
  NOR2_X1 U6902 ( .A1(n7443), .A2(n6197), .ZN(n6200) );
  OAI22_X1 U6903 ( .A1(n6198), .A2(n7450), .B1(n7420), .B2(n6451), .ZN(n6199)
         );
  AOI211_X1 U6904 ( .C1(n6202), .C2(n6201), .A(n6200), .B(n6199), .ZN(n6206)
         );
  AOI21_X1 U6905 ( .B1(n6204), .B2(n6310), .A(n6203), .ZN(n6640) );
  NAND2_X1 U6906 ( .A1(n6640), .A2(n7473), .ZN(n6205) );
  OAI211_X1 U6907 ( .C1(n6379), .C2(n7437), .A(n6206), .B(n6205), .ZN(U2803)
         );
  OAI21_X1 U6908 ( .B1(n6207), .B2(n6209), .A(n6208), .ZN(n6466) );
  AOI21_X1 U6909 ( .B1(n6210), .B2(n6324), .A(n3760), .ZN(n6654) );
  INV_X1 U6910 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6318) );
  INV_X1 U6911 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U6912 ( .A1(n6465), .A2(n7450), .ZN(n6211) );
  AOI21_X1 U6913 ( .B1(n7475), .B2(n6469), .A(n6211), .ZN(n6212) );
  OAI21_X1 U6914 ( .B1(n7443), .B2(n6318), .A(n6212), .ZN(n6217) );
  INV_X1 U6915 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U6916 ( .A1(n7470), .A2(n6213), .ZN(n6227) );
  NOR2_X1 U6917 ( .A1(n7230), .A2(n6227), .ZN(n7462) );
  AOI21_X1 U6918 ( .B1(REIP_REG_21__SCAN_IN), .B2(n7462), .A(
        REIP_REG_22__SCAN_IN), .ZN(n6215) );
  INV_X1 U6919 ( .A(n7375), .ZN(n6214) );
  AOI211_X1 U6920 ( .C1(n7469), .C2(n7426), .A(n6215), .B(n6214), .ZN(n6216)
         );
  AOI211_X1 U6921 ( .C1(n6654), .C2(n7473), .A(n6217), .B(n6216), .ZN(n6218)
         );
  OAI21_X1 U6922 ( .B1(n6466), .B2(n7437), .A(n6218), .ZN(U2805) );
  AND2_X1 U6923 ( .A1(n6330), .A2(n6219), .ZN(n6221) );
  AND2_X1 U6924 ( .A1(n3724), .A2(n6222), .ZN(n6223) );
  OR2_X1 U6925 ( .A1(n6322), .A2(n6223), .ZN(n6669) );
  INV_X1 U6926 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6481) );
  INV_X1 U6927 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6326) );
  OAI22_X1 U6928 ( .A1(n6481), .A2(n7450), .B1(n6326), .B2(n7443), .ZN(n6224)
         );
  AOI21_X1 U6929 ( .B1(n7475), .B2(n6485), .A(n6224), .ZN(n6230) );
  INV_X1 U6930 ( .A(n6225), .ZN(n6226) );
  OAI21_X1 U6931 ( .B1(n7446), .B2(n6226), .A(n7426), .ZN(n7460) );
  NAND2_X1 U6932 ( .A1(n6227), .A2(n7230), .ZN(n6228) );
  NAND2_X1 U6933 ( .A1(n7460), .A2(n6228), .ZN(n6229) );
  OAI211_X1 U6934 ( .C1(n6669), .C2(n7467), .A(n6230), .B(n6229), .ZN(n6231)
         );
  INV_X1 U6935 ( .A(n6231), .ZN(n6232) );
  OAI21_X1 U6936 ( .B1(n6482), .B2(n7437), .A(n6232), .ZN(U2807) );
  OAI21_X1 U6937 ( .B1(n3708), .B2(n4503), .A(n6234), .ZN(n6508) );
  OAI21_X1 U6938 ( .B1(n6235), .B2(n7376), .A(n7375), .ZN(n6267) );
  AOI21_X1 U6939 ( .B1(n7472), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7423), 
        .ZN(n6238) );
  NOR2_X1 U6940 ( .A1(n6235), .A2(n7388), .ZN(n7424) );
  OAI211_X1 U6941 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n7424), .B(n6236), .ZN(n6237) );
  OAI211_X1 U6942 ( .C1(n6267), .C2(n7223), .A(n6238), .B(n6237), .ZN(n6246)
         );
  INV_X1 U6943 ( .A(n6250), .ZN(n6240) );
  OAI21_X1 U6944 ( .B1(n6259), .B2(n6240), .A(n6239), .ZN(n6241) );
  AND2_X1 U6945 ( .A1(n6241), .A2(n6345), .ZN(n7331) );
  INV_X1 U6946 ( .A(n7331), .ZN(n6244) );
  INV_X1 U6947 ( .A(n6242), .ZN(n6505) );
  AOI22_X1 U6948 ( .A1(n7471), .A2(EBX_REG_16__SCAN_IN), .B1(n7475), .B2(n6505), .ZN(n6243) );
  OAI21_X1 U6949 ( .B1(n6244), .B2(n7467), .A(n6243), .ZN(n6245) );
  NOR2_X1 U6950 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  OAI21_X1 U6951 ( .B1(n6508), .B2(n7437), .A(n6247), .ZN(U2811) );
  AOI21_X1 U6952 ( .B1(n6249), .B2(n6248), .A(n3708), .ZN(n7286) );
  INV_X1 U6953 ( .A(n7286), .ZN(n6388) );
  XNOR2_X1 U6954 ( .A(n6259), .B(n6250), .ZN(n7283) );
  INV_X1 U6955 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6515) );
  AOI21_X1 U6956 ( .B1(n7475), .B2(n6512), .A(n7423), .ZN(n6251) );
  OAI21_X1 U6957 ( .B1(n7450), .B2(n6515), .A(n6251), .ZN(n6254) );
  AOI22_X1 U6958 ( .A1(EBX_REG_15__SCAN_IN), .A2(n7471), .B1(n7424), .B2(n7221), .ZN(n6252) );
  OAI21_X1 U6959 ( .B1(n7221), .B2(n6267), .A(n6252), .ZN(n6253) );
  AOI211_X1 U6960 ( .C1(n7473), .C2(n7283), .A(n6254), .B(n6253), .ZN(n6255)
         );
  OAI21_X1 U6961 ( .B1(n6388), .B2(n7437), .A(n6255), .ZN(U2812) );
  OAI21_X1 U6962 ( .B1(n6257), .B2(n6256), .A(n6248), .ZN(n6522) );
  OR2_X1 U6963 ( .A1(n6277), .A2(n6258), .ZN(n6260) );
  AND2_X1 U6964 ( .A1(n6260), .A2(n6259), .ZN(n6722) );
  INV_X1 U6965 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6356) );
  INV_X1 U6966 ( .A(n6525), .ZN(n6263) );
  OAI21_X1 U6967 ( .B1(n7450), .B2(n6261), .A(n7448), .ZN(n6262) );
  AOI21_X1 U6968 ( .B1(n7475), .B2(n6263), .A(n6262), .ZN(n6264) );
  OAI21_X1 U6969 ( .B1(n7443), .B2(n6356), .A(n6264), .ZN(n6271) );
  INV_X1 U6970 ( .A(n6265), .ZN(n6266) );
  NOR2_X1 U6971 ( .A1(n6266), .A2(n6281), .ZN(n6269) );
  INV_X1 U6972 ( .A(n6267), .ZN(n6268) );
  MUX2_X1 U6973 ( .A(n6269), .B(n6268), .S(REIP_REG_14__SCAN_IN), .Z(n6270) );
  AOI211_X1 U6974 ( .C1(n6722), .C2(n7473), .A(n6271), .B(n6270), .ZN(n6272)
         );
  OAI21_X1 U6975 ( .B1(n6522), .B2(n7437), .A(n6272), .ZN(U2813) );
  XOR2_X1 U6976 ( .A(n6274), .B(n6273), .Z(n6535) );
  INV_X1 U6977 ( .A(n6535), .ZN(n6392) );
  INV_X1 U6978 ( .A(n6532), .ZN(n6287) );
  NOR2_X1 U6979 ( .A1(n3722), .A2(n6275), .ZN(n6276) );
  OR2_X1 U6980 ( .A1(n6277), .A2(n6276), .ZN(n6743) );
  NAND2_X1 U6981 ( .A1(n6282), .A2(n7375), .ZN(n7407) );
  NAND2_X1 U6982 ( .A1(n7407), .A2(n6278), .ZN(n7415) );
  INV_X1 U6983 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6279) );
  OAI22_X1 U6984 ( .A1(n6279), .A2(n7450), .B1(n6358), .B2(n7443), .ZN(n6280)
         );
  AOI211_X1 U6985 ( .C1(REIP_REG_13__SCAN_IN), .C2(n7415), .A(n7423), .B(n6280), .ZN(n6285) );
  NOR2_X1 U6986 ( .A1(n6282), .A2(n6281), .ZN(n7417) );
  OAI211_X1 U6987 ( .C1(REIP_REG_12__SCAN_IN), .C2(REIP_REG_13__SCAN_IN), .A(
        n7417), .B(n6283), .ZN(n6284) );
  OAI211_X1 U6988 ( .C1(n6743), .C2(n7467), .A(n6285), .B(n6284), .ZN(n6286)
         );
  AOI21_X1 U6989 ( .B1(n7475), .B2(n6287), .A(n6286), .ZN(n6288) );
  OAI21_X1 U6990 ( .B1(n6392), .B2(n7437), .A(n6288), .ZN(U2814) );
  NAND2_X1 U6991 ( .A1(n6289), .A2(n7370), .ZN(n6299) );
  AOI22_X1 U6992 ( .A1(EBX_REG_2__SCAN_IN), .A2(n7471), .B1(n7473), .B2(n6290), 
        .ZN(n6291) );
  OAI21_X1 U6993 ( .B1(n7426), .B2(n7199), .A(n6291), .ZN(n6294) );
  NOR2_X1 U6994 ( .A1(n7420), .A2(n6292), .ZN(n6293) );
  AOI211_X1 U6995 ( .C1(n7472), .C2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6294), 
        .B(n6293), .ZN(n6298) );
  NAND2_X1 U6996 ( .A1(n7358), .A2(n3665), .ZN(n6297) );
  OAI211_X1 U6997 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n7470), .B(n6295), .ZN(n6296) );
  NAND4_X1 U6998 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(U2825)
         );
  OAI22_X1 U6999 ( .A1(n6578), .A2(n6359), .B1(n6300), .B2(n6352), .ZN(U2828)
         );
  AOI22_X1 U7000 ( .A1(n6598), .A2(n7284), .B1(EBX_REG_29__SCAN_IN), .B2(n6353), .ZN(n6301) );
  OAI21_X1 U7001 ( .B1(n6366), .B2(n6355), .A(n6301), .ZN(U2830) );
  AOI22_X1 U7002 ( .A1(n6606), .A2(n7284), .B1(n6353), .B2(EBX_REG_28__SCAN_IN), .ZN(n6302) );
  OAI21_X1 U7003 ( .B1(n6369), .B2(n6355), .A(n6302), .ZN(U2831) );
  OAI222_X1 U7004 ( .A1(n6303), .A2(n6352), .B1(n6359), .B2(n6612), .C1(n6419), 
        .C2(n6355), .ZN(U2832) );
  INV_X1 U7005 ( .A(n6624), .ZN(n6304) );
  OAI222_X1 U7006 ( .A1(n6305), .A2(n6352), .B1(n6359), .B2(n6304), .C1(n6426), 
        .C2(n6355), .ZN(U2833) );
  AOI22_X1 U7007 ( .A1(n6632), .A2(n7284), .B1(n6353), .B2(EBX_REG_25__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7008 ( .B1(n6376), .B2(n6355), .A(n6306), .ZN(U2834) );
  INV_X1 U7009 ( .A(n6640), .ZN(n6307) );
  OAI222_X1 U7010 ( .A1(n6355), .A2(n6379), .B1(n6352), .B2(n6197), .C1(n6307), 
        .C2(n6359), .ZN(U2835) );
  AOI21_X1 U7011 ( .B1(n6309), .B2(n6208), .A(n6193), .ZN(n7582) );
  INV_X1 U7012 ( .A(n7582), .ZN(n6316) );
  INV_X1 U7013 ( .A(n6310), .ZN(n6311) );
  AOI21_X1 U7014 ( .B1(n6313), .B2(n6312), .A(n6311), .ZN(n7474) );
  INV_X1 U7015 ( .A(n7474), .ZN(n6314) );
  OAI222_X1 U7016 ( .A1(n6355), .A2(n6316), .B1(n6352), .B2(n6315), .C1(n6314), 
        .C2(n6359), .ZN(U2836) );
  INV_X1 U7017 ( .A(n6654), .ZN(n6317) );
  OAI222_X1 U7018 ( .A1(n6318), .A2(n6352), .B1(n6359), .B2(n6317), .C1(n6466), 
        .C2(n6355), .ZN(U2837) );
  INV_X1 U7019 ( .A(n6207), .ZN(n6319) );
  OAI21_X1 U7020 ( .B1(n6320), .B2(n6220), .A(n6319), .ZN(n7463) );
  INV_X1 U7021 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6325) );
  OR2_X1 U7022 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  NAND2_X1 U7023 ( .A1(n6324), .A2(n6323), .ZN(n7468) );
  OAI222_X1 U7024 ( .A1(n6355), .A2(n7463), .B1(n6352), .B2(n6325), .C1(n7468), 
        .C2(n6359), .ZN(U2838) );
  OAI22_X1 U7025 ( .A1(n6669), .A2(n6359), .B1(n6326), .B2(n6352), .ZN(n6327)
         );
  INV_X1 U7026 ( .A(n6327), .ZN(n6328) );
  OAI21_X1 U7027 ( .B1(n6482), .B2(n6355), .A(n6328), .ZN(U2839) );
  INV_X1 U7028 ( .A(n6330), .ZN(n6331) );
  AOI21_X1 U7029 ( .B1(n6332), .B2(n6329), .A(n6331), .ZN(n7574) );
  INV_X1 U7030 ( .A(n7574), .ZN(n6336) );
  INV_X1 U7031 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6335) );
  OR2_X1 U7032 ( .A1(n6341), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7033 ( .A1(n3724), .A2(n6334), .ZN(n7457) );
  OAI222_X1 U7034 ( .A1(n6355), .A2(n6336), .B1(n6352), .B2(n6335), .C1(n7457), 
        .C2(n6359), .ZN(U2840) );
  OAI21_X1 U7035 ( .B1(n6337), .B2(n6338), .A(n6329), .ZN(n7438) );
  NOR2_X1 U7036 ( .A1(n6346), .A2(n6339), .ZN(n6340) );
  OR2_X1 U7037 ( .A1(n6341), .A2(n6340), .ZN(n7436) );
  OAI22_X1 U7038 ( .A1(n7436), .A2(n6359), .B1(n7444), .B2(n6352), .ZN(n6342)
         );
  INV_X1 U7039 ( .A(n6342), .ZN(n6343) );
  OAI21_X1 U7040 ( .B1(n7438), .B2(n6355), .A(n6343), .ZN(U2841) );
  AND2_X1 U7041 ( .A1(n6345), .A2(n6344), .ZN(n6347) );
  OR2_X1 U7042 ( .A1(n6347), .A2(n6346), .ZN(n7431) );
  AND2_X1 U7043 ( .A1(n6234), .A2(n6348), .ZN(n6349) );
  NOR2_X1 U7044 ( .A1(n6337), .A2(n6349), .ZN(n7571) );
  INV_X1 U7045 ( .A(n7571), .ZN(n6350) );
  OAI222_X1 U7046 ( .A1(n6359), .A2(n7431), .B1(n6352), .B2(n6351), .C1(n6355), 
        .C2(n6350), .ZN(U2842) );
  AOI22_X1 U7047 ( .A1(n7331), .A2(n7284), .B1(n6353), .B2(EBX_REG_16__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U7048 ( .B1(n6508), .B2(n6355), .A(n6354), .ZN(U2843) );
  INV_X1 U7049 ( .A(n6722), .ZN(n6357) );
  OAI222_X1 U7050 ( .A1(n6357), .A2(n6359), .B1(n6356), .B2(n6352), .C1(n6522), 
        .C2(n6355), .ZN(U2845) );
  OAI22_X1 U7051 ( .A1(n6743), .A2(n6359), .B1(n6358), .B2(n6352), .ZN(n6360)
         );
  AOI21_X1 U7052 ( .B1(n6535), .B2(n7285), .A(n6360), .ZN(n6361) );
  INV_X1 U7053 ( .A(n6361), .ZN(U2846) );
  NAND3_X1 U7054 ( .A1(n6404), .A2(n3901), .A3(n6391), .ZN(n6363) );
  AOI22_X1 U7055 ( .A1(n7580), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7583), .ZN(n6362) );
  NAND2_X1 U7056 ( .A1(n6363), .A2(n6362), .ZN(U2860) );
  AOI22_X1 U7057 ( .A1(n7580), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n7583), .ZN(n6365) );
  NAND2_X1 U7058 ( .A1(n7584), .A2(DATAI_13_), .ZN(n6364) );
  OAI211_X1 U7059 ( .C1(n6366), .C2(n7570), .A(n6365), .B(n6364), .ZN(U2862)
         );
  AOI22_X1 U7060 ( .A1(n7580), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n7583), .ZN(n6368) );
  NAND2_X1 U7061 ( .A1(n7584), .A2(DATAI_12_), .ZN(n6367) );
  OAI211_X1 U7062 ( .C1(n6369), .C2(n7570), .A(n6368), .B(n6367), .ZN(U2863)
         );
  AOI22_X1 U7063 ( .A1(n7580), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n7583), .ZN(n6371) );
  NAND2_X1 U7064 ( .A1(n7584), .A2(DATAI_11_), .ZN(n6370) );
  OAI211_X1 U7065 ( .C1(n6419), .C2(n7570), .A(n6371), .B(n6370), .ZN(U2864)
         );
  AOI22_X1 U7066 ( .A1(n7580), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n7583), .ZN(n6373) );
  NAND2_X1 U7067 ( .A1(n7584), .A2(DATAI_10_), .ZN(n6372) );
  OAI211_X1 U7068 ( .C1(n6426), .C2(n7570), .A(n6373), .B(n6372), .ZN(U2865)
         );
  AOI22_X1 U7069 ( .A1(n7580), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n7583), .ZN(n6375) );
  NAND2_X1 U7070 ( .A1(n7584), .A2(DATAI_9_), .ZN(n6374) );
  OAI211_X1 U7071 ( .C1(n6376), .C2(n7570), .A(n6375), .B(n6374), .ZN(U2866)
         );
  AOI22_X1 U7072 ( .A1(n7580), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7583), .ZN(n6378) );
  NAND2_X1 U7073 ( .A1(n7584), .A2(DATAI_8_), .ZN(n6377) );
  OAI211_X1 U7074 ( .C1(n6379), .C2(n7570), .A(n6378), .B(n6377), .ZN(U2867)
         );
  AOI22_X1 U7075 ( .A1(n7580), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7583), .ZN(n6381) );
  NAND2_X1 U7076 ( .A1(n7584), .A2(DATAI_6_), .ZN(n6380) );
  OAI211_X1 U7077 ( .C1(n6466), .C2(n7570), .A(n6381), .B(n6380), .ZN(U2869)
         );
  AOI22_X1 U7078 ( .A1(n7580), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n7583), .ZN(n6383) );
  NAND2_X1 U7079 ( .A1(n7584), .A2(DATAI_4_), .ZN(n6382) );
  OAI211_X1 U7080 ( .C1(n6482), .C2(n7570), .A(n6383), .B(n6382), .ZN(U2871)
         );
  AOI22_X1 U7081 ( .A1(n7580), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n7583), .ZN(n6385) );
  NAND2_X1 U7082 ( .A1(n7584), .A2(DATAI_2_), .ZN(n6384) );
  OAI211_X1 U7083 ( .C1(n7438), .C2(n7570), .A(n6385), .B(n6384), .ZN(U2873)
         );
  AOI22_X1 U7084 ( .A1(n7580), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n7583), .ZN(n6387) );
  NAND2_X1 U7085 ( .A1(n7584), .A2(DATAI_0_), .ZN(n6386) );
  OAI211_X1 U7086 ( .C1(n6508), .C2(n7570), .A(n6387), .B(n6386), .ZN(U2875)
         );
  INV_X1 U7087 ( .A(DATAI_15_), .ZN(n6389) );
  INV_X1 U7088 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7197) );
  OAI222_X1 U7089 ( .A1(n6389), .A2(n6394), .B1(n6391), .B2(n7197), .C1(n7570), 
        .C2(n6388), .ZN(U2876) );
  INV_X1 U7090 ( .A(DATAI_14_), .ZN(n6390) );
  OAI222_X1 U7091 ( .A1(n6394), .A2(n6390), .B1(n6391), .B2(n4993), .C1(n7570), 
        .C2(n6522), .ZN(U2877) );
  INV_X1 U7092 ( .A(DATAI_13_), .ZN(n6393) );
  OAI222_X1 U7093 ( .A1(n6394), .A2(n6393), .B1(n7570), .B2(n6392), .C1(n7191), 
        .C2(n6391), .ZN(U2878) );
  NAND3_X1 U7094 ( .A1(n6593), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U7095 ( .A1(n3783), .A2(n6574), .ZN(n6398) );
  NOR2_X1 U7096 ( .A1(n6395), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6396)
         );
  AOI22_X1 U7097 ( .A1(n6399), .A2(n6398), .B1(n6397), .B2(n6396), .ZN(n6400)
         );
  XOR2_X1 U7098 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n6400), .Z(n6582) );
  AND2_X1 U7099 ( .A1(n6546), .A2(REIP_REG_31__SCAN_IN), .ZN(n6576) );
  AOI21_X1 U7100 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6576), 
        .ZN(n6401) );
  OAI21_X1 U7101 ( .B1(n7294), .B2(n6402), .A(n6401), .ZN(n6403) );
  INV_X1 U7102 ( .A(n6408), .ZN(n6410) );
  AND2_X1 U7103 ( .A1(n6546), .A2(REIP_REG_28__SCAN_IN), .ZN(n6605) );
  AOI21_X1 U7104 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6605), 
        .ZN(n6409) );
  OAI21_X1 U7105 ( .B1(n7294), .B2(n6410), .A(n6409), .ZN(n6411) );
  AOI21_X1 U7106 ( .B1(n6412), .B2(n6534), .A(n6411), .ZN(n6413) );
  OAI21_X1 U7107 ( .B1(n6609), .B2(n7482), .A(n6413), .ZN(U2958) );
  AND2_X1 U7108 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6618) );
  MUX2_X1 U7109 ( .A(n3783), .B(n6618), .S(n3686), .Z(n6415) );
  OAI21_X1 U7110 ( .B1(n6622), .B2(n6697), .A(n6415), .ZN(n6417) );
  XNOR2_X1 U7111 ( .A(n6417), .B(n6416), .ZN(n6617) );
  NAND2_X1 U7112 ( .A1(n6546), .A2(REIP_REG_27__SCAN_IN), .ZN(n6610) );
  OAI21_X1 U7113 ( .B1(n6516), .B2(n6418), .A(n6610), .ZN(n6421) );
  NOR2_X1 U7114 ( .A1(n6419), .A2(n6509), .ZN(n6420) );
  OAI21_X1 U7115 ( .B1(n6617), .B2(n7482), .A(n6423), .ZN(U2959) );
  XNOR2_X1 U7116 ( .A(n3783), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6424)
         );
  NAND2_X1 U7117 ( .A1(n6546), .A2(REIP_REG_26__SCAN_IN), .ZN(n6621) );
  OAI21_X1 U7118 ( .B1(n6516), .B2(n6425), .A(n6621), .ZN(n6428) );
  NOR2_X1 U7119 ( .A1(n6426), .A2(n6509), .ZN(n6427) );
  OAI21_X1 U7120 ( .B1(n6626), .B2(n7482), .A(n6430), .ZN(U2960) );
  AOI21_X1 U7122 ( .B1(n6434), .B2(n6432), .A(n6433), .ZN(n6634) );
  NAND2_X1 U7123 ( .A1(n7330), .A2(REIP_REG_25__SCAN_IN), .ZN(n6629) );
  INV_X1 U7124 ( .A(n6629), .ZN(n6435) );
  AOI21_X1 U7125 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6435), 
        .ZN(n6436) );
  OAI21_X1 U7126 ( .B1(n7294), .B2(n6437), .A(n6436), .ZN(n6438) );
  AOI21_X1 U7127 ( .B1(n6439), .B2(n6534), .A(n6438), .ZN(n6440) );
  OAI21_X1 U7128 ( .B1(n6634), .B2(n7482), .A(n6440), .ZN(U2961) );
  XNOR2_X1 U7129 ( .A(n3783), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6488)
         );
  INV_X1 U7130 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6668) );
  XNOR2_X1 U7131 ( .A(n3783), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6472)
         );
  NOR2_X1 U7132 ( .A1(n6473), .A2(n6472), .ZN(n6471) );
  NAND3_X1 U7133 ( .A1(n6697), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6448) );
  INV_X1 U7134 ( .A(n6445), .ZN(n6447) );
  NAND3_X1 U7135 ( .A1(n6447), .A2(n3783), .A3(n6446), .ZN(n6455) );
  OAI22_X1 U7136 ( .A1(n6464), .A2(n6448), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6455), .ZN(n6449) );
  XNOR2_X1 U7137 ( .A(n6449), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6642)
         );
  NAND2_X1 U7138 ( .A1(n7330), .A2(REIP_REG_24__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U7139 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6450)
         );
  OAI211_X1 U7140 ( .C1(n7294), .C2(n6451), .A(n6636), .B(n6450), .ZN(n6452)
         );
  AOI21_X1 U7141 ( .B1(n6453), .B2(n6534), .A(n6452), .ZN(n6454) );
  OAI21_X1 U7142 ( .B1(n6642), .B2(n7482), .A(n6454), .ZN(U2962) );
  NAND3_X1 U7143 ( .A1(n6697), .A2(n6570), .A3(n6565), .ZN(n6456) );
  OAI21_X1 U7144 ( .B1(n3682), .B2(n6456), .A(n6455), .ZN(n6458) );
  XNOR2_X1 U7145 ( .A(n6458), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6648)
         );
  NAND2_X1 U7146 ( .A1(n6513), .A2(n7476), .ZN(n6459) );
  NAND2_X1 U7147 ( .A1(n7330), .A2(REIP_REG_23__SCAN_IN), .ZN(n6643) );
  OAI211_X1 U7148 ( .C1(n6516), .C2(n6460), .A(n6459), .B(n6643), .ZN(n6461)
         );
  AOI21_X1 U7149 ( .B1(n7582), .B2(n6534), .A(n6461), .ZN(n6462) );
  OAI21_X1 U7150 ( .B1(n6648), .B2(n7482), .A(n6462), .ZN(U2963) );
  XNOR2_X1 U7151 ( .A(n3783), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6463)
         );
  XNOR2_X1 U7152 ( .A(n6464), .B(n6463), .ZN(n6656) );
  NAND2_X1 U7153 ( .A1(n7330), .A2(REIP_REG_22__SCAN_IN), .ZN(n6650) );
  OAI21_X1 U7154 ( .B1(n6516), .B2(n6465), .A(n6650), .ZN(n6468) );
  NOR2_X1 U7155 ( .A1(n6466), .A2(n6509), .ZN(n6467) );
  AOI211_X1 U7156 ( .C1(n6513), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6470)
         );
  OAI21_X1 U7157 ( .B1(n6656), .B2(n7482), .A(n6470), .ZN(U2964) );
  INV_X1 U7158 ( .A(n6471), .ZN(n6658) );
  NAND2_X1 U7159 ( .A1(n6473), .A2(n6472), .ZN(n6657) );
  NAND3_X1 U7160 ( .A1(n6658), .A2(n7290), .A3(n6657), .ZN(n6478) );
  INV_X1 U7161 ( .A(n6474), .ZN(n7464) );
  NAND2_X1 U7162 ( .A1(n7330), .A2(REIP_REG_21__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U7163 ( .B1(n6516), .B2(n6475), .A(n6660), .ZN(n6476) );
  AOI21_X1 U7164 ( .B1(n7464), .B2(n6513), .A(n6476), .ZN(n6477) );
  OAI211_X1 U7165 ( .C1(n6509), .C2(n7463), .A(n6478), .B(n6477), .ZN(U2965)
         );
  NAND2_X1 U7166 ( .A1(n6697), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6479) );
  MUX2_X1 U7167 ( .A(n6479), .B(n6697), .S(n6487), .Z(n6480) );
  XOR2_X1 U7168 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(n6480), .Z(n6674) );
  NAND2_X1 U7169 ( .A1(n7330), .A2(REIP_REG_20__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7170 ( .B1(n6516), .B2(n6481), .A(n6667), .ZN(n6484) );
  NOR2_X1 U7171 ( .A1(n6482), .A2(n6509), .ZN(n6483) );
  AOI211_X1 U7172 ( .C1(n6513), .C2(n6485), .A(n6484), .B(n6483), .ZN(n6486)
         );
  OAI21_X1 U7173 ( .B1(n6674), .B2(n7482), .A(n6486), .ZN(U2966) );
  AOI21_X1 U7174 ( .B1(n6441), .B2(n6488), .A(n6487), .ZN(n6682) );
  INV_X1 U7175 ( .A(n7447), .ZN(n6490) );
  NAND2_X1 U7176 ( .A1(n7330), .A2(REIP_REG_19__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7177 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6489)
         );
  OAI211_X1 U7178 ( .C1(n7294), .C2(n6490), .A(n6675), .B(n6489), .ZN(n6491)
         );
  AOI21_X1 U7179 ( .B1(n7574), .B2(n6534), .A(n6491), .ZN(n6492) );
  OAI21_X1 U7180 ( .B1(n6682), .B2(n7482), .A(n6492), .ZN(U2967) );
  NAND2_X1 U7181 ( .A1(n6493), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6496) );
  AOI21_X1 U7182 ( .B1(n3783), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6493), 
        .ZN(n6699) );
  INV_X1 U7183 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7184 ( .A1(n6699), .A2(n6494), .ZN(n6495) );
  MUX2_X1 U7185 ( .A(n6496), .B(n6495), .S(n3783), .Z(n6497) );
  XOR2_X1 U7186 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n6497), .Z(n6696) );
  NAND2_X1 U7187 ( .A1(n7330), .A2(REIP_REG_18__SCAN_IN), .ZN(n6692) );
  OAI21_X1 U7188 ( .B1(n6516), .B2(n7434), .A(n6692), .ZN(n6499) );
  NOR2_X1 U7189 ( .A1(n7438), .A2(n6509), .ZN(n6498) );
  AOI211_X1 U7190 ( .C1(n6513), .C2(n7440), .A(n6499), .B(n6498), .ZN(n6500)
         );
  OAI21_X1 U7191 ( .B1(n6696), .B2(n7482), .A(n6500), .ZN(U2968) );
  XNOR2_X1 U7192 ( .A(n6697), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6502)
         );
  XNOR2_X1 U7193 ( .A(n6501), .B(n6502), .ZN(n7333) );
  NAND2_X1 U7194 ( .A1(n7333), .A2(n7290), .ZN(n6507) );
  OAI22_X1 U7195 ( .A1(n6516), .A2(n6503), .B1(n6759), .B2(n7223), .ZN(n6504)
         );
  AOI21_X1 U7196 ( .B1(n6513), .B2(n6505), .A(n6504), .ZN(n6506) );
  OAI211_X1 U7197 ( .C1(n6509), .C2(n6508), .A(n6507), .B(n6506), .ZN(U2970)
         );
  XNOR2_X1 U7198 ( .A(n6511), .B(n6510), .ZN(n6718) );
  NAND2_X1 U7199 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  NAND2_X1 U7200 ( .A1(n7330), .A2(REIP_REG_15__SCAN_IN), .ZN(n6713) );
  OAI211_X1 U7201 ( .C1(n6516), .C2(n6515), .A(n6514), .B(n6713), .ZN(n6517)
         );
  AOI21_X1 U7202 ( .B1(n7286), .B2(n6534), .A(n6517), .ZN(n6518) );
  OAI21_X1 U7203 ( .B1(n6718), .B2(n7482), .A(n6518), .ZN(U2971) );
  OAI21_X1 U7204 ( .B1(n6521), .B2(n6520), .A(n6519), .ZN(n6736) );
  INV_X1 U7205 ( .A(n6522), .ZN(n6527) );
  INV_X1 U7206 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6523) );
  NOR2_X1 U7207 ( .A1(n6759), .A2(n6523), .ZN(n6721) );
  AOI21_X1 U7208 ( .B1(n7289), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6721), 
        .ZN(n6524) );
  OAI21_X1 U7209 ( .B1(n7294), .B2(n6525), .A(n6524), .ZN(n6526) );
  AOI21_X1 U7210 ( .B1(n6527), .B2(n6534), .A(n6526), .ZN(n6528) );
  OAI21_X1 U7211 ( .B1(n6736), .B2(n7482), .A(n6528), .ZN(U2972) );
  XOR2_X1 U7212 ( .A(n3693), .B(n6529), .Z(n6748) );
  NAND2_X1 U7213 ( .A1(n7330), .A2(REIP_REG_13__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U7214 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6531)
         );
  OAI211_X1 U7215 ( .C1(n7294), .C2(n6532), .A(n6742), .B(n6531), .ZN(n6533)
         );
  AOI21_X1 U7216 ( .B1(n6535), .B2(n6534), .A(n6533), .ZN(n6536) );
  OAI21_X1 U7217 ( .B1(n6748), .B2(n7482), .A(n6536), .ZN(U2973) );
  XNOR2_X1 U7218 ( .A(n6537), .B(n6538), .ZN(n6758) );
  INV_X1 U7219 ( .A(n6539), .ZN(n7410) );
  AOI22_X1 U7220 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6546), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6540) );
  OAI21_X1 U7221 ( .B1(n7294), .B2(n7408), .A(n6540), .ZN(n6541) );
  AOI21_X1 U7222 ( .B1(n7410), .B2(n6534), .A(n6541), .ZN(n6542) );
  OAI21_X1 U7223 ( .B1(n6758), .B2(n7482), .A(n6542), .ZN(U2974) );
  XNOR2_X1 U7224 ( .A(n6544), .B(n6543), .ZN(n6766) );
  INV_X1 U7225 ( .A(n6545), .ZN(n7401) );
  AOI22_X1 U7226 ( .A1(n7289), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6546), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U7227 ( .B1(n7294), .B2(n7401), .A(n6547), .ZN(n6548) );
  AOI21_X1 U7228 ( .B1(n6549), .B2(n6534), .A(n6548), .ZN(n6550) );
  OAI21_X1 U7229 ( .B1(n6766), .B2(n7482), .A(n6550), .ZN(U2975) );
  INV_X1 U7230 ( .A(n6574), .ZN(n6569) );
  NOR3_X1 U7231 ( .A1(n6552), .A2(n6551), .A3(n7320), .ZN(n6557) );
  NAND2_X1 U7232 ( .A1(n6553), .A2(n6557), .ZN(n6685) );
  INV_X1 U7233 ( .A(n6685), .ZN(n6725) );
  INV_X1 U7234 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U7235 ( .A1(n6753), .A2(n6752), .ZN(n6724) );
  NAND2_X1 U7236 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6724), .ZN(n6719) );
  NOR2_X1 U7237 ( .A1(n6712), .A2(n6719), .ZN(n6711) );
  NAND3_X1 U7238 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6711), .ZN(n6701) );
  INV_X1 U7239 ( .A(n6554), .ZN(n6555) );
  NOR2_X1 U7240 ( .A1(n6701), .A2(n6555), .ZN(n6558) );
  NAND2_X1 U7241 ( .A1(n6725), .A2(n6558), .ZN(n6559) );
  AND2_X1 U7242 ( .A1(n6557), .A2(n6556), .ZN(n6723) );
  NAND2_X1 U7243 ( .A1(n6723), .A2(n6558), .ZN(n6561) );
  OAI22_X1 U7244 ( .A1(n6741), .A2(n6559), .B1(n6683), .B2(n6561), .ZN(n6680)
         );
  NAND2_X1 U7245 ( .A1(n6680), .A2(n6565), .ZN(n6659) );
  OR2_X1 U7246 ( .A1(n6659), .A2(n6570), .ZN(n6652) );
  INV_X1 U7247 ( .A(n6559), .ZN(n6560) );
  OR2_X1 U7248 ( .A1(n6727), .A2(n6560), .ZN(n6564) );
  NAND2_X1 U7249 ( .A1(n6731), .A2(n6561), .ZN(n6562) );
  AND3_X1 U7250 ( .A1(n6564), .A2(n6563), .A3(n6562), .ZN(n6676) );
  NAND2_X1 U7251 ( .A1(n6687), .A2(n6443), .ZN(n6566) );
  AND2_X1 U7252 ( .A1(n6676), .A2(n6566), .ZN(n6661) );
  NAND2_X1 U7253 ( .A1(n6652), .A2(n6661), .ZN(n6649) );
  AOI21_X1 U7254 ( .B1(n6741), .B2(n6683), .A(n6572), .ZN(n6567) );
  NOR2_X1 U7255 ( .A1(n6649), .A2(n6567), .ZN(n6638) );
  OAI21_X1 U7256 ( .B1(n6710), .B2(n6618), .A(n6638), .ZN(n6615) );
  INV_X1 U7257 ( .A(n6615), .ZN(n6568) );
  OAI21_X1 U7258 ( .B1(n6710), .B2(n6569), .A(n6568), .ZN(n6577) );
  INV_X1 U7259 ( .A(n6570), .ZN(n6571) );
  INV_X1 U7260 ( .A(n6572), .ZN(n6573) );
  NOR2_X1 U7261 ( .A1(n6645), .A2(n6573), .ZN(n6627) );
  INV_X1 U7262 ( .A(n6603), .ZN(n6611) );
  NOR3_X1 U7263 ( .A1(n6611), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6574), 
        .ZN(n6575) );
  AOI211_X1 U7264 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n6577), .A(n6576), .B(n6575), .ZN(n6581) );
  INV_X1 U7265 ( .A(n6578), .ZN(n6579) );
  NAND2_X1 U7266 ( .A1(n6579), .A2(n7332), .ZN(n6580) );
  OAI211_X1 U7267 ( .C1(n6582), .C2(n6765), .A(n6581), .B(n6580), .ZN(U2987)
         );
  AOI211_X1 U7268 ( .C1(n6687), .C2(n6602), .A(n6584), .B(n6615), .ZN(n6596)
         );
  INV_X1 U7269 ( .A(n6638), .ZN(n6585) );
  OAI21_X1 U7270 ( .B1(n6585), .B2(n6687), .A(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n6589) );
  INV_X1 U7271 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6586) );
  NAND4_X1 U7272 ( .A1(n6603), .A2(n6593), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n6586), .ZN(n6588) );
  OAI211_X1 U7273 ( .C1(n6596), .C2(n6589), .A(n6588), .B(n6587), .ZN(n6590)
         );
  AOI21_X1 U7274 ( .B1(n6591), .B2(n7332), .A(n6590), .ZN(n6592) );
  OAI21_X1 U7275 ( .B1(n6583), .B2(n6765), .A(n6592), .ZN(U2988) );
  AOI21_X1 U7276 ( .B1(n6603), .B2(n6593), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n6595) );
  OAI21_X1 U7277 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(n6597) );
  AOI21_X1 U7278 ( .B1(n6598), .B2(n7332), .A(n6597), .ZN(n6599) );
  OAI21_X1 U7279 ( .B1(n6600), .B2(n6765), .A(n6599), .ZN(U2989) );
  AND3_X1 U7280 ( .A1(n6603), .A2(n6602), .A3(n6601), .ZN(n6604) );
  AOI211_X1 U7281 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n6615), .A(n6605), .B(n6604), .ZN(n6608) );
  NAND2_X1 U7282 ( .A1(n6606), .A2(n7332), .ZN(n6607) );
  OAI211_X1 U7283 ( .C1(n6609), .C2(n6765), .A(n6608), .B(n6607), .ZN(U2990)
         );
  OAI21_X1 U7284 ( .B1(n6611), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6610), 
        .ZN(n6614) );
  NOR2_X1 U7285 ( .A1(n6612), .A2(n7342), .ZN(n6613) );
  AOI211_X1 U7286 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n6615), .A(n6614), .B(n6613), .ZN(n6616) );
  OAI21_X1 U7287 ( .B1(n6617), .B2(n6765), .A(n6616), .ZN(U2991) );
  INV_X1 U7288 ( .A(n6618), .ZN(n6619) );
  OAI211_X1 U7289 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6627), .B(n6619), .ZN(n6620) );
  OAI211_X1 U7290 ( .C1(n6638), .C2(n6622), .A(n6621), .B(n6620), .ZN(n6623)
         );
  AOI21_X1 U7291 ( .B1(n6624), .B2(n7332), .A(n6623), .ZN(n6625) );
  OAI21_X1 U7292 ( .B1(n6626), .B2(n6765), .A(n6625), .ZN(U2992) );
  NAND2_X1 U7293 ( .A1(n6627), .A2(n6630), .ZN(n6628) );
  OAI211_X1 U7294 ( .C1(n6638), .C2(n6630), .A(n6629), .B(n6628), .ZN(n6631)
         );
  AOI21_X1 U7295 ( .B1(n6632), .B2(n7332), .A(n6631), .ZN(n6633) );
  OAI21_X1 U7296 ( .B1(n6634), .B2(n6765), .A(n6633), .ZN(U2993) );
  INV_X1 U7297 ( .A(n6645), .ZN(n6635) );
  AOI21_X1 U7298 ( .B1(n6635), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6637) );
  OAI21_X1 U7299 ( .B1(n6638), .B2(n6637), .A(n6636), .ZN(n6639) );
  AOI21_X1 U7300 ( .B1(n6640), .B2(n7332), .A(n6639), .ZN(n6641) );
  OAI21_X1 U7301 ( .B1(n6642), .B2(n6765), .A(n6641), .ZN(U2994) );
  NAND2_X1 U7302 ( .A1(n6649), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6644) );
  OAI211_X1 U7303 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6646) );
  AOI21_X1 U7304 ( .B1(n7474), .B2(n7332), .A(n6646), .ZN(n6647) );
  OAI21_X1 U7305 ( .B1(n6648), .B2(n6765), .A(n6647), .ZN(U2995) );
  INV_X1 U7306 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U7307 ( .A1(n6649), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6651) );
  OAI211_X1 U7308 ( .C1(n6652), .C2(n6663), .A(n6651), .B(n6650), .ZN(n6653)
         );
  AOI21_X1 U7309 ( .B1(n6654), .B2(n7332), .A(n6653), .ZN(n6655) );
  OAI21_X1 U7310 ( .B1(n6656), .B2(n6765), .A(n6655), .ZN(U2996) );
  NAND3_X1 U7311 ( .A1(n6658), .A2(n7344), .A3(n6657), .ZN(n6666) );
  INV_X1 U7312 ( .A(n6659), .ZN(n6664) );
  OAI21_X1 U7313 ( .B1(n6661), .B2(n6663), .A(n6660), .ZN(n6662) );
  AOI21_X1 U7314 ( .B1(n6664), .B2(n6663), .A(n6662), .ZN(n6665) );
  OAI211_X1 U7315 ( .C1(n7342), .C2(n7468), .A(n6666), .B(n6665), .ZN(U2997)
         );
  XOR2_X1 U7316 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .B(
        INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n6672) );
  OAI21_X1 U7317 ( .B1(n6676), .B2(n6668), .A(n6667), .ZN(n6671) );
  NOR2_X1 U7318 ( .A1(n6669), .A2(n7342), .ZN(n6670) );
  AOI211_X1 U7319 ( .C1(n6672), .C2(n6680), .A(n6671), .B(n6670), .ZN(n6673)
         );
  OAI21_X1 U7320 ( .B1(n6674), .B2(n6765), .A(n6673), .ZN(U2998) );
  INV_X1 U7321 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U7322 ( .B1(n6676), .B2(n6679), .A(n6675), .ZN(n6678) );
  NOR2_X1 U7323 ( .A1(n7457), .A2(n7342), .ZN(n6677) );
  AOI211_X1 U7324 ( .C1(n6680), .C2(n6679), .A(n6678), .B(n6677), .ZN(n6681)
         );
  OAI21_X1 U7325 ( .B1(n6682), .B2(n6765), .A(n6681), .ZN(U2999) );
  OAI21_X1 U7326 ( .B1(n6741), .B2(n6685), .A(n6683), .ZN(n6751) );
  INV_X1 U7327 ( .A(n6751), .ZN(n6688) );
  INV_X1 U7328 ( .A(n6727), .ZN(n6686) );
  NOR2_X1 U7329 ( .A1(n6723), .A2(n6683), .ZN(n6684) );
  AOI211_X1 U7330 ( .C1(n6686), .C2(n6685), .A(n6684), .B(n6729), .ZN(n6709)
         );
  INV_X1 U7331 ( .A(n6709), .ZN(n6763) );
  AOI21_X1 U7332 ( .B1(n6687), .B2(n6701), .A(n6763), .ZN(n6700) );
  OAI21_X1 U7333 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6688), .A(n6700), 
        .ZN(n6694) );
  NAND2_X1 U7334 ( .A1(n6751), .A2(n6723), .ZN(n6760) );
  INV_X1 U7335 ( .A(n6760), .ZN(n6703) );
  INV_X1 U7336 ( .A(n6701), .ZN(n6690) );
  INV_X1 U7337 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6689) );
  NAND4_X1 U7338 ( .A1(n6703), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6690), .A4(n6689), .ZN(n6691) );
  OAI211_X1 U7339 ( .C1(n7436), .C2(n7342), .A(n6692), .B(n6691), .ZN(n6693)
         );
  AOI21_X1 U7340 ( .B1(n6694), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6693), 
        .ZN(n6695) );
  OAI21_X1 U7341 ( .B1(n6696), .B2(n6765), .A(n6695), .ZN(U3000) );
  XNOR2_X1 U7342 ( .A(n6697), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6698)
         );
  XNOR2_X1 U7343 ( .A(n6699), .B(n6698), .ZN(n7291) );
  INV_X1 U7344 ( .A(n7291), .ZN(n6708) );
  INV_X1 U7345 ( .A(n6700), .ZN(n6706) );
  NOR2_X1 U7346 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6701), .ZN(n6702)
         );
  AOI22_X1 U7347 ( .A1(n6703), .A2(n6702), .B1(n7330), .B2(
        REIP_REG_17__SCAN_IN), .ZN(n6704) );
  OAI21_X1 U7348 ( .B1(n7431), .B2(n7342), .A(n6704), .ZN(n6705) );
  AOI21_X1 U7349 ( .B1(n6706), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6705), 
        .ZN(n6707) );
  OAI21_X1 U7350 ( .B1(n6708), .B2(n6765), .A(n6707), .ZN(U3001) );
  OAI21_X1 U7351 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(n7329) );
  INV_X1 U7352 ( .A(n7329), .ZN(n6715) );
  NOR3_X1 U7353 ( .A1(n6760), .A2(n6719), .A3(n6712), .ZN(n7334) );
  NAND2_X1 U7354 ( .A1(n7334), .A2(n4223), .ZN(n6714) );
  OAI211_X1 U7355 ( .C1(n4223), .C2(n6715), .A(n6714), .B(n6713), .ZN(n6716)
         );
  AOI21_X1 U7356 ( .B1(n7283), .B2(n7332), .A(n6716), .ZN(n6717) );
  OAI21_X1 U7357 ( .B1(n6718), .B2(n6765), .A(n6717), .ZN(U3003) );
  NOR3_X1 U7358 ( .A1(n6760), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6719), 
        .ZN(n6720) );
  AOI211_X1 U7359 ( .C1(n6722), .C2(n7332), .A(n6721), .B(n6720), .ZN(n6735)
         );
  NAND3_X1 U7360 ( .A1(n6725), .A2(n6724), .A3(n6730), .ZN(n6740) );
  NAND2_X1 U7361 ( .A1(n6724), .A2(n6723), .ZN(n6739) );
  AND2_X1 U7362 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  OAI22_X1 U7363 ( .A1(n6727), .A2(n6726), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n7348), .ZN(n6728) );
  AOI211_X1 U7364 ( .C1(n6731), .C2(n6739), .A(n6729), .B(n6728), .ZN(n6737)
         );
  NAND2_X1 U7365 ( .A1(n6731), .A2(n6730), .ZN(n6738) );
  OAI211_X1 U7366 ( .C1(n6732), .C2(n6740), .A(n6737), .B(n6738), .ZN(n6733)
         );
  NAND2_X1 U7367 ( .A1(n6733), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6734) );
  OAI211_X1 U7368 ( .C1(n6736), .C2(n6765), .A(n6735), .B(n6734), .ZN(U3004)
         );
  INV_X1 U7369 ( .A(n6737), .ZN(n6746) );
  OAI22_X1 U7370 ( .A1(n6741), .A2(n6740), .B1(n6739), .B2(n6738), .ZN(n6745)
         );
  OAI21_X1 U7371 ( .B1(n6743), .B2(n7342), .A(n6742), .ZN(n6744) );
  AOI211_X1 U7372 ( .C1(n6746), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6745), .B(n6744), .ZN(n6747) );
  OAI21_X1 U7373 ( .B1(n6748), .B2(n6765), .A(n6747), .ZN(U3005) );
  AOI21_X1 U7374 ( .B1(n6750), .B2(n6749), .A(n3722), .ZN(n7411) );
  NOR3_X1 U7375 ( .A1(n6760), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n6752), 
        .ZN(n6756) );
  INV_X1 U7376 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7416) );
  AOI21_X1 U7377 ( .B1(n6752), .B2(n6751), .A(n6763), .ZN(n6754) );
  OAI22_X1 U7378 ( .A1(n6759), .A2(n7416), .B1(n6754), .B2(n6753), .ZN(n6755)
         );
  AOI211_X1 U7379 ( .C1(n7411), .C2(n7332), .A(n6756), .B(n6755), .ZN(n6757)
         );
  OAI21_X1 U7380 ( .B1(n6758), .B2(n6765), .A(n6757), .ZN(U3006) );
  NOR2_X1 U7381 ( .A1(n7399), .A2(n7342), .ZN(n6762) );
  INV_X1 U7382 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7215) );
  OAI22_X1 U7383 ( .A1(n6760), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .B1(n7215), .B2(n6759), .ZN(n6761) );
  AOI211_X1 U7384 ( .C1(n6763), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6762), .B(n6761), .ZN(n6764) );
  OAI21_X1 U7385 ( .B1(n6766), .B2(n6765), .A(n6764), .ZN(U3007) );
  INV_X1 U7386 ( .A(n6767), .ZN(n6769) );
  OAI22_X1 U7387 ( .A1(n6769), .A2(n7486), .B1(n6768), .B2(n7543), .ZN(n6770)
         );
  MUX2_X1 U7388 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6770), .S(n7491), 
        .Z(U3456) );
  XNOR2_X1 U7389 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n6772) );
  XNOR2_X1 U7390 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .ZN(n6771) );
  NAND2_X1 U7391 ( .A1(n6772), .A2(n6771), .ZN(n6844) );
  INV_X1 U7392 ( .A(n6844), .ZN(n6849) );
  XOR2_X1 U7393 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n6848) );
  XOR2_X1 U7394 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .Z(n6847) );
  XOR2_X1 U7395 ( .A(DATAI_31_), .B(keyinput_0), .Z(n6775) );
  XOR2_X1 U7396 ( .A(DATAI_30_), .B(keyinput_1), .Z(n6774) );
  XNOR2_X1 U7397 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n6773) );
  AOI21_X1 U7398 ( .B1(n6775), .B2(n6774), .A(n6773), .ZN(n6778) );
  XOR2_X1 U7399 ( .A(DATAI_28_), .B(keyinput_3), .Z(n6777) );
  XNOR2_X1 U7400 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n6776) );
  NOR3_X1 U7401 ( .A1(n6778), .A2(n6777), .A3(n6776), .ZN(n6781) );
  XOR2_X1 U7402 ( .A(DATAI_26_), .B(keyinput_5), .Z(n6780) );
  XOR2_X1 U7403 ( .A(DATAI_25_), .B(keyinput_6), .Z(n6779) );
  OAI21_X1 U7404 ( .B1(n6781), .B2(n6780), .A(n6779), .ZN(n6785) );
  XOR2_X1 U7405 ( .A(DATAI_22_), .B(keyinput_9), .Z(n6784) );
  XNOR2_X1 U7406 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n6783) );
  XNOR2_X1 U7407 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n6782) );
  NAND4_X1 U7408 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6788)
         );
  XOR2_X1 U7409 ( .A(DATAI_20_), .B(keyinput_11), .Z(n6787) );
  XNOR2_X1 U7410 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n6786) );
  NAND3_X1 U7411 ( .A1(n6788), .A2(n6787), .A3(n6786), .ZN(n6791) );
  XNOR2_X1 U7412 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n6790) );
  XOR2_X1 U7413 ( .A(DATAI_18_), .B(keyinput_13), .Z(n6789) );
  AOI21_X1 U7414 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6795) );
  XNOR2_X1 U7415 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n6794) );
  XOR2_X1 U7416 ( .A(DATAI_16_), .B(keyinput_15), .Z(n6793) );
  XNOR2_X1 U7417 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n6792) );
  OAI211_X1 U7418 ( .C1(n6795), .C2(n6794), .A(n6793), .B(n6792), .ZN(n6798)
         );
  XNOR2_X1 U7419 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n6797) );
  XOR2_X1 U7420 ( .A(DATAI_13_), .B(keyinput_18), .Z(n6796) );
  AOI21_X1 U7421 ( .B1(n6798), .B2(n6797), .A(n6796), .ZN(n6802) );
  XNOR2_X1 U7422 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n6801) );
  XOR2_X1 U7423 ( .A(DATAI_10_), .B(keyinput_21), .Z(n6800) );
  XNOR2_X1 U7424 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n6799) );
  OAI211_X1 U7425 ( .C1(n6802), .C2(n6801), .A(n6800), .B(n6799), .ZN(n6805)
         );
  XOR2_X1 U7426 ( .A(DATAI_9_), .B(keyinput_22), .Z(n6804) );
  XOR2_X1 U7427 ( .A(DATAI_8_), .B(keyinput_23), .Z(n6803) );
  NAND3_X1 U7428 ( .A1(n6805), .A2(n6804), .A3(n6803), .ZN(n6808) );
  XOR2_X1 U7429 ( .A(DATAI_6_), .B(keyinput_25), .Z(n6807) );
  XOR2_X1 U7430 ( .A(DATAI_7_), .B(keyinput_24), .Z(n6806) );
  NAND3_X1 U7431 ( .A1(n6808), .A2(n6807), .A3(n6806), .ZN(n6811) );
  XNOR2_X1 U7432 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n6810) );
  XNOR2_X1 U7433 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n6809) );
  AOI21_X1 U7434 ( .B1(n6811), .B2(n6810), .A(n6809), .ZN(n6814) );
  XOR2_X1 U7435 ( .A(DATAI_3_), .B(keyinput_28), .Z(n6813) );
  XNOR2_X1 U7436 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n6812) );
  NOR3_X1 U7437 ( .A1(n6814), .A2(n6813), .A3(n6812), .ZN(n6828) );
  XOR2_X1 U7438 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_37), .Z(n6818) );
  XOR2_X1 U7439 ( .A(BS16_N), .B(keyinput_34), .Z(n6817) );
  XOR2_X1 U7440 ( .A(NA_N), .B(keyinput_33), .Z(n6816) );
  XOR2_X1 U7441 ( .A(HOLD), .B(keyinput_36), .Z(n6815) );
  NOR4_X1 U7442 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6825)
         );
  XOR2_X1 U7443 ( .A(DATAI_1_), .B(keyinput_30), .Z(n6824) );
  XOR2_X1 U7444 ( .A(DATAI_0_), .B(keyinput_31), .Z(n6821) );
  XOR2_X1 U7445 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_38), .Z(n6820) );
  XNOR2_X1 U7446 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_32), .ZN(n6819) );
  NOR3_X1 U7447 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(n6823) );
  XNOR2_X1 U7448 ( .A(READY_N), .B(keyinput_35), .ZN(n6822) );
  NAND4_X1 U7449 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .ZN(n6827)
         );
  INV_X1 U7450 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n7296) );
  XNOR2_X1 U7451 ( .A(n7296), .B(keyinput_39), .ZN(n6826) );
  OAI21_X1 U7452 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n6831) );
  INV_X1 U7453 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7567) );
  XNOR2_X1 U7454 ( .A(n7567), .B(keyinput_40), .ZN(n6830) );
  XNOR2_X1 U7455 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n6829) );
  AOI21_X1 U7456 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(n6834) );
  XOR2_X1 U7457 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_42), .Z(n6833)
         );
  XNOR2_X1 U7458 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_43), .ZN(n6832) );
  NOR3_X1 U7459 ( .A1(n6834), .A2(n6833), .A3(n6832), .ZN(n6838) );
  XOR2_X1 U7460 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_45), .Z(n6837) );
  XOR2_X1 U7461 ( .A(MORE_REG_SCAN_IN), .B(keyinput_44), .Z(n6836) );
  XNOR2_X1 U7462 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_46), .ZN(n6835) );
  NOR4_X1 U7463 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n6842)
         );
  XOR2_X1 U7464 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_47), .Z(n6841) );
  XNOR2_X1 U7465 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_49), .ZN(n6840)
         );
  XNOR2_X1 U7466 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_48), .ZN(n6839)
         );
  NOR4_X1 U7467 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6845)
         );
  XNOR2_X1 U7468 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_50), .ZN(n6843)
         );
  NOR3_X1 U7469 ( .A1(n6845), .A2(n6844), .A3(n6843), .ZN(n6846) );
  AOI211_X1 U7470 ( .C1(n6849), .C2(n6848), .A(n6847), .B(n6846), .ZN(n6852)
         );
  XNOR2_X1 U7471 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .ZN(n6851) );
  XNOR2_X1 U7472 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n6850) );
  NOR3_X1 U7473 ( .A1(n6852), .A2(n6851), .A3(n6850), .ZN(n6854) );
  XOR2_X1 U7474 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .Z(n6853) );
  NOR2_X1 U7475 ( .A1(n6854), .A2(n6853), .ZN(n6862) );
  INV_X1 U7476 ( .A(keyinput_59), .ZN(n6855) );
  XNOR2_X1 U7477 ( .A(n6855), .B(REIP_REG_23__SCAN_IN), .ZN(n6859) );
  XNOR2_X1 U7478 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n6858) );
  XNOR2_X1 U7479 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .ZN(n6857) );
  XNOR2_X1 U7480 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n6856) );
  NAND4_X1 U7481 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n6861)
         );
  XNOR2_X1 U7482 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n6860) );
  OAI21_X1 U7483 ( .B1(n6862), .B2(n6861), .A(n6860), .ZN(n6865) );
  XOR2_X1 U7484 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .Z(n6864) );
  XNOR2_X1 U7485 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .ZN(n6863) );
  AOI21_X1 U7486 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6868) );
  XNOR2_X1 U7487 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_65), .ZN(n6867) );
  XOR2_X1 U7488 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n6866) );
  OAI21_X1 U7489 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6872) );
  INV_X1 U7490 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7253) );
  XNOR2_X1 U7491 ( .A(n7253), .B(keyinput_67), .ZN(n6871) );
  INV_X1 U7492 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7266) );
  XNOR2_X1 U7493 ( .A(n7266), .B(keyinput_68), .ZN(n6870) );
  XNOR2_X1 U7494 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_69), .ZN(n6869) );
  AOI211_X1 U7495 ( .C1(n6872), .C2(n6871), .A(n6870), .B(n6869), .ZN(n6876)
         );
  INV_X1 U7496 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7274) );
  XNOR2_X1 U7497 ( .A(n7274), .B(keyinput_70), .ZN(n6875) );
  INV_X1 U7498 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7247) );
  XNOR2_X1 U7499 ( .A(n7247), .B(keyinput_72), .ZN(n6874) );
  XNOR2_X1 U7500 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_71), .ZN(n6873) );
  OAI211_X1 U7501 ( .C1(n6876), .C2(n6875), .A(n6874), .B(n6873), .ZN(n6879)
         );
  INV_X1 U7502 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7243) );
  XNOR2_X1 U7503 ( .A(n7243), .B(keyinput_74), .ZN(n6878) );
  XNOR2_X1 U7504 ( .A(ADDRESS_REG_27__SCAN_IN), .B(keyinput_73), .ZN(n6877) );
  NAND3_X1 U7505 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(n6882) );
  XNOR2_X1 U7506 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_76), .ZN(n6881) );
  XNOR2_X1 U7507 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_75), .ZN(n6880) );
  NAND3_X1 U7508 ( .A1(n6882), .A2(n6881), .A3(n6880), .ZN(n6885) );
  XNOR2_X1 U7509 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_77), .ZN(n6884) );
  XNOR2_X1 U7510 ( .A(ADDRESS_REG_22__SCAN_IN), .B(keyinput_78), .ZN(n6883) );
  AOI21_X1 U7511 ( .B1(n6885), .B2(n6884), .A(n6883), .ZN(n6888) );
  XNOR2_X1 U7512 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_79), .ZN(n6887) );
  XNOR2_X1 U7513 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_80), .ZN(n6886) );
  OAI21_X1 U7514 ( .B1(n6888), .B2(n6887), .A(n6886), .ZN(n6891) );
  INV_X1 U7515 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7229) );
  XNOR2_X1 U7516 ( .A(n7229), .B(keyinput_81), .ZN(n6890) );
  XNOR2_X1 U7517 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_82), .ZN(n6889) );
  NAND3_X1 U7518 ( .A1(n6891), .A2(n6890), .A3(n6889), .ZN(n6894) );
  XNOR2_X1 U7519 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_83), .ZN(n6893) );
  XNOR2_X1 U7520 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_84), .ZN(n6892) );
  NAND3_X1 U7521 ( .A1(n6894), .A2(n6893), .A3(n6892), .ZN(n6901) );
  XNOR2_X1 U7522 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_85), .ZN(n6900) );
  XOR2_X1 U7523 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_89), .Z(n6898) );
  XOR2_X1 U7524 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_88), .Z(n6897) );
  XOR2_X1 U7525 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_86), .Z(n6896) );
  XOR2_X1 U7526 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_87), .Z(n6895) );
  NAND4_X1 U7527 ( .A1(n6898), .A2(n6897), .A3(n6896), .A4(n6895), .ZN(n6899)
         );
  AOI21_X1 U7528 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(n6905) );
  INV_X1 U7529 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7214) );
  XNOR2_X1 U7530 ( .A(n7214), .B(keyinput_90), .ZN(n6904) );
  INV_X1 U7531 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7212) );
  XNOR2_X1 U7532 ( .A(n7212), .B(keyinput_91), .ZN(n6903) );
  INV_X1 U7533 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7211) );
  XNOR2_X1 U7534 ( .A(n7211), .B(keyinput_92), .ZN(n6902) );
  NOR4_X1 U7535 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6908)
         );
  INV_X1 U7536 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7208) );
  XNOR2_X1 U7537 ( .A(n7208), .B(keyinput_93), .ZN(n6907) );
  INV_X1 U7538 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7207) );
  XNOR2_X1 U7539 ( .A(n7207), .B(keyinput_94), .ZN(n6906) );
  NOR3_X1 U7540 ( .A1(n6908), .A2(n6907), .A3(n6906), .ZN(n6911) );
  INV_X1 U7541 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7205) );
  XNOR2_X1 U7542 ( .A(n7205), .B(keyinput_96), .ZN(n6910) );
  XNOR2_X1 U7543 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n6909) );
  NOR3_X1 U7544 ( .A1(n6911), .A2(n6910), .A3(n6909), .ZN(n6915) );
  INV_X1 U7545 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7200) );
  XNOR2_X1 U7546 ( .A(n7200), .B(keyinput_99), .ZN(n6914) );
  INV_X1 U7547 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7202) );
  XNOR2_X1 U7548 ( .A(n7202), .B(keyinput_98), .ZN(n6913) );
  XNOR2_X1 U7549 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_97), .ZN(n6912) );
  NOR4_X1 U7550 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(n6920)
         );
  INV_X1 U7551 ( .A(keyinput_101), .ZN(n6916) );
  XNOR2_X1 U7552 ( .A(n6916), .B(STATE_REG_2__SCAN_IN), .ZN(n6919) );
  XNOR2_X1 U7553 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .ZN(n6918) );
  XNOR2_X1 U7554 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_100), .ZN(n6917) );
  NOR4_X1 U7555 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6923)
         );
  XNOR2_X1 U7556 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .ZN(n6922) );
  XNOR2_X1 U7557 ( .A(n7103), .B(keyinput_104), .ZN(n6921) );
  OAI21_X1 U7558 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(n6929) );
  XOR2_X1 U7559 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .Z(n6925) );
  XNOR2_X1 U7560 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_106), .ZN(n6924)
         );
  NOR2_X1 U7561 ( .A1(n6925), .A2(n6924), .ZN(n6928) );
  INV_X1 U7562 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7153) );
  XNOR2_X1 U7563 ( .A(n7153), .B(keyinput_107), .ZN(n6927) );
  XNOR2_X1 U7564 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_108), .ZN(n6926)
         );
  AOI211_X1 U7565 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n6926), .ZN(n6932)
         );
  INV_X1 U7566 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7154) );
  XNOR2_X1 U7567 ( .A(n7154), .B(keyinput_109), .ZN(n6931) );
  INV_X1 U7568 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7155) );
  XNOR2_X1 U7569 ( .A(n7155), .B(keyinput_110), .ZN(n6930) );
  OAI21_X1 U7570 ( .B1(n6932), .B2(n6931), .A(n6930), .ZN(n6936) );
  XNOR2_X1 U7571 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_111), .ZN(n6935)
         );
  INV_X1 U7572 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7158) );
  XNOR2_X1 U7573 ( .A(n7158), .B(keyinput_113), .ZN(n6934) );
  INV_X1 U7574 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7157) );
  XNOR2_X1 U7575 ( .A(n7157), .B(keyinput_112), .ZN(n6933) );
  AOI211_X1 U7576 ( .C1(n6936), .C2(n6935), .A(n6934), .B(n6933), .ZN(n6939)
         );
  INV_X1 U7577 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7160) );
  XNOR2_X1 U7578 ( .A(n7160), .B(keyinput_115), .ZN(n6938) );
  XNOR2_X1 U7579 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_114), .ZN(n6937)
         );
  NOR3_X1 U7580 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(n6942) );
  INV_X1 U7581 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7161) );
  XNOR2_X1 U7582 ( .A(n7161), .B(keyinput_116), .ZN(n6941) );
  INV_X1 U7583 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7162) );
  XNOR2_X1 U7584 ( .A(n7162), .B(keyinput_117), .ZN(n6940) );
  OAI21_X1 U7585 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(n6945) );
  INV_X1 U7586 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7163) );
  XNOR2_X1 U7587 ( .A(n7163), .B(keyinput_118), .ZN(n6944) );
  INV_X1 U7588 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7164) );
  XNOR2_X1 U7589 ( .A(n7164), .B(keyinput_119), .ZN(n6943) );
  AOI21_X1 U7590 ( .B1(n6945), .B2(n6944), .A(n6943), .ZN(n6949) );
  INV_X1 U7591 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7165) );
  XNOR2_X1 U7592 ( .A(n7165), .B(keyinput_120), .ZN(n6948) );
  INV_X1 U7593 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7167) );
  XNOR2_X1 U7594 ( .A(n7167), .B(keyinput_122), .ZN(n6947) );
  XNOR2_X1 U7595 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_121), .ZN(n6946)
         );
  OAI211_X1 U7596 ( .C1(n6949), .C2(n6948), .A(n6947), .B(n6946), .ZN(n6952)
         );
  INV_X1 U7597 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7168) );
  XNOR2_X1 U7598 ( .A(n7168), .B(keyinput_123), .ZN(n6951) );
  INV_X1 U7599 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7169) );
  XNOR2_X1 U7600 ( .A(n7169), .B(keyinput_124), .ZN(n6950) );
  NAND3_X1 U7601 ( .A1(n6952), .A2(n6951), .A3(n6950), .ZN(n6955) );
  XOR2_X1 U7602 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .Z(n6954)
         );
  XOR2_X1 U7603 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_126), .Z(n6953)
         );
  NAND3_X1 U7604 ( .A1(n6955), .A2(n6954), .A3(n6953), .ZN(n7142) );
  XNOR2_X1 U7605 ( .A(keyinput_255), .B(keyinput_127), .ZN(n7141) );
  XOR2_X1 U7606 ( .A(DATAI_31_), .B(keyinput_128), .Z(n6958) );
  XOR2_X1 U7607 ( .A(DATAI_30_), .B(keyinput_129), .Z(n6957) );
  XOR2_X1 U7608 ( .A(DATAI_29_), .B(keyinput_130), .Z(n6956) );
  AOI21_X1 U7609 ( .B1(n6958), .B2(n6957), .A(n6956), .ZN(n6961) );
  XOR2_X1 U7610 ( .A(DATAI_27_), .B(keyinput_132), .Z(n6960) );
  XNOR2_X1 U7611 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n6959) );
  NOR3_X1 U7612 ( .A1(n6961), .A2(n6960), .A3(n6959), .ZN(n6964) );
  XOR2_X1 U7613 ( .A(DATAI_26_), .B(keyinput_133), .Z(n6963) );
  XOR2_X1 U7614 ( .A(DATAI_25_), .B(keyinput_134), .Z(n6962) );
  OAI21_X1 U7615 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6968) );
  XOR2_X1 U7616 ( .A(DATAI_23_), .B(keyinput_136), .Z(n6967) );
  XNOR2_X1 U7617 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n6966) );
  XNOR2_X1 U7618 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n6965) );
  NAND4_X1 U7619 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n6971)
         );
  XOR2_X1 U7620 ( .A(DATAI_20_), .B(keyinput_139), .Z(n6970) );
  XOR2_X1 U7621 ( .A(DATAI_21_), .B(keyinput_138), .Z(n6969) );
  NAND3_X1 U7622 ( .A1(n6971), .A2(n6970), .A3(n6969), .ZN(n6974) );
  XNOR2_X1 U7623 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n6973) );
  XNOR2_X1 U7624 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n6972) );
  AOI21_X1 U7625 ( .B1(n6974), .B2(n6973), .A(n6972), .ZN(n6978) );
  XNOR2_X1 U7626 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n6977) );
  XOR2_X1 U7627 ( .A(DATAI_15_), .B(keyinput_144), .Z(n6976) );
  XOR2_X1 U7628 ( .A(DATAI_16_), .B(keyinput_143), .Z(n6975) );
  OAI211_X1 U7629 ( .C1(n6978), .C2(n6977), .A(n6976), .B(n6975), .ZN(n6981)
         );
  XNOR2_X1 U7630 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n6980) );
  XNOR2_X1 U7631 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n6979) );
  AOI21_X1 U7632 ( .B1(n6981), .B2(n6980), .A(n6979), .ZN(n6985) );
  XNOR2_X1 U7633 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n6984) );
  XOR2_X1 U7634 ( .A(DATAI_10_), .B(keyinput_149), .Z(n6983) );
  XNOR2_X1 U7635 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n6982) );
  OAI211_X1 U7636 ( .C1(n6985), .C2(n6984), .A(n6983), .B(n6982), .ZN(n6988)
         );
  XOR2_X1 U7637 ( .A(DATAI_9_), .B(keyinput_150), .Z(n6987) );
  XOR2_X1 U7638 ( .A(DATAI_8_), .B(keyinput_151), .Z(n6986) );
  NAND3_X1 U7639 ( .A1(n6988), .A2(n6987), .A3(n6986), .ZN(n6991) );
  XNOR2_X1 U7640 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n6990) );
  XNOR2_X1 U7641 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n6989) );
  NAND3_X1 U7642 ( .A1(n6991), .A2(n6990), .A3(n6989), .ZN(n6994) );
  XNOR2_X1 U7643 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n6993) );
  XOR2_X1 U7644 ( .A(DATAI_4_), .B(keyinput_155), .Z(n6992) );
  AOI21_X1 U7645 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n6997) );
  XOR2_X1 U7646 ( .A(DATAI_3_), .B(keyinput_156), .Z(n6996) );
  XOR2_X1 U7647 ( .A(DATAI_2_), .B(keyinput_157), .Z(n6995) );
  NOR3_X1 U7648 ( .A1(n6997), .A2(n6996), .A3(n6995), .ZN(n7011) );
  XOR2_X1 U7649 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .Z(n7001) );
  XOR2_X1 U7650 ( .A(DATAI_0_), .B(keyinput_159), .Z(n7000) );
  XOR2_X1 U7651 ( .A(DATAI_1_), .B(keyinput_158), .Z(n6999) );
  XNOR2_X1 U7652 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_166), .ZN(n6998) );
  NOR4_X1 U7653 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7008)
         );
  XOR2_X1 U7654 ( .A(HOLD), .B(keyinput_164), .Z(n7007) );
  XOR2_X1 U7655 ( .A(NA_N), .B(keyinput_161), .Z(n7006) );
  XOR2_X1 U7656 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .Z(n7004) );
  XNOR2_X1 U7657 ( .A(n7516), .B(keyinput_163), .ZN(n7003) );
  XNOR2_X1 U7658 ( .A(BS16_N), .B(keyinput_162), .ZN(n7002) );
  NOR3_X1 U7659 ( .A1(n7004), .A2(n7003), .A3(n7002), .ZN(n7005) );
  NAND4_X1 U7660 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), .ZN(n7010)
         );
  XNOR2_X1 U7661 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_167), .ZN(n7009) );
  OAI21_X1 U7662 ( .B1(n7011), .B2(n7010), .A(n7009), .ZN(n7014) );
  XNOR2_X1 U7663 ( .A(n7567), .B(keyinput_168), .ZN(n7013) );
  INV_X1 U7664 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7300) );
  XNOR2_X1 U7665 ( .A(n7300), .B(keyinput_169), .ZN(n7012) );
  AOI21_X1 U7666 ( .B1(n7014), .B2(n7013), .A(n7012), .ZN(n7017) );
  XOR2_X1 U7667 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .Z(n7016)
         );
  XNOR2_X1 U7668 ( .A(n7303), .B(keyinput_171), .ZN(n7015) );
  NOR3_X1 U7669 ( .A1(n7017), .A2(n7016), .A3(n7015), .ZN(n7021) );
  XOR2_X1 U7670 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .Z(n7020) );
  XNOR2_X1 U7671 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .ZN(n7019) );
  XNOR2_X1 U7672 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .ZN(n7018) );
  NOR4_X1 U7673 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7025)
         );
  XOR2_X1 U7674 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_177), .Z(n7024)
         );
  XNOR2_X1 U7675 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_176), .ZN(n7023)
         );
  XNOR2_X1 U7676 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_175), .ZN(n7022)
         );
  NOR4_X1 U7677 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(n7028)
         );
  INV_X1 U7678 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7254) );
  XNOR2_X1 U7679 ( .A(n7254), .B(keyinput_178), .ZN(n7027) );
  XNOR2_X1 U7680 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n7026) );
  OAI21_X1 U7681 ( .B1(n7028), .B2(n7027), .A(n7026), .ZN(n7031) );
  XOR2_X1 U7682 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .Z(n7030) );
  XNOR2_X1 U7683 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .ZN(n7029) );
  NAND3_X1 U7684 ( .A1(n7031), .A2(n7030), .A3(n7029), .ZN(n7035) );
  XNOR2_X1 U7685 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .ZN(n7034) );
  XNOR2_X1 U7686 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .ZN(n7033) );
  XNOR2_X1 U7687 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n7032) );
  AOI211_X1 U7688 ( .C1(n7035), .C2(n7034), .A(n7033), .B(n7032), .ZN(n7042)
         );
  XOR2_X1 U7689 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .Z(n7041) );
  XOR2_X1 U7690 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .Z(n7039) );
  XOR2_X1 U7691 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .Z(n7038) );
  XNOR2_X1 U7692 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n7037) );
  XNOR2_X1 U7693 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .ZN(n7036) );
  NOR4_X1 U7694 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7040)
         );
  OAI21_X1 U7695 ( .B1(n7042), .B2(n7041), .A(n7040), .ZN(n7045) );
  XOR2_X1 U7696 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .Z(n7044) );
  XOR2_X1 U7697 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n7043) );
  AOI21_X1 U7698 ( .B1(n7045), .B2(n7044), .A(n7043), .ZN(n7048) );
  XOR2_X1 U7699 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .Z(n7047) );
  XNOR2_X1 U7700 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .ZN(n7046) );
  OAI21_X1 U7701 ( .B1(n7048), .B2(n7047), .A(n7046), .ZN(n7051) );
  XOR2_X1 U7702 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .Z(n7050) );
  XNOR2_X1 U7703 ( .A(n7253), .B(keyinput_195), .ZN(n7049) );
  AOI21_X1 U7704 ( .B1(n7051), .B2(n7050), .A(n7049), .ZN(n7054) );
  XNOR2_X1 U7705 ( .A(n7266), .B(keyinput_196), .ZN(n7053) );
  XNOR2_X1 U7706 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_197), .ZN(n7052) );
  NOR3_X1 U7707 ( .A1(n7054), .A2(n7053), .A3(n7052), .ZN(n7058) );
  XNOR2_X1 U7708 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_198), .ZN(n7057) );
  INV_X1 U7709 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7250) );
  XNOR2_X1 U7710 ( .A(n7250), .B(keyinput_199), .ZN(n7056) );
  XNOR2_X1 U7711 ( .A(ADDRESS_REG_28__SCAN_IN), .B(keyinput_200), .ZN(n7055)
         );
  OAI211_X1 U7712 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n7055), .ZN(n7061)
         );
  XNOR2_X1 U7713 ( .A(ADDRESS_REG_27__SCAN_IN), .B(keyinput_201), .ZN(n7060)
         );
  XNOR2_X1 U7714 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_202), .ZN(n7059)
         );
  NAND3_X1 U7715 ( .A1(n7061), .A2(n7060), .A3(n7059), .ZN(n7064) );
  INV_X1 U7716 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7238) );
  XNOR2_X1 U7717 ( .A(n7238), .B(keyinput_204), .ZN(n7063) );
  XNOR2_X1 U7718 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_203), .ZN(n7062)
         );
  NAND3_X1 U7719 ( .A1(n7064), .A2(n7063), .A3(n7062), .ZN(n7067) );
  XNOR2_X1 U7720 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_205), .ZN(n7066)
         );
  INV_X1 U7721 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7235) );
  XNOR2_X1 U7722 ( .A(n7235), .B(keyinput_206), .ZN(n7065) );
  AOI21_X1 U7723 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7070) );
  INV_X1 U7724 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7233) );
  XNOR2_X1 U7725 ( .A(n7233), .B(keyinput_207), .ZN(n7069) );
  XNOR2_X1 U7726 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_208), .ZN(n7068)
         );
  OAI21_X1 U7727 ( .B1(n7070), .B2(n7069), .A(n7068), .ZN(n7073) );
  XNOR2_X1 U7728 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_210), .ZN(n7072)
         );
  XNOR2_X1 U7729 ( .A(ADDRESS_REG_19__SCAN_IN), .B(keyinput_209), .ZN(n7071)
         );
  NAND3_X1 U7730 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7076) );
  XNOR2_X1 U7731 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_211), .ZN(n7075)
         );
  XNOR2_X1 U7732 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_212), .ZN(n7074)
         );
  NAND3_X1 U7733 ( .A1(n7076), .A2(n7075), .A3(n7074), .ZN(n7083) );
  XNOR2_X1 U7734 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_213), .ZN(n7082)
         );
  XOR2_X1 U7735 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_217), .Z(n7080) );
  XOR2_X1 U7736 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_215), .Z(n7079) );
  XOR2_X1 U7737 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_214), .Z(n7078) );
  XOR2_X1 U7738 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .Z(n7077) );
  NAND4_X1 U7739 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(n7081)
         );
  AOI21_X1 U7740 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7087) );
  XNOR2_X1 U7741 ( .A(n7211), .B(keyinput_220), .ZN(n7086) );
  XNOR2_X1 U7742 ( .A(n7214), .B(keyinput_218), .ZN(n7085) );
  XNOR2_X1 U7743 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n7084) );
  NOR4_X1 U7744 ( .A1(n7087), .A2(n7086), .A3(n7085), .A4(n7084), .ZN(n7090)
         );
  XNOR2_X1 U7745 ( .A(n7208), .B(keyinput_221), .ZN(n7089) );
  XNOR2_X1 U7746 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_222), .ZN(n7088) );
  NOR3_X1 U7747 ( .A1(n7090), .A2(n7089), .A3(n7088), .ZN(n7093) );
  INV_X1 U7748 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7206) );
  XNOR2_X1 U7749 ( .A(n7206), .B(keyinput_223), .ZN(n7092) );
  XNOR2_X1 U7750 ( .A(n7205), .B(keyinput_224), .ZN(n7091) );
  NOR3_X1 U7751 ( .A1(n7093), .A2(n7092), .A3(n7091), .ZN(n7097) );
  INV_X1 U7752 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7204) );
  XNOR2_X1 U7753 ( .A(n7204), .B(keyinput_225), .ZN(n7096) );
  XNOR2_X1 U7754 ( .A(n7202), .B(keyinput_226), .ZN(n7095) );
  XNOR2_X1 U7755 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_227), .ZN(n7094) );
  NOR4_X1 U7756 ( .A1(n7097), .A2(n7096), .A3(n7095), .A4(n7094), .ZN(n7102)
         );
  XNOR2_X1 U7757 ( .A(n7098), .B(keyinput_230), .ZN(n7101) );
  XOR2_X1 U7758 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_229), .Z(n7100) );
  XNOR2_X1 U7759 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_228), .ZN(n7099) );
  NOR4_X1 U7760 ( .A1(n7102), .A2(n7101), .A3(n7100), .A4(n7099), .ZN(n7106)
         );
  XNOR2_X1 U7761 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_231), .ZN(n7105) );
  XNOR2_X1 U7762 ( .A(n7103), .B(keyinput_232), .ZN(n7104) );
  OAI21_X1 U7763 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7109) );
  XOR2_X1 U7764 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_234), .Z(n7108) );
  XNOR2_X1 U7765 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .ZN(n7107)
         );
  NAND3_X1 U7766 ( .A1(n7109), .A2(n7108), .A3(n7107), .ZN(n7112) );
  XNOR2_X1 U7767 ( .A(n7153), .B(keyinput_235), .ZN(n7111) );
  XOR2_X1 U7768 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_236), .Z(n7110) );
  NAND3_X1 U7769 ( .A1(n7112), .A2(n7111), .A3(n7110), .ZN(n7115) );
  XNOR2_X1 U7770 ( .A(n7154), .B(keyinput_237), .ZN(n7114) );
  XNOR2_X1 U7771 ( .A(DATAWIDTH_REG_6__SCAN_IN), .B(keyinput_238), .ZN(n7113)
         );
  AOI21_X1 U7772 ( .B1(n7115), .B2(n7114), .A(n7113), .ZN(n7119) );
  XNOR2_X1 U7773 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_239), .ZN(n7118)
         );
  XNOR2_X1 U7774 ( .A(n7158), .B(keyinput_241), .ZN(n7117) );
  XNOR2_X1 U7775 ( .A(n7157), .B(keyinput_240), .ZN(n7116) );
  OAI211_X1 U7776 ( .C1(n7119), .C2(n7118), .A(n7117), .B(n7116), .ZN(n7122)
         );
  XNOR2_X1 U7777 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_242), .ZN(n7121)
         );
  XNOR2_X1 U7778 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_243), .ZN(n7120)
         );
  NAND3_X1 U7779 ( .A1(n7122), .A2(n7121), .A3(n7120), .ZN(n7125) );
  XNOR2_X1 U7780 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_244), .ZN(n7124)
         );
  XNOR2_X1 U7781 ( .A(n7162), .B(keyinput_245), .ZN(n7123) );
  AOI21_X1 U7782 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7128) );
  XNOR2_X1 U7783 ( .A(n7163), .B(keyinput_246), .ZN(n7127) );
  XNOR2_X1 U7784 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_247), .ZN(n7126)
         );
  OAI21_X1 U7785 ( .B1(n7128), .B2(n7127), .A(n7126), .ZN(n7132) );
  XNOR2_X1 U7786 ( .A(n7165), .B(keyinput_248), .ZN(n7131) );
  INV_X1 U7787 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7166) );
  XNOR2_X1 U7788 ( .A(n7166), .B(keyinput_249), .ZN(n7130) );
  XNOR2_X1 U7789 ( .A(n7167), .B(keyinput_250), .ZN(n7129) );
  AOI211_X1 U7790 ( .C1(n7132), .C2(n7131), .A(n7130), .B(n7129), .ZN(n7135)
         );
  XNOR2_X1 U7791 ( .A(n7168), .B(keyinput_251), .ZN(n7134) );
  XNOR2_X1 U7792 ( .A(n7169), .B(keyinput_252), .ZN(n7133) );
  NOR3_X1 U7793 ( .A1(n7135), .A2(n7134), .A3(n7133), .ZN(n7138) );
  XNOR2_X1 U7794 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_254), .ZN(n7137)
         );
  XNOR2_X1 U7795 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_253), .ZN(n7136)
         );
  NOR3_X1 U7796 ( .A1(n7138), .A2(n7137), .A3(n7136), .ZN(n7140) );
  XOR2_X1 U7797 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .Z(n7139)
         );
  AOI211_X1 U7798 ( .C1(n7142), .C2(n7141), .A(n7140), .B(n7139), .ZN(n7152)
         );
  AOI22_X1 U7799 ( .A1(n7691), .A2(n7145), .B1(n7144), .B2(n7143), .ZN(n7146)
         );
  OAI21_X1 U7800 ( .B1(n7147), .B2(n7674), .A(n7146), .ZN(n7149) );
  NOR2_X1 U7801 ( .A1(n7740), .A2(n7680), .ZN(n7148) );
  AOI211_X1 U7802 ( .C1(INSTQUEUE_REG_0__6__SCAN_IN), .C2(n7150), .A(n7149), 
        .B(n7148), .ZN(n7151) );
  XNOR2_X1 U7803 ( .A(n7152), .B(n7151), .ZN(U3026) );
  AND2_X1 U7804 ( .A1(n7171), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  NOR2_X1 U7805 ( .A1(n7170), .A2(n7153), .ZN(U3179) );
  AND2_X1 U7806 ( .A1(n7171), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  NOR2_X1 U7807 ( .A1(n7170), .A2(n7154), .ZN(U3177) );
  NOR2_X1 U7808 ( .A1(n7170), .A2(n7155), .ZN(U3176) );
  INV_X1 U7809 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7156) );
  NOR2_X1 U7810 ( .A1(n7170), .A2(n7156), .ZN(U3175) );
  NOR2_X1 U7811 ( .A1(n7170), .A2(n7157), .ZN(U3174) );
  NOR2_X1 U7812 ( .A1(n7170), .A2(n7158), .ZN(U3173) );
  INV_X1 U7813 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7159) );
  NOR2_X1 U7814 ( .A1(n7170), .A2(n7159), .ZN(U3172) );
  NOR2_X1 U7815 ( .A1(n7170), .A2(n7160), .ZN(U3171) );
  NOR2_X1 U7816 ( .A1(n7170), .A2(n7161), .ZN(U3170) );
  NOR2_X1 U7817 ( .A1(n7170), .A2(n7162), .ZN(U3169) );
  NOR2_X1 U7818 ( .A1(n7170), .A2(n7163), .ZN(U3168) );
  NOR2_X1 U7819 ( .A1(n7170), .A2(n7164), .ZN(U3167) );
  NOR2_X1 U7820 ( .A1(n7170), .A2(n7165), .ZN(U3166) );
  NOR2_X1 U7821 ( .A1(n7170), .A2(n7166), .ZN(U3165) );
  NOR2_X1 U7822 ( .A1(n7170), .A2(n7167), .ZN(U3164) );
  NOR2_X1 U7823 ( .A1(n7170), .A2(n7168), .ZN(U3163) );
  NOR2_X1 U7824 ( .A1(n7170), .A2(n7169), .ZN(U3162) );
  AND2_X1 U7825 ( .A1(n7171), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7826 ( .A1(n7171), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U7827 ( .A1(n7171), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7828 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7171), .ZN(U3158) );
  AND2_X1 U7829 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7171), .ZN(U3157) );
  AND2_X1 U7830 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7171), .ZN(U3156) );
  AND2_X1 U7831 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7171), .ZN(U3155) );
  AND2_X1 U7832 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7171), .ZN(U3154) );
  AND2_X1 U7833 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7171), .ZN(U3153) );
  AND2_X1 U7834 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7171), .ZN(U3152) );
  AND2_X1 U7835 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7171), .ZN(U3151) );
  AND2_X1 U7836 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n7551), .ZN(U3019)
         );
  AND2_X1 U7837 ( .A1(n7172), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7838 ( .A1(n7182), .A2(LWORD_REG_0__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n7173) );
  OAI21_X1 U7839 ( .B1(n7174), .B2(n7196), .A(n7173), .ZN(U2923) );
  AOI22_X1 U7840 ( .A1(n7182), .A2(LWORD_REG_1__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7175) );
  OAI21_X1 U7841 ( .B1(n4991), .B2(n7196), .A(n7175), .ZN(U2922) );
  AOI22_X1 U7842 ( .A1(n7182), .A2(LWORD_REG_2__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n7176) );
  OAI21_X1 U7843 ( .B1(n5003), .B2(n7196), .A(n7176), .ZN(U2921) );
  AOI22_X1 U7844 ( .A1(n7182), .A2(LWORD_REG_3__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7177) );
  OAI21_X1 U7845 ( .B1(n5033), .B2(n7196), .A(n7177), .ZN(U2920) );
  AOI22_X1 U7846 ( .A1(n7182), .A2(LWORD_REG_4__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7178) );
  OAI21_X1 U7847 ( .B1(n7179), .B2(n7196), .A(n7178), .ZN(U2919) );
  AOI22_X1 U7848 ( .A1(n7182), .A2(LWORD_REG_5__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7180) );
  OAI21_X1 U7849 ( .B1(n7181), .B2(n7196), .A(n7180), .ZN(U2918) );
  AOI22_X1 U7850 ( .A1(n7182), .A2(LWORD_REG_6__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7183) );
  OAI21_X1 U7851 ( .B1(n4864), .B2(n7196), .A(n7183), .ZN(U2917) );
  AOI22_X1 U7852 ( .A1(n7182), .A2(LWORD_REG_7__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7184) );
  OAI21_X1 U7853 ( .B1(n5028), .B2(n7196), .A(n7184), .ZN(U2916) );
  AOI22_X1 U7854 ( .A1(n7182), .A2(LWORD_REG_8__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7185) );
  OAI21_X1 U7855 ( .B1(n5045), .B2(n7196), .A(n7185), .ZN(U2915) );
  AOI22_X1 U7856 ( .A1(n7182), .A2(LWORD_REG_9__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7186) );
  OAI21_X1 U7857 ( .B1(n5018), .B2(n7196), .A(n7186), .ZN(U2914) );
  AOI22_X1 U7858 ( .A1(n7182), .A2(LWORD_REG_10__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7187) );
  OAI21_X1 U7859 ( .B1(n5025), .B2(n7196), .A(n7187), .ZN(U2913) );
  AOI22_X1 U7860 ( .A1(n7182), .A2(LWORD_REG_11__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7188) );
  OAI21_X1 U7861 ( .B1(n5022), .B2(n7196), .A(n7188), .ZN(U2912) );
  AOI22_X1 U7862 ( .A1(n7182), .A2(LWORD_REG_12__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7189) );
  OAI21_X1 U7863 ( .B1(n5039), .B2(n7196), .A(n7189), .ZN(U2911) );
  AOI22_X1 U7864 ( .A1(n7182), .A2(LWORD_REG_13__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7190) );
  OAI21_X1 U7865 ( .B1(n7191), .B2(n7196), .A(n7190), .ZN(U2910) );
  AOI22_X1 U7866 ( .A1(n7182), .A2(LWORD_REG_14__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U7867 ( .B1(n4993), .B2(n7196), .A(n7192), .ZN(U2909) );
  AOI22_X1 U7868 ( .A1(n7182), .A2(LWORD_REG_15__SCAN_IN), .B1(n7193), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7195) );
  OAI21_X1 U7869 ( .B1(n7197), .B2(n7196), .A(n7195), .ZN(U2908) );
  INV_X1 U7870 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7198) );
  OAI222_X1 U7871 ( .A1(n7242), .A2(n7199), .B1(n7198), .B2(n7569), .C1(n7350), 
        .C2(n7252), .ZN(U3184) );
  OAI222_X1 U7872 ( .A1(n7242), .A2(n7201), .B1(n7200), .B2(n7569), .C1(n7199), 
        .C2(n7252), .ZN(U3185) );
  OAI222_X1 U7873 ( .A1(n7242), .A2(n7203), .B1(n7202), .B2(n7569), .C1(n7201), 
        .C2(n7252), .ZN(U3186) );
  OAI222_X1 U7874 ( .A1(n7242), .A2(n7366), .B1(n7204), .B2(n7569), .C1(n7203), 
        .C2(n7252), .ZN(U3187) );
  OAI222_X1 U7875 ( .A1(n7242), .A2(n7387), .B1(n7205), .B2(n7569), .C1(n7366), 
        .C2(n7252), .ZN(U3188) );
  INV_X1 U7876 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7386) );
  OAI222_X1 U7877 ( .A1(n7242), .A2(n7386), .B1(n7206), .B2(n7569), .C1(n7387), 
        .C2(n7252), .ZN(U3189) );
  OAI222_X1 U7878 ( .A1(n7242), .A2(n7209), .B1(n7207), .B2(n7569), .C1(n7386), 
        .C2(n7252), .ZN(U3190) );
  OAI222_X1 U7879 ( .A1(n7252), .A2(n7209), .B1(n7208), .B2(n7569), .C1(n7210), 
        .C2(n7242), .ZN(U3191) );
  OAI222_X1 U7880 ( .A1(n7242), .A2(n7213), .B1(n7211), .B2(n7569), .C1(n7210), 
        .C2(n7252), .ZN(U3192) );
  OAI222_X1 U7881 ( .A1(n7252), .A2(n7213), .B1(n7212), .B2(n7569), .C1(n7215), 
        .C2(n7242), .ZN(U3193) );
  OAI222_X1 U7882 ( .A1(n7252), .A2(n7215), .B1(n7214), .B2(n7569), .C1(n7416), 
        .C2(n7242), .ZN(U3194) );
  INV_X1 U7883 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7217) );
  INV_X1 U7884 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7216) );
  OAI222_X1 U7885 ( .A1(n7242), .A2(n7217), .B1(n7216), .B2(n7569), .C1(n7416), 
        .C2(n7252), .ZN(U3195) );
  INV_X1 U7886 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7218) );
  OAI222_X1 U7887 ( .A1(n7242), .A2(n6523), .B1(n7218), .B2(n7569), .C1(n7217), 
        .C2(n7252), .ZN(U3196) );
  INV_X1 U7888 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7219) );
  OAI222_X1 U7889 ( .A1(n7252), .A2(n6523), .B1(n7219), .B2(n7569), .C1(n7221), 
        .C2(n7242), .ZN(U3197) );
  INV_X1 U7890 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7220) );
  OAI222_X1 U7891 ( .A1(n7252), .A2(n7221), .B1(n7220), .B2(n7569), .C1(n7223), 
        .C2(n7242), .ZN(U3198) );
  INV_X1 U7892 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7222) );
  OAI222_X1 U7893 ( .A1(n7252), .A2(n7223), .B1(n7222), .B2(n7569), .C1(n7433), 
        .C2(n7242), .ZN(U3199) );
  INV_X1 U7894 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7224) );
  INV_X1 U7895 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7226) );
  OAI222_X1 U7896 ( .A1(n7252), .A2(n7433), .B1(n7224), .B2(n7569), .C1(n7226), 
        .C2(n7242), .ZN(U3200) );
  INV_X1 U7897 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7225) );
  OAI222_X1 U7898 ( .A1(n7252), .A2(n7226), .B1(n7225), .B2(n7569), .C1(n7228), 
        .C2(n7242), .ZN(U3201) );
  INV_X1 U7899 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7227) );
  OAI222_X1 U7900 ( .A1(n7252), .A2(n7228), .B1(n7227), .B2(n7569), .C1(n7230), 
        .C2(n7242), .ZN(U3202) );
  OAI222_X1 U7901 ( .A1(n7252), .A2(n7230), .B1(n7229), .B2(n7569), .C1(n7461), 
        .C2(n7242), .ZN(U3203) );
  INV_X1 U7902 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7231) );
  OAI222_X1 U7903 ( .A1(n7252), .A2(n7461), .B1(n7231), .B2(n7569), .C1(n7232), 
        .C2(n7242), .ZN(U3204) );
  INV_X1 U7904 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7234) );
  OAI222_X1 U7905 ( .A1(n7242), .A2(n7234), .B1(n7233), .B2(n7569), .C1(n7232), 
        .C2(n7252), .ZN(U3205) );
  OAI222_X1 U7906 ( .A1(n7242), .A2(n7237), .B1(n7235), .B2(n7569), .C1(n7234), 
        .C2(n7252), .ZN(U3206) );
  INV_X1 U7907 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7236) );
  OAI222_X1 U7908 ( .A1(n7252), .A2(n7237), .B1(n7236), .B2(n7569), .C1(n7239), 
        .C2(n7242), .ZN(U3207) );
  OAI222_X1 U7909 ( .A1(n7252), .A2(n7239), .B1(n7238), .B2(n7569), .C1(n7240), 
        .C2(n7242), .ZN(U3208) );
  INV_X1 U7910 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7241) );
  OAI222_X1 U7911 ( .A1(n7242), .A2(n7244), .B1(n7241), .B2(n7569), .C1(n7240), 
        .C2(n7252), .ZN(U3209) );
  INV_X1 U7912 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7246) );
  OAI222_X1 U7913 ( .A1(n7252), .A2(n7244), .B1(n7243), .B2(n7569), .C1(n7246), 
        .C2(n7242), .ZN(U3210) );
  INV_X1 U7914 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7245) );
  OAI222_X1 U7915 ( .A1(n7252), .A2(n7246), .B1(n7245), .B2(n7569), .C1(n7248), 
        .C2(n7242), .ZN(U3211) );
  OAI222_X1 U7916 ( .A1(n7252), .A2(n7248), .B1(n7247), .B2(n7569), .C1(n7251), 
        .C2(n7242), .ZN(U3212) );
  INV_X1 U7917 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7249) );
  OAI222_X1 U7918 ( .A1(n7252), .A2(n7251), .B1(n7250), .B2(n7569), .C1(n7249), 
        .C2(n7242), .ZN(U3213) );
  AOI22_X1 U7919 ( .A1(n7569), .A2(n7254), .B1(n7253), .B2(n7566), .ZN(U3445)
         );
  AOI221_X1 U7920 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7265) );
  NOR4_X1 U7921 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n7258) );
  NOR4_X1 U7922 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n7257) );
  NOR4_X1 U7923 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(DATAWIDTH_REG_21__SCAN_IN), .ZN(
        n7256) );
  NOR4_X1 U7924 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7255) );
  NAND4_X1 U7925 ( .A1(n7258), .A2(n7257), .A3(n7256), .A4(n7255), .ZN(n7264)
         );
  NOR4_X1 U7926 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7262)
         );
  AOI211_X1 U7927 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_11__SCAN_IN), .B(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n7261) );
  NOR4_X1 U7928 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7260)
         );
  NOR4_X1 U7929 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n7259) );
  NAND4_X1 U7930 ( .A1(n7262), .A2(n7261), .A3(n7260), .A4(n7259), .ZN(n7263)
         );
  NOR2_X1 U7931 ( .A1(n7264), .A2(n7263), .ZN(n7277) );
  MUX2_X1 U7932 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7265), .S(n7277), .Z(
        U2795) );
  INV_X1 U7933 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7269) );
  AOI22_X1 U7934 ( .A1(n7569), .A2(n7269), .B1(n7266), .B2(n7566), .ZN(U3446)
         );
  AOI21_X1 U7935 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7267) );
  OAI221_X1 U7936 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7267), .C1(n7350), .C2(
        REIP_REG_0__SCAN_IN), .A(n7277), .ZN(n7268) );
  OAI21_X1 U7937 ( .B1(n7277), .B2(n7269), .A(n7268), .ZN(U3468) );
  OAI22_X1 U7938 ( .A1(n7566), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n7569), .ZN(n7270) );
  INV_X1 U7939 ( .A(n7270), .ZN(U3447) );
  INV_X1 U7940 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7273) );
  NOR3_X1 U7941 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7271) );
  OAI21_X1 U7942 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7271), .A(n7277), .ZN(n7272)
         );
  OAI21_X1 U7943 ( .B1(n7277), .B2(n7273), .A(n7272), .ZN(U2794) );
  INV_X1 U7944 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7276) );
  AOI22_X1 U7945 ( .A1(n7569), .A2(n7276), .B1(n7274), .B2(n7566), .ZN(U3448)
         );
  OAI21_X1 U7946 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .A(
        n7277), .ZN(n7275) );
  OAI21_X1 U7947 ( .B1(n7277), .B2(n7276), .A(n7275), .ZN(U3469) );
  INV_X1 U7948 ( .A(n7355), .ZN(n7279) );
  AOI22_X1 U7949 ( .A1(n7279), .A2(n7285), .B1(n7284), .B2(n7278), .ZN(n7280)
         );
  OAI21_X1 U7950 ( .B1(n6352), .B2(n7361), .A(n7280), .ZN(U2858) );
  INV_X1 U7951 ( .A(EBX_REG_12__SCAN_IN), .ZN(n7282) );
  AOI22_X1 U7952 ( .A1(n7410), .A2(n7285), .B1(n7284), .B2(n7411), .ZN(n7281)
         );
  OAI21_X1 U7953 ( .B1(n6352), .B2(n7282), .A(n7281), .ZN(U2847) );
  AOI22_X1 U7954 ( .A1(n7286), .A2(n7285), .B1(n7284), .B2(n7283), .ZN(n7287)
         );
  OAI21_X1 U7955 ( .B1(n6352), .B2(n7288), .A(n7287), .ZN(U2844) );
  AOI22_X1 U7956 ( .A1(REIP_REG_17__SCAN_IN), .A2(n7330), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n7289), .ZN(n7293) );
  AOI22_X1 U7957 ( .A1(n7291), .A2(n7290), .B1(n6534), .B2(n7571), .ZN(n7292)
         );
  OAI211_X1 U7958 ( .C1(n7421), .C2(n7294), .A(n7293), .B(n7292), .ZN(U2969)
         );
  NOR2_X1 U7959 ( .A1(n7295), .A2(n7546), .ZN(n7297) );
  OAI22_X1 U7960 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7527), .B1(n7297), .B2(
        n7296), .ZN(U2790) );
  OAI21_X1 U7961 ( .B1(STATE_REG_1__SCAN_IN), .B2(n7562), .A(n7298), .ZN(n7299) );
  AOI22_X1 U7962 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7569), .B1(n7300), .B2(
        n7299), .ZN(U2791) );
  INV_X1 U7963 ( .A(n7301), .ZN(n7302) );
  AOI211_X1 U7964 ( .C1(n7304), .C2(n7303), .A(n7522), .B(n7302), .ZN(n7305)
         );
  OAI21_X1 U7965 ( .B1(n7305), .B2(n3966), .A(n7542), .ZN(n7309) );
  OAI211_X1 U7966 ( .C1(READY_N), .C2(n7517), .A(n7307), .B(n7306), .ZN(n7308)
         );
  MUX2_X1 U7967 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n7309), .S(n7308), .Z(
        U3472) );
  NOR2_X1 U7968 ( .A1(n7310), .A2(n4161), .ZN(n7314) );
  OAI21_X1 U7969 ( .B1(n7342), .B2(n7312), .A(n7311), .ZN(n7313) );
  AOI211_X1 U7970 ( .C1(n7315), .C2(n7344), .A(n7314), .B(n7313), .ZN(n7319)
         );
  OAI211_X1 U7971 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7317), .B(n7316), .ZN(n7318) );
  NAND2_X1 U7972 ( .A1(n7319), .A2(n7318), .ZN(U3014) );
  OAI21_X1 U7973 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n7320), .ZN(n7327) );
  AOI22_X1 U7974 ( .A1(n7321), .A2(n7332), .B1(n7330), .B2(REIP_REG_8__SCAN_IN), .ZN(n7322) );
  OAI21_X1 U7975 ( .B1(n7323), .B2(n4216), .A(n7322), .ZN(n7324) );
  AOI21_X1 U7976 ( .B1(n7325), .B2(n7344), .A(n7324), .ZN(n7326) );
  OAI21_X1 U7977 ( .B1(n7328), .B2(n7327), .A(n7326), .ZN(U3010) );
  AOI22_X1 U7978 ( .A1(REIP_REG_16__SCAN_IN), .A2(n7330), .B1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n7329), .ZN(n7338) );
  AOI22_X1 U7979 ( .A1(n7333), .A2(n7344), .B1(n7332), .B2(n7331), .ZN(n7337)
         );
  OAI221_X1 U7980 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n7335), .C2(n4223), .A(n7334), 
        .ZN(n7336) );
  NAND3_X1 U7981 ( .A1(n7338), .A2(n7337), .A3(n7336), .ZN(U3002) );
  OAI211_X1 U7982 ( .C1(n7342), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7343)
         );
  AOI21_X1 U7983 ( .B1(n7345), .B2(n7344), .A(n7343), .ZN(n7346) );
  OAI221_X1 U7984 ( .B1(n7349), .B2(n7348), .C1(n7349), .C2(n7347), .A(n7346), 
        .ZN(U3018) );
  AOI22_X1 U7985 ( .A1(n7473), .A2(n7351), .B1(n7470), .B2(n7350), .ZN(n7360)
         );
  AOI22_X1 U7986 ( .A1(n7472), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7352), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n7353) );
  OAI21_X1 U7987 ( .B1(n7420), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n7353), 
        .ZN(n7357) );
  NOR2_X1 U7988 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  AOI211_X1 U7989 ( .C1(n7358), .C2(n4054), .A(n7357), .B(n7356), .ZN(n7359)
         );
  OAI211_X1 U7990 ( .C1(n7361), .C2(n7443), .A(n7360), .B(n7359), .ZN(U2826)
         );
  OAI22_X1 U7991 ( .A1(n7363), .A2(n7443), .B1(n7467), .B2(n7362), .ZN(n7364)
         );
  AOI211_X1 U7992 ( .C1(n7472), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n7423), 
        .B(n7364), .ZN(n7373) );
  AND2_X1 U7993 ( .A1(n7375), .A2(n7376), .ZN(n7369) );
  INV_X1 U7994 ( .A(n7365), .ZN(n7367) );
  OAI21_X1 U7995 ( .B1(n7446), .B2(n7367), .A(n7366), .ZN(n7368) );
  AOI22_X1 U7996 ( .A1(n7371), .A2(n7370), .B1(n7369), .B2(n7368), .ZN(n7372)
         );
  OAI211_X1 U7997 ( .C1(n7374), .C2(n7420), .A(n7373), .B(n7372), .ZN(U2822)
         );
  OAI21_X1 U7998 ( .B1(n7387), .B2(n7376), .A(n7375), .ZN(n7385) );
  AOI21_X1 U7999 ( .B1(n7388), .B2(n7387), .A(n7385), .ZN(n7381) );
  AOI22_X1 U8000 ( .A1(EBX_REG_6__SCAN_IN), .A2(n7471), .B1(n7473), .B2(n7377), 
        .ZN(n7378) );
  OAI211_X1 U8001 ( .C1(n7450), .C2(n7379), .A(n7378), .B(n7448), .ZN(n7380)
         );
  AOI211_X1 U8002 ( .C1(n7382), .C2(n7477), .A(n7381), .B(n7380), .ZN(n7383)
         );
  OAI21_X1 U8003 ( .B1(n7384), .B2(n7420), .A(n7383), .ZN(U2821) );
  AOI22_X1 U8004 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7472), .B1(
        EBX_REG_7__SCAN_IN), .B2(n7471), .ZN(n7393) );
  OAI21_X1 U8005 ( .B1(n7386), .B2(n7385), .A(n7448), .ZN(n7390) );
  NOR3_X1 U8006 ( .A1(n7388), .A2(REIP_REG_7__SCAN_IN), .A3(n7387), .ZN(n7389)
         );
  AOI211_X1 U8007 ( .C1(n7391), .C2(n7473), .A(n7390), .B(n7389), .ZN(n7392)
         );
  OAI211_X1 U8008 ( .C1(n7394), .C2(n7437), .A(n7393), .B(n7392), .ZN(n7395)
         );
  INV_X1 U8009 ( .A(n7395), .ZN(n7396) );
  OAI21_X1 U8010 ( .B1(n7397), .B2(n7420), .A(n7396), .ZN(U2820) );
  AOI22_X1 U8011 ( .A1(EBX_REG_11__SCAN_IN), .A2(n7471), .B1(
        REIP_REG_11__SCAN_IN), .B2(n7415), .ZN(n7398) );
  OAI21_X1 U8012 ( .B1(n7467), .B2(n7399), .A(n7398), .ZN(n7400) );
  AOI211_X1 U8013 ( .C1(n7472), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7423), 
        .B(n7400), .ZN(n7405) );
  OAI22_X1 U8014 ( .A1(n7402), .A2(n7437), .B1(n7420), .B2(n7401), .ZN(n7403)
         );
  INV_X1 U8015 ( .A(n7403), .ZN(n7404) );
  OAI211_X1 U8016 ( .C1(n7407), .C2(n7406), .A(n7405), .B(n7404), .ZN(U2816)
         );
  INV_X1 U8017 ( .A(n7408), .ZN(n7409) );
  AOI22_X1 U8018 ( .A1(n7410), .A2(n7477), .B1(n7475), .B2(n7409), .ZN(n7419)
         );
  AOI22_X1 U8019 ( .A1(EBX_REG_12__SCAN_IN), .A2(n7471), .B1(n7473), .B2(n7411), .ZN(n7412) );
  OAI211_X1 U8020 ( .C1(n7450), .C2(n7413), .A(n7412), .B(n7448), .ZN(n7414)
         );
  AOI221_X1 U8021 ( .B1(n7417), .B2(n7416), .C1(n7415), .C2(
        REIP_REG_12__SCAN_IN), .A(n7414), .ZN(n7418) );
  NAND2_X1 U8022 ( .A1(n7419), .A2(n7418), .ZN(U2815) );
  OAI22_X1 U8023 ( .A1(n4521), .A2(n7450), .B1(n7421), .B2(n7420), .ZN(n7422)
         );
  AOI211_X1 U8024 ( .C1(n7471), .C2(EBX_REG_17__SCAN_IN), .A(n7423), .B(n7422), 
        .ZN(n7430) );
  NAND2_X1 U8025 ( .A1(n7425), .A2(n7424), .ZN(n7432) );
  NAND2_X1 U8026 ( .A1(n7433), .A2(n7432), .ZN(n7428) );
  OAI21_X1 U8027 ( .B1(n7446), .B2(n7427), .A(n7426), .ZN(n7453) );
  AOI22_X1 U8028 ( .A1(n7571), .A2(n7477), .B1(n7428), .B2(n7453), .ZN(n7429)
         );
  OAI211_X1 U8029 ( .C1(n7431), .C2(n7467), .A(n7430), .B(n7429), .ZN(U2810)
         );
  NOR3_X1 U8030 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7433), .A3(n7432), .ZN(n7454) );
  OAI21_X1 U8031 ( .B1(n7450), .B2(n7434), .A(n7448), .ZN(n7435) );
  AOI211_X1 U8032 ( .C1(REIP_REG_18__SCAN_IN), .C2(n7453), .A(n7454), .B(n7435), .ZN(n7442) );
  OAI22_X1 U8033 ( .A1(n7438), .A2(n7437), .B1(n7436), .B2(n7467), .ZN(n7439)
         );
  AOI21_X1 U8034 ( .B1(n7440), .B2(n7475), .A(n7439), .ZN(n7441) );
  OAI211_X1 U8035 ( .C1(n7444), .C2(n7443), .A(n7442), .B(n7441), .ZN(U2809)
         );
  NOR3_X1 U8036 ( .A1(n7446), .A2(REIP_REG_19__SCAN_IN), .A3(n7445), .ZN(n7452) );
  AOI22_X1 U8037 ( .A1(n7447), .A2(n7475), .B1(EBX_REG_19__SCAN_IN), .B2(n7471), .ZN(n7449) );
  OAI211_X1 U8038 ( .C1(n7450), .C2(n4558), .A(n7449), .B(n7448), .ZN(n7451)
         );
  AOI211_X1 U8039 ( .C1(n7574), .C2(n7477), .A(n7452), .B(n7451), .ZN(n7456)
         );
  OAI21_X1 U8040 ( .B1(n7454), .B2(n7453), .A(REIP_REG_19__SCAN_IN), .ZN(n7455) );
  OAI211_X1 U8041 ( .C1(n7467), .C2(n7457), .A(n7456), .B(n7455), .ZN(U2808)
         );
  AOI22_X1 U8042 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n7472), .B1(
        EBX_REG_21__SCAN_IN), .B2(n7471), .ZN(n7458) );
  INV_X1 U8043 ( .A(n7458), .ZN(n7459) );
  AOI221_X1 U8044 ( .B1(n7462), .B2(n7461), .C1(n7460), .C2(
        REIP_REG_21__SCAN_IN), .A(n7459), .ZN(n7466) );
  INV_X1 U8045 ( .A(n7463), .ZN(n7577) );
  AOI22_X1 U8046 ( .A1(n7577), .A2(n7477), .B1(n7464), .B2(n7475), .ZN(n7465)
         );
  OAI211_X1 U8047 ( .C1(n7468), .C2(n7467), .A(n7466), .B(n7465), .ZN(U2806)
         );
  AOI21_X1 U8048 ( .B1(n7470), .B2(n7469), .A(REIP_REG_23__SCAN_IN), .ZN(n7480) );
  AOI22_X1 U8049 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n7472), .B1(
        EBX_REG_23__SCAN_IN), .B2(n7471), .ZN(n7479) );
  AOI222_X1 U8050 ( .A1(n7582), .A2(n7477), .B1(n7476), .B2(n7475), .C1(n7474), 
        .C2(n7473), .ZN(n7478) );
  OAI211_X1 U8051 ( .C1(n7481), .C2(n7480), .A(n7479), .B(n7478), .ZN(U2804)
         );
  OAI21_X1 U8052 ( .B1(n7484), .B2(n7483), .A(n7482), .ZN(U2793) );
  NOR3_X1 U8053 ( .A1(n7486), .A2(n7485), .A3(n3692), .ZN(n7487) );
  NAND2_X1 U8054 ( .A1(n7488), .A2(n7487), .ZN(n7489) );
  OAI21_X1 U8055 ( .B1(n7491), .B2(n7490), .A(n7489), .ZN(U3455) );
  INV_X1 U8056 ( .A(n7492), .ZN(n7514) );
  INV_X1 U8057 ( .A(n7502), .ZN(n7504) );
  NOR3_X1 U8058 ( .A1(n7494), .A2(n7493), .A3(n7557), .ZN(n7498) );
  NAND2_X1 U8059 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7498), .ZN(n7500) );
  INV_X1 U8060 ( .A(n7495), .ZN(n7497) );
  OAI22_X1 U8061 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7498), .B1(n7497), .B2(n7496), .ZN(n7499) );
  OAI211_X1 U8062 ( .C1(n7502), .C2(n7501), .A(n7500), .B(n7499), .ZN(n7503)
         );
  OAI21_X1 U8063 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7504), .A(n7503), 
        .ZN(n7507) );
  AOI222_X1 U8064 ( .A1(n7507), .A2(n7506), .B1(n7507), .B2(n7505), .C1(n7506), 
        .C2(n7505), .ZN(n7511) );
  OAI21_X1 U8065 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n7508), 
        .ZN(n7510) );
  OAI211_X1 U8066 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7511), .A(n7510), .B(n7509), .ZN(n7512) );
  OAI22_X1 U8067 ( .A1(n7535), .A2(n7546), .B1(n7517), .B2(n7516), .ZN(n7518)
         );
  OAI21_X1 U8068 ( .B1(n7520), .B2(n7519), .A(n7518), .ZN(n7541) );
  INV_X1 U8069 ( .A(n7541), .ZN(n7521) );
  AOI21_X1 U8070 ( .B1(READY_N), .B2(n7522), .A(n7521), .ZN(n7538) );
  INV_X1 U8071 ( .A(n7538), .ZN(n7526) );
  INV_X1 U8072 ( .A(n7523), .ZN(n7524) );
  AOI21_X1 U8073 ( .B1(n7526), .B2(n7525), .A(n7524), .ZN(n7530) );
  OAI21_X1 U8074 ( .B1(READY_N), .B2(n7527), .A(n7546), .ZN(n7528) );
  NAND2_X1 U8075 ( .A1(n7541), .A2(n7528), .ZN(n7529) );
  OAI211_X1 U8076 ( .C1(n7536), .C2(n7541), .A(n7530), .B(n7529), .ZN(U3149)
         );
  INV_X1 U8077 ( .A(n7531), .ZN(n7532) );
  OAI211_X1 U8078 ( .C1(n7534), .C2(n7541), .A(n7533), .B(n7532), .ZN(U3453)
         );
  INV_X1 U8079 ( .A(n7535), .ZN(n7547) );
  OR2_X1 U8080 ( .A1(n7537), .A2(n7536), .ZN(n7550) );
  AOI21_X1 U8081 ( .B1(n7538), .B2(n7550), .A(n3966), .ZN(n7540) );
  NOR2_X1 U8082 ( .A1(n7540), .A2(n7539), .ZN(n7545) );
  OAI211_X1 U8083 ( .C1(n7543), .C2(n7542), .A(n3966), .B(n7541), .ZN(n7544)
         );
  OAI211_X1 U8084 ( .C1(n7547), .C2(n7546), .A(n7545), .B(n7544), .ZN(U3148)
         );
  OAI22_X1 U8085 ( .A1(n7551), .A2(n7550), .B1(n7549), .B2(n7548), .ZN(n7552)
         );
  AOI21_X1 U8086 ( .B1(n7554), .B2(n7553), .A(n7552), .ZN(n7555) );
  OAI21_X1 U8087 ( .B1(n7557), .B2(n7556), .A(n7555), .ZN(U3465) );
  AOI211_X1 U8088 ( .C1(HOLD), .C2(STATE_REG_1__SCAN_IN), .A(n7559), .B(n7558), 
        .ZN(n7565) );
  INV_X1 U8089 ( .A(n7560), .ZN(n7563) );
  AOI21_X1 U8090 ( .B1(n7563), .B2(n7562), .A(n7561), .ZN(n7564) );
  OAI21_X1 U8091 ( .B1(n7569), .B2(n7565), .A(n7564), .ZN(U3181) );
  AOI22_X1 U8092 ( .A1(n7569), .A2(n7568), .B1(n7567), .B2(n7566), .ZN(U3473)
         );
  INV_X1 U8093 ( .A(n7570), .ZN(n7581) );
  AOI22_X1 U8094 ( .A1(n7571), .A2(n7581), .B1(n7580), .B2(DATAI_17_), .ZN(
        n7573) );
  AOI22_X1 U8095 ( .A1(n7584), .A2(DATAI_1_), .B1(n7583), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U8096 ( .A1(n7573), .A2(n7572), .ZN(U2874) );
  AOI22_X1 U8097 ( .A1(n7574), .A2(n7581), .B1(n7580), .B2(DATAI_19_), .ZN(
        n7576) );
  AOI22_X1 U8098 ( .A1(n7584), .A2(DATAI_3_), .B1(n7583), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U8099 ( .A1(n7576), .A2(n7575), .ZN(U2872) );
  AOI22_X1 U8100 ( .A1(n7577), .A2(n7581), .B1(n7580), .B2(DATAI_21_), .ZN(
        n7579) );
  AOI22_X1 U8101 ( .A1(n7584), .A2(DATAI_5_), .B1(n7583), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U8102 ( .A1(n7579), .A2(n7578), .ZN(U2870) );
  AOI22_X1 U8103 ( .A1(n7582), .A2(n7581), .B1(n7580), .B2(DATAI_23_), .ZN(
        n7586) );
  AOI22_X1 U8104 ( .A1(n7584), .A2(DATAI_7_), .B1(n7583), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U8105 ( .A1(n7586), .A2(n7585), .ZN(U2868) );
  OAI22_X1 U8106 ( .A1(n7699), .A2(n7597), .B1(n7601), .B2(n7698), .ZN(n7587)
         );
  INV_X1 U8107 ( .A(n7587), .ZN(n7589) );
  AOI22_X1 U8108 ( .A1(n7702), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7605), 
        .B2(n7701), .ZN(n7588) );
  OAI211_X1 U8109 ( .C1(n7705), .C2(n7608), .A(n7589), .B(n7588), .ZN(U3108)
         );
  AOI22_X1 U8110 ( .A1(n7716), .A2(n7605), .B1(n7594), .B2(n7657), .ZN(n7591)
         );
  AOI22_X1 U8111 ( .A1(n7710), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7603), 
        .B2(n7701), .ZN(n7590) );
  OAI211_X1 U8112 ( .C1(n7713), .C2(n7608), .A(n7591), .B(n7590), .ZN(U3100)
         );
  AOI22_X1 U8113 ( .A1(n7715), .A2(n7605), .B1(n7594), .B2(n7714), .ZN(n7593)
         );
  AOI22_X1 U8114 ( .A1(n7717), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7603), 
        .B2(n7716), .ZN(n7592) );
  OAI211_X1 U8115 ( .C1(n7720), .C2(n7608), .A(n7593), .B(n7592), .ZN(U3092)
         );
  AOI22_X1 U8116 ( .A1(n7722), .A2(n7605), .B1(n7594), .B2(n7721), .ZN(n7596)
         );
  AOI22_X1 U8117 ( .A1(n7724), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n7603), 
        .B2(n7723), .ZN(n7595) );
  OAI211_X1 U8118 ( .C1(n7727), .C2(n7608), .A(n7596), .B(n7595), .ZN(U3060)
         );
  OAI22_X1 U8119 ( .A1(n7643), .A2(n7597), .B1(n7601), .B2(n7619), .ZN(n7598)
         );
  INV_X1 U8120 ( .A(n7598), .ZN(n7600) );
  AOI22_X1 U8121 ( .A1(n7733), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n7605), 
        .B2(n7731), .ZN(n7599) );
  OAI211_X1 U8122 ( .C1(n7736), .C2(n7608), .A(n7600), .B(n7599), .ZN(U3044)
         );
  NOR2_X1 U8123 ( .A1(n7601), .A2(n7737), .ZN(n7602) );
  AOI21_X1 U8124 ( .B1(n7742), .B2(n7603), .A(n7602), .ZN(n7607) );
  INV_X1 U8125 ( .A(n7604), .ZN(n7744) );
  AOI22_X1 U8126 ( .A1(n7744), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n7694), 
        .B2(n7605), .ZN(n7606) );
  OAI211_X1 U8127 ( .C1(n7748), .C2(n7608), .A(n7607), .B(n7606), .ZN(U3028)
         );
  OAI22_X1 U8128 ( .A1(n7699), .A2(n7620), .B1(n7625), .B2(n7698), .ZN(n7609)
         );
  INV_X1 U8129 ( .A(n7609), .ZN(n7611) );
  AOI22_X1 U8130 ( .A1(n7702), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7622), 
        .B2(n7701), .ZN(n7610) );
  OAI211_X1 U8131 ( .C1(n7705), .C2(n7631), .A(n7611), .B(n7610), .ZN(U3109)
         );
  AOI22_X1 U8132 ( .A1(n7716), .A2(n7622), .B1(n7616), .B2(n7657), .ZN(n7613)
         );
  AOI22_X1 U8133 ( .A1(n7710), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7628), 
        .B2(n7701), .ZN(n7612) );
  OAI211_X1 U8134 ( .C1(n7713), .C2(n7631), .A(n7613), .B(n7612), .ZN(U3101)
         );
  AOI22_X1 U8135 ( .A1(n7715), .A2(n7622), .B1(n7616), .B2(n7714), .ZN(n7615)
         );
  AOI22_X1 U8136 ( .A1(n7717), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7628), 
        .B2(n7716), .ZN(n7614) );
  OAI211_X1 U8137 ( .C1(n7720), .C2(n7631), .A(n7615), .B(n7614), .ZN(U3093)
         );
  AOI22_X1 U8138 ( .A1(n7722), .A2(n7622), .B1(n7616), .B2(n7721), .ZN(n7618)
         );
  AOI22_X1 U8139 ( .A1(n7724), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n7628), 
        .B2(n7723), .ZN(n7617) );
  OAI211_X1 U8140 ( .C1(n7727), .C2(n7631), .A(n7618), .B(n7617), .ZN(U3061)
         );
  OAI22_X1 U8141 ( .A1(n7643), .A2(n7620), .B1(n7625), .B2(n7619), .ZN(n7621)
         );
  INV_X1 U8142 ( .A(n7621), .ZN(n7624) );
  AOI22_X1 U8143 ( .A1(n7733), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n7622), 
        .B2(n7731), .ZN(n7623) );
  OAI211_X1 U8144 ( .C1(n7736), .C2(n7631), .A(n7624), .B(n7623), .ZN(U3045)
         );
  OAI22_X1 U8145 ( .A1(n7740), .A2(n7626), .B1(n7625), .B2(n7737), .ZN(n7627)
         );
  INV_X1 U8146 ( .A(n7627), .ZN(n7630) );
  AOI22_X1 U8147 ( .A1(n7744), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n7628), 
        .B2(n7742), .ZN(n7629) );
  OAI211_X1 U8148 ( .C1(n7748), .C2(n7631), .A(n7630), .B(n7629), .ZN(U3029)
         );
  OAI22_X1 U8149 ( .A1(n7708), .A2(n7632), .B1(n7646), .B2(n7698), .ZN(n7633)
         );
  INV_X1 U8150 ( .A(n7633), .ZN(n7635) );
  AOI22_X1 U8151 ( .A1(n7702), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7648), 
        .B2(n7676), .ZN(n7634) );
  OAI211_X1 U8152 ( .C1(n7705), .C2(n7652), .A(n7635), .B(n7634), .ZN(U3110)
         );
  AOI22_X1 U8153 ( .A1(n7716), .A2(n7649), .B1(n7642), .B2(n7657), .ZN(n7637)
         );
  AOI22_X1 U8154 ( .A1(n7710), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7648), 
        .B2(n7701), .ZN(n7636) );
  OAI211_X1 U8155 ( .C1(n7713), .C2(n7652), .A(n7637), .B(n7636), .ZN(U3102)
         );
  AOI22_X1 U8156 ( .A1(n7715), .A2(n7649), .B1(n7642), .B2(n7714), .ZN(n7639)
         );
  AOI22_X1 U8157 ( .A1(n7717), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7648), 
        .B2(n7716), .ZN(n7638) );
  OAI211_X1 U8158 ( .C1(n7720), .C2(n7652), .A(n7639), .B(n7638), .ZN(U3094)
         );
  AOI22_X1 U8159 ( .A1(n7723), .A2(n7648), .B1(n7642), .B2(n7721), .ZN(n7641)
         );
  AOI22_X1 U8160 ( .A1(n7724), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n7649), 
        .B2(n7722), .ZN(n7640) );
  OAI211_X1 U8161 ( .C1(n7727), .C2(n7652), .A(n7641), .B(n7640), .ZN(U3062)
         );
  AOI22_X1 U8162 ( .A1(n7731), .A2(n7649), .B1(n7642), .B2(n7728), .ZN(n7645)
         );
  INV_X1 U8163 ( .A(n7643), .ZN(n7732) );
  AOI22_X1 U8164 ( .A1(n7733), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n7648), 
        .B2(n7732), .ZN(n7644) );
  OAI211_X1 U8165 ( .C1(n7736), .C2(n7652), .A(n7645), .B(n7644), .ZN(U3046)
         );
  NOR2_X1 U8166 ( .A1(n7646), .A2(n7737), .ZN(n7647) );
  AOI21_X1 U8167 ( .B1(n7742), .B2(n7648), .A(n7647), .ZN(n7651) );
  AOI22_X1 U8168 ( .A1(n7744), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n7694), 
        .B2(n7649), .ZN(n7650) );
  OAI211_X1 U8169 ( .C1(n7748), .C2(n7652), .A(n7651), .B(n7650), .ZN(U3030)
         );
  OAI22_X1 U8170 ( .A1(n7699), .A2(n7653), .B1(n7667), .B2(n7698), .ZN(n7654)
         );
  INV_X1 U8171 ( .A(n7654), .ZN(n7656) );
  AOI22_X1 U8172 ( .A1(n7702), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7670), 
        .B2(n7701), .ZN(n7655) );
  OAI211_X1 U8173 ( .C1(n7705), .C2(n7673), .A(n7656), .B(n7655), .ZN(U3112)
         );
  AOI22_X1 U8174 ( .A1(n7716), .A2(n7670), .B1(n7664), .B2(n7657), .ZN(n7659)
         );
  AOI22_X1 U8175 ( .A1(n7710), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7669), 
        .B2(n7701), .ZN(n7658) );
  OAI211_X1 U8176 ( .C1(n7713), .C2(n7673), .A(n7659), .B(n7658), .ZN(U3104)
         );
  AOI22_X1 U8177 ( .A1(n7716), .A2(n7669), .B1(n7664), .B2(n7714), .ZN(n7661)
         );
  AOI22_X1 U8178 ( .A1(n7717), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7715), 
        .B2(n7670), .ZN(n7660) );
  OAI211_X1 U8179 ( .C1(n7720), .C2(n7673), .A(n7661), .B(n7660), .ZN(U3096)
         );
  AOI22_X1 U8180 ( .A1(n7722), .A2(n7670), .B1(n7664), .B2(n7721), .ZN(n7663)
         );
  AOI22_X1 U8181 ( .A1(n7724), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n7669), 
        .B2(n7723), .ZN(n7662) );
  OAI211_X1 U8182 ( .C1(n7727), .C2(n7673), .A(n7663), .B(n7662), .ZN(U3064)
         );
  AOI22_X1 U8183 ( .A1(n7731), .A2(n7670), .B1(n7664), .B2(n7728), .ZN(n7666)
         );
  AOI22_X1 U8184 ( .A1(n7733), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n7669), 
        .B2(n7732), .ZN(n7665) );
  OAI211_X1 U8185 ( .C1(n7736), .C2(n7673), .A(n7666), .B(n7665), .ZN(U3048)
         );
  NOR2_X1 U8186 ( .A1(n7667), .A2(n7737), .ZN(n7668) );
  AOI21_X1 U8187 ( .B1(n7742), .B2(n7669), .A(n7668), .ZN(n7672) );
  AOI22_X1 U8188 ( .A1(n7744), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n7694), 
        .B2(n7670), .ZN(n7671) );
  OAI211_X1 U8189 ( .C1(n7748), .C2(n7673), .A(n7672), .B(n7671), .ZN(U3032)
         );
  OAI22_X1 U8190 ( .A1(n7708), .A2(n7674), .B1(n7679), .B2(n7698), .ZN(n7675)
         );
  INV_X1 U8191 ( .A(n7675), .ZN(n7678) );
  AOI22_X1 U8192 ( .A1(n7702), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7692), 
        .B2(n7676), .ZN(n7677) );
  OAI211_X1 U8193 ( .C1(n7705), .C2(n7697), .A(n7678), .B(n7677), .ZN(U3114)
         );
  OAI22_X1 U8194 ( .A1(n7708), .A2(n7680), .B1(n7679), .B2(n7706), .ZN(n7681)
         );
  INV_X1 U8195 ( .A(n7681), .ZN(n7683) );
  AOI22_X1 U8196 ( .A1(n7710), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7693), 
        .B2(n7716), .ZN(n7682) );
  OAI211_X1 U8197 ( .C1(n7713), .C2(n7697), .A(n7683), .B(n7682), .ZN(U3106)
         );
  AOI22_X1 U8198 ( .A1(n7715), .A2(n7693), .B1(n7691), .B2(n7714), .ZN(n7685)
         );
  AOI22_X1 U8199 ( .A1(n7717), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7692), 
        .B2(n7716), .ZN(n7684) );
  OAI211_X1 U8200 ( .C1(n7720), .C2(n7697), .A(n7685), .B(n7684), .ZN(U3098)
         );
  AOI22_X1 U8201 ( .A1(n7722), .A2(n7693), .B1(n7691), .B2(n7721), .ZN(n7687)
         );
  AOI22_X1 U8202 ( .A1(n7724), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n7692), 
        .B2(n7723), .ZN(n7686) );
  OAI211_X1 U8203 ( .C1(n7727), .C2(n7697), .A(n7687), .B(n7686), .ZN(U3066)
         );
  AOI22_X1 U8204 ( .A1(n7731), .A2(n7693), .B1(n7691), .B2(n7728), .ZN(n7689)
         );
  AOI22_X1 U8205 ( .A1(n7733), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n7692), 
        .B2(n7732), .ZN(n7688) );
  OAI211_X1 U8206 ( .C1(n7736), .C2(n7697), .A(n7689), .B(n7688), .ZN(U3050)
         );
  INV_X1 U8207 ( .A(n7737), .ZN(n7690) );
  AOI22_X1 U8208 ( .A1(n7742), .A2(n7692), .B1(n7691), .B2(n7690), .ZN(n7696)
         );
  AOI22_X1 U8209 ( .A1(n7744), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n7694), 
        .B2(n7693), .ZN(n7695) );
  OAI211_X1 U8210 ( .C1(n7748), .C2(n7697), .A(n7696), .B(n7695), .ZN(U3034)
         );
  OAI22_X1 U8211 ( .A1(n7699), .A2(n7707), .B1(n7738), .B2(n7698), .ZN(n7700)
         );
  INV_X1 U8212 ( .A(n7700), .ZN(n7704) );
  AOI22_X1 U8213 ( .A1(n7702), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7730), 
        .B2(n7701), .ZN(n7703) );
  OAI211_X1 U8214 ( .C1(n7705), .C2(n7747), .A(n7704), .B(n7703), .ZN(U3115)
         );
  OAI22_X1 U8215 ( .A1(n7708), .A2(n7707), .B1(n7738), .B2(n7706), .ZN(n7709)
         );
  INV_X1 U8216 ( .A(n7709), .ZN(n7712) );
  AOI22_X1 U8217 ( .A1(n7710), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7730), 
        .B2(n7716), .ZN(n7711) );
  OAI211_X1 U8218 ( .C1(n7713), .C2(n7747), .A(n7712), .B(n7711), .ZN(U3107)
         );
  AOI22_X1 U8219 ( .A1(n7715), .A2(n7730), .B1(n7729), .B2(n7714), .ZN(n7719)
         );
  AOI22_X1 U8220 ( .A1(n7717), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7743), 
        .B2(n7716), .ZN(n7718) );
  OAI211_X1 U8221 ( .C1(n7720), .C2(n7747), .A(n7719), .B(n7718), .ZN(U3099)
         );
  AOI22_X1 U8222 ( .A1(n7722), .A2(n7730), .B1(n7729), .B2(n7721), .ZN(n7726)
         );
  AOI22_X1 U8223 ( .A1(n7724), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7743), 
        .B2(n7723), .ZN(n7725) );
  OAI211_X1 U8224 ( .C1(n7727), .C2(n7747), .A(n7726), .B(n7725), .ZN(U3067)
         );
  AOI22_X1 U8225 ( .A1(n7731), .A2(n7730), .B1(n7729), .B2(n7728), .ZN(n7735)
         );
  AOI22_X1 U8226 ( .A1(n7733), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n7743), 
        .B2(n7732), .ZN(n7734) );
  OAI211_X1 U8227 ( .C1(n7736), .C2(n7747), .A(n7735), .B(n7734), .ZN(U3051)
         );
  OAI22_X1 U8228 ( .A1(n7740), .A2(n7739), .B1(n7738), .B2(n7737), .ZN(n7741)
         );
  INV_X1 U8229 ( .A(n7741), .ZN(n7746) );
  AOI22_X1 U8230 ( .A1(n7744), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n7743), 
        .B2(n7742), .ZN(n7745) );
  OAI211_X1 U8231 ( .C1(n7748), .C2(n7747), .A(n7746), .B(n7745), .ZN(U3035)
         );
  OR2_X1 U3864 ( .A1(n6582), .A2(n7482), .ZN(n3685) );
  NAND2_X1 U3779 ( .A1(n6142), .A2(n6143), .ZN(n4817) );
  CLKBUF_X1 U3878 ( .A(n3905), .Z(n5225) );
  INV_X1 U3892 ( .A(n6018), .ZN(n6113) );
  CLKBUF_X1 U4298 ( .A(n7172), .Z(n7193) );
  CLKBUF_X1 U5425 ( .A(n6431), .Z(n6432) );
  CLKBUF_X1 U5426 ( .A(n6530), .Z(n3693) );
  INV_X2 U5488 ( .A(n7517), .ZN(n7182) );
endmodule

